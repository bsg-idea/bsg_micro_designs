

module top
(
  clk_i,
  reset_i,
  ready_o,
  v_i,
  data_i,
  v_o,
  data_o,
  ready_i
);

  input [63:0] data_i;
  output [499:0] v_o;
  output [31999:0] data_o;
  input [499:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output ready_o;

  bsg_front_side_bus_hop_in
  wrapper
  (
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .ready_i(ready_i),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p64_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [63:0] w_data_i;
  input [0:0] r_addr_i;
  output [63:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [63:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [127:0] mem;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[127] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[126] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[125] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[124] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[123] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[122] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[121] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[120] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[119] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[118] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[117] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[116] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[115] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[114] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[113] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[112] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[111] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[110] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[109] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[108] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[107] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[106] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[105] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[104] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[103] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[102] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[101] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[100] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[99] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[98] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[97] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[96] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[95] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[94] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[93] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[92] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[91] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[90] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[89] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[88] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[87] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[86] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[85] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[84] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[83] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[82] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[81] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[80] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[79] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[78] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[77] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[76] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[75] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[74] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[73] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[72] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[71] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[70] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[69] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[68] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[67] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[66] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[65] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[64] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[127:64] } <= { w_data_i[63:0] };
    end 
    if(N7) begin
      { mem[63:0] } <= { w_data_i[63:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p64_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [63:0] w_data_i;
  input [0:0] r_addr_i;
  output [63:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [63:0] r_data_o;

  bsg_mem_1r1w_synth_width_p64_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p64
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [63:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [63:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p64_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_front_side_bus_hop_in
(
  clk_i,
  reset_i,
  ready_o,
  v_i,
  data_i,
  v_o,
  data_o,
  ready_i
);

  input [63:0] data_i;
  output [499:0] v_o;
  output [31999:0] data_o;
  input [499:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output ready_o;
  wire [499:0] v_o,sent_n;
  wire [31999:0] data_o;
  wire ready_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
  N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,
  N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,
  N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,
  N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,
  N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,
  N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,
  N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,
  N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,
  N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
  N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,
  N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,
  N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,fifo_v,fifo_yumi,
  N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,
  N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,
  N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,
  N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,
  N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,
  N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,
  N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,
  N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,
  N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,
  N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,
  N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,
  N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,
  N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,
  N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,
  N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,
  N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,
  N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,
  N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,
  N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,
  N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,
  N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,
  N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,
  N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,
  N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,
  N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,
  N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,
  N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
  N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,
  N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,
  N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,
  N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,
  N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,
  N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,
  N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,
  N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,
  N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,
  N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,
  N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,
  N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,
  N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
  N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,
  N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,
  N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,
  N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,
  N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,
  N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,
  N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,
  N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,
  N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,
  N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,
  N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,
  N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,
  N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,
  N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,
  N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,
  N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,
  N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,
  N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,
  N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,
  N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,
  N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,
  N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,
  N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,
  N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,
  N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,
  N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,
  N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,
  N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,
  N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,
  N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,
  N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,
  N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,
  N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,
  N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,
  N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,
  N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,
  N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,
  N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,
  N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,
  N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,
  N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,
  N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,
  N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,
  N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,
  N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,
  N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,
  N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,
  N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,
  N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,
  N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,
  N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,
  N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,
  N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,
  N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,
  N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,
  N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,
  N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,
  N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,
  N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,
  N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,
  N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,
  N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,
  N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,
  N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,
  N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,
  N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,
  N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,
  N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,
  N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,
  N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,
  N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,
  N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,
  N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,
  N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,
  N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,
  N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,
  N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,
  N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,
  N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,
  N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,
  N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,
  N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,
  N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,
  N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,
  N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,
  N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,
  N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,
  N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,
  N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,
  N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,
  N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,
  N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,
  N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,
  N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,
  N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,
  N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,
  N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,
  N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,
  N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,
  N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,
  N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,
  N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,
  N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,
  N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,
  N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,
  N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,
  N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,
  N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,
  N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
  N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,
  N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,
  N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,
  N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,
  N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,
  N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,
  N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,
  N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,
  N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,
  N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,
  N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,
  N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,
  N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,
  N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,
  N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,
  N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,
  N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,
  N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,
  N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,
  N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,
  N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,
  N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,
  N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,
  N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,
  N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,
  N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,
  N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,
  N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,
  N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,
  N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,
  N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,
  N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,
  N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,
  N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,
  N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,
  N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,
  N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,
  N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,
  N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,
  N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,
  N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,
  N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,
  N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,
  N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,
  N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,
  N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,
  N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,
  N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,
  N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,
  N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,
  N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,
  N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,
  N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,
  N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,
  N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,
  N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,
  N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,
  N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,
  N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,
  N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,
  N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,
  N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,
  N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,
  N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,
  N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,
  N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,
  N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,
  N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,
  N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,
  N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,
  N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,
  N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,
  N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,
  N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,
  N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,
  N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,
  N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,
  N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,
  N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,
  N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,
  N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,
  N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,
  N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,
  N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,
  N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,
  N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,
  N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,
  N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,
  N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,
  N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,
  N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,
  N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,
  N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,
  N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,
  N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,
  N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,
  N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,
  N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,
  N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,
  N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,
  N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,
  N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,
  N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,
  N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,
  N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,
  N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,
  N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,
  N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,
  N4927,N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,
  N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,
  N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,
  N4967,N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,
  N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,
  N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,
  N5007,N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,
  N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,
  N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,
  N5047,N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,
  N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,
  N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,
  N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,
  N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,
  N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,
  N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,
  N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,
  N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,
  N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,
  N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,
  N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,
  N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,
  N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,
  N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,
  N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,
  N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,
  N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,
  N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,
  N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,
  N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,
  N5327,N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,
  N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,
  N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,
  N5367,N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,
  N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,
  N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,
  N5407,N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,
  N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,
  N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,
  N5447,N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,
  N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,
  N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,
  N5487,N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,
  N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,
  N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,
  N5527,N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,
  N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,
  N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,
  N5567,N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,
  N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,
  N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,
  N5607,N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,
  N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,
  N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,
  N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,
  N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,
  N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,
  N5687,N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,
  N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,
  N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,
  N5727,N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,
  N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,
  N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,
  N5767,N5768,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,
  N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,
  N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,
  N5807,N5808,N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,
  N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,
  N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,
  N5847,N5848,N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,
  N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,
  N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,
  N5887,N5888,N5889,N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,
  N5900,N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,
  N5914,N5915,N5916,N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,
  N5927,N5928,N5929,N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,
  N5940,N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,
  N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,
  N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,
  N5980,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,
  N5994,N5995,N5996,N5997;
  reg [499:0] sent_r;
  assign data_o[127] = data_o[63];
  assign data_o[191] = data_o[63];
  assign data_o[255] = data_o[63];
  assign data_o[319] = data_o[63];
  assign data_o[383] = data_o[63];
  assign data_o[447] = data_o[63];
  assign data_o[511] = data_o[63];
  assign data_o[575] = data_o[63];
  assign data_o[639] = data_o[63];
  assign data_o[703] = data_o[63];
  assign data_o[767] = data_o[63];
  assign data_o[831] = data_o[63];
  assign data_o[895] = data_o[63];
  assign data_o[959] = data_o[63];
  assign data_o[1023] = data_o[63];
  assign data_o[1087] = data_o[63];
  assign data_o[1151] = data_o[63];
  assign data_o[1215] = data_o[63];
  assign data_o[1279] = data_o[63];
  assign data_o[1343] = data_o[63];
  assign data_o[1407] = data_o[63];
  assign data_o[1471] = data_o[63];
  assign data_o[1535] = data_o[63];
  assign data_o[1599] = data_o[63];
  assign data_o[1663] = data_o[63];
  assign data_o[1727] = data_o[63];
  assign data_o[1791] = data_o[63];
  assign data_o[1855] = data_o[63];
  assign data_o[1919] = data_o[63];
  assign data_o[1983] = data_o[63];
  assign data_o[2047] = data_o[63];
  assign data_o[2111] = data_o[63];
  assign data_o[2175] = data_o[63];
  assign data_o[2239] = data_o[63];
  assign data_o[2303] = data_o[63];
  assign data_o[2367] = data_o[63];
  assign data_o[2431] = data_o[63];
  assign data_o[2495] = data_o[63];
  assign data_o[2559] = data_o[63];
  assign data_o[2623] = data_o[63];
  assign data_o[2687] = data_o[63];
  assign data_o[2751] = data_o[63];
  assign data_o[2815] = data_o[63];
  assign data_o[2879] = data_o[63];
  assign data_o[2943] = data_o[63];
  assign data_o[3007] = data_o[63];
  assign data_o[3071] = data_o[63];
  assign data_o[3135] = data_o[63];
  assign data_o[3199] = data_o[63];
  assign data_o[3263] = data_o[63];
  assign data_o[3327] = data_o[63];
  assign data_o[3391] = data_o[63];
  assign data_o[3455] = data_o[63];
  assign data_o[3519] = data_o[63];
  assign data_o[3583] = data_o[63];
  assign data_o[3647] = data_o[63];
  assign data_o[3711] = data_o[63];
  assign data_o[3775] = data_o[63];
  assign data_o[3839] = data_o[63];
  assign data_o[3903] = data_o[63];
  assign data_o[3967] = data_o[63];
  assign data_o[4031] = data_o[63];
  assign data_o[4095] = data_o[63];
  assign data_o[4159] = data_o[63];
  assign data_o[4223] = data_o[63];
  assign data_o[4287] = data_o[63];
  assign data_o[4351] = data_o[63];
  assign data_o[4415] = data_o[63];
  assign data_o[4479] = data_o[63];
  assign data_o[4543] = data_o[63];
  assign data_o[4607] = data_o[63];
  assign data_o[4671] = data_o[63];
  assign data_o[4735] = data_o[63];
  assign data_o[4799] = data_o[63];
  assign data_o[4863] = data_o[63];
  assign data_o[4927] = data_o[63];
  assign data_o[4991] = data_o[63];
  assign data_o[5055] = data_o[63];
  assign data_o[5119] = data_o[63];
  assign data_o[5183] = data_o[63];
  assign data_o[5247] = data_o[63];
  assign data_o[5311] = data_o[63];
  assign data_o[5375] = data_o[63];
  assign data_o[5439] = data_o[63];
  assign data_o[5503] = data_o[63];
  assign data_o[5567] = data_o[63];
  assign data_o[5631] = data_o[63];
  assign data_o[5695] = data_o[63];
  assign data_o[5759] = data_o[63];
  assign data_o[5823] = data_o[63];
  assign data_o[5887] = data_o[63];
  assign data_o[5951] = data_o[63];
  assign data_o[6015] = data_o[63];
  assign data_o[6079] = data_o[63];
  assign data_o[6143] = data_o[63];
  assign data_o[6207] = data_o[63];
  assign data_o[6271] = data_o[63];
  assign data_o[6335] = data_o[63];
  assign data_o[6399] = data_o[63];
  assign data_o[6463] = data_o[63];
  assign data_o[6527] = data_o[63];
  assign data_o[6591] = data_o[63];
  assign data_o[6655] = data_o[63];
  assign data_o[6719] = data_o[63];
  assign data_o[6783] = data_o[63];
  assign data_o[6847] = data_o[63];
  assign data_o[6911] = data_o[63];
  assign data_o[6975] = data_o[63];
  assign data_o[7039] = data_o[63];
  assign data_o[7103] = data_o[63];
  assign data_o[7167] = data_o[63];
  assign data_o[7231] = data_o[63];
  assign data_o[7295] = data_o[63];
  assign data_o[7359] = data_o[63];
  assign data_o[7423] = data_o[63];
  assign data_o[7487] = data_o[63];
  assign data_o[7551] = data_o[63];
  assign data_o[7615] = data_o[63];
  assign data_o[7679] = data_o[63];
  assign data_o[7743] = data_o[63];
  assign data_o[7807] = data_o[63];
  assign data_o[7871] = data_o[63];
  assign data_o[7935] = data_o[63];
  assign data_o[7999] = data_o[63];
  assign data_o[8063] = data_o[63];
  assign data_o[8127] = data_o[63];
  assign data_o[8191] = data_o[63];
  assign data_o[8255] = data_o[63];
  assign data_o[8319] = data_o[63];
  assign data_o[8383] = data_o[63];
  assign data_o[8447] = data_o[63];
  assign data_o[8511] = data_o[63];
  assign data_o[8575] = data_o[63];
  assign data_o[8639] = data_o[63];
  assign data_o[8703] = data_o[63];
  assign data_o[8767] = data_o[63];
  assign data_o[8831] = data_o[63];
  assign data_o[8895] = data_o[63];
  assign data_o[8959] = data_o[63];
  assign data_o[9023] = data_o[63];
  assign data_o[9087] = data_o[63];
  assign data_o[9151] = data_o[63];
  assign data_o[9215] = data_o[63];
  assign data_o[9279] = data_o[63];
  assign data_o[9343] = data_o[63];
  assign data_o[9407] = data_o[63];
  assign data_o[9471] = data_o[63];
  assign data_o[9535] = data_o[63];
  assign data_o[9599] = data_o[63];
  assign data_o[9663] = data_o[63];
  assign data_o[9727] = data_o[63];
  assign data_o[9791] = data_o[63];
  assign data_o[9855] = data_o[63];
  assign data_o[9919] = data_o[63];
  assign data_o[9983] = data_o[63];
  assign data_o[10047] = data_o[63];
  assign data_o[10111] = data_o[63];
  assign data_o[10175] = data_o[63];
  assign data_o[10239] = data_o[63];
  assign data_o[10303] = data_o[63];
  assign data_o[10367] = data_o[63];
  assign data_o[10431] = data_o[63];
  assign data_o[10495] = data_o[63];
  assign data_o[10559] = data_o[63];
  assign data_o[10623] = data_o[63];
  assign data_o[10687] = data_o[63];
  assign data_o[10751] = data_o[63];
  assign data_o[10815] = data_o[63];
  assign data_o[10879] = data_o[63];
  assign data_o[10943] = data_o[63];
  assign data_o[11007] = data_o[63];
  assign data_o[11071] = data_o[63];
  assign data_o[11135] = data_o[63];
  assign data_o[11199] = data_o[63];
  assign data_o[11263] = data_o[63];
  assign data_o[11327] = data_o[63];
  assign data_o[11391] = data_o[63];
  assign data_o[11455] = data_o[63];
  assign data_o[11519] = data_o[63];
  assign data_o[11583] = data_o[63];
  assign data_o[11647] = data_o[63];
  assign data_o[11711] = data_o[63];
  assign data_o[11775] = data_o[63];
  assign data_o[11839] = data_o[63];
  assign data_o[11903] = data_o[63];
  assign data_o[11967] = data_o[63];
  assign data_o[12031] = data_o[63];
  assign data_o[12095] = data_o[63];
  assign data_o[12159] = data_o[63];
  assign data_o[12223] = data_o[63];
  assign data_o[12287] = data_o[63];
  assign data_o[12351] = data_o[63];
  assign data_o[12415] = data_o[63];
  assign data_o[12479] = data_o[63];
  assign data_o[12543] = data_o[63];
  assign data_o[12607] = data_o[63];
  assign data_o[12671] = data_o[63];
  assign data_o[12735] = data_o[63];
  assign data_o[12799] = data_o[63];
  assign data_o[12863] = data_o[63];
  assign data_o[12927] = data_o[63];
  assign data_o[12991] = data_o[63];
  assign data_o[13055] = data_o[63];
  assign data_o[13119] = data_o[63];
  assign data_o[13183] = data_o[63];
  assign data_o[13247] = data_o[63];
  assign data_o[13311] = data_o[63];
  assign data_o[13375] = data_o[63];
  assign data_o[13439] = data_o[63];
  assign data_o[13503] = data_o[63];
  assign data_o[13567] = data_o[63];
  assign data_o[13631] = data_o[63];
  assign data_o[13695] = data_o[63];
  assign data_o[13759] = data_o[63];
  assign data_o[13823] = data_o[63];
  assign data_o[13887] = data_o[63];
  assign data_o[13951] = data_o[63];
  assign data_o[14015] = data_o[63];
  assign data_o[14079] = data_o[63];
  assign data_o[14143] = data_o[63];
  assign data_o[14207] = data_o[63];
  assign data_o[14271] = data_o[63];
  assign data_o[14335] = data_o[63];
  assign data_o[14399] = data_o[63];
  assign data_o[14463] = data_o[63];
  assign data_o[14527] = data_o[63];
  assign data_o[14591] = data_o[63];
  assign data_o[14655] = data_o[63];
  assign data_o[14719] = data_o[63];
  assign data_o[14783] = data_o[63];
  assign data_o[14847] = data_o[63];
  assign data_o[14911] = data_o[63];
  assign data_o[14975] = data_o[63];
  assign data_o[15039] = data_o[63];
  assign data_o[15103] = data_o[63];
  assign data_o[15167] = data_o[63];
  assign data_o[15231] = data_o[63];
  assign data_o[15295] = data_o[63];
  assign data_o[15359] = data_o[63];
  assign data_o[15423] = data_o[63];
  assign data_o[15487] = data_o[63];
  assign data_o[15551] = data_o[63];
  assign data_o[15615] = data_o[63];
  assign data_o[15679] = data_o[63];
  assign data_o[15743] = data_o[63];
  assign data_o[15807] = data_o[63];
  assign data_o[15871] = data_o[63];
  assign data_o[15935] = data_o[63];
  assign data_o[15999] = data_o[63];
  assign data_o[16063] = data_o[63];
  assign data_o[16127] = data_o[63];
  assign data_o[16191] = data_o[63];
  assign data_o[16255] = data_o[63];
  assign data_o[16319] = data_o[63];
  assign data_o[16383] = data_o[63];
  assign data_o[16447] = data_o[63];
  assign data_o[16511] = data_o[63];
  assign data_o[16575] = data_o[63];
  assign data_o[16639] = data_o[63];
  assign data_o[16703] = data_o[63];
  assign data_o[16767] = data_o[63];
  assign data_o[16831] = data_o[63];
  assign data_o[16895] = data_o[63];
  assign data_o[16959] = data_o[63];
  assign data_o[17023] = data_o[63];
  assign data_o[17087] = data_o[63];
  assign data_o[17151] = data_o[63];
  assign data_o[17215] = data_o[63];
  assign data_o[17279] = data_o[63];
  assign data_o[17343] = data_o[63];
  assign data_o[17407] = data_o[63];
  assign data_o[17471] = data_o[63];
  assign data_o[17535] = data_o[63];
  assign data_o[17599] = data_o[63];
  assign data_o[17663] = data_o[63];
  assign data_o[17727] = data_o[63];
  assign data_o[17791] = data_o[63];
  assign data_o[17855] = data_o[63];
  assign data_o[17919] = data_o[63];
  assign data_o[17983] = data_o[63];
  assign data_o[18047] = data_o[63];
  assign data_o[18111] = data_o[63];
  assign data_o[18175] = data_o[63];
  assign data_o[18239] = data_o[63];
  assign data_o[18303] = data_o[63];
  assign data_o[18367] = data_o[63];
  assign data_o[18431] = data_o[63];
  assign data_o[18495] = data_o[63];
  assign data_o[18559] = data_o[63];
  assign data_o[18623] = data_o[63];
  assign data_o[18687] = data_o[63];
  assign data_o[18751] = data_o[63];
  assign data_o[18815] = data_o[63];
  assign data_o[18879] = data_o[63];
  assign data_o[18943] = data_o[63];
  assign data_o[19007] = data_o[63];
  assign data_o[19071] = data_o[63];
  assign data_o[19135] = data_o[63];
  assign data_o[19199] = data_o[63];
  assign data_o[19263] = data_o[63];
  assign data_o[19327] = data_o[63];
  assign data_o[19391] = data_o[63];
  assign data_o[19455] = data_o[63];
  assign data_o[19519] = data_o[63];
  assign data_o[19583] = data_o[63];
  assign data_o[19647] = data_o[63];
  assign data_o[19711] = data_o[63];
  assign data_o[19775] = data_o[63];
  assign data_o[19839] = data_o[63];
  assign data_o[19903] = data_o[63];
  assign data_o[19967] = data_o[63];
  assign data_o[20031] = data_o[63];
  assign data_o[20095] = data_o[63];
  assign data_o[20159] = data_o[63];
  assign data_o[20223] = data_o[63];
  assign data_o[20287] = data_o[63];
  assign data_o[20351] = data_o[63];
  assign data_o[20415] = data_o[63];
  assign data_o[20479] = data_o[63];
  assign data_o[20543] = data_o[63];
  assign data_o[20607] = data_o[63];
  assign data_o[20671] = data_o[63];
  assign data_o[20735] = data_o[63];
  assign data_o[20799] = data_o[63];
  assign data_o[20863] = data_o[63];
  assign data_o[20927] = data_o[63];
  assign data_o[20991] = data_o[63];
  assign data_o[21055] = data_o[63];
  assign data_o[21119] = data_o[63];
  assign data_o[21183] = data_o[63];
  assign data_o[21247] = data_o[63];
  assign data_o[21311] = data_o[63];
  assign data_o[21375] = data_o[63];
  assign data_o[21439] = data_o[63];
  assign data_o[21503] = data_o[63];
  assign data_o[21567] = data_o[63];
  assign data_o[21631] = data_o[63];
  assign data_o[21695] = data_o[63];
  assign data_o[21759] = data_o[63];
  assign data_o[21823] = data_o[63];
  assign data_o[21887] = data_o[63];
  assign data_o[21951] = data_o[63];
  assign data_o[22015] = data_o[63];
  assign data_o[22079] = data_o[63];
  assign data_o[22143] = data_o[63];
  assign data_o[22207] = data_o[63];
  assign data_o[22271] = data_o[63];
  assign data_o[22335] = data_o[63];
  assign data_o[22399] = data_o[63];
  assign data_o[22463] = data_o[63];
  assign data_o[22527] = data_o[63];
  assign data_o[22591] = data_o[63];
  assign data_o[22655] = data_o[63];
  assign data_o[22719] = data_o[63];
  assign data_o[22783] = data_o[63];
  assign data_o[22847] = data_o[63];
  assign data_o[22911] = data_o[63];
  assign data_o[22975] = data_o[63];
  assign data_o[23039] = data_o[63];
  assign data_o[23103] = data_o[63];
  assign data_o[23167] = data_o[63];
  assign data_o[23231] = data_o[63];
  assign data_o[23295] = data_o[63];
  assign data_o[23359] = data_o[63];
  assign data_o[23423] = data_o[63];
  assign data_o[23487] = data_o[63];
  assign data_o[23551] = data_o[63];
  assign data_o[23615] = data_o[63];
  assign data_o[23679] = data_o[63];
  assign data_o[23743] = data_o[63];
  assign data_o[23807] = data_o[63];
  assign data_o[23871] = data_o[63];
  assign data_o[23935] = data_o[63];
  assign data_o[23999] = data_o[63];
  assign data_o[24063] = data_o[63];
  assign data_o[24127] = data_o[63];
  assign data_o[24191] = data_o[63];
  assign data_o[24255] = data_o[63];
  assign data_o[24319] = data_o[63];
  assign data_o[24383] = data_o[63];
  assign data_o[24447] = data_o[63];
  assign data_o[24511] = data_o[63];
  assign data_o[24575] = data_o[63];
  assign data_o[24639] = data_o[63];
  assign data_o[24703] = data_o[63];
  assign data_o[24767] = data_o[63];
  assign data_o[24831] = data_o[63];
  assign data_o[24895] = data_o[63];
  assign data_o[24959] = data_o[63];
  assign data_o[25023] = data_o[63];
  assign data_o[25087] = data_o[63];
  assign data_o[25151] = data_o[63];
  assign data_o[25215] = data_o[63];
  assign data_o[25279] = data_o[63];
  assign data_o[25343] = data_o[63];
  assign data_o[25407] = data_o[63];
  assign data_o[25471] = data_o[63];
  assign data_o[25535] = data_o[63];
  assign data_o[25599] = data_o[63];
  assign data_o[25663] = data_o[63];
  assign data_o[25727] = data_o[63];
  assign data_o[25791] = data_o[63];
  assign data_o[25855] = data_o[63];
  assign data_o[25919] = data_o[63];
  assign data_o[25983] = data_o[63];
  assign data_o[26047] = data_o[63];
  assign data_o[26111] = data_o[63];
  assign data_o[26175] = data_o[63];
  assign data_o[26239] = data_o[63];
  assign data_o[26303] = data_o[63];
  assign data_o[26367] = data_o[63];
  assign data_o[26431] = data_o[63];
  assign data_o[26495] = data_o[63];
  assign data_o[26559] = data_o[63];
  assign data_o[26623] = data_o[63];
  assign data_o[26687] = data_o[63];
  assign data_o[26751] = data_o[63];
  assign data_o[26815] = data_o[63];
  assign data_o[26879] = data_o[63];
  assign data_o[26943] = data_o[63];
  assign data_o[27007] = data_o[63];
  assign data_o[27071] = data_o[63];
  assign data_o[27135] = data_o[63];
  assign data_o[27199] = data_o[63];
  assign data_o[27263] = data_o[63];
  assign data_o[27327] = data_o[63];
  assign data_o[27391] = data_o[63];
  assign data_o[27455] = data_o[63];
  assign data_o[27519] = data_o[63];
  assign data_o[27583] = data_o[63];
  assign data_o[27647] = data_o[63];
  assign data_o[27711] = data_o[63];
  assign data_o[27775] = data_o[63];
  assign data_o[27839] = data_o[63];
  assign data_o[27903] = data_o[63];
  assign data_o[27967] = data_o[63];
  assign data_o[28031] = data_o[63];
  assign data_o[28095] = data_o[63];
  assign data_o[28159] = data_o[63];
  assign data_o[28223] = data_o[63];
  assign data_o[28287] = data_o[63];
  assign data_o[28351] = data_o[63];
  assign data_o[28415] = data_o[63];
  assign data_o[28479] = data_o[63];
  assign data_o[28543] = data_o[63];
  assign data_o[28607] = data_o[63];
  assign data_o[28671] = data_o[63];
  assign data_o[28735] = data_o[63];
  assign data_o[28799] = data_o[63];
  assign data_o[28863] = data_o[63];
  assign data_o[28927] = data_o[63];
  assign data_o[28991] = data_o[63];
  assign data_o[29055] = data_o[63];
  assign data_o[29119] = data_o[63];
  assign data_o[29183] = data_o[63];
  assign data_o[29247] = data_o[63];
  assign data_o[29311] = data_o[63];
  assign data_o[29375] = data_o[63];
  assign data_o[29439] = data_o[63];
  assign data_o[29503] = data_o[63];
  assign data_o[29567] = data_o[63];
  assign data_o[29631] = data_o[63];
  assign data_o[29695] = data_o[63];
  assign data_o[29759] = data_o[63];
  assign data_o[29823] = data_o[63];
  assign data_o[29887] = data_o[63];
  assign data_o[29951] = data_o[63];
  assign data_o[30015] = data_o[63];
  assign data_o[30079] = data_o[63];
  assign data_o[30143] = data_o[63];
  assign data_o[30207] = data_o[63];
  assign data_o[30271] = data_o[63];
  assign data_o[30335] = data_o[63];
  assign data_o[30399] = data_o[63];
  assign data_o[30463] = data_o[63];
  assign data_o[30527] = data_o[63];
  assign data_o[30591] = data_o[63];
  assign data_o[30655] = data_o[63];
  assign data_o[30719] = data_o[63];
  assign data_o[30783] = data_o[63];
  assign data_o[30847] = data_o[63];
  assign data_o[30911] = data_o[63];
  assign data_o[30975] = data_o[63];
  assign data_o[31039] = data_o[63];
  assign data_o[31103] = data_o[63];
  assign data_o[31167] = data_o[63];
  assign data_o[31231] = data_o[63];
  assign data_o[31295] = data_o[63];
  assign data_o[31359] = data_o[63];
  assign data_o[31423] = data_o[63];
  assign data_o[31487] = data_o[63];
  assign data_o[31551] = data_o[63];
  assign data_o[31615] = data_o[63];
  assign data_o[31679] = data_o[63];
  assign data_o[31743] = data_o[63];
  assign data_o[31807] = data_o[63];
  assign data_o[31871] = data_o[63];
  assign data_o[31935] = data_o[63];
  assign data_o[31999] = data_o[63];
  assign data_o[126] = data_o[62];
  assign data_o[190] = data_o[62];
  assign data_o[254] = data_o[62];
  assign data_o[318] = data_o[62];
  assign data_o[382] = data_o[62];
  assign data_o[446] = data_o[62];
  assign data_o[510] = data_o[62];
  assign data_o[574] = data_o[62];
  assign data_o[638] = data_o[62];
  assign data_o[702] = data_o[62];
  assign data_o[766] = data_o[62];
  assign data_o[830] = data_o[62];
  assign data_o[894] = data_o[62];
  assign data_o[958] = data_o[62];
  assign data_o[1022] = data_o[62];
  assign data_o[1086] = data_o[62];
  assign data_o[1150] = data_o[62];
  assign data_o[1214] = data_o[62];
  assign data_o[1278] = data_o[62];
  assign data_o[1342] = data_o[62];
  assign data_o[1406] = data_o[62];
  assign data_o[1470] = data_o[62];
  assign data_o[1534] = data_o[62];
  assign data_o[1598] = data_o[62];
  assign data_o[1662] = data_o[62];
  assign data_o[1726] = data_o[62];
  assign data_o[1790] = data_o[62];
  assign data_o[1854] = data_o[62];
  assign data_o[1918] = data_o[62];
  assign data_o[1982] = data_o[62];
  assign data_o[2046] = data_o[62];
  assign data_o[2110] = data_o[62];
  assign data_o[2174] = data_o[62];
  assign data_o[2238] = data_o[62];
  assign data_o[2302] = data_o[62];
  assign data_o[2366] = data_o[62];
  assign data_o[2430] = data_o[62];
  assign data_o[2494] = data_o[62];
  assign data_o[2558] = data_o[62];
  assign data_o[2622] = data_o[62];
  assign data_o[2686] = data_o[62];
  assign data_o[2750] = data_o[62];
  assign data_o[2814] = data_o[62];
  assign data_o[2878] = data_o[62];
  assign data_o[2942] = data_o[62];
  assign data_o[3006] = data_o[62];
  assign data_o[3070] = data_o[62];
  assign data_o[3134] = data_o[62];
  assign data_o[3198] = data_o[62];
  assign data_o[3262] = data_o[62];
  assign data_o[3326] = data_o[62];
  assign data_o[3390] = data_o[62];
  assign data_o[3454] = data_o[62];
  assign data_o[3518] = data_o[62];
  assign data_o[3582] = data_o[62];
  assign data_o[3646] = data_o[62];
  assign data_o[3710] = data_o[62];
  assign data_o[3774] = data_o[62];
  assign data_o[3838] = data_o[62];
  assign data_o[3902] = data_o[62];
  assign data_o[3966] = data_o[62];
  assign data_o[4030] = data_o[62];
  assign data_o[4094] = data_o[62];
  assign data_o[4158] = data_o[62];
  assign data_o[4222] = data_o[62];
  assign data_o[4286] = data_o[62];
  assign data_o[4350] = data_o[62];
  assign data_o[4414] = data_o[62];
  assign data_o[4478] = data_o[62];
  assign data_o[4542] = data_o[62];
  assign data_o[4606] = data_o[62];
  assign data_o[4670] = data_o[62];
  assign data_o[4734] = data_o[62];
  assign data_o[4798] = data_o[62];
  assign data_o[4862] = data_o[62];
  assign data_o[4926] = data_o[62];
  assign data_o[4990] = data_o[62];
  assign data_o[5054] = data_o[62];
  assign data_o[5118] = data_o[62];
  assign data_o[5182] = data_o[62];
  assign data_o[5246] = data_o[62];
  assign data_o[5310] = data_o[62];
  assign data_o[5374] = data_o[62];
  assign data_o[5438] = data_o[62];
  assign data_o[5502] = data_o[62];
  assign data_o[5566] = data_o[62];
  assign data_o[5630] = data_o[62];
  assign data_o[5694] = data_o[62];
  assign data_o[5758] = data_o[62];
  assign data_o[5822] = data_o[62];
  assign data_o[5886] = data_o[62];
  assign data_o[5950] = data_o[62];
  assign data_o[6014] = data_o[62];
  assign data_o[6078] = data_o[62];
  assign data_o[6142] = data_o[62];
  assign data_o[6206] = data_o[62];
  assign data_o[6270] = data_o[62];
  assign data_o[6334] = data_o[62];
  assign data_o[6398] = data_o[62];
  assign data_o[6462] = data_o[62];
  assign data_o[6526] = data_o[62];
  assign data_o[6590] = data_o[62];
  assign data_o[6654] = data_o[62];
  assign data_o[6718] = data_o[62];
  assign data_o[6782] = data_o[62];
  assign data_o[6846] = data_o[62];
  assign data_o[6910] = data_o[62];
  assign data_o[6974] = data_o[62];
  assign data_o[7038] = data_o[62];
  assign data_o[7102] = data_o[62];
  assign data_o[7166] = data_o[62];
  assign data_o[7230] = data_o[62];
  assign data_o[7294] = data_o[62];
  assign data_o[7358] = data_o[62];
  assign data_o[7422] = data_o[62];
  assign data_o[7486] = data_o[62];
  assign data_o[7550] = data_o[62];
  assign data_o[7614] = data_o[62];
  assign data_o[7678] = data_o[62];
  assign data_o[7742] = data_o[62];
  assign data_o[7806] = data_o[62];
  assign data_o[7870] = data_o[62];
  assign data_o[7934] = data_o[62];
  assign data_o[7998] = data_o[62];
  assign data_o[8062] = data_o[62];
  assign data_o[8126] = data_o[62];
  assign data_o[8190] = data_o[62];
  assign data_o[8254] = data_o[62];
  assign data_o[8318] = data_o[62];
  assign data_o[8382] = data_o[62];
  assign data_o[8446] = data_o[62];
  assign data_o[8510] = data_o[62];
  assign data_o[8574] = data_o[62];
  assign data_o[8638] = data_o[62];
  assign data_o[8702] = data_o[62];
  assign data_o[8766] = data_o[62];
  assign data_o[8830] = data_o[62];
  assign data_o[8894] = data_o[62];
  assign data_o[8958] = data_o[62];
  assign data_o[9022] = data_o[62];
  assign data_o[9086] = data_o[62];
  assign data_o[9150] = data_o[62];
  assign data_o[9214] = data_o[62];
  assign data_o[9278] = data_o[62];
  assign data_o[9342] = data_o[62];
  assign data_o[9406] = data_o[62];
  assign data_o[9470] = data_o[62];
  assign data_o[9534] = data_o[62];
  assign data_o[9598] = data_o[62];
  assign data_o[9662] = data_o[62];
  assign data_o[9726] = data_o[62];
  assign data_o[9790] = data_o[62];
  assign data_o[9854] = data_o[62];
  assign data_o[9918] = data_o[62];
  assign data_o[9982] = data_o[62];
  assign data_o[10046] = data_o[62];
  assign data_o[10110] = data_o[62];
  assign data_o[10174] = data_o[62];
  assign data_o[10238] = data_o[62];
  assign data_o[10302] = data_o[62];
  assign data_o[10366] = data_o[62];
  assign data_o[10430] = data_o[62];
  assign data_o[10494] = data_o[62];
  assign data_o[10558] = data_o[62];
  assign data_o[10622] = data_o[62];
  assign data_o[10686] = data_o[62];
  assign data_o[10750] = data_o[62];
  assign data_o[10814] = data_o[62];
  assign data_o[10878] = data_o[62];
  assign data_o[10942] = data_o[62];
  assign data_o[11006] = data_o[62];
  assign data_o[11070] = data_o[62];
  assign data_o[11134] = data_o[62];
  assign data_o[11198] = data_o[62];
  assign data_o[11262] = data_o[62];
  assign data_o[11326] = data_o[62];
  assign data_o[11390] = data_o[62];
  assign data_o[11454] = data_o[62];
  assign data_o[11518] = data_o[62];
  assign data_o[11582] = data_o[62];
  assign data_o[11646] = data_o[62];
  assign data_o[11710] = data_o[62];
  assign data_o[11774] = data_o[62];
  assign data_o[11838] = data_o[62];
  assign data_o[11902] = data_o[62];
  assign data_o[11966] = data_o[62];
  assign data_o[12030] = data_o[62];
  assign data_o[12094] = data_o[62];
  assign data_o[12158] = data_o[62];
  assign data_o[12222] = data_o[62];
  assign data_o[12286] = data_o[62];
  assign data_o[12350] = data_o[62];
  assign data_o[12414] = data_o[62];
  assign data_o[12478] = data_o[62];
  assign data_o[12542] = data_o[62];
  assign data_o[12606] = data_o[62];
  assign data_o[12670] = data_o[62];
  assign data_o[12734] = data_o[62];
  assign data_o[12798] = data_o[62];
  assign data_o[12862] = data_o[62];
  assign data_o[12926] = data_o[62];
  assign data_o[12990] = data_o[62];
  assign data_o[13054] = data_o[62];
  assign data_o[13118] = data_o[62];
  assign data_o[13182] = data_o[62];
  assign data_o[13246] = data_o[62];
  assign data_o[13310] = data_o[62];
  assign data_o[13374] = data_o[62];
  assign data_o[13438] = data_o[62];
  assign data_o[13502] = data_o[62];
  assign data_o[13566] = data_o[62];
  assign data_o[13630] = data_o[62];
  assign data_o[13694] = data_o[62];
  assign data_o[13758] = data_o[62];
  assign data_o[13822] = data_o[62];
  assign data_o[13886] = data_o[62];
  assign data_o[13950] = data_o[62];
  assign data_o[14014] = data_o[62];
  assign data_o[14078] = data_o[62];
  assign data_o[14142] = data_o[62];
  assign data_o[14206] = data_o[62];
  assign data_o[14270] = data_o[62];
  assign data_o[14334] = data_o[62];
  assign data_o[14398] = data_o[62];
  assign data_o[14462] = data_o[62];
  assign data_o[14526] = data_o[62];
  assign data_o[14590] = data_o[62];
  assign data_o[14654] = data_o[62];
  assign data_o[14718] = data_o[62];
  assign data_o[14782] = data_o[62];
  assign data_o[14846] = data_o[62];
  assign data_o[14910] = data_o[62];
  assign data_o[14974] = data_o[62];
  assign data_o[15038] = data_o[62];
  assign data_o[15102] = data_o[62];
  assign data_o[15166] = data_o[62];
  assign data_o[15230] = data_o[62];
  assign data_o[15294] = data_o[62];
  assign data_o[15358] = data_o[62];
  assign data_o[15422] = data_o[62];
  assign data_o[15486] = data_o[62];
  assign data_o[15550] = data_o[62];
  assign data_o[15614] = data_o[62];
  assign data_o[15678] = data_o[62];
  assign data_o[15742] = data_o[62];
  assign data_o[15806] = data_o[62];
  assign data_o[15870] = data_o[62];
  assign data_o[15934] = data_o[62];
  assign data_o[15998] = data_o[62];
  assign data_o[16062] = data_o[62];
  assign data_o[16126] = data_o[62];
  assign data_o[16190] = data_o[62];
  assign data_o[16254] = data_o[62];
  assign data_o[16318] = data_o[62];
  assign data_o[16382] = data_o[62];
  assign data_o[16446] = data_o[62];
  assign data_o[16510] = data_o[62];
  assign data_o[16574] = data_o[62];
  assign data_o[16638] = data_o[62];
  assign data_o[16702] = data_o[62];
  assign data_o[16766] = data_o[62];
  assign data_o[16830] = data_o[62];
  assign data_o[16894] = data_o[62];
  assign data_o[16958] = data_o[62];
  assign data_o[17022] = data_o[62];
  assign data_o[17086] = data_o[62];
  assign data_o[17150] = data_o[62];
  assign data_o[17214] = data_o[62];
  assign data_o[17278] = data_o[62];
  assign data_o[17342] = data_o[62];
  assign data_o[17406] = data_o[62];
  assign data_o[17470] = data_o[62];
  assign data_o[17534] = data_o[62];
  assign data_o[17598] = data_o[62];
  assign data_o[17662] = data_o[62];
  assign data_o[17726] = data_o[62];
  assign data_o[17790] = data_o[62];
  assign data_o[17854] = data_o[62];
  assign data_o[17918] = data_o[62];
  assign data_o[17982] = data_o[62];
  assign data_o[18046] = data_o[62];
  assign data_o[18110] = data_o[62];
  assign data_o[18174] = data_o[62];
  assign data_o[18238] = data_o[62];
  assign data_o[18302] = data_o[62];
  assign data_o[18366] = data_o[62];
  assign data_o[18430] = data_o[62];
  assign data_o[18494] = data_o[62];
  assign data_o[18558] = data_o[62];
  assign data_o[18622] = data_o[62];
  assign data_o[18686] = data_o[62];
  assign data_o[18750] = data_o[62];
  assign data_o[18814] = data_o[62];
  assign data_o[18878] = data_o[62];
  assign data_o[18942] = data_o[62];
  assign data_o[19006] = data_o[62];
  assign data_o[19070] = data_o[62];
  assign data_o[19134] = data_o[62];
  assign data_o[19198] = data_o[62];
  assign data_o[19262] = data_o[62];
  assign data_o[19326] = data_o[62];
  assign data_o[19390] = data_o[62];
  assign data_o[19454] = data_o[62];
  assign data_o[19518] = data_o[62];
  assign data_o[19582] = data_o[62];
  assign data_o[19646] = data_o[62];
  assign data_o[19710] = data_o[62];
  assign data_o[19774] = data_o[62];
  assign data_o[19838] = data_o[62];
  assign data_o[19902] = data_o[62];
  assign data_o[19966] = data_o[62];
  assign data_o[20030] = data_o[62];
  assign data_o[20094] = data_o[62];
  assign data_o[20158] = data_o[62];
  assign data_o[20222] = data_o[62];
  assign data_o[20286] = data_o[62];
  assign data_o[20350] = data_o[62];
  assign data_o[20414] = data_o[62];
  assign data_o[20478] = data_o[62];
  assign data_o[20542] = data_o[62];
  assign data_o[20606] = data_o[62];
  assign data_o[20670] = data_o[62];
  assign data_o[20734] = data_o[62];
  assign data_o[20798] = data_o[62];
  assign data_o[20862] = data_o[62];
  assign data_o[20926] = data_o[62];
  assign data_o[20990] = data_o[62];
  assign data_o[21054] = data_o[62];
  assign data_o[21118] = data_o[62];
  assign data_o[21182] = data_o[62];
  assign data_o[21246] = data_o[62];
  assign data_o[21310] = data_o[62];
  assign data_o[21374] = data_o[62];
  assign data_o[21438] = data_o[62];
  assign data_o[21502] = data_o[62];
  assign data_o[21566] = data_o[62];
  assign data_o[21630] = data_o[62];
  assign data_o[21694] = data_o[62];
  assign data_o[21758] = data_o[62];
  assign data_o[21822] = data_o[62];
  assign data_o[21886] = data_o[62];
  assign data_o[21950] = data_o[62];
  assign data_o[22014] = data_o[62];
  assign data_o[22078] = data_o[62];
  assign data_o[22142] = data_o[62];
  assign data_o[22206] = data_o[62];
  assign data_o[22270] = data_o[62];
  assign data_o[22334] = data_o[62];
  assign data_o[22398] = data_o[62];
  assign data_o[22462] = data_o[62];
  assign data_o[22526] = data_o[62];
  assign data_o[22590] = data_o[62];
  assign data_o[22654] = data_o[62];
  assign data_o[22718] = data_o[62];
  assign data_o[22782] = data_o[62];
  assign data_o[22846] = data_o[62];
  assign data_o[22910] = data_o[62];
  assign data_o[22974] = data_o[62];
  assign data_o[23038] = data_o[62];
  assign data_o[23102] = data_o[62];
  assign data_o[23166] = data_o[62];
  assign data_o[23230] = data_o[62];
  assign data_o[23294] = data_o[62];
  assign data_o[23358] = data_o[62];
  assign data_o[23422] = data_o[62];
  assign data_o[23486] = data_o[62];
  assign data_o[23550] = data_o[62];
  assign data_o[23614] = data_o[62];
  assign data_o[23678] = data_o[62];
  assign data_o[23742] = data_o[62];
  assign data_o[23806] = data_o[62];
  assign data_o[23870] = data_o[62];
  assign data_o[23934] = data_o[62];
  assign data_o[23998] = data_o[62];
  assign data_o[24062] = data_o[62];
  assign data_o[24126] = data_o[62];
  assign data_o[24190] = data_o[62];
  assign data_o[24254] = data_o[62];
  assign data_o[24318] = data_o[62];
  assign data_o[24382] = data_o[62];
  assign data_o[24446] = data_o[62];
  assign data_o[24510] = data_o[62];
  assign data_o[24574] = data_o[62];
  assign data_o[24638] = data_o[62];
  assign data_o[24702] = data_o[62];
  assign data_o[24766] = data_o[62];
  assign data_o[24830] = data_o[62];
  assign data_o[24894] = data_o[62];
  assign data_o[24958] = data_o[62];
  assign data_o[25022] = data_o[62];
  assign data_o[25086] = data_o[62];
  assign data_o[25150] = data_o[62];
  assign data_o[25214] = data_o[62];
  assign data_o[25278] = data_o[62];
  assign data_o[25342] = data_o[62];
  assign data_o[25406] = data_o[62];
  assign data_o[25470] = data_o[62];
  assign data_o[25534] = data_o[62];
  assign data_o[25598] = data_o[62];
  assign data_o[25662] = data_o[62];
  assign data_o[25726] = data_o[62];
  assign data_o[25790] = data_o[62];
  assign data_o[25854] = data_o[62];
  assign data_o[25918] = data_o[62];
  assign data_o[25982] = data_o[62];
  assign data_o[26046] = data_o[62];
  assign data_o[26110] = data_o[62];
  assign data_o[26174] = data_o[62];
  assign data_o[26238] = data_o[62];
  assign data_o[26302] = data_o[62];
  assign data_o[26366] = data_o[62];
  assign data_o[26430] = data_o[62];
  assign data_o[26494] = data_o[62];
  assign data_o[26558] = data_o[62];
  assign data_o[26622] = data_o[62];
  assign data_o[26686] = data_o[62];
  assign data_o[26750] = data_o[62];
  assign data_o[26814] = data_o[62];
  assign data_o[26878] = data_o[62];
  assign data_o[26942] = data_o[62];
  assign data_o[27006] = data_o[62];
  assign data_o[27070] = data_o[62];
  assign data_o[27134] = data_o[62];
  assign data_o[27198] = data_o[62];
  assign data_o[27262] = data_o[62];
  assign data_o[27326] = data_o[62];
  assign data_o[27390] = data_o[62];
  assign data_o[27454] = data_o[62];
  assign data_o[27518] = data_o[62];
  assign data_o[27582] = data_o[62];
  assign data_o[27646] = data_o[62];
  assign data_o[27710] = data_o[62];
  assign data_o[27774] = data_o[62];
  assign data_o[27838] = data_o[62];
  assign data_o[27902] = data_o[62];
  assign data_o[27966] = data_o[62];
  assign data_o[28030] = data_o[62];
  assign data_o[28094] = data_o[62];
  assign data_o[28158] = data_o[62];
  assign data_o[28222] = data_o[62];
  assign data_o[28286] = data_o[62];
  assign data_o[28350] = data_o[62];
  assign data_o[28414] = data_o[62];
  assign data_o[28478] = data_o[62];
  assign data_o[28542] = data_o[62];
  assign data_o[28606] = data_o[62];
  assign data_o[28670] = data_o[62];
  assign data_o[28734] = data_o[62];
  assign data_o[28798] = data_o[62];
  assign data_o[28862] = data_o[62];
  assign data_o[28926] = data_o[62];
  assign data_o[28990] = data_o[62];
  assign data_o[29054] = data_o[62];
  assign data_o[29118] = data_o[62];
  assign data_o[29182] = data_o[62];
  assign data_o[29246] = data_o[62];
  assign data_o[29310] = data_o[62];
  assign data_o[29374] = data_o[62];
  assign data_o[29438] = data_o[62];
  assign data_o[29502] = data_o[62];
  assign data_o[29566] = data_o[62];
  assign data_o[29630] = data_o[62];
  assign data_o[29694] = data_o[62];
  assign data_o[29758] = data_o[62];
  assign data_o[29822] = data_o[62];
  assign data_o[29886] = data_o[62];
  assign data_o[29950] = data_o[62];
  assign data_o[30014] = data_o[62];
  assign data_o[30078] = data_o[62];
  assign data_o[30142] = data_o[62];
  assign data_o[30206] = data_o[62];
  assign data_o[30270] = data_o[62];
  assign data_o[30334] = data_o[62];
  assign data_o[30398] = data_o[62];
  assign data_o[30462] = data_o[62];
  assign data_o[30526] = data_o[62];
  assign data_o[30590] = data_o[62];
  assign data_o[30654] = data_o[62];
  assign data_o[30718] = data_o[62];
  assign data_o[30782] = data_o[62];
  assign data_o[30846] = data_o[62];
  assign data_o[30910] = data_o[62];
  assign data_o[30974] = data_o[62];
  assign data_o[31038] = data_o[62];
  assign data_o[31102] = data_o[62];
  assign data_o[31166] = data_o[62];
  assign data_o[31230] = data_o[62];
  assign data_o[31294] = data_o[62];
  assign data_o[31358] = data_o[62];
  assign data_o[31422] = data_o[62];
  assign data_o[31486] = data_o[62];
  assign data_o[31550] = data_o[62];
  assign data_o[31614] = data_o[62];
  assign data_o[31678] = data_o[62];
  assign data_o[31742] = data_o[62];
  assign data_o[31806] = data_o[62];
  assign data_o[31870] = data_o[62];
  assign data_o[31934] = data_o[62];
  assign data_o[31998] = data_o[62];
  assign data_o[125] = data_o[61];
  assign data_o[189] = data_o[61];
  assign data_o[253] = data_o[61];
  assign data_o[317] = data_o[61];
  assign data_o[381] = data_o[61];
  assign data_o[445] = data_o[61];
  assign data_o[509] = data_o[61];
  assign data_o[573] = data_o[61];
  assign data_o[637] = data_o[61];
  assign data_o[701] = data_o[61];
  assign data_o[765] = data_o[61];
  assign data_o[829] = data_o[61];
  assign data_o[893] = data_o[61];
  assign data_o[957] = data_o[61];
  assign data_o[1021] = data_o[61];
  assign data_o[1085] = data_o[61];
  assign data_o[1149] = data_o[61];
  assign data_o[1213] = data_o[61];
  assign data_o[1277] = data_o[61];
  assign data_o[1341] = data_o[61];
  assign data_o[1405] = data_o[61];
  assign data_o[1469] = data_o[61];
  assign data_o[1533] = data_o[61];
  assign data_o[1597] = data_o[61];
  assign data_o[1661] = data_o[61];
  assign data_o[1725] = data_o[61];
  assign data_o[1789] = data_o[61];
  assign data_o[1853] = data_o[61];
  assign data_o[1917] = data_o[61];
  assign data_o[1981] = data_o[61];
  assign data_o[2045] = data_o[61];
  assign data_o[2109] = data_o[61];
  assign data_o[2173] = data_o[61];
  assign data_o[2237] = data_o[61];
  assign data_o[2301] = data_o[61];
  assign data_o[2365] = data_o[61];
  assign data_o[2429] = data_o[61];
  assign data_o[2493] = data_o[61];
  assign data_o[2557] = data_o[61];
  assign data_o[2621] = data_o[61];
  assign data_o[2685] = data_o[61];
  assign data_o[2749] = data_o[61];
  assign data_o[2813] = data_o[61];
  assign data_o[2877] = data_o[61];
  assign data_o[2941] = data_o[61];
  assign data_o[3005] = data_o[61];
  assign data_o[3069] = data_o[61];
  assign data_o[3133] = data_o[61];
  assign data_o[3197] = data_o[61];
  assign data_o[3261] = data_o[61];
  assign data_o[3325] = data_o[61];
  assign data_o[3389] = data_o[61];
  assign data_o[3453] = data_o[61];
  assign data_o[3517] = data_o[61];
  assign data_o[3581] = data_o[61];
  assign data_o[3645] = data_o[61];
  assign data_o[3709] = data_o[61];
  assign data_o[3773] = data_o[61];
  assign data_o[3837] = data_o[61];
  assign data_o[3901] = data_o[61];
  assign data_o[3965] = data_o[61];
  assign data_o[4029] = data_o[61];
  assign data_o[4093] = data_o[61];
  assign data_o[4157] = data_o[61];
  assign data_o[4221] = data_o[61];
  assign data_o[4285] = data_o[61];
  assign data_o[4349] = data_o[61];
  assign data_o[4413] = data_o[61];
  assign data_o[4477] = data_o[61];
  assign data_o[4541] = data_o[61];
  assign data_o[4605] = data_o[61];
  assign data_o[4669] = data_o[61];
  assign data_o[4733] = data_o[61];
  assign data_o[4797] = data_o[61];
  assign data_o[4861] = data_o[61];
  assign data_o[4925] = data_o[61];
  assign data_o[4989] = data_o[61];
  assign data_o[5053] = data_o[61];
  assign data_o[5117] = data_o[61];
  assign data_o[5181] = data_o[61];
  assign data_o[5245] = data_o[61];
  assign data_o[5309] = data_o[61];
  assign data_o[5373] = data_o[61];
  assign data_o[5437] = data_o[61];
  assign data_o[5501] = data_o[61];
  assign data_o[5565] = data_o[61];
  assign data_o[5629] = data_o[61];
  assign data_o[5693] = data_o[61];
  assign data_o[5757] = data_o[61];
  assign data_o[5821] = data_o[61];
  assign data_o[5885] = data_o[61];
  assign data_o[5949] = data_o[61];
  assign data_o[6013] = data_o[61];
  assign data_o[6077] = data_o[61];
  assign data_o[6141] = data_o[61];
  assign data_o[6205] = data_o[61];
  assign data_o[6269] = data_o[61];
  assign data_o[6333] = data_o[61];
  assign data_o[6397] = data_o[61];
  assign data_o[6461] = data_o[61];
  assign data_o[6525] = data_o[61];
  assign data_o[6589] = data_o[61];
  assign data_o[6653] = data_o[61];
  assign data_o[6717] = data_o[61];
  assign data_o[6781] = data_o[61];
  assign data_o[6845] = data_o[61];
  assign data_o[6909] = data_o[61];
  assign data_o[6973] = data_o[61];
  assign data_o[7037] = data_o[61];
  assign data_o[7101] = data_o[61];
  assign data_o[7165] = data_o[61];
  assign data_o[7229] = data_o[61];
  assign data_o[7293] = data_o[61];
  assign data_o[7357] = data_o[61];
  assign data_o[7421] = data_o[61];
  assign data_o[7485] = data_o[61];
  assign data_o[7549] = data_o[61];
  assign data_o[7613] = data_o[61];
  assign data_o[7677] = data_o[61];
  assign data_o[7741] = data_o[61];
  assign data_o[7805] = data_o[61];
  assign data_o[7869] = data_o[61];
  assign data_o[7933] = data_o[61];
  assign data_o[7997] = data_o[61];
  assign data_o[8061] = data_o[61];
  assign data_o[8125] = data_o[61];
  assign data_o[8189] = data_o[61];
  assign data_o[8253] = data_o[61];
  assign data_o[8317] = data_o[61];
  assign data_o[8381] = data_o[61];
  assign data_o[8445] = data_o[61];
  assign data_o[8509] = data_o[61];
  assign data_o[8573] = data_o[61];
  assign data_o[8637] = data_o[61];
  assign data_o[8701] = data_o[61];
  assign data_o[8765] = data_o[61];
  assign data_o[8829] = data_o[61];
  assign data_o[8893] = data_o[61];
  assign data_o[8957] = data_o[61];
  assign data_o[9021] = data_o[61];
  assign data_o[9085] = data_o[61];
  assign data_o[9149] = data_o[61];
  assign data_o[9213] = data_o[61];
  assign data_o[9277] = data_o[61];
  assign data_o[9341] = data_o[61];
  assign data_o[9405] = data_o[61];
  assign data_o[9469] = data_o[61];
  assign data_o[9533] = data_o[61];
  assign data_o[9597] = data_o[61];
  assign data_o[9661] = data_o[61];
  assign data_o[9725] = data_o[61];
  assign data_o[9789] = data_o[61];
  assign data_o[9853] = data_o[61];
  assign data_o[9917] = data_o[61];
  assign data_o[9981] = data_o[61];
  assign data_o[10045] = data_o[61];
  assign data_o[10109] = data_o[61];
  assign data_o[10173] = data_o[61];
  assign data_o[10237] = data_o[61];
  assign data_o[10301] = data_o[61];
  assign data_o[10365] = data_o[61];
  assign data_o[10429] = data_o[61];
  assign data_o[10493] = data_o[61];
  assign data_o[10557] = data_o[61];
  assign data_o[10621] = data_o[61];
  assign data_o[10685] = data_o[61];
  assign data_o[10749] = data_o[61];
  assign data_o[10813] = data_o[61];
  assign data_o[10877] = data_o[61];
  assign data_o[10941] = data_o[61];
  assign data_o[11005] = data_o[61];
  assign data_o[11069] = data_o[61];
  assign data_o[11133] = data_o[61];
  assign data_o[11197] = data_o[61];
  assign data_o[11261] = data_o[61];
  assign data_o[11325] = data_o[61];
  assign data_o[11389] = data_o[61];
  assign data_o[11453] = data_o[61];
  assign data_o[11517] = data_o[61];
  assign data_o[11581] = data_o[61];
  assign data_o[11645] = data_o[61];
  assign data_o[11709] = data_o[61];
  assign data_o[11773] = data_o[61];
  assign data_o[11837] = data_o[61];
  assign data_o[11901] = data_o[61];
  assign data_o[11965] = data_o[61];
  assign data_o[12029] = data_o[61];
  assign data_o[12093] = data_o[61];
  assign data_o[12157] = data_o[61];
  assign data_o[12221] = data_o[61];
  assign data_o[12285] = data_o[61];
  assign data_o[12349] = data_o[61];
  assign data_o[12413] = data_o[61];
  assign data_o[12477] = data_o[61];
  assign data_o[12541] = data_o[61];
  assign data_o[12605] = data_o[61];
  assign data_o[12669] = data_o[61];
  assign data_o[12733] = data_o[61];
  assign data_o[12797] = data_o[61];
  assign data_o[12861] = data_o[61];
  assign data_o[12925] = data_o[61];
  assign data_o[12989] = data_o[61];
  assign data_o[13053] = data_o[61];
  assign data_o[13117] = data_o[61];
  assign data_o[13181] = data_o[61];
  assign data_o[13245] = data_o[61];
  assign data_o[13309] = data_o[61];
  assign data_o[13373] = data_o[61];
  assign data_o[13437] = data_o[61];
  assign data_o[13501] = data_o[61];
  assign data_o[13565] = data_o[61];
  assign data_o[13629] = data_o[61];
  assign data_o[13693] = data_o[61];
  assign data_o[13757] = data_o[61];
  assign data_o[13821] = data_o[61];
  assign data_o[13885] = data_o[61];
  assign data_o[13949] = data_o[61];
  assign data_o[14013] = data_o[61];
  assign data_o[14077] = data_o[61];
  assign data_o[14141] = data_o[61];
  assign data_o[14205] = data_o[61];
  assign data_o[14269] = data_o[61];
  assign data_o[14333] = data_o[61];
  assign data_o[14397] = data_o[61];
  assign data_o[14461] = data_o[61];
  assign data_o[14525] = data_o[61];
  assign data_o[14589] = data_o[61];
  assign data_o[14653] = data_o[61];
  assign data_o[14717] = data_o[61];
  assign data_o[14781] = data_o[61];
  assign data_o[14845] = data_o[61];
  assign data_o[14909] = data_o[61];
  assign data_o[14973] = data_o[61];
  assign data_o[15037] = data_o[61];
  assign data_o[15101] = data_o[61];
  assign data_o[15165] = data_o[61];
  assign data_o[15229] = data_o[61];
  assign data_o[15293] = data_o[61];
  assign data_o[15357] = data_o[61];
  assign data_o[15421] = data_o[61];
  assign data_o[15485] = data_o[61];
  assign data_o[15549] = data_o[61];
  assign data_o[15613] = data_o[61];
  assign data_o[15677] = data_o[61];
  assign data_o[15741] = data_o[61];
  assign data_o[15805] = data_o[61];
  assign data_o[15869] = data_o[61];
  assign data_o[15933] = data_o[61];
  assign data_o[15997] = data_o[61];
  assign data_o[16061] = data_o[61];
  assign data_o[16125] = data_o[61];
  assign data_o[16189] = data_o[61];
  assign data_o[16253] = data_o[61];
  assign data_o[16317] = data_o[61];
  assign data_o[16381] = data_o[61];
  assign data_o[16445] = data_o[61];
  assign data_o[16509] = data_o[61];
  assign data_o[16573] = data_o[61];
  assign data_o[16637] = data_o[61];
  assign data_o[16701] = data_o[61];
  assign data_o[16765] = data_o[61];
  assign data_o[16829] = data_o[61];
  assign data_o[16893] = data_o[61];
  assign data_o[16957] = data_o[61];
  assign data_o[17021] = data_o[61];
  assign data_o[17085] = data_o[61];
  assign data_o[17149] = data_o[61];
  assign data_o[17213] = data_o[61];
  assign data_o[17277] = data_o[61];
  assign data_o[17341] = data_o[61];
  assign data_o[17405] = data_o[61];
  assign data_o[17469] = data_o[61];
  assign data_o[17533] = data_o[61];
  assign data_o[17597] = data_o[61];
  assign data_o[17661] = data_o[61];
  assign data_o[17725] = data_o[61];
  assign data_o[17789] = data_o[61];
  assign data_o[17853] = data_o[61];
  assign data_o[17917] = data_o[61];
  assign data_o[17981] = data_o[61];
  assign data_o[18045] = data_o[61];
  assign data_o[18109] = data_o[61];
  assign data_o[18173] = data_o[61];
  assign data_o[18237] = data_o[61];
  assign data_o[18301] = data_o[61];
  assign data_o[18365] = data_o[61];
  assign data_o[18429] = data_o[61];
  assign data_o[18493] = data_o[61];
  assign data_o[18557] = data_o[61];
  assign data_o[18621] = data_o[61];
  assign data_o[18685] = data_o[61];
  assign data_o[18749] = data_o[61];
  assign data_o[18813] = data_o[61];
  assign data_o[18877] = data_o[61];
  assign data_o[18941] = data_o[61];
  assign data_o[19005] = data_o[61];
  assign data_o[19069] = data_o[61];
  assign data_o[19133] = data_o[61];
  assign data_o[19197] = data_o[61];
  assign data_o[19261] = data_o[61];
  assign data_o[19325] = data_o[61];
  assign data_o[19389] = data_o[61];
  assign data_o[19453] = data_o[61];
  assign data_o[19517] = data_o[61];
  assign data_o[19581] = data_o[61];
  assign data_o[19645] = data_o[61];
  assign data_o[19709] = data_o[61];
  assign data_o[19773] = data_o[61];
  assign data_o[19837] = data_o[61];
  assign data_o[19901] = data_o[61];
  assign data_o[19965] = data_o[61];
  assign data_o[20029] = data_o[61];
  assign data_o[20093] = data_o[61];
  assign data_o[20157] = data_o[61];
  assign data_o[20221] = data_o[61];
  assign data_o[20285] = data_o[61];
  assign data_o[20349] = data_o[61];
  assign data_o[20413] = data_o[61];
  assign data_o[20477] = data_o[61];
  assign data_o[20541] = data_o[61];
  assign data_o[20605] = data_o[61];
  assign data_o[20669] = data_o[61];
  assign data_o[20733] = data_o[61];
  assign data_o[20797] = data_o[61];
  assign data_o[20861] = data_o[61];
  assign data_o[20925] = data_o[61];
  assign data_o[20989] = data_o[61];
  assign data_o[21053] = data_o[61];
  assign data_o[21117] = data_o[61];
  assign data_o[21181] = data_o[61];
  assign data_o[21245] = data_o[61];
  assign data_o[21309] = data_o[61];
  assign data_o[21373] = data_o[61];
  assign data_o[21437] = data_o[61];
  assign data_o[21501] = data_o[61];
  assign data_o[21565] = data_o[61];
  assign data_o[21629] = data_o[61];
  assign data_o[21693] = data_o[61];
  assign data_o[21757] = data_o[61];
  assign data_o[21821] = data_o[61];
  assign data_o[21885] = data_o[61];
  assign data_o[21949] = data_o[61];
  assign data_o[22013] = data_o[61];
  assign data_o[22077] = data_o[61];
  assign data_o[22141] = data_o[61];
  assign data_o[22205] = data_o[61];
  assign data_o[22269] = data_o[61];
  assign data_o[22333] = data_o[61];
  assign data_o[22397] = data_o[61];
  assign data_o[22461] = data_o[61];
  assign data_o[22525] = data_o[61];
  assign data_o[22589] = data_o[61];
  assign data_o[22653] = data_o[61];
  assign data_o[22717] = data_o[61];
  assign data_o[22781] = data_o[61];
  assign data_o[22845] = data_o[61];
  assign data_o[22909] = data_o[61];
  assign data_o[22973] = data_o[61];
  assign data_o[23037] = data_o[61];
  assign data_o[23101] = data_o[61];
  assign data_o[23165] = data_o[61];
  assign data_o[23229] = data_o[61];
  assign data_o[23293] = data_o[61];
  assign data_o[23357] = data_o[61];
  assign data_o[23421] = data_o[61];
  assign data_o[23485] = data_o[61];
  assign data_o[23549] = data_o[61];
  assign data_o[23613] = data_o[61];
  assign data_o[23677] = data_o[61];
  assign data_o[23741] = data_o[61];
  assign data_o[23805] = data_o[61];
  assign data_o[23869] = data_o[61];
  assign data_o[23933] = data_o[61];
  assign data_o[23997] = data_o[61];
  assign data_o[24061] = data_o[61];
  assign data_o[24125] = data_o[61];
  assign data_o[24189] = data_o[61];
  assign data_o[24253] = data_o[61];
  assign data_o[24317] = data_o[61];
  assign data_o[24381] = data_o[61];
  assign data_o[24445] = data_o[61];
  assign data_o[24509] = data_o[61];
  assign data_o[24573] = data_o[61];
  assign data_o[24637] = data_o[61];
  assign data_o[24701] = data_o[61];
  assign data_o[24765] = data_o[61];
  assign data_o[24829] = data_o[61];
  assign data_o[24893] = data_o[61];
  assign data_o[24957] = data_o[61];
  assign data_o[25021] = data_o[61];
  assign data_o[25085] = data_o[61];
  assign data_o[25149] = data_o[61];
  assign data_o[25213] = data_o[61];
  assign data_o[25277] = data_o[61];
  assign data_o[25341] = data_o[61];
  assign data_o[25405] = data_o[61];
  assign data_o[25469] = data_o[61];
  assign data_o[25533] = data_o[61];
  assign data_o[25597] = data_o[61];
  assign data_o[25661] = data_o[61];
  assign data_o[25725] = data_o[61];
  assign data_o[25789] = data_o[61];
  assign data_o[25853] = data_o[61];
  assign data_o[25917] = data_o[61];
  assign data_o[25981] = data_o[61];
  assign data_o[26045] = data_o[61];
  assign data_o[26109] = data_o[61];
  assign data_o[26173] = data_o[61];
  assign data_o[26237] = data_o[61];
  assign data_o[26301] = data_o[61];
  assign data_o[26365] = data_o[61];
  assign data_o[26429] = data_o[61];
  assign data_o[26493] = data_o[61];
  assign data_o[26557] = data_o[61];
  assign data_o[26621] = data_o[61];
  assign data_o[26685] = data_o[61];
  assign data_o[26749] = data_o[61];
  assign data_o[26813] = data_o[61];
  assign data_o[26877] = data_o[61];
  assign data_o[26941] = data_o[61];
  assign data_o[27005] = data_o[61];
  assign data_o[27069] = data_o[61];
  assign data_o[27133] = data_o[61];
  assign data_o[27197] = data_o[61];
  assign data_o[27261] = data_o[61];
  assign data_o[27325] = data_o[61];
  assign data_o[27389] = data_o[61];
  assign data_o[27453] = data_o[61];
  assign data_o[27517] = data_o[61];
  assign data_o[27581] = data_o[61];
  assign data_o[27645] = data_o[61];
  assign data_o[27709] = data_o[61];
  assign data_o[27773] = data_o[61];
  assign data_o[27837] = data_o[61];
  assign data_o[27901] = data_o[61];
  assign data_o[27965] = data_o[61];
  assign data_o[28029] = data_o[61];
  assign data_o[28093] = data_o[61];
  assign data_o[28157] = data_o[61];
  assign data_o[28221] = data_o[61];
  assign data_o[28285] = data_o[61];
  assign data_o[28349] = data_o[61];
  assign data_o[28413] = data_o[61];
  assign data_o[28477] = data_o[61];
  assign data_o[28541] = data_o[61];
  assign data_o[28605] = data_o[61];
  assign data_o[28669] = data_o[61];
  assign data_o[28733] = data_o[61];
  assign data_o[28797] = data_o[61];
  assign data_o[28861] = data_o[61];
  assign data_o[28925] = data_o[61];
  assign data_o[28989] = data_o[61];
  assign data_o[29053] = data_o[61];
  assign data_o[29117] = data_o[61];
  assign data_o[29181] = data_o[61];
  assign data_o[29245] = data_o[61];
  assign data_o[29309] = data_o[61];
  assign data_o[29373] = data_o[61];
  assign data_o[29437] = data_o[61];
  assign data_o[29501] = data_o[61];
  assign data_o[29565] = data_o[61];
  assign data_o[29629] = data_o[61];
  assign data_o[29693] = data_o[61];
  assign data_o[29757] = data_o[61];
  assign data_o[29821] = data_o[61];
  assign data_o[29885] = data_o[61];
  assign data_o[29949] = data_o[61];
  assign data_o[30013] = data_o[61];
  assign data_o[30077] = data_o[61];
  assign data_o[30141] = data_o[61];
  assign data_o[30205] = data_o[61];
  assign data_o[30269] = data_o[61];
  assign data_o[30333] = data_o[61];
  assign data_o[30397] = data_o[61];
  assign data_o[30461] = data_o[61];
  assign data_o[30525] = data_o[61];
  assign data_o[30589] = data_o[61];
  assign data_o[30653] = data_o[61];
  assign data_o[30717] = data_o[61];
  assign data_o[30781] = data_o[61];
  assign data_o[30845] = data_o[61];
  assign data_o[30909] = data_o[61];
  assign data_o[30973] = data_o[61];
  assign data_o[31037] = data_o[61];
  assign data_o[31101] = data_o[61];
  assign data_o[31165] = data_o[61];
  assign data_o[31229] = data_o[61];
  assign data_o[31293] = data_o[61];
  assign data_o[31357] = data_o[61];
  assign data_o[31421] = data_o[61];
  assign data_o[31485] = data_o[61];
  assign data_o[31549] = data_o[61];
  assign data_o[31613] = data_o[61];
  assign data_o[31677] = data_o[61];
  assign data_o[31741] = data_o[61];
  assign data_o[31805] = data_o[61];
  assign data_o[31869] = data_o[61];
  assign data_o[31933] = data_o[61];
  assign data_o[31997] = data_o[61];
  assign data_o[124] = data_o[60];
  assign data_o[188] = data_o[60];
  assign data_o[252] = data_o[60];
  assign data_o[316] = data_o[60];
  assign data_o[380] = data_o[60];
  assign data_o[444] = data_o[60];
  assign data_o[508] = data_o[60];
  assign data_o[572] = data_o[60];
  assign data_o[636] = data_o[60];
  assign data_o[700] = data_o[60];
  assign data_o[764] = data_o[60];
  assign data_o[828] = data_o[60];
  assign data_o[892] = data_o[60];
  assign data_o[956] = data_o[60];
  assign data_o[1020] = data_o[60];
  assign data_o[1084] = data_o[60];
  assign data_o[1148] = data_o[60];
  assign data_o[1212] = data_o[60];
  assign data_o[1276] = data_o[60];
  assign data_o[1340] = data_o[60];
  assign data_o[1404] = data_o[60];
  assign data_o[1468] = data_o[60];
  assign data_o[1532] = data_o[60];
  assign data_o[1596] = data_o[60];
  assign data_o[1660] = data_o[60];
  assign data_o[1724] = data_o[60];
  assign data_o[1788] = data_o[60];
  assign data_o[1852] = data_o[60];
  assign data_o[1916] = data_o[60];
  assign data_o[1980] = data_o[60];
  assign data_o[2044] = data_o[60];
  assign data_o[2108] = data_o[60];
  assign data_o[2172] = data_o[60];
  assign data_o[2236] = data_o[60];
  assign data_o[2300] = data_o[60];
  assign data_o[2364] = data_o[60];
  assign data_o[2428] = data_o[60];
  assign data_o[2492] = data_o[60];
  assign data_o[2556] = data_o[60];
  assign data_o[2620] = data_o[60];
  assign data_o[2684] = data_o[60];
  assign data_o[2748] = data_o[60];
  assign data_o[2812] = data_o[60];
  assign data_o[2876] = data_o[60];
  assign data_o[2940] = data_o[60];
  assign data_o[3004] = data_o[60];
  assign data_o[3068] = data_o[60];
  assign data_o[3132] = data_o[60];
  assign data_o[3196] = data_o[60];
  assign data_o[3260] = data_o[60];
  assign data_o[3324] = data_o[60];
  assign data_o[3388] = data_o[60];
  assign data_o[3452] = data_o[60];
  assign data_o[3516] = data_o[60];
  assign data_o[3580] = data_o[60];
  assign data_o[3644] = data_o[60];
  assign data_o[3708] = data_o[60];
  assign data_o[3772] = data_o[60];
  assign data_o[3836] = data_o[60];
  assign data_o[3900] = data_o[60];
  assign data_o[3964] = data_o[60];
  assign data_o[4028] = data_o[60];
  assign data_o[4092] = data_o[60];
  assign data_o[4156] = data_o[60];
  assign data_o[4220] = data_o[60];
  assign data_o[4284] = data_o[60];
  assign data_o[4348] = data_o[60];
  assign data_o[4412] = data_o[60];
  assign data_o[4476] = data_o[60];
  assign data_o[4540] = data_o[60];
  assign data_o[4604] = data_o[60];
  assign data_o[4668] = data_o[60];
  assign data_o[4732] = data_o[60];
  assign data_o[4796] = data_o[60];
  assign data_o[4860] = data_o[60];
  assign data_o[4924] = data_o[60];
  assign data_o[4988] = data_o[60];
  assign data_o[5052] = data_o[60];
  assign data_o[5116] = data_o[60];
  assign data_o[5180] = data_o[60];
  assign data_o[5244] = data_o[60];
  assign data_o[5308] = data_o[60];
  assign data_o[5372] = data_o[60];
  assign data_o[5436] = data_o[60];
  assign data_o[5500] = data_o[60];
  assign data_o[5564] = data_o[60];
  assign data_o[5628] = data_o[60];
  assign data_o[5692] = data_o[60];
  assign data_o[5756] = data_o[60];
  assign data_o[5820] = data_o[60];
  assign data_o[5884] = data_o[60];
  assign data_o[5948] = data_o[60];
  assign data_o[6012] = data_o[60];
  assign data_o[6076] = data_o[60];
  assign data_o[6140] = data_o[60];
  assign data_o[6204] = data_o[60];
  assign data_o[6268] = data_o[60];
  assign data_o[6332] = data_o[60];
  assign data_o[6396] = data_o[60];
  assign data_o[6460] = data_o[60];
  assign data_o[6524] = data_o[60];
  assign data_o[6588] = data_o[60];
  assign data_o[6652] = data_o[60];
  assign data_o[6716] = data_o[60];
  assign data_o[6780] = data_o[60];
  assign data_o[6844] = data_o[60];
  assign data_o[6908] = data_o[60];
  assign data_o[6972] = data_o[60];
  assign data_o[7036] = data_o[60];
  assign data_o[7100] = data_o[60];
  assign data_o[7164] = data_o[60];
  assign data_o[7228] = data_o[60];
  assign data_o[7292] = data_o[60];
  assign data_o[7356] = data_o[60];
  assign data_o[7420] = data_o[60];
  assign data_o[7484] = data_o[60];
  assign data_o[7548] = data_o[60];
  assign data_o[7612] = data_o[60];
  assign data_o[7676] = data_o[60];
  assign data_o[7740] = data_o[60];
  assign data_o[7804] = data_o[60];
  assign data_o[7868] = data_o[60];
  assign data_o[7932] = data_o[60];
  assign data_o[7996] = data_o[60];
  assign data_o[8060] = data_o[60];
  assign data_o[8124] = data_o[60];
  assign data_o[8188] = data_o[60];
  assign data_o[8252] = data_o[60];
  assign data_o[8316] = data_o[60];
  assign data_o[8380] = data_o[60];
  assign data_o[8444] = data_o[60];
  assign data_o[8508] = data_o[60];
  assign data_o[8572] = data_o[60];
  assign data_o[8636] = data_o[60];
  assign data_o[8700] = data_o[60];
  assign data_o[8764] = data_o[60];
  assign data_o[8828] = data_o[60];
  assign data_o[8892] = data_o[60];
  assign data_o[8956] = data_o[60];
  assign data_o[9020] = data_o[60];
  assign data_o[9084] = data_o[60];
  assign data_o[9148] = data_o[60];
  assign data_o[9212] = data_o[60];
  assign data_o[9276] = data_o[60];
  assign data_o[9340] = data_o[60];
  assign data_o[9404] = data_o[60];
  assign data_o[9468] = data_o[60];
  assign data_o[9532] = data_o[60];
  assign data_o[9596] = data_o[60];
  assign data_o[9660] = data_o[60];
  assign data_o[9724] = data_o[60];
  assign data_o[9788] = data_o[60];
  assign data_o[9852] = data_o[60];
  assign data_o[9916] = data_o[60];
  assign data_o[9980] = data_o[60];
  assign data_o[10044] = data_o[60];
  assign data_o[10108] = data_o[60];
  assign data_o[10172] = data_o[60];
  assign data_o[10236] = data_o[60];
  assign data_o[10300] = data_o[60];
  assign data_o[10364] = data_o[60];
  assign data_o[10428] = data_o[60];
  assign data_o[10492] = data_o[60];
  assign data_o[10556] = data_o[60];
  assign data_o[10620] = data_o[60];
  assign data_o[10684] = data_o[60];
  assign data_o[10748] = data_o[60];
  assign data_o[10812] = data_o[60];
  assign data_o[10876] = data_o[60];
  assign data_o[10940] = data_o[60];
  assign data_o[11004] = data_o[60];
  assign data_o[11068] = data_o[60];
  assign data_o[11132] = data_o[60];
  assign data_o[11196] = data_o[60];
  assign data_o[11260] = data_o[60];
  assign data_o[11324] = data_o[60];
  assign data_o[11388] = data_o[60];
  assign data_o[11452] = data_o[60];
  assign data_o[11516] = data_o[60];
  assign data_o[11580] = data_o[60];
  assign data_o[11644] = data_o[60];
  assign data_o[11708] = data_o[60];
  assign data_o[11772] = data_o[60];
  assign data_o[11836] = data_o[60];
  assign data_o[11900] = data_o[60];
  assign data_o[11964] = data_o[60];
  assign data_o[12028] = data_o[60];
  assign data_o[12092] = data_o[60];
  assign data_o[12156] = data_o[60];
  assign data_o[12220] = data_o[60];
  assign data_o[12284] = data_o[60];
  assign data_o[12348] = data_o[60];
  assign data_o[12412] = data_o[60];
  assign data_o[12476] = data_o[60];
  assign data_o[12540] = data_o[60];
  assign data_o[12604] = data_o[60];
  assign data_o[12668] = data_o[60];
  assign data_o[12732] = data_o[60];
  assign data_o[12796] = data_o[60];
  assign data_o[12860] = data_o[60];
  assign data_o[12924] = data_o[60];
  assign data_o[12988] = data_o[60];
  assign data_o[13052] = data_o[60];
  assign data_o[13116] = data_o[60];
  assign data_o[13180] = data_o[60];
  assign data_o[13244] = data_o[60];
  assign data_o[13308] = data_o[60];
  assign data_o[13372] = data_o[60];
  assign data_o[13436] = data_o[60];
  assign data_o[13500] = data_o[60];
  assign data_o[13564] = data_o[60];
  assign data_o[13628] = data_o[60];
  assign data_o[13692] = data_o[60];
  assign data_o[13756] = data_o[60];
  assign data_o[13820] = data_o[60];
  assign data_o[13884] = data_o[60];
  assign data_o[13948] = data_o[60];
  assign data_o[14012] = data_o[60];
  assign data_o[14076] = data_o[60];
  assign data_o[14140] = data_o[60];
  assign data_o[14204] = data_o[60];
  assign data_o[14268] = data_o[60];
  assign data_o[14332] = data_o[60];
  assign data_o[14396] = data_o[60];
  assign data_o[14460] = data_o[60];
  assign data_o[14524] = data_o[60];
  assign data_o[14588] = data_o[60];
  assign data_o[14652] = data_o[60];
  assign data_o[14716] = data_o[60];
  assign data_o[14780] = data_o[60];
  assign data_o[14844] = data_o[60];
  assign data_o[14908] = data_o[60];
  assign data_o[14972] = data_o[60];
  assign data_o[15036] = data_o[60];
  assign data_o[15100] = data_o[60];
  assign data_o[15164] = data_o[60];
  assign data_o[15228] = data_o[60];
  assign data_o[15292] = data_o[60];
  assign data_o[15356] = data_o[60];
  assign data_o[15420] = data_o[60];
  assign data_o[15484] = data_o[60];
  assign data_o[15548] = data_o[60];
  assign data_o[15612] = data_o[60];
  assign data_o[15676] = data_o[60];
  assign data_o[15740] = data_o[60];
  assign data_o[15804] = data_o[60];
  assign data_o[15868] = data_o[60];
  assign data_o[15932] = data_o[60];
  assign data_o[15996] = data_o[60];
  assign data_o[16060] = data_o[60];
  assign data_o[16124] = data_o[60];
  assign data_o[16188] = data_o[60];
  assign data_o[16252] = data_o[60];
  assign data_o[16316] = data_o[60];
  assign data_o[16380] = data_o[60];
  assign data_o[16444] = data_o[60];
  assign data_o[16508] = data_o[60];
  assign data_o[16572] = data_o[60];
  assign data_o[16636] = data_o[60];
  assign data_o[16700] = data_o[60];
  assign data_o[16764] = data_o[60];
  assign data_o[16828] = data_o[60];
  assign data_o[16892] = data_o[60];
  assign data_o[16956] = data_o[60];
  assign data_o[17020] = data_o[60];
  assign data_o[17084] = data_o[60];
  assign data_o[17148] = data_o[60];
  assign data_o[17212] = data_o[60];
  assign data_o[17276] = data_o[60];
  assign data_o[17340] = data_o[60];
  assign data_o[17404] = data_o[60];
  assign data_o[17468] = data_o[60];
  assign data_o[17532] = data_o[60];
  assign data_o[17596] = data_o[60];
  assign data_o[17660] = data_o[60];
  assign data_o[17724] = data_o[60];
  assign data_o[17788] = data_o[60];
  assign data_o[17852] = data_o[60];
  assign data_o[17916] = data_o[60];
  assign data_o[17980] = data_o[60];
  assign data_o[18044] = data_o[60];
  assign data_o[18108] = data_o[60];
  assign data_o[18172] = data_o[60];
  assign data_o[18236] = data_o[60];
  assign data_o[18300] = data_o[60];
  assign data_o[18364] = data_o[60];
  assign data_o[18428] = data_o[60];
  assign data_o[18492] = data_o[60];
  assign data_o[18556] = data_o[60];
  assign data_o[18620] = data_o[60];
  assign data_o[18684] = data_o[60];
  assign data_o[18748] = data_o[60];
  assign data_o[18812] = data_o[60];
  assign data_o[18876] = data_o[60];
  assign data_o[18940] = data_o[60];
  assign data_o[19004] = data_o[60];
  assign data_o[19068] = data_o[60];
  assign data_o[19132] = data_o[60];
  assign data_o[19196] = data_o[60];
  assign data_o[19260] = data_o[60];
  assign data_o[19324] = data_o[60];
  assign data_o[19388] = data_o[60];
  assign data_o[19452] = data_o[60];
  assign data_o[19516] = data_o[60];
  assign data_o[19580] = data_o[60];
  assign data_o[19644] = data_o[60];
  assign data_o[19708] = data_o[60];
  assign data_o[19772] = data_o[60];
  assign data_o[19836] = data_o[60];
  assign data_o[19900] = data_o[60];
  assign data_o[19964] = data_o[60];
  assign data_o[20028] = data_o[60];
  assign data_o[20092] = data_o[60];
  assign data_o[20156] = data_o[60];
  assign data_o[20220] = data_o[60];
  assign data_o[20284] = data_o[60];
  assign data_o[20348] = data_o[60];
  assign data_o[20412] = data_o[60];
  assign data_o[20476] = data_o[60];
  assign data_o[20540] = data_o[60];
  assign data_o[20604] = data_o[60];
  assign data_o[20668] = data_o[60];
  assign data_o[20732] = data_o[60];
  assign data_o[20796] = data_o[60];
  assign data_o[20860] = data_o[60];
  assign data_o[20924] = data_o[60];
  assign data_o[20988] = data_o[60];
  assign data_o[21052] = data_o[60];
  assign data_o[21116] = data_o[60];
  assign data_o[21180] = data_o[60];
  assign data_o[21244] = data_o[60];
  assign data_o[21308] = data_o[60];
  assign data_o[21372] = data_o[60];
  assign data_o[21436] = data_o[60];
  assign data_o[21500] = data_o[60];
  assign data_o[21564] = data_o[60];
  assign data_o[21628] = data_o[60];
  assign data_o[21692] = data_o[60];
  assign data_o[21756] = data_o[60];
  assign data_o[21820] = data_o[60];
  assign data_o[21884] = data_o[60];
  assign data_o[21948] = data_o[60];
  assign data_o[22012] = data_o[60];
  assign data_o[22076] = data_o[60];
  assign data_o[22140] = data_o[60];
  assign data_o[22204] = data_o[60];
  assign data_o[22268] = data_o[60];
  assign data_o[22332] = data_o[60];
  assign data_o[22396] = data_o[60];
  assign data_o[22460] = data_o[60];
  assign data_o[22524] = data_o[60];
  assign data_o[22588] = data_o[60];
  assign data_o[22652] = data_o[60];
  assign data_o[22716] = data_o[60];
  assign data_o[22780] = data_o[60];
  assign data_o[22844] = data_o[60];
  assign data_o[22908] = data_o[60];
  assign data_o[22972] = data_o[60];
  assign data_o[23036] = data_o[60];
  assign data_o[23100] = data_o[60];
  assign data_o[23164] = data_o[60];
  assign data_o[23228] = data_o[60];
  assign data_o[23292] = data_o[60];
  assign data_o[23356] = data_o[60];
  assign data_o[23420] = data_o[60];
  assign data_o[23484] = data_o[60];
  assign data_o[23548] = data_o[60];
  assign data_o[23612] = data_o[60];
  assign data_o[23676] = data_o[60];
  assign data_o[23740] = data_o[60];
  assign data_o[23804] = data_o[60];
  assign data_o[23868] = data_o[60];
  assign data_o[23932] = data_o[60];
  assign data_o[23996] = data_o[60];
  assign data_o[24060] = data_o[60];
  assign data_o[24124] = data_o[60];
  assign data_o[24188] = data_o[60];
  assign data_o[24252] = data_o[60];
  assign data_o[24316] = data_o[60];
  assign data_o[24380] = data_o[60];
  assign data_o[24444] = data_o[60];
  assign data_o[24508] = data_o[60];
  assign data_o[24572] = data_o[60];
  assign data_o[24636] = data_o[60];
  assign data_o[24700] = data_o[60];
  assign data_o[24764] = data_o[60];
  assign data_o[24828] = data_o[60];
  assign data_o[24892] = data_o[60];
  assign data_o[24956] = data_o[60];
  assign data_o[25020] = data_o[60];
  assign data_o[25084] = data_o[60];
  assign data_o[25148] = data_o[60];
  assign data_o[25212] = data_o[60];
  assign data_o[25276] = data_o[60];
  assign data_o[25340] = data_o[60];
  assign data_o[25404] = data_o[60];
  assign data_o[25468] = data_o[60];
  assign data_o[25532] = data_o[60];
  assign data_o[25596] = data_o[60];
  assign data_o[25660] = data_o[60];
  assign data_o[25724] = data_o[60];
  assign data_o[25788] = data_o[60];
  assign data_o[25852] = data_o[60];
  assign data_o[25916] = data_o[60];
  assign data_o[25980] = data_o[60];
  assign data_o[26044] = data_o[60];
  assign data_o[26108] = data_o[60];
  assign data_o[26172] = data_o[60];
  assign data_o[26236] = data_o[60];
  assign data_o[26300] = data_o[60];
  assign data_o[26364] = data_o[60];
  assign data_o[26428] = data_o[60];
  assign data_o[26492] = data_o[60];
  assign data_o[26556] = data_o[60];
  assign data_o[26620] = data_o[60];
  assign data_o[26684] = data_o[60];
  assign data_o[26748] = data_o[60];
  assign data_o[26812] = data_o[60];
  assign data_o[26876] = data_o[60];
  assign data_o[26940] = data_o[60];
  assign data_o[27004] = data_o[60];
  assign data_o[27068] = data_o[60];
  assign data_o[27132] = data_o[60];
  assign data_o[27196] = data_o[60];
  assign data_o[27260] = data_o[60];
  assign data_o[27324] = data_o[60];
  assign data_o[27388] = data_o[60];
  assign data_o[27452] = data_o[60];
  assign data_o[27516] = data_o[60];
  assign data_o[27580] = data_o[60];
  assign data_o[27644] = data_o[60];
  assign data_o[27708] = data_o[60];
  assign data_o[27772] = data_o[60];
  assign data_o[27836] = data_o[60];
  assign data_o[27900] = data_o[60];
  assign data_o[27964] = data_o[60];
  assign data_o[28028] = data_o[60];
  assign data_o[28092] = data_o[60];
  assign data_o[28156] = data_o[60];
  assign data_o[28220] = data_o[60];
  assign data_o[28284] = data_o[60];
  assign data_o[28348] = data_o[60];
  assign data_o[28412] = data_o[60];
  assign data_o[28476] = data_o[60];
  assign data_o[28540] = data_o[60];
  assign data_o[28604] = data_o[60];
  assign data_o[28668] = data_o[60];
  assign data_o[28732] = data_o[60];
  assign data_o[28796] = data_o[60];
  assign data_o[28860] = data_o[60];
  assign data_o[28924] = data_o[60];
  assign data_o[28988] = data_o[60];
  assign data_o[29052] = data_o[60];
  assign data_o[29116] = data_o[60];
  assign data_o[29180] = data_o[60];
  assign data_o[29244] = data_o[60];
  assign data_o[29308] = data_o[60];
  assign data_o[29372] = data_o[60];
  assign data_o[29436] = data_o[60];
  assign data_o[29500] = data_o[60];
  assign data_o[29564] = data_o[60];
  assign data_o[29628] = data_o[60];
  assign data_o[29692] = data_o[60];
  assign data_o[29756] = data_o[60];
  assign data_o[29820] = data_o[60];
  assign data_o[29884] = data_o[60];
  assign data_o[29948] = data_o[60];
  assign data_o[30012] = data_o[60];
  assign data_o[30076] = data_o[60];
  assign data_o[30140] = data_o[60];
  assign data_o[30204] = data_o[60];
  assign data_o[30268] = data_o[60];
  assign data_o[30332] = data_o[60];
  assign data_o[30396] = data_o[60];
  assign data_o[30460] = data_o[60];
  assign data_o[30524] = data_o[60];
  assign data_o[30588] = data_o[60];
  assign data_o[30652] = data_o[60];
  assign data_o[30716] = data_o[60];
  assign data_o[30780] = data_o[60];
  assign data_o[30844] = data_o[60];
  assign data_o[30908] = data_o[60];
  assign data_o[30972] = data_o[60];
  assign data_o[31036] = data_o[60];
  assign data_o[31100] = data_o[60];
  assign data_o[31164] = data_o[60];
  assign data_o[31228] = data_o[60];
  assign data_o[31292] = data_o[60];
  assign data_o[31356] = data_o[60];
  assign data_o[31420] = data_o[60];
  assign data_o[31484] = data_o[60];
  assign data_o[31548] = data_o[60];
  assign data_o[31612] = data_o[60];
  assign data_o[31676] = data_o[60];
  assign data_o[31740] = data_o[60];
  assign data_o[31804] = data_o[60];
  assign data_o[31868] = data_o[60];
  assign data_o[31932] = data_o[60];
  assign data_o[31996] = data_o[60];
  assign data_o[123] = data_o[59];
  assign data_o[187] = data_o[59];
  assign data_o[251] = data_o[59];
  assign data_o[315] = data_o[59];
  assign data_o[379] = data_o[59];
  assign data_o[443] = data_o[59];
  assign data_o[507] = data_o[59];
  assign data_o[571] = data_o[59];
  assign data_o[635] = data_o[59];
  assign data_o[699] = data_o[59];
  assign data_o[763] = data_o[59];
  assign data_o[827] = data_o[59];
  assign data_o[891] = data_o[59];
  assign data_o[955] = data_o[59];
  assign data_o[1019] = data_o[59];
  assign data_o[1083] = data_o[59];
  assign data_o[1147] = data_o[59];
  assign data_o[1211] = data_o[59];
  assign data_o[1275] = data_o[59];
  assign data_o[1339] = data_o[59];
  assign data_o[1403] = data_o[59];
  assign data_o[1467] = data_o[59];
  assign data_o[1531] = data_o[59];
  assign data_o[1595] = data_o[59];
  assign data_o[1659] = data_o[59];
  assign data_o[1723] = data_o[59];
  assign data_o[1787] = data_o[59];
  assign data_o[1851] = data_o[59];
  assign data_o[1915] = data_o[59];
  assign data_o[1979] = data_o[59];
  assign data_o[2043] = data_o[59];
  assign data_o[2107] = data_o[59];
  assign data_o[2171] = data_o[59];
  assign data_o[2235] = data_o[59];
  assign data_o[2299] = data_o[59];
  assign data_o[2363] = data_o[59];
  assign data_o[2427] = data_o[59];
  assign data_o[2491] = data_o[59];
  assign data_o[2555] = data_o[59];
  assign data_o[2619] = data_o[59];
  assign data_o[2683] = data_o[59];
  assign data_o[2747] = data_o[59];
  assign data_o[2811] = data_o[59];
  assign data_o[2875] = data_o[59];
  assign data_o[2939] = data_o[59];
  assign data_o[3003] = data_o[59];
  assign data_o[3067] = data_o[59];
  assign data_o[3131] = data_o[59];
  assign data_o[3195] = data_o[59];
  assign data_o[3259] = data_o[59];
  assign data_o[3323] = data_o[59];
  assign data_o[3387] = data_o[59];
  assign data_o[3451] = data_o[59];
  assign data_o[3515] = data_o[59];
  assign data_o[3579] = data_o[59];
  assign data_o[3643] = data_o[59];
  assign data_o[3707] = data_o[59];
  assign data_o[3771] = data_o[59];
  assign data_o[3835] = data_o[59];
  assign data_o[3899] = data_o[59];
  assign data_o[3963] = data_o[59];
  assign data_o[4027] = data_o[59];
  assign data_o[4091] = data_o[59];
  assign data_o[4155] = data_o[59];
  assign data_o[4219] = data_o[59];
  assign data_o[4283] = data_o[59];
  assign data_o[4347] = data_o[59];
  assign data_o[4411] = data_o[59];
  assign data_o[4475] = data_o[59];
  assign data_o[4539] = data_o[59];
  assign data_o[4603] = data_o[59];
  assign data_o[4667] = data_o[59];
  assign data_o[4731] = data_o[59];
  assign data_o[4795] = data_o[59];
  assign data_o[4859] = data_o[59];
  assign data_o[4923] = data_o[59];
  assign data_o[4987] = data_o[59];
  assign data_o[5051] = data_o[59];
  assign data_o[5115] = data_o[59];
  assign data_o[5179] = data_o[59];
  assign data_o[5243] = data_o[59];
  assign data_o[5307] = data_o[59];
  assign data_o[5371] = data_o[59];
  assign data_o[5435] = data_o[59];
  assign data_o[5499] = data_o[59];
  assign data_o[5563] = data_o[59];
  assign data_o[5627] = data_o[59];
  assign data_o[5691] = data_o[59];
  assign data_o[5755] = data_o[59];
  assign data_o[5819] = data_o[59];
  assign data_o[5883] = data_o[59];
  assign data_o[5947] = data_o[59];
  assign data_o[6011] = data_o[59];
  assign data_o[6075] = data_o[59];
  assign data_o[6139] = data_o[59];
  assign data_o[6203] = data_o[59];
  assign data_o[6267] = data_o[59];
  assign data_o[6331] = data_o[59];
  assign data_o[6395] = data_o[59];
  assign data_o[6459] = data_o[59];
  assign data_o[6523] = data_o[59];
  assign data_o[6587] = data_o[59];
  assign data_o[6651] = data_o[59];
  assign data_o[6715] = data_o[59];
  assign data_o[6779] = data_o[59];
  assign data_o[6843] = data_o[59];
  assign data_o[6907] = data_o[59];
  assign data_o[6971] = data_o[59];
  assign data_o[7035] = data_o[59];
  assign data_o[7099] = data_o[59];
  assign data_o[7163] = data_o[59];
  assign data_o[7227] = data_o[59];
  assign data_o[7291] = data_o[59];
  assign data_o[7355] = data_o[59];
  assign data_o[7419] = data_o[59];
  assign data_o[7483] = data_o[59];
  assign data_o[7547] = data_o[59];
  assign data_o[7611] = data_o[59];
  assign data_o[7675] = data_o[59];
  assign data_o[7739] = data_o[59];
  assign data_o[7803] = data_o[59];
  assign data_o[7867] = data_o[59];
  assign data_o[7931] = data_o[59];
  assign data_o[7995] = data_o[59];
  assign data_o[8059] = data_o[59];
  assign data_o[8123] = data_o[59];
  assign data_o[8187] = data_o[59];
  assign data_o[8251] = data_o[59];
  assign data_o[8315] = data_o[59];
  assign data_o[8379] = data_o[59];
  assign data_o[8443] = data_o[59];
  assign data_o[8507] = data_o[59];
  assign data_o[8571] = data_o[59];
  assign data_o[8635] = data_o[59];
  assign data_o[8699] = data_o[59];
  assign data_o[8763] = data_o[59];
  assign data_o[8827] = data_o[59];
  assign data_o[8891] = data_o[59];
  assign data_o[8955] = data_o[59];
  assign data_o[9019] = data_o[59];
  assign data_o[9083] = data_o[59];
  assign data_o[9147] = data_o[59];
  assign data_o[9211] = data_o[59];
  assign data_o[9275] = data_o[59];
  assign data_o[9339] = data_o[59];
  assign data_o[9403] = data_o[59];
  assign data_o[9467] = data_o[59];
  assign data_o[9531] = data_o[59];
  assign data_o[9595] = data_o[59];
  assign data_o[9659] = data_o[59];
  assign data_o[9723] = data_o[59];
  assign data_o[9787] = data_o[59];
  assign data_o[9851] = data_o[59];
  assign data_o[9915] = data_o[59];
  assign data_o[9979] = data_o[59];
  assign data_o[10043] = data_o[59];
  assign data_o[10107] = data_o[59];
  assign data_o[10171] = data_o[59];
  assign data_o[10235] = data_o[59];
  assign data_o[10299] = data_o[59];
  assign data_o[10363] = data_o[59];
  assign data_o[10427] = data_o[59];
  assign data_o[10491] = data_o[59];
  assign data_o[10555] = data_o[59];
  assign data_o[10619] = data_o[59];
  assign data_o[10683] = data_o[59];
  assign data_o[10747] = data_o[59];
  assign data_o[10811] = data_o[59];
  assign data_o[10875] = data_o[59];
  assign data_o[10939] = data_o[59];
  assign data_o[11003] = data_o[59];
  assign data_o[11067] = data_o[59];
  assign data_o[11131] = data_o[59];
  assign data_o[11195] = data_o[59];
  assign data_o[11259] = data_o[59];
  assign data_o[11323] = data_o[59];
  assign data_o[11387] = data_o[59];
  assign data_o[11451] = data_o[59];
  assign data_o[11515] = data_o[59];
  assign data_o[11579] = data_o[59];
  assign data_o[11643] = data_o[59];
  assign data_o[11707] = data_o[59];
  assign data_o[11771] = data_o[59];
  assign data_o[11835] = data_o[59];
  assign data_o[11899] = data_o[59];
  assign data_o[11963] = data_o[59];
  assign data_o[12027] = data_o[59];
  assign data_o[12091] = data_o[59];
  assign data_o[12155] = data_o[59];
  assign data_o[12219] = data_o[59];
  assign data_o[12283] = data_o[59];
  assign data_o[12347] = data_o[59];
  assign data_o[12411] = data_o[59];
  assign data_o[12475] = data_o[59];
  assign data_o[12539] = data_o[59];
  assign data_o[12603] = data_o[59];
  assign data_o[12667] = data_o[59];
  assign data_o[12731] = data_o[59];
  assign data_o[12795] = data_o[59];
  assign data_o[12859] = data_o[59];
  assign data_o[12923] = data_o[59];
  assign data_o[12987] = data_o[59];
  assign data_o[13051] = data_o[59];
  assign data_o[13115] = data_o[59];
  assign data_o[13179] = data_o[59];
  assign data_o[13243] = data_o[59];
  assign data_o[13307] = data_o[59];
  assign data_o[13371] = data_o[59];
  assign data_o[13435] = data_o[59];
  assign data_o[13499] = data_o[59];
  assign data_o[13563] = data_o[59];
  assign data_o[13627] = data_o[59];
  assign data_o[13691] = data_o[59];
  assign data_o[13755] = data_o[59];
  assign data_o[13819] = data_o[59];
  assign data_o[13883] = data_o[59];
  assign data_o[13947] = data_o[59];
  assign data_o[14011] = data_o[59];
  assign data_o[14075] = data_o[59];
  assign data_o[14139] = data_o[59];
  assign data_o[14203] = data_o[59];
  assign data_o[14267] = data_o[59];
  assign data_o[14331] = data_o[59];
  assign data_o[14395] = data_o[59];
  assign data_o[14459] = data_o[59];
  assign data_o[14523] = data_o[59];
  assign data_o[14587] = data_o[59];
  assign data_o[14651] = data_o[59];
  assign data_o[14715] = data_o[59];
  assign data_o[14779] = data_o[59];
  assign data_o[14843] = data_o[59];
  assign data_o[14907] = data_o[59];
  assign data_o[14971] = data_o[59];
  assign data_o[15035] = data_o[59];
  assign data_o[15099] = data_o[59];
  assign data_o[15163] = data_o[59];
  assign data_o[15227] = data_o[59];
  assign data_o[15291] = data_o[59];
  assign data_o[15355] = data_o[59];
  assign data_o[15419] = data_o[59];
  assign data_o[15483] = data_o[59];
  assign data_o[15547] = data_o[59];
  assign data_o[15611] = data_o[59];
  assign data_o[15675] = data_o[59];
  assign data_o[15739] = data_o[59];
  assign data_o[15803] = data_o[59];
  assign data_o[15867] = data_o[59];
  assign data_o[15931] = data_o[59];
  assign data_o[15995] = data_o[59];
  assign data_o[16059] = data_o[59];
  assign data_o[16123] = data_o[59];
  assign data_o[16187] = data_o[59];
  assign data_o[16251] = data_o[59];
  assign data_o[16315] = data_o[59];
  assign data_o[16379] = data_o[59];
  assign data_o[16443] = data_o[59];
  assign data_o[16507] = data_o[59];
  assign data_o[16571] = data_o[59];
  assign data_o[16635] = data_o[59];
  assign data_o[16699] = data_o[59];
  assign data_o[16763] = data_o[59];
  assign data_o[16827] = data_o[59];
  assign data_o[16891] = data_o[59];
  assign data_o[16955] = data_o[59];
  assign data_o[17019] = data_o[59];
  assign data_o[17083] = data_o[59];
  assign data_o[17147] = data_o[59];
  assign data_o[17211] = data_o[59];
  assign data_o[17275] = data_o[59];
  assign data_o[17339] = data_o[59];
  assign data_o[17403] = data_o[59];
  assign data_o[17467] = data_o[59];
  assign data_o[17531] = data_o[59];
  assign data_o[17595] = data_o[59];
  assign data_o[17659] = data_o[59];
  assign data_o[17723] = data_o[59];
  assign data_o[17787] = data_o[59];
  assign data_o[17851] = data_o[59];
  assign data_o[17915] = data_o[59];
  assign data_o[17979] = data_o[59];
  assign data_o[18043] = data_o[59];
  assign data_o[18107] = data_o[59];
  assign data_o[18171] = data_o[59];
  assign data_o[18235] = data_o[59];
  assign data_o[18299] = data_o[59];
  assign data_o[18363] = data_o[59];
  assign data_o[18427] = data_o[59];
  assign data_o[18491] = data_o[59];
  assign data_o[18555] = data_o[59];
  assign data_o[18619] = data_o[59];
  assign data_o[18683] = data_o[59];
  assign data_o[18747] = data_o[59];
  assign data_o[18811] = data_o[59];
  assign data_o[18875] = data_o[59];
  assign data_o[18939] = data_o[59];
  assign data_o[19003] = data_o[59];
  assign data_o[19067] = data_o[59];
  assign data_o[19131] = data_o[59];
  assign data_o[19195] = data_o[59];
  assign data_o[19259] = data_o[59];
  assign data_o[19323] = data_o[59];
  assign data_o[19387] = data_o[59];
  assign data_o[19451] = data_o[59];
  assign data_o[19515] = data_o[59];
  assign data_o[19579] = data_o[59];
  assign data_o[19643] = data_o[59];
  assign data_o[19707] = data_o[59];
  assign data_o[19771] = data_o[59];
  assign data_o[19835] = data_o[59];
  assign data_o[19899] = data_o[59];
  assign data_o[19963] = data_o[59];
  assign data_o[20027] = data_o[59];
  assign data_o[20091] = data_o[59];
  assign data_o[20155] = data_o[59];
  assign data_o[20219] = data_o[59];
  assign data_o[20283] = data_o[59];
  assign data_o[20347] = data_o[59];
  assign data_o[20411] = data_o[59];
  assign data_o[20475] = data_o[59];
  assign data_o[20539] = data_o[59];
  assign data_o[20603] = data_o[59];
  assign data_o[20667] = data_o[59];
  assign data_o[20731] = data_o[59];
  assign data_o[20795] = data_o[59];
  assign data_o[20859] = data_o[59];
  assign data_o[20923] = data_o[59];
  assign data_o[20987] = data_o[59];
  assign data_o[21051] = data_o[59];
  assign data_o[21115] = data_o[59];
  assign data_o[21179] = data_o[59];
  assign data_o[21243] = data_o[59];
  assign data_o[21307] = data_o[59];
  assign data_o[21371] = data_o[59];
  assign data_o[21435] = data_o[59];
  assign data_o[21499] = data_o[59];
  assign data_o[21563] = data_o[59];
  assign data_o[21627] = data_o[59];
  assign data_o[21691] = data_o[59];
  assign data_o[21755] = data_o[59];
  assign data_o[21819] = data_o[59];
  assign data_o[21883] = data_o[59];
  assign data_o[21947] = data_o[59];
  assign data_o[22011] = data_o[59];
  assign data_o[22075] = data_o[59];
  assign data_o[22139] = data_o[59];
  assign data_o[22203] = data_o[59];
  assign data_o[22267] = data_o[59];
  assign data_o[22331] = data_o[59];
  assign data_o[22395] = data_o[59];
  assign data_o[22459] = data_o[59];
  assign data_o[22523] = data_o[59];
  assign data_o[22587] = data_o[59];
  assign data_o[22651] = data_o[59];
  assign data_o[22715] = data_o[59];
  assign data_o[22779] = data_o[59];
  assign data_o[22843] = data_o[59];
  assign data_o[22907] = data_o[59];
  assign data_o[22971] = data_o[59];
  assign data_o[23035] = data_o[59];
  assign data_o[23099] = data_o[59];
  assign data_o[23163] = data_o[59];
  assign data_o[23227] = data_o[59];
  assign data_o[23291] = data_o[59];
  assign data_o[23355] = data_o[59];
  assign data_o[23419] = data_o[59];
  assign data_o[23483] = data_o[59];
  assign data_o[23547] = data_o[59];
  assign data_o[23611] = data_o[59];
  assign data_o[23675] = data_o[59];
  assign data_o[23739] = data_o[59];
  assign data_o[23803] = data_o[59];
  assign data_o[23867] = data_o[59];
  assign data_o[23931] = data_o[59];
  assign data_o[23995] = data_o[59];
  assign data_o[24059] = data_o[59];
  assign data_o[24123] = data_o[59];
  assign data_o[24187] = data_o[59];
  assign data_o[24251] = data_o[59];
  assign data_o[24315] = data_o[59];
  assign data_o[24379] = data_o[59];
  assign data_o[24443] = data_o[59];
  assign data_o[24507] = data_o[59];
  assign data_o[24571] = data_o[59];
  assign data_o[24635] = data_o[59];
  assign data_o[24699] = data_o[59];
  assign data_o[24763] = data_o[59];
  assign data_o[24827] = data_o[59];
  assign data_o[24891] = data_o[59];
  assign data_o[24955] = data_o[59];
  assign data_o[25019] = data_o[59];
  assign data_o[25083] = data_o[59];
  assign data_o[25147] = data_o[59];
  assign data_o[25211] = data_o[59];
  assign data_o[25275] = data_o[59];
  assign data_o[25339] = data_o[59];
  assign data_o[25403] = data_o[59];
  assign data_o[25467] = data_o[59];
  assign data_o[25531] = data_o[59];
  assign data_o[25595] = data_o[59];
  assign data_o[25659] = data_o[59];
  assign data_o[25723] = data_o[59];
  assign data_o[25787] = data_o[59];
  assign data_o[25851] = data_o[59];
  assign data_o[25915] = data_o[59];
  assign data_o[25979] = data_o[59];
  assign data_o[26043] = data_o[59];
  assign data_o[26107] = data_o[59];
  assign data_o[26171] = data_o[59];
  assign data_o[26235] = data_o[59];
  assign data_o[26299] = data_o[59];
  assign data_o[26363] = data_o[59];
  assign data_o[26427] = data_o[59];
  assign data_o[26491] = data_o[59];
  assign data_o[26555] = data_o[59];
  assign data_o[26619] = data_o[59];
  assign data_o[26683] = data_o[59];
  assign data_o[26747] = data_o[59];
  assign data_o[26811] = data_o[59];
  assign data_o[26875] = data_o[59];
  assign data_o[26939] = data_o[59];
  assign data_o[27003] = data_o[59];
  assign data_o[27067] = data_o[59];
  assign data_o[27131] = data_o[59];
  assign data_o[27195] = data_o[59];
  assign data_o[27259] = data_o[59];
  assign data_o[27323] = data_o[59];
  assign data_o[27387] = data_o[59];
  assign data_o[27451] = data_o[59];
  assign data_o[27515] = data_o[59];
  assign data_o[27579] = data_o[59];
  assign data_o[27643] = data_o[59];
  assign data_o[27707] = data_o[59];
  assign data_o[27771] = data_o[59];
  assign data_o[27835] = data_o[59];
  assign data_o[27899] = data_o[59];
  assign data_o[27963] = data_o[59];
  assign data_o[28027] = data_o[59];
  assign data_o[28091] = data_o[59];
  assign data_o[28155] = data_o[59];
  assign data_o[28219] = data_o[59];
  assign data_o[28283] = data_o[59];
  assign data_o[28347] = data_o[59];
  assign data_o[28411] = data_o[59];
  assign data_o[28475] = data_o[59];
  assign data_o[28539] = data_o[59];
  assign data_o[28603] = data_o[59];
  assign data_o[28667] = data_o[59];
  assign data_o[28731] = data_o[59];
  assign data_o[28795] = data_o[59];
  assign data_o[28859] = data_o[59];
  assign data_o[28923] = data_o[59];
  assign data_o[28987] = data_o[59];
  assign data_o[29051] = data_o[59];
  assign data_o[29115] = data_o[59];
  assign data_o[29179] = data_o[59];
  assign data_o[29243] = data_o[59];
  assign data_o[29307] = data_o[59];
  assign data_o[29371] = data_o[59];
  assign data_o[29435] = data_o[59];
  assign data_o[29499] = data_o[59];
  assign data_o[29563] = data_o[59];
  assign data_o[29627] = data_o[59];
  assign data_o[29691] = data_o[59];
  assign data_o[29755] = data_o[59];
  assign data_o[29819] = data_o[59];
  assign data_o[29883] = data_o[59];
  assign data_o[29947] = data_o[59];
  assign data_o[30011] = data_o[59];
  assign data_o[30075] = data_o[59];
  assign data_o[30139] = data_o[59];
  assign data_o[30203] = data_o[59];
  assign data_o[30267] = data_o[59];
  assign data_o[30331] = data_o[59];
  assign data_o[30395] = data_o[59];
  assign data_o[30459] = data_o[59];
  assign data_o[30523] = data_o[59];
  assign data_o[30587] = data_o[59];
  assign data_o[30651] = data_o[59];
  assign data_o[30715] = data_o[59];
  assign data_o[30779] = data_o[59];
  assign data_o[30843] = data_o[59];
  assign data_o[30907] = data_o[59];
  assign data_o[30971] = data_o[59];
  assign data_o[31035] = data_o[59];
  assign data_o[31099] = data_o[59];
  assign data_o[31163] = data_o[59];
  assign data_o[31227] = data_o[59];
  assign data_o[31291] = data_o[59];
  assign data_o[31355] = data_o[59];
  assign data_o[31419] = data_o[59];
  assign data_o[31483] = data_o[59];
  assign data_o[31547] = data_o[59];
  assign data_o[31611] = data_o[59];
  assign data_o[31675] = data_o[59];
  assign data_o[31739] = data_o[59];
  assign data_o[31803] = data_o[59];
  assign data_o[31867] = data_o[59];
  assign data_o[31931] = data_o[59];
  assign data_o[31995] = data_o[59];
  assign data_o[122] = data_o[58];
  assign data_o[186] = data_o[58];
  assign data_o[250] = data_o[58];
  assign data_o[314] = data_o[58];
  assign data_o[378] = data_o[58];
  assign data_o[442] = data_o[58];
  assign data_o[506] = data_o[58];
  assign data_o[570] = data_o[58];
  assign data_o[634] = data_o[58];
  assign data_o[698] = data_o[58];
  assign data_o[762] = data_o[58];
  assign data_o[826] = data_o[58];
  assign data_o[890] = data_o[58];
  assign data_o[954] = data_o[58];
  assign data_o[1018] = data_o[58];
  assign data_o[1082] = data_o[58];
  assign data_o[1146] = data_o[58];
  assign data_o[1210] = data_o[58];
  assign data_o[1274] = data_o[58];
  assign data_o[1338] = data_o[58];
  assign data_o[1402] = data_o[58];
  assign data_o[1466] = data_o[58];
  assign data_o[1530] = data_o[58];
  assign data_o[1594] = data_o[58];
  assign data_o[1658] = data_o[58];
  assign data_o[1722] = data_o[58];
  assign data_o[1786] = data_o[58];
  assign data_o[1850] = data_o[58];
  assign data_o[1914] = data_o[58];
  assign data_o[1978] = data_o[58];
  assign data_o[2042] = data_o[58];
  assign data_o[2106] = data_o[58];
  assign data_o[2170] = data_o[58];
  assign data_o[2234] = data_o[58];
  assign data_o[2298] = data_o[58];
  assign data_o[2362] = data_o[58];
  assign data_o[2426] = data_o[58];
  assign data_o[2490] = data_o[58];
  assign data_o[2554] = data_o[58];
  assign data_o[2618] = data_o[58];
  assign data_o[2682] = data_o[58];
  assign data_o[2746] = data_o[58];
  assign data_o[2810] = data_o[58];
  assign data_o[2874] = data_o[58];
  assign data_o[2938] = data_o[58];
  assign data_o[3002] = data_o[58];
  assign data_o[3066] = data_o[58];
  assign data_o[3130] = data_o[58];
  assign data_o[3194] = data_o[58];
  assign data_o[3258] = data_o[58];
  assign data_o[3322] = data_o[58];
  assign data_o[3386] = data_o[58];
  assign data_o[3450] = data_o[58];
  assign data_o[3514] = data_o[58];
  assign data_o[3578] = data_o[58];
  assign data_o[3642] = data_o[58];
  assign data_o[3706] = data_o[58];
  assign data_o[3770] = data_o[58];
  assign data_o[3834] = data_o[58];
  assign data_o[3898] = data_o[58];
  assign data_o[3962] = data_o[58];
  assign data_o[4026] = data_o[58];
  assign data_o[4090] = data_o[58];
  assign data_o[4154] = data_o[58];
  assign data_o[4218] = data_o[58];
  assign data_o[4282] = data_o[58];
  assign data_o[4346] = data_o[58];
  assign data_o[4410] = data_o[58];
  assign data_o[4474] = data_o[58];
  assign data_o[4538] = data_o[58];
  assign data_o[4602] = data_o[58];
  assign data_o[4666] = data_o[58];
  assign data_o[4730] = data_o[58];
  assign data_o[4794] = data_o[58];
  assign data_o[4858] = data_o[58];
  assign data_o[4922] = data_o[58];
  assign data_o[4986] = data_o[58];
  assign data_o[5050] = data_o[58];
  assign data_o[5114] = data_o[58];
  assign data_o[5178] = data_o[58];
  assign data_o[5242] = data_o[58];
  assign data_o[5306] = data_o[58];
  assign data_o[5370] = data_o[58];
  assign data_o[5434] = data_o[58];
  assign data_o[5498] = data_o[58];
  assign data_o[5562] = data_o[58];
  assign data_o[5626] = data_o[58];
  assign data_o[5690] = data_o[58];
  assign data_o[5754] = data_o[58];
  assign data_o[5818] = data_o[58];
  assign data_o[5882] = data_o[58];
  assign data_o[5946] = data_o[58];
  assign data_o[6010] = data_o[58];
  assign data_o[6074] = data_o[58];
  assign data_o[6138] = data_o[58];
  assign data_o[6202] = data_o[58];
  assign data_o[6266] = data_o[58];
  assign data_o[6330] = data_o[58];
  assign data_o[6394] = data_o[58];
  assign data_o[6458] = data_o[58];
  assign data_o[6522] = data_o[58];
  assign data_o[6586] = data_o[58];
  assign data_o[6650] = data_o[58];
  assign data_o[6714] = data_o[58];
  assign data_o[6778] = data_o[58];
  assign data_o[6842] = data_o[58];
  assign data_o[6906] = data_o[58];
  assign data_o[6970] = data_o[58];
  assign data_o[7034] = data_o[58];
  assign data_o[7098] = data_o[58];
  assign data_o[7162] = data_o[58];
  assign data_o[7226] = data_o[58];
  assign data_o[7290] = data_o[58];
  assign data_o[7354] = data_o[58];
  assign data_o[7418] = data_o[58];
  assign data_o[7482] = data_o[58];
  assign data_o[7546] = data_o[58];
  assign data_o[7610] = data_o[58];
  assign data_o[7674] = data_o[58];
  assign data_o[7738] = data_o[58];
  assign data_o[7802] = data_o[58];
  assign data_o[7866] = data_o[58];
  assign data_o[7930] = data_o[58];
  assign data_o[7994] = data_o[58];
  assign data_o[8058] = data_o[58];
  assign data_o[8122] = data_o[58];
  assign data_o[8186] = data_o[58];
  assign data_o[8250] = data_o[58];
  assign data_o[8314] = data_o[58];
  assign data_o[8378] = data_o[58];
  assign data_o[8442] = data_o[58];
  assign data_o[8506] = data_o[58];
  assign data_o[8570] = data_o[58];
  assign data_o[8634] = data_o[58];
  assign data_o[8698] = data_o[58];
  assign data_o[8762] = data_o[58];
  assign data_o[8826] = data_o[58];
  assign data_o[8890] = data_o[58];
  assign data_o[8954] = data_o[58];
  assign data_o[9018] = data_o[58];
  assign data_o[9082] = data_o[58];
  assign data_o[9146] = data_o[58];
  assign data_o[9210] = data_o[58];
  assign data_o[9274] = data_o[58];
  assign data_o[9338] = data_o[58];
  assign data_o[9402] = data_o[58];
  assign data_o[9466] = data_o[58];
  assign data_o[9530] = data_o[58];
  assign data_o[9594] = data_o[58];
  assign data_o[9658] = data_o[58];
  assign data_o[9722] = data_o[58];
  assign data_o[9786] = data_o[58];
  assign data_o[9850] = data_o[58];
  assign data_o[9914] = data_o[58];
  assign data_o[9978] = data_o[58];
  assign data_o[10042] = data_o[58];
  assign data_o[10106] = data_o[58];
  assign data_o[10170] = data_o[58];
  assign data_o[10234] = data_o[58];
  assign data_o[10298] = data_o[58];
  assign data_o[10362] = data_o[58];
  assign data_o[10426] = data_o[58];
  assign data_o[10490] = data_o[58];
  assign data_o[10554] = data_o[58];
  assign data_o[10618] = data_o[58];
  assign data_o[10682] = data_o[58];
  assign data_o[10746] = data_o[58];
  assign data_o[10810] = data_o[58];
  assign data_o[10874] = data_o[58];
  assign data_o[10938] = data_o[58];
  assign data_o[11002] = data_o[58];
  assign data_o[11066] = data_o[58];
  assign data_o[11130] = data_o[58];
  assign data_o[11194] = data_o[58];
  assign data_o[11258] = data_o[58];
  assign data_o[11322] = data_o[58];
  assign data_o[11386] = data_o[58];
  assign data_o[11450] = data_o[58];
  assign data_o[11514] = data_o[58];
  assign data_o[11578] = data_o[58];
  assign data_o[11642] = data_o[58];
  assign data_o[11706] = data_o[58];
  assign data_o[11770] = data_o[58];
  assign data_o[11834] = data_o[58];
  assign data_o[11898] = data_o[58];
  assign data_o[11962] = data_o[58];
  assign data_o[12026] = data_o[58];
  assign data_o[12090] = data_o[58];
  assign data_o[12154] = data_o[58];
  assign data_o[12218] = data_o[58];
  assign data_o[12282] = data_o[58];
  assign data_o[12346] = data_o[58];
  assign data_o[12410] = data_o[58];
  assign data_o[12474] = data_o[58];
  assign data_o[12538] = data_o[58];
  assign data_o[12602] = data_o[58];
  assign data_o[12666] = data_o[58];
  assign data_o[12730] = data_o[58];
  assign data_o[12794] = data_o[58];
  assign data_o[12858] = data_o[58];
  assign data_o[12922] = data_o[58];
  assign data_o[12986] = data_o[58];
  assign data_o[13050] = data_o[58];
  assign data_o[13114] = data_o[58];
  assign data_o[13178] = data_o[58];
  assign data_o[13242] = data_o[58];
  assign data_o[13306] = data_o[58];
  assign data_o[13370] = data_o[58];
  assign data_o[13434] = data_o[58];
  assign data_o[13498] = data_o[58];
  assign data_o[13562] = data_o[58];
  assign data_o[13626] = data_o[58];
  assign data_o[13690] = data_o[58];
  assign data_o[13754] = data_o[58];
  assign data_o[13818] = data_o[58];
  assign data_o[13882] = data_o[58];
  assign data_o[13946] = data_o[58];
  assign data_o[14010] = data_o[58];
  assign data_o[14074] = data_o[58];
  assign data_o[14138] = data_o[58];
  assign data_o[14202] = data_o[58];
  assign data_o[14266] = data_o[58];
  assign data_o[14330] = data_o[58];
  assign data_o[14394] = data_o[58];
  assign data_o[14458] = data_o[58];
  assign data_o[14522] = data_o[58];
  assign data_o[14586] = data_o[58];
  assign data_o[14650] = data_o[58];
  assign data_o[14714] = data_o[58];
  assign data_o[14778] = data_o[58];
  assign data_o[14842] = data_o[58];
  assign data_o[14906] = data_o[58];
  assign data_o[14970] = data_o[58];
  assign data_o[15034] = data_o[58];
  assign data_o[15098] = data_o[58];
  assign data_o[15162] = data_o[58];
  assign data_o[15226] = data_o[58];
  assign data_o[15290] = data_o[58];
  assign data_o[15354] = data_o[58];
  assign data_o[15418] = data_o[58];
  assign data_o[15482] = data_o[58];
  assign data_o[15546] = data_o[58];
  assign data_o[15610] = data_o[58];
  assign data_o[15674] = data_o[58];
  assign data_o[15738] = data_o[58];
  assign data_o[15802] = data_o[58];
  assign data_o[15866] = data_o[58];
  assign data_o[15930] = data_o[58];
  assign data_o[15994] = data_o[58];
  assign data_o[16058] = data_o[58];
  assign data_o[16122] = data_o[58];
  assign data_o[16186] = data_o[58];
  assign data_o[16250] = data_o[58];
  assign data_o[16314] = data_o[58];
  assign data_o[16378] = data_o[58];
  assign data_o[16442] = data_o[58];
  assign data_o[16506] = data_o[58];
  assign data_o[16570] = data_o[58];
  assign data_o[16634] = data_o[58];
  assign data_o[16698] = data_o[58];
  assign data_o[16762] = data_o[58];
  assign data_o[16826] = data_o[58];
  assign data_o[16890] = data_o[58];
  assign data_o[16954] = data_o[58];
  assign data_o[17018] = data_o[58];
  assign data_o[17082] = data_o[58];
  assign data_o[17146] = data_o[58];
  assign data_o[17210] = data_o[58];
  assign data_o[17274] = data_o[58];
  assign data_o[17338] = data_o[58];
  assign data_o[17402] = data_o[58];
  assign data_o[17466] = data_o[58];
  assign data_o[17530] = data_o[58];
  assign data_o[17594] = data_o[58];
  assign data_o[17658] = data_o[58];
  assign data_o[17722] = data_o[58];
  assign data_o[17786] = data_o[58];
  assign data_o[17850] = data_o[58];
  assign data_o[17914] = data_o[58];
  assign data_o[17978] = data_o[58];
  assign data_o[18042] = data_o[58];
  assign data_o[18106] = data_o[58];
  assign data_o[18170] = data_o[58];
  assign data_o[18234] = data_o[58];
  assign data_o[18298] = data_o[58];
  assign data_o[18362] = data_o[58];
  assign data_o[18426] = data_o[58];
  assign data_o[18490] = data_o[58];
  assign data_o[18554] = data_o[58];
  assign data_o[18618] = data_o[58];
  assign data_o[18682] = data_o[58];
  assign data_o[18746] = data_o[58];
  assign data_o[18810] = data_o[58];
  assign data_o[18874] = data_o[58];
  assign data_o[18938] = data_o[58];
  assign data_o[19002] = data_o[58];
  assign data_o[19066] = data_o[58];
  assign data_o[19130] = data_o[58];
  assign data_o[19194] = data_o[58];
  assign data_o[19258] = data_o[58];
  assign data_o[19322] = data_o[58];
  assign data_o[19386] = data_o[58];
  assign data_o[19450] = data_o[58];
  assign data_o[19514] = data_o[58];
  assign data_o[19578] = data_o[58];
  assign data_o[19642] = data_o[58];
  assign data_o[19706] = data_o[58];
  assign data_o[19770] = data_o[58];
  assign data_o[19834] = data_o[58];
  assign data_o[19898] = data_o[58];
  assign data_o[19962] = data_o[58];
  assign data_o[20026] = data_o[58];
  assign data_o[20090] = data_o[58];
  assign data_o[20154] = data_o[58];
  assign data_o[20218] = data_o[58];
  assign data_o[20282] = data_o[58];
  assign data_o[20346] = data_o[58];
  assign data_o[20410] = data_o[58];
  assign data_o[20474] = data_o[58];
  assign data_o[20538] = data_o[58];
  assign data_o[20602] = data_o[58];
  assign data_o[20666] = data_o[58];
  assign data_o[20730] = data_o[58];
  assign data_o[20794] = data_o[58];
  assign data_o[20858] = data_o[58];
  assign data_o[20922] = data_o[58];
  assign data_o[20986] = data_o[58];
  assign data_o[21050] = data_o[58];
  assign data_o[21114] = data_o[58];
  assign data_o[21178] = data_o[58];
  assign data_o[21242] = data_o[58];
  assign data_o[21306] = data_o[58];
  assign data_o[21370] = data_o[58];
  assign data_o[21434] = data_o[58];
  assign data_o[21498] = data_o[58];
  assign data_o[21562] = data_o[58];
  assign data_o[21626] = data_o[58];
  assign data_o[21690] = data_o[58];
  assign data_o[21754] = data_o[58];
  assign data_o[21818] = data_o[58];
  assign data_o[21882] = data_o[58];
  assign data_o[21946] = data_o[58];
  assign data_o[22010] = data_o[58];
  assign data_o[22074] = data_o[58];
  assign data_o[22138] = data_o[58];
  assign data_o[22202] = data_o[58];
  assign data_o[22266] = data_o[58];
  assign data_o[22330] = data_o[58];
  assign data_o[22394] = data_o[58];
  assign data_o[22458] = data_o[58];
  assign data_o[22522] = data_o[58];
  assign data_o[22586] = data_o[58];
  assign data_o[22650] = data_o[58];
  assign data_o[22714] = data_o[58];
  assign data_o[22778] = data_o[58];
  assign data_o[22842] = data_o[58];
  assign data_o[22906] = data_o[58];
  assign data_o[22970] = data_o[58];
  assign data_o[23034] = data_o[58];
  assign data_o[23098] = data_o[58];
  assign data_o[23162] = data_o[58];
  assign data_o[23226] = data_o[58];
  assign data_o[23290] = data_o[58];
  assign data_o[23354] = data_o[58];
  assign data_o[23418] = data_o[58];
  assign data_o[23482] = data_o[58];
  assign data_o[23546] = data_o[58];
  assign data_o[23610] = data_o[58];
  assign data_o[23674] = data_o[58];
  assign data_o[23738] = data_o[58];
  assign data_o[23802] = data_o[58];
  assign data_o[23866] = data_o[58];
  assign data_o[23930] = data_o[58];
  assign data_o[23994] = data_o[58];
  assign data_o[24058] = data_o[58];
  assign data_o[24122] = data_o[58];
  assign data_o[24186] = data_o[58];
  assign data_o[24250] = data_o[58];
  assign data_o[24314] = data_o[58];
  assign data_o[24378] = data_o[58];
  assign data_o[24442] = data_o[58];
  assign data_o[24506] = data_o[58];
  assign data_o[24570] = data_o[58];
  assign data_o[24634] = data_o[58];
  assign data_o[24698] = data_o[58];
  assign data_o[24762] = data_o[58];
  assign data_o[24826] = data_o[58];
  assign data_o[24890] = data_o[58];
  assign data_o[24954] = data_o[58];
  assign data_o[25018] = data_o[58];
  assign data_o[25082] = data_o[58];
  assign data_o[25146] = data_o[58];
  assign data_o[25210] = data_o[58];
  assign data_o[25274] = data_o[58];
  assign data_o[25338] = data_o[58];
  assign data_o[25402] = data_o[58];
  assign data_o[25466] = data_o[58];
  assign data_o[25530] = data_o[58];
  assign data_o[25594] = data_o[58];
  assign data_o[25658] = data_o[58];
  assign data_o[25722] = data_o[58];
  assign data_o[25786] = data_o[58];
  assign data_o[25850] = data_o[58];
  assign data_o[25914] = data_o[58];
  assign data_o[25978] = data_o[58];
  assign data_o[26042] = data_o[58];
  assign data_o[26106] = data_o[58];
  assign data_o[26170] = data_o[58];
  assign data_o[26234] = data_o[58];
  assign data_o[26298] = data_o[58];
  assign data_o[26362] = data_o[58];
  assign data_o[26426] = data_o[58];
  assign data_o[26490] = data_o[58];
  assign data_o[26554] = data_o[58];
  assign data_o[26618] = data_o[58];
  assign data_o[26682] = data_o[58];
  assign data_o[26746] = data_o[58];
  assign data_o[26810] = data_o[58];
  assign data_o[26874] = data_o[58];
  assign data_o[26938] = data_o[58];
  assign data_o[27002] = data_o[58];
  assign data_o[27066] = data_o[58];
  assign data_o[27130] = data_o[58];
  assign data_o[27194] = data_o[58];
  assign data_o[27258] = data_o[58];
  assign data_o[27322] = data_o[58];
  assign data_o[27386] = data_o[58];
  assign data_o[27450] = data_o[58];
  assign data_o[27514] = data_o[58];
  assign data_o[27578] = data_o[58];
  assign data_o[27642] = data_o[58];
  assign data_o[27706] = data_o[58];
  assign data_o[27770] = data_o[58];
  assign data_o[27834] = data_o[58];
  assign data_o[27898] = data_o[58];
  assign data_o[27962] = data_o[58];
  assign data_o[28026] = data_o[58];
  assign data_o[28090] = data_o[58];
  assign data_o[28154] = data_o[58];
  assign data_o[28218] = data_o[58];
  assign data_o[28282] = data_o[58];
  assign data_o[28346] = data_o[58];
  assign data_o[28410] = data_o[58];
  assign data_o[28474] = data_o[58];
  assign data_o[28538] = data_o[58];
  assign data_o[28602] = data_o[58];
  assign data_o[28666] = data_o[58];
  assign data_o[28730] = data_o[58];
  assign data_o[28794] = data_o[58];
  assign data_o[28858] = data_o[58];
  assign data_o[28922] = data_o[58];
  assign data_o[28986] = data_o[58];
  assign data_o[29050] = data_o[58];
  assign data_o[29114] = data_o[58];
  assign data_o[29178] = data_o[58];
  assign data_o[29242] = data_o[58];
  assign data_o[29306] = data_o[58];
  assign data_o[29370] = data_o[58];
  assign data_o[29434] = data_o[58];
  assign data_o[29498] = data_o[58];
  assign data_o[29562] = data_o[58];
  assign data_o[29626] = data_o[58];
  assign data_o[29690] = data_o[58];
  assign data_o[29754] = data_o[58];
  assign data_o[29818] = data_o[58];
  assign data_o[29882] = data_o[58];
  assign data_o[29946] = data_o[58];
  assign data_o[30010] = data_o[58];
  assign data_o[30074] = data_o[58];
  assign data_o[30138] = data_o[58];
  assign data_o[30202] = data_o[58];
  assign data_o[30266] = data_o[58];
  assign data_o[30330] = data_o[58];
  assign data_o[30394] = data_o[58];
  assign data_o[30458] = data_o[58];
  assign data_o[30522] = data_o[58];
  assign data_o[30586] = data_o[58];
  assign data_o[30650] = data_o[58];
  assign data_o[30714] = data_o[58];
  assign data_o[30778] = data_o[58];
  assign data_o[30842] = data_o[58];
  assign data_o[30906] = data_o[58];
  assign data_o[30970] = data_o[58];
  assign data_o[31034] = data_o[58];
  assign data_o[31098] = data_o[58];
  assign data_o[31162] = data_o[58];
  assign data_o[31226] = data_o[58];
  assign data_o[31290] = data_o[58];
  assign data_o[31354] = data_o[58];
  assign data_o[31418] = data_o[58];
  assign data_o[31482] = data_o[58];
  assign data_o[31546] = data_o[58];
  assign data_o[31610] = data_o[58];
  assign data_o[31674] = data_o[58];
  assign data_o[31738] = data_o[58];
  assign data_o[31802] = data_o[58];
  assign data_o[31866] = data_o[58];
  assign data_o[31930] = data_o[58];
  assign data_o[31994] = data_o[58];
  assign data_o[121] = data_o[57];
  assign data_o[185] = data_o[57];
  assign data_o[249] = data_o[57];
  assign data_o[313] = data_o[57];
  assign data_o[377] = data_o[57];
  assign data_o[441] = data_o[57];
  assign data_o[505] = data_o[57];
  assign data_o[569] = data_o[57];
  assign data_o[633] = data_o[57];
  assign data_o[697] = data_o[57];
  assign data_o[761] = data_o[57];
  assign data_o[825] = data_o[57];
  assign data_o[889] = data_o[57];
  assign data_o[953] = data_o[57];
  assign data_o[1017] = data_o[57];
  assign data_o[1081] = data_o[57];
  assign data_o[1145] = data_o[57];
  assign data_o[1209] = data_o[57];
  assign data_o[1273] = data_o[57];
  assign data_o[1337] = data_o[57];
  assign data_o[1401] = data_o[57];
  assign data_o[1465] = data_o[57];
  assign data_o[1529] = data_o[57];
  assign data_o[1593] = data_o[57];
  assign data_o[1657] = data_o[57];
  assign data_o[1721] = data_o[57];
  assign data_o[1785] = data_o[57];
  assign data_o[1849] = data_o[57];
  assign data_o[1913] = data_o[57];
  assign data_o[1977] = data_o[57];
  assign data_o[2041] = data_o[57];
  assign data_o[2105] = data_o[57];
  assign data_o[2169] = data_o[57];
  assign data_o[2233] = data_o[57];
  assign data_o[2297] = data_o[57];
  assign data_o[2361] = data_o[57];
  assign data_o[2425] = data_o[57];
  assign data_o[2489] = data_o[57];
  assign data_o[2553] = data_o[57];
  assign data_o[2617] = data_o[57];
  assign data_o[2681] = data_o[57];
  assign data_o[2745] = data_o[57];
  assign data_o[2809] = data_o[57];
  assign data_o[2873] = data_o[57];
  assign data_o[2937] = data_o[57];
  assign data_o[3001] = data_o[57];
  assign data_o[3065] = data_o[57];
  assign data_o[3129] = data_o[57];
  assign data_o[3193] = data_o[57];
  assign data_o[3257] = data_o[57];
  assign data_o[3321] = data_o[57];
  assign data_o[3385] = data_o[57];
  assign data_o[3449] = data_o[57];
  assign data_o[3513] = data_o[57];
  assign data_o[3577] = data_o[57];
  assign data_o[3641] = data_o[57];
  assign data_o[3705] = data_o[57];
  assign data_o[3769] = data_o[57];
  assign data_o[3833] = data_o[57];
  assign data_o[3897] = data_o[57];
  assign data_o[3961] = data_o[57];
  assign data_o[4025] = data_o[57];
  assign data_o[4089] = data_o[57];
  assign data_o[4153] = data_o[57];
  assign data_o[4217] = data_o[57];
  assign data_o[4281] = data_o[57];
  assign data_o[4345] = data_o[57];
  assign data_o[4409] = data_o[57];
  assign data_o[4473] = data_o[57];
  assign data_o[4537] = data_o[57];
  assign data_o[4601] = data_o[57];
  assign data_o[4665] = data_o[57];
  assign data_o[4729] = data_o[57];
  assign data_o[4793] = data_o[57];
  assign data_o[4857] = data_o[57];
  assign data_o[4921] = data_o[57];
  assign data_o[4985] = data_o[57];
  assign data_o[5049] = data_o[57];
  assign data_o[5113] = data_o[57];
  assign data_o[5177] = data_o[57];
  assign data_o[5241] = data_o[57];
  assign data_o[5305] = data_o[57];
  assign data_o[5369] = data_o[57];
  assign data_o[5433] = data_o[57];
  assign data_o[5497] = data_o[57];
  assign data_o[5561] = data_o[57];
  assign data_o[5625] = data_o[57];
  assign data_o[5689] = data_o[57];
  assign data_o[5753] = data_o[57];
  assign data_o[5817] = data_o[57];
  assign data_o[5881] = data_o[57];
  assign data_o[5945] = data_o[57];
  assign data_o[6009] = data_o[57];
  assign data_o[6073] = data_o[57];
  assign data_o[6137] = data_o[57];
  assign data_o[6201] = data_o[57];
  assign data_o[6265] = data_o[57];
  assign data_o[6329] = data_o[57];
  assign data_o[6393] = data_o[57];
  assign data_o[6457] = data_o[57];
  assign data_o[6521] = data_o[57];
  assign data_o[6585] = data_o[57];
  assign data_o[6649] = data_o[57];
  assign data_o[6713] = data_o[57];
  assign data_o[6777] = data_o[57];
  assign data_o[6841] = data_o[57];
  assign data_o[6905] = data_o[57];
  assign data_o[6969] = data_o[57];
  assign data_o[7033] = data_o[57];
  assign data_o[7097] = data_o[57];
  assign data_o[7161] = data_o[57];
  assign data_o[7225] = data_o[57];
  assign data_o[7289] = data_o[57];
  assign data_o[7353] = data_o[57];
  assign data_o[7417] = data_o[57];
  assign data_o[7481] = data_o[57];
  assign data_o[7545] = data_o[57];
  assign data_o[7609] = data_o[57];
  assign data_o[7673] = data_o[57];
  assign data_o[7737] = data_o[57];
  assign data_o[7801] = data_o[57];
  assign data_o[7865] = data_o[57];
  assign data_o[7929] = data_o[57];
  assign data_o[7993] = data_o[57];
  assign data_o[8057] = data_o[57];
  assign data_o[8121] = data_o[57];
  assign data_o[8185] = data_o[57];
  assign data_o[8249] = data_o[57];
  assign data_o[8313] = data_o[57];
  assign data_o[8377] = data_o[57];
  assign data_o[8441] = data_o[57];
  assign data_o[8505] = data_o[57];
  assign data_o[8569] = data_o[57];
  assign data_o[8633] = data_o[57];
  assign data_o[8697] = data_o[57];
  assign data_o[8761] = data_o[57];
  assign data_o[8825] = data_o[57];
  assign data_o[8889] = data_o[57];
  assign data_o[8953] = data_o[57];
  assign data_o[9017] = data_o[57];
  assign data_o[9081] = data_o[57];
  assign data_o[9145] = data_o[57];
  assign data_o[9209] = data_o[57];
  assign data_o[9273] = data_o[57];
  assign data_o[9337] = data_o[57];
  assign data_o[9401] = data_o[57];
  assign data_o[9465] = data_o[57];
  assign data_o[9529] = data_o[57];
  assign data_o[9593] = data_o[57];
  assign data_o[9657] = data_o[57];
  assign data_o[9721] = data_o[57];
  assign data_o[9785] = data_o[57];
  assign data_o[9849] = data_o[57];
  assign data_o[9913] = data_o[57];
  assign data_o[9977] = data_o[57];
  assign data_o[10041] = data_o[57];
  assign data_o[10105] = data_o[57];
  assign data_o[10169] = data_o[57];
  assign data_o[10233] = data_o[57];
  assign data_o[10297] = data_o[57];
  assign data_o[10361] = data_o[57];
  assign data_o[10425] = data_o[57];
  assign data_o[10489] = data_o[57];
  assign data_o[10553] = data_o[57];
  assign data_o[10617] = data_o[57];
  assign data_o[10681] = data_o[57];
  assign data_o[10745] = data_o[57];
  assign data_o[10809] = data_o[57];
  assign data_o[10873] = data_o[57];
  assign data_o[10937] = data_o[57];
  assign data_o[11001] = data_o[57];
  assign data_o[11065] = data_o[57];
  assign data_o[11129] = data_o[57];
  assign data_o[11193] = data_o[57];
  assign data_o[11257] = data_o[57];
  assign data_o[11321] = data_o[57];
  assign data_o[11385] = data_o[57];
  assign data_o[11449] = data_o[57];
  assign data_o[11513] = data_o[57];
  assign data_o[11577] = data_o[57];
  assign data_o[11641] = data_o[57];
  assign data_o[11705] = data_o[57];
  assign data_o[11769] = data_o[57];
  assign data_o[11833] = data_o[57];
  assign data_o[11897] = data_o[57];
  assign data_o[11961] = data_o[57];
  assign data_o[12025] = data_o[57];
  assign data_o[12089] = data_o[57];
  assign data_o[12153] = data_o[57];
  assign data_o[12217] = data_o[57];
  assign data_o[12281] = data_o[57];
  assign data_o[12345] = data_o[57];
  assign data_o[12409] = data_o[57];
  assign data_o[12473] = data_o[57];
  assign data_o[12537] = data_o[57];
  assign data_o[12601] = data_o[57];
  assign data_o[12665] = data_o[57];
  assign data_o[12729] = data_o[57];
  assign data_o[12793] = data_o[57];
  assign data_o[12857] = data_o[57];
  assign data_o[12921] = data_o[57];
  assign data_o[12985] = data_o[57];
  assign data_o[13049] = data_o[57];
  assign data_o[13113] = data_o[57];
  assign data_o[13177] = data_o[57];
  assign data_o[13241] = data_o[57];
  assign data_o[13305] = data_o[57];
  assign data_o[13369] = data_o[57];
  assign data_o[13433] = data_o[57];
  assign data_o[13497] = data_o[57];
  assign data_o[13561] = data_o[57];
  assign data_o[13625] = data_o[57];
  assign data_o[13689] = data_o[57];
  assign data_o[13753] = data_o[57];
  assign data_o[13817] = data_o[57];
  assign data_o[13881] = data_o[57];
  assign data_o[13945] = data_o[57];
  assign data_o[14009] = data_o[57];
  assign data_o[14073] = data_o[57];
  assign data_o[14137] = data_o[57];
  assign data_o[14201] = data_o[57];
  assign data_o[14265] = data_o[57];
  assign data_o[14329] = data_o[57];
  assign data_o[14393] = data_o[57];
  assign data_o[14457] = data_o[57];
  assign data_o[14521] = data_o[57];
  assign data_o[14585] = data_o[57];
  assign data_o[14649] = data_o[57];
  assign data_o[14713] = data_o[57];
  assign data_o[14777] = data_o[57];
  assign data_o[14841] = data_o[57];
  assign data_o[14905] = data_o[57];
  assign data_o[14969] = data_o[57];
  assign data_o[15033] = data_o[57];
  assign data_o[15097] = data_o[57];
  assign data_o[15161] = data_o[57];
  assign data_o[15225] = data_o[57];
  assign data_o[15289] = data_o[57];
  assign data_o[15353] = data_o[57];
  assign data_o[15417] = data_o[57];
  assign data_o[15481] = data_o[57];
  assign data_o[15545] = data_o[57];
  assign data_o[15609] = data_o[57];
  assign data_o[15673] = data_o[57];
  assign data_o[15737] = data_o[57];
  assign data_o[15801] = data_o[57];
  assign data_o[15865] = data_o[57];
  assign data_o[15929] = data_o[57];
  assign data_o[15993] = data_o[57];
  assign data_o[16057] = data_o[57];
  assign data_o[16121] = data_o[57];
  assign data_o[16185] = data_o[57];
  assign data_o[16249] = data_o[57];
  assign data_o[16313] = data_o[57];
  assign data_o[16377] = data_o[57];
  assign data_o[16441] = data_o[57];
  assign data_o[16505] = data_o[57];
  assign data_o[16569] = data_o[57];
  assign data_o[16633] = data_o[57];
  assign data_o[16697] = data_o[57];
  assign data_o[16761] = data_o[57];
  assign data_o[16825] = data_o[57];
  assign data_o[16889] = data_o[57];
  assign data_o[16953] = data_o[57];
  assign data_o[17017] = data_o[57];
  assign data_o[17081] = data_o[57];
  assign data_o[17145] = data_o[57];
  assign data_o[17209] = data_o[57];
  assign data_o[17273] = data_o[57];
  assign data_o[17337] = data_o[57];
  assign data_o[17401] = data_o[57];
  assign data_o[17465] = data_o[57];
  assign data_o[17529] = data_o[57];
  assign data_o[17593] = data_o[57];
  assign data_o[17657] = data_o[57];
  assign data_o[17721] = data_o[57];
  assign data_o[17785] = data_o[57];
  assign data_o[17849] = data_o[57];
  assign data_o[17913] = data_o[57];
  assign data_o[17977] = data_o[57];
  assign data_o[18041] = data_o[57];
  assign data_o[18105] = data_o[57];
  assign data_o[18169] = data_o[57];
  assign data_o[18233] = data_o[57];
  assign data_o[18297] = data_o[57];
  assign data_o[18361] = data_o[57];
  assign data_o[18425] = data_o[57];
  assign data_o[18489] = data_o[57];
  assign data_o[18553] = data_o[57];
  assign data_o[18617] = data_o[57];
  assign data_o[18681] = data_o[57];
  assign data_o[18745] = data_o[57];
  assign data_o[18809] = data_o[57];
  assign data_o[18873] = data_o[57];
  assign data_o[18937] = data_o[57];
  assign data_o[19001] = data_o[57];
  assign data_o[19065] = data_o[57];
  assign data_o[19129] = data_o[57];
  assign data_o[19193] = data_o[57];
  assign data_o[19257] = data_o[57];
  assign data_o[19321] = data_o[57];
  assign data_o[19385] = data_o[57];
  assign data_o[19449] = data_o[57];
  assign data_o[19513] = data_o[57];
  assign data_o[19577] = data_o[57];
  assign data_o[19641] = data_o[57];
  assign data_o[19705] = data_o[57];
  assign data_o[19769] = data_o[57];
  assign data_o[19833] = data_o[57];
  assign data_o[19897] = data_o[57];
  assign data_o[19961] = data_o[57];
  assign data_o[20025] = data_o[57];
  assign data_o[20089] = data_o[57];
  assign data_o[20153] = data_o[57];
  assign data_o[20217] = data_o[57];
  assign data_o[20281] = data_o[57];
  assign data_o[20345] = data_o[57];
  assign data_o[20409] = data_o[57];
  assign data_o[20473] = data_o[57];
  assign data_o[20537] = data_o[57];
  assign data_o[20601] = data_o[57];
  assign data_o[20665] = data_o[57];
  assign data_o[20729] = data_o[57];
  assign data_o[20793] = data_o[57];
  assign data_o[20857] = data_o[57];
  assign data_o[20921] = data_o[57];
  assign data_o[20985] = data_o[57];
  assign data_o[21049] = data_o[57];
  assign data_o[21113] = data_o[57];
  assign data_o[21177] = data_o[57];
  assign data_o[21241] = data_o[57];
  assign data_o[21305] = data_o[57];
  assign data_o[21369] = data_o[57];
  assign data_o[21433] = data_o[57];
  assign data_o[21497] = data_o[57];
  assign data_o[21561] = data_o[57];
  assign data_o[21625] = data_o[57];
  assign data_o[21689] = data_o[57];
  assign data_o[21753] = data_o[57];
  assign data_o[21817] = data_o[57];
  assign data_o[21881] = data_o[57];
  assign data_o[21945] = data_o[57];
  assign data_o[22009] = data_o[57];
  assign data_o[22073] = data_o[57];
  assign data_o[22137] = data_o[57];
  assign data_o[22201] = data_o[57];
  assign data_o[22265] = data_o[57];
  assign data_o[22329] = data_o[57];
  assign data_o[22393] = data_o[57];
  assign data_o[22457] = data_o[57];
  assign data_o[22521] = data_o[57];
  assign data_o[22585] = data_o[57];
  assign data_o[22649] = data_o[57];
  assign data_o[22713] = data_o[57];
  assign data_o[22777] = data_o[57];
  assign data_o[22841] = data_o[57];
  assign data_o[22905] = data_o[57];
  assign data_o[22969] = data_o[57];
  assign data_o[23033] = data_o[57];
  assign data_o[23097] = data_o[57];
  assign data_o[23161] = data_o[57];
  assign data_o[23225] = data_o[57];
  assign data_o[23289] = data_o[57];
  assign data_o[23353] = data_o[57];
  assign data_o[23417] = data_o[57];
  assign data_o[23481] = data_o[57];
  assign data_o[23545] = data_o[57];
  assign data_o[23609] = data_o[57];
  assign data_o[23673] = data_o[57];
  assign data_o[23737] = data_o[57];
  assign data_o[23801] = data_o[57];
  assign data_o[23865] = data_o[57];
  assign data_o[23929] = data_o[57];
  assign data_o[23993] = data_o[57];
  assign data_o[24057] = data_o[57];
  assign data_o[24121] = data_o[57];
  assign data_o[24185] = data_o[57];
  assign data_o[24249] = data_o[57];
  assign data_o[24313] = data_o[57];
  assign data_o[24377] = data_o[57];
  assign data_o[24441] = data_o[57];
  assign data_o[24505] = data_o[57];
  assign data_o[24569] = data_o[57];
  assign data_o[24633] = data_o[57];
  assign data_o[24697] = data_o[57];
  assign data_o[24761] = data_o[57];
  assign data_o[24825] = data_o[57];
  assign data_o[24889] = data_o[57];
  assign data_o[24953] = data_o[57];
  assign data_o[25017] = data_o[57];
  assign data_o[25081] = data_o[57];
  assign data_o[25145] = data_o[57];
  assign data_o[25209] = data_o[57];
  assign data_o[25273] = data_o[57];
  assign data_o[25337] = data_o[57];
  assign data_o[25401] = data_o[57];
  assign data_o[25465] = data_o[57];
  assign data_o[25529] = data_o[57];
  assign data_o[25593] = data_o[57];
  assign data_o[25657] = data_o[57];
  assign data_o[25721] = data_o[57];
  assign data_o[25785] = data_o[57];
  assign data_o[25849] = data_o[57];
  assign data_o[25913] = data_o[57];
  assign data_o[25977] = data_o[57];
  assign data_o[26041] = data_o[57];
  assign data_o[26105] = data_o[57];
  assign data_o[26169] = data_o[57];
  assign data_o[26233] = data_o[57];
  assign data_o[26297] = data_o[57];
  assign data_o[26361] = data_o[57];
  assign data_o[26425] = data_o[57];
  assign data_o[26489] = data_o[57];
  assign data_o[26553] = data_o[57];
  assign data_o[26617] = data_o[57];
  assign data_o[26681] = data_o[57];
  assign data_o[26745] = data_o[57];
  assign data_o[26809] = data_o[57];
  assign data_o[26873] = data_o[57];
  assign data_o[26937] = data_o[57];
  assign data_o[27001] = data_o[57];
  assign data_o[27065] = data_o[57];
  assign data_o[27129] = data_o[57];
  assign data_o[27193] = data_o[57];
  assign data_o[27257] = data_o[57];
  assign data_o[27321] = data_o[57];
  assign data_o[27385] = data_o[57];
  assign data_o[27449] = data_o[57];
  assign data_o[27513] = data_o[57];
  assign data_o[27577] = data_o[57];
  assign data_o[27641] = data_o[57];
  assign data_o[27705] = data_o[57];
  assign data_o[27769] = data_o[57];
  assign data_o[27833] = data_o[57];
  assign data_o[27897] = data_o[57];
  assign data_o[27961] = data_o[57];
  assign data_o[28025] = data_o[57];
  assign data_o[28089] = data_o[57];
  assign data_o[28153] = data_o[57];
  assign data_o[28217] = data_o[57];
  assign data_o[28281] = data_o[57];
  assign data_o[28345] = data_o[57];
  assign data_o[28409] = data_o[57];
  assign data_o[28473] = data_o[57];
  assign data_o[28537] = data_o[57];
  assign data_o[28601] = data_o[57];
  assign data_o[28665] = data_o[57];
  assign data_o[28729] = data_o[57];
  assign data_o[28793] = data_o[57];
  assign data_o[28857] = data_o[57];
  assign data_o[28921] = data_o[57];
  assign data_o[28985] = data_o[57];
  assign data_o[29049] = data_o[57];
  assign data_o[29113] = data_o[57];
  assign data_o[29177] = data_o[57];
  assign data_o[29241] = data_o[57];
  assign data_o[29305] = data_o[57];
  assign data_o[29369] = data_o[57];
  assign data_o[29433] = data_o[57];
  assign data_o[29497] = data_o[57];
  assign data_o[29561] = data_o[57];
  assign data_o[29625] = data_o[57];
  assign data_o[29689] = data_o[57];
  assign data_o[29753] = data_o[57];
  assign data_o[29817] = data_o[57];
  assign data_o[29881] = data_o[57];
  assign data_o[29945] = data_o[57];
  assign data_o[30009] = data_o[57];
  assign data_o[30073] = data_o[57];
  assign data_o[30137] = data_o[57];
  assign data_o[30201] = data_o[57];
  assign data_o[30265] = data_o[57];
  assign data_o[30329] = data_o[57];
  assign data_o[30393] = data_o[57];
  assign data_o[30457] = data_o[57];
  assign data_o[30521] = data_o[57];
  assign data_o[30585] = data_o[57];
  assign data_o[30649] = data_o[57];
  assign data_o[30713] = data_o[57];
  assign data_o[30777] = data_o[57];
  assign data_o[30841] = data_o[57];
  assign data_o[30905] = data_o[57];
  assign data_o[30969] = data_o[57];
  assign data_o[31033] = data_o[57];
  assign data_o[31097] = data_o[57];
  assign data_o[31161] = data_o[57];
  assign data_o[31225] = data_o[57];
  assign data_o[31289] = data_o[57];
  assign data_o[31353] = data_o[57];
  assign data_o[31417] = data_o[57];
  assign data_o[31481] = data_o[57];
  assign data_o[31545] = data_o[57];
  assign data_o[31609] = data_o[57];
  assign data_o[31673] = data_o[57];
  assign data_o[31737] = data_o[57];
  assign data_o[31801] = data_o[57];
  assign data_o[31865] = data_o[57];
  assign data_o[31929] = data_o[57];
  assign data_o[31993] = data_o[57];
  assign data_o[120] = data_o[56];
  assign data_o[184] = data_o[56];
  assign data_o[248] = data_o[56];
  assign data_o[312] = data_o[56];
  assign data_o[376] = data_o[56];
  assign data_o[440] = data_o[56];
  assign data_o[504] = data_o[56];
  assign data_o[568] = data_o[56];
  assign data_o[632] = data_o[56];
  assign data_o[696] = data_o[56];
  assign data_o[760] = data_o[56];
  assign data_o[824] = data_o[56];
  assign data_o[888] = data_o[56];
  assign data_o[952] = data_o[56];
  assign data_o[1016] = data_o[56];
  assign data_o[1080] = data_o[56];
  assign data_o[1144] = data_o[56];
  assign data_o[1208] = data_o[56];
  assign data_o[1272] = data_o[56];
  assign data_o[1336] = data_o[56];
  assign data_o[1400] = data_o[56];
  assign data_o[1464] = data_o[56];
  assign data_o[1528] = data_o[56];
  assign data_o[1592] = data_o[56];
  assign data_o[1656] = data_o[56];
  assign data_o[1720] = data_o[56];
  assign data_o[1784] = data_o[56];
  assign data_o[1848] = data_o[56];
  assign data_o[1912] = data_o[56];
  assign data_o[1976] = data_o[56];
  assign data_o[2040] = data_o[56];
  assign data_o[2104] = data_o[56];
  assign data_o[2168] = data_o[56];
  assign data_o[2232] = data_o[56];
  assign data_o[2296] = data_o[56];
  assign data_o[2360] = data_o[56];
  assign data_o[2424] = data_o[56];
  assign data_o[2488] = data_o[56];
  assign data_o[2552] = data_o[56];
  assign data_o[2616] = data_o[56];
  assign data_o[2680] = data_o[56];
  assign data_o[2744] = data_o[56];
  assign data_o[2808] = data_o[56];
  assign data_o[2872] = data_o[56];
  assign data_o[2936] = data_o[56];
  assign data_o[3000] = data_o[56];
  assign data_o[3064] = data_o[56];
  assign data_o[3128] = data_o[56];
  assign data_o[3192] = data_o[56];
  assign data_o[3256] = data_o[56];
  assign data_o[3320] = data_o[56];
  assign data_o[3384] = data_o[56];
  assign data_o[3448] = data_o[56];
  assign data_o[3512] = data_o[56];
  assign data_o[3576] = data_o[56];
  assign data_o[3640] = data_o[56];
  assign data_o[3704] = data_o[56];
  assign data_o[3768] = data_o[56];
  assign data_o[3832] = data_o[56];
  assign data_o[3896] = data_o[56];
  assign data_o[3960] = data_o[56];
  assign data_o[4024] = data_o[56];
  assign data_o[4088] = data_o[56];
  assign data_o[4152] = data_o[56];
  assign data_o[4216] = data_o[56];
  assign data_o[4280] = data_o[56];
  assign data_o[4344] = data_o[56];
  assign data_o[4408] = data_o[56];
  assign data_o[4472] = data_o[56];
  assign data_o[4536] = data_o[56];
  assign data_o[4600] = data_o[56];
  assign data_o[4664] = data_o[56];
  assign data_o[4728] = data_o[56];
  assign data_o[4792] = data_o[56];
  assign data_o[4856] = data_o[56];
  assign data_o[4920] = data_o[56];
  assign data_o[4984] = data_o[56];
  assign data_o[5048] = data_o[56];
  assign data_o[5112] = data_o[56];
  assign data_o[5176] = data_o[56];
  assign data_o[5240] = data_o[56];
  assign data_o[5304] = data_o[56];
  assign data_o[5368] = data_o[56];
  assign data_o[5432] = data_o[56];
  assign data_o[5496] = data_o[56];
  assign data_o[5560] = data_o[56];
  assign data_o[5624] = data_o[56];
  assign data_o[5688] = data_o[56];
  assign data_o[5752] = data_o[56];
  assign data_o[5816] = data_o[56];
  assign data_o[5880] = data_o[56];
  assign data_o[5944] = data_o[56];
  assign data_o[6008] = data_o[56];
  assign data_o[6072] = data_o[56];
  assign data_o[6136] = data_o[56];
  assign data_o[6200] = data_o[56];
  assign data_o[6264] = data_o[56];
  assign data_o[6328] = data_o[56];
  assign data_o[6392] = data_o[56];
  assign data_o[6456] = data_o[56];
  assign data_o[6520] = data_o[56];
  assign data_o[6584] = data_o[56];
  assign data_o[6648] = data_o[56];
  assign data_o[6712] = data_o[56];
  assign data_o[6776] = data_o[56];
  assign data_o[6840] = data_o[56];
  assign data_o[6904] = data_o[56];
  assign data_o[6968] = data_o[56];
  assign data_o[7032] = data_o[56];
  assign data_o[7096] = data_o[56];
  assign data_o[7160] = data_o[56];
  assign data_o[7224] = data_o[56];
  assign data_o[7288] = data_o[56];
  assign data_o[7352] = data_o[56];
  assign data_o[7416] = data_o[56];
  assign data_o[7480] = data_o[56];
  assign data_o[7544] = data_o[56];
  assign data_o[7608] = data_o[56];
  assign data_o[7672] = data_o[56];
  assign data_o[7736] = data_o[56];
  assign data_o[7800] = data_o[56];
  assign data_o[7864] = data_o[56];
  assign data_o[7928] = data_o[56];
  assign data_o[7992] = data_o[56];
  assign data_o[8056] = data_o[56];
  assign data_o[8120] = data_o[56];
  assign data_o[8184] = data_o[56];
  assign data_o[8248] = data_o[56];
  assign data_o[8312] = data_o[56];
  assign data_o[8376] = data_o[56];
  assign data_o[8440] = data_o[56];
  assign data_o[8504] = data_o[56];
  assign data_o[8568] = data_o[56];
  assign data_o[8632] = data_o[56];
  assign data_o[8696] = data_o[56];
  assign data_o[8760] = data_o[56];
  assign data_o[8824] = data_o[56];
  assign data_o[8888] = data_o[56];
  assign data_o[8952] = data_o[56];
  assign data_o[9016] = data_o[56];
  assign data_o[9080] = data_o[56];
  assign data_o[9144] = data_o[56];
  assign data_o[9208] = data_o[56];
  assign data_o[9272] = data_o[56];
  assign data_o[9336] = data_o[56];
  assign data_o[9400] = data_o[56];
  assign data_o[9464] = data_o[56];
  assign data_o[9528] = data_o[56];
  assign data_o[9592] = data_o[56];
  assign data_o[9656] = data_o[56];
  assign data_o[9720] = data_o[56];
  assign data_o[9784] = data_o[56];
  assign data_o[9848] = data_o[56];
  assign data_o[9912] = data_o[56];
  assign data_o[9976] = data_o[56];
  assign data_o[10040] = data_o[56];
  assign data_o[10104] = data_o[56];
  assign data_o[10168] = data_o[56];
  assign data_o[10232] = data_o[56];
  assign data_o[10296] = data_o[56];
  assign data_o[10360] = data_o[56];
  assign data_o[10424] = data_o[56];
  assign data_o[10488] = data_o[56];
  assign data_o[10552] = data_o[56];
  assign data_o[10616] = data_o[56];
  assign data_o[10680] = data_o[56];
  assign data_o[10744] = data_o[56];
  assign data_o[10808] = data_o[56];
  assign data_o[10872] = data_o[56];
  assign data_o[10936] = data_o[56];
  assign data_o[11000] = data_o[56];
  assign data_o[11064] = data_o[56];
  assign data_o[11128] = data_o[56];
  assign data_o[11192] = data_o[56];
  assign data_o[11256] = data_o[56];
  assign data_o[11320] = data_o[56];
  assign data_o[11384] = data_o[56];
  assign data_o[11448] = data_o[56];
  assign data_o[11512] = data_o[56];
  assign data_o[11576] = data_o[56];
  assign data_o[11640] = data_o[56];
  assign data_o[11704] = data_o[56];
  assign data_o[11768] = data_o[56];
  assign data_o[11832] = data_o[56];
  assign data_o[11896] = data_o[56];
  assign data_o[11960] = data_o[56];
  assign data_o[12024] = data_o[56];
  assign data_o[12088] = data_o[56];
  assign data_o[12152] = data_o[56];
  assign data_o[12216] = data_o[56];
  assign data_o[12280] = data_o[56];
  assign data_o[12344] = data_o[56];
  assign data_o[12408] = data_o[56];
  assign data_o[12472] = data_o[56];
  assign data_o[12536] = data_o[56];
  assign data_o[12600] = data_o[56];
  assign data_o[12664] = data_o[56];
  assign data_o[12728] = data_o[56];
  assign data_o[12792] = data_o[56];
  assign data_o[12856] = data_o[56];
  assign data_o[12920] = data_o[56];
  assign data_o[12984] = data_o[56];
  assign data_o[13048] = data_o[56];
  assign data_o[13112] = data_o[56];
  assign data_o[13176] = data_o[56];
  assign data_o[13240] = data_o[56];
  assign data_o[13304] = data_o[56];
  assign data_o[13368] = data_o[56];
  assign data_o[13432] = data_o[56];
  assign data_o[13496] = data_o[56];
  assign data_o[13560] = data_o[56];
  assign data_o[13624] = data_o[56];
  assign data_o[13688] = data_o[56];
  assign data_o[13752] = data_o[56];
  assign data_o[13816] = data_o[56];
  assign data_o[13880] = data_o[56];
  assign data_o[13944] = data_o[56];
  assign data_o[14008] = data_o[56];
  assign data_o[14072] = data_o[56];
  assign data_o[14136] = data_o[56];
  assign data_o[14200] = data_o[56];
  assign data_o[14264] = data_o[56];
  assign data_o[14328] = data_o[56];
  assign data_o[14392] = data_o[56];
  assign data_o[14456] = data_o[56];
  assign data_o[14520] = data_o[56];
  assign data_o[14584] = data_o[56];
  assign data_o[14648] = data_o[56];
  assign data_o[14712] = data_o[56];
  assign data_o[14776] = data_o[56];
  assign data_o[14840] = data_o[56];
  assign data_o[14904] = data_o[56];
  assign data_o[14968] = data_o[56];
  assign data_o[15032] = data_o[56];
  assign data_o[15096] = data_o[56];
  assign data_o[15160] = data_o[56];
  assign data_o[15224] = data_o[56];
  assign data_o[15288] = data_o[56];
  assign data_o[15352] = data_o[56];
  assign data_o[15416] = data_o[56];
  assign data_o[15480] = data_o[56];
  assign data_o[15544] = data_o[56];
  assign data_o[15608] = data_o[56];
  assign data_o[15672] = data_o[56];
  assign data_o[15736] = data_o[56];
  assign data_o[15800] = data_o[56];
  assign data_o[15864] = data_o[56];
  assign data_o[15928] = data_o[56];
  assign data_o[15992] = data_o[56];
  assign data_o[16056] = data_o[56];
  assign data_o[16120] = data_o[56];
  assign data_o[16184] = data_o[56];
  assign data_o[16248] = data_o[56];
  assign data_o[16312] = data_o[56];
  assign data_o[16376] = data_o[56];
  assign data_o[16440] = data_o[56];
  assign data_o[16504] = data_o[56];
  assign data_o[16568] = data_o[56];
  assign data_o[16632] = data_o[56];
  assign data_o[16696] = data_o[56];
  assign data_o[16760] = data_o[56];
  assign data_o[16824] = data_o[56];
  assign data_o[16888] = data_o[56];
  assign data_o[16952] = data_o[56];
  assign data_o[17016] = data_o[56];
  assign data_o[17080] = data_o[56];
  assign data_o[17144] = data_o[56];
  assign data_o[17208] = data_o[56];
  assign data_o[17272] = data_o[56];
  assign data_o[17336] = data_o[56];
  assign data_o[17400] = data_o[56];
  assign data_o[17464] = data_o[56];
  assign data_o[17528] = data_o[56];
  assign data_o[17592] = data_o[56];
  assign data_o[17656] = data_o[56];
  assign data_o[17720] = data_o[56];
  assign data_o[17784] = data_o[56];
  assign data_o[17848] = data_o[56];
  assign data_o[17912] = data_o[56];
  assign data_o[17976] = data_o[56];
  assign data_o[18040] = data_o[56];
  assign data_o[18104] = data_o[56];
  assign data_o[18168] = data_o[56];
  assign data_o[18232] = data_o[56];
  assign data_o[18296] = data_o[56];
  assign data_o[18360] = data_o[56];
  assign data_o[18424] = data_o[56];
  assign data_o[18488] = data_o[56];
  assign data_o[18552] = data_o[56];
  assign data_o[18616] = data_o[56];
  assign data_o[18680] = data_o[56];
  assign data_o[18744] = data_o[56];
  assign data_o[18808] = data_o[56];
  assign data_o[18872] = data_o[56];
  assign data_o[18936] = data_o[56];
  assign data_o[19000] = data_o[56];
  assign data_o[19064] = data_o[56];
  assign data_o[19128] = data_o[56];
  assign data_o[19192] = data_o[56];
  assign data_o[19256] = data_o[56];
  assign data_o[19320] = data_o[56];
  assign data_o[19384] = data_o[56];
  assign data_o[19448] = data_o[56];
  assign data_o[19512] = data_o[56];
  assign data_o[19576] = data_o[56];
  assign data_o[19640] = data_o[56];
  assign data_o[19704] = data_o[56];
  assign data_o[19768] = data_o[56];
  assign data_o[19832] = data_o[56];
  assign data_o[19896] = data_o[56];
  assign data_o[19960] = data_o[56];
  assign data_o[20024] = data_o[56];
  assign data_o[20088] = data_o[56];
  assign data_o[20152] = data_o[56];
  assign data_o[20216] = data_o[56];
  assign data_o[20280] = data_o[56];
  assign data_o[20344] = data_o[56];
  assign data_o[20408] = data_o[56];
  assign data_o[20472] = data_o[56];
  assign data_o[20536] = data_o[56];
  assign data_o[20600] = data_o[56];
  assign data_o[20664] = data_o[56];
  assign data_o[20728] = data_o[56];
  assign data_o[20792] = data_o[56];
  assign data_o[20856] = data_o[56];
  assign data_o[20920] = data_o[56];
  assign data_o[20984] = data_o[56];
  assign data_o[21048] = data_o[56];
  assign data_o[21112] = data_o[56];
  assign data_o[21176] = data_o[56];
  assign data_o[21240] = data_o[56];
  assign data_o[21304] = data_o[56];
  assign data_o[21368] = data_o[56];
  assign data_o[21432] = data_o[56];
  assign data_o[21496] = data_o[56];
  assign data_o[21560] = data_o[56];
  assign data_o[21624] = data_o[56];
  assign data_o[21688] = data_o[56];
  assign data_o[21752] = data_o[56];
  assign data_o[21816] = data_o[56];
  assign data_o[21880] = data_o[56];
  assign data_o[21944] = data_o[56];
  assign data_o[22008] = data_o[56];
  assign data_o[22072] = data_o[56];
  assign data_o[22136] = data_o[56];
  assign data_o[22200] = data_o[56];
  assign data_o[22264] = data_o[56];
  assign data_o[22328] = data_o[56];
  assign data_o[22392] = data_o[56];
  assign data_o[22456] = data_o[56];
  assign data_o[22520] = data_o[56];
  assign data_o[22584] = data_o[56];
  assign data_o[22648] = data_o[56];
  assign data_o[22712] = data_o[56];
  assign data_o[22776] = data_o[56];
  assign data_o[22840] = data_o[56];
  assign data_o[22904] = data_o[56];
  assign data_o[22968] = data_o[56];
  assign data_o[23032] = data_o[56];
  assign data_o[23096] = data_o[56];
  assign data_o[23160] = data_o[56];
  assign data_o[23224] = data_o[56];
  assign data_o[23288] = data_o[56];
  assign data_o[23352] = data_o[56];
  assign data_o[23416] = data_o[56];
  assign data_o[23480] = data_o[56];
  assign data_o[23544] = data_o[56];
  assign data_o[23608] = data_o[56];
  assign data_o[23672] = data_o[56];
  assign data_o[23736] = data_o[56];
  assign data_o[23800] = data_o[56];
  assign data_o[23864] = data_o[56];
  assign data_o[23928] = data_o[56];
  assign data_o[23992] = data_o[56];
  assign data_o[24056] = data_o[56];
  assign data_o[24120] = data_o[56];
  assign data_o[24184] = data_o[56];
  assign data_o[24248] = data_o[56];
  assign data_o[24312] = data_o[56];
  assign data_o[24376] = data_o[56];
  assign data_o[24440] = data_o[56];
  assign data_o[24504] = data_o[56];
  assign data_o[24568] = data_o[56];
  assign data_o[24632] = data_o[56];
  assign data_o[24696] = data_o[56];
  assign data_o[24760] = data_o[56];
  assign data_o[24824] = data_o[56];
  assign data_o[24888] = data_o[56];
  assign data_o[24952] = data_o[56];
  assign data_o[25016] = data_o[56];
  assign data_o[25080] = data_o[56];
  assign data_o[25144] = data_o[56];
  assign data_o[25208] = data_o[56];
  assign data_o[25272] = data_o[56];
  assign data_o[25336] = data_o[56];
  assign data_o[25400] = data_o[56];
  assign data_o[25464] = data_o[56];
  assign data_o[25528] = data_o[56];
  assign data_o[25592] = data_o[56];
  assign data_o[25656] = data_o[56];
  assign data_o[25720] = data_o[56];
  assign data_o[25784] = data_o[56];
  assign data_o[25848] = data_o[56];
  assign data_o[25912] = data_o[56];
  assign data_o[25976] = data_o[56];
  assign data_o[26040] = data_o[56];
  assign data_o[26104] = data_o[56];
  assign data_o[26168] = data_o[56];
  assign data_o[26232] = data_o[56];
  assign data_o[26296] = data_o[56];
  assign data_o[26360] = data_o[56];
  assign data_o[26424] = data_o[56];
  assign data_o[26488] = data_o[56];
  assign data_o[26552] = data_o[56];
  assign data_o[26616] = data_o[56];
  assign data_o[26680] = data_o[56];
  assign data_o[26744] = data_o[56];
  assign data_o[26808] = data_o[56];
  assign data_o[26872] = data_o[56];
  assign data_o[26936] = data_o[56];
  assign data_o[27000] = data_o[56];
  assign data_o[27064] = data_o[56];
  assign data_o[27128] = data_o[56];
  assign data_o[27192] = data_o[56];
  assign data_o[27256] = data_o[56];
  assign data_o[27320] = data_o[56];
  assign data_o[27384] = data_o[56];
  assign data_o[27448] = data_o[56];
  assign data_o[27512] = data_o[56];
  assign data_o[27576] = data_o[56];
  assign data_o[27640] = data_o[56];
  assign data_o[27704] = data_o[56];
  assign data_o[27768] = data_o[56];
  assign data_o[27832] = data_o[56];
  assign data_o[27896] = data_o[56];
  assign data_o[27960] = data_o[56];
  assign data_o[28024] = data_o[56];
  assign data_o[28088] = data_o[56];
  assign data_o[28152] = data_o[56];
  assign data_o[28216] = data_o[56];
  assign data_o[28280] = data_o[56];
  assign data_o[28344] = data_o[56];
  assign data_o[28408] = data_o[56];
  assign data_o[28472] = data_o[56];
  assign data_o[28536] = data_o[56];
  assign data_o[28600] = data_o[56];
  assign data_o[28664] = data_o[56];
  assign data_o[28728] = data_o[56];
  assign data_o[28792] = data_o[56];
  assign data_o[28856] = data_o[56];
  assign data_o[28920] = data_o[56];
  assign data_o[28984] = data_o[56];
  assign data_o[29048] = data_o[56];
  assign data_o[29112] = data_o[56];
  assign data_o[29176] = data_o[56];
  assign data_o[29240] = data_o[56];
  assign data_o[29304] = data_o[56];
  assign data_o[29368] = data_o[56];
  assign data_o[29432] = data_o[56];
  assign data_o[29496] = data_o[56];
  assign data_o[29560] = data_o[56];
  assign data_o[29624] = data_o[56];
  assign data_o[29688] = data_o[56];
  assign data_o[29752] = data_o[56];
  assign data_o[29816] = data_o[56];
  assign data_o[29880] = data_o[56];
  assign data_o[29944] = data_o[56];
  assign data_o[30008] = data_o[56];
  assign data_o[30072] = data_o[56];
  assign data_o[30136] = data_o[56];
  assign data_o[30200] = data_o[56];
  assign data_o[30264] = data_o[56];
  assign data_o[30328] = data_o[56];
  assign data_o[30392] = data_o[56];
  assign data_o[30456] = data_o[56];
  assign data_o[30520] = data_o[56];
  assign data_o[30584] = data_o[56];
  assign data_o[30648] = data_o[56];
  assign data_o[30712] = data_o[56];
  assign data_o[30776] = data_o[56];
  assign data_o[30840] = data_o[56];
  assign data_o[30904] = data_o[56];
  assign data_o[30968] = data_o[56];
  assign data_o[31032] = data_o[56];
  assign data_o[31096] = data_o[56];
  assign data_o[31160] = data_o[56];
  assign data_o[31224] = data_o[56];
  assign data_o[31288] = data_o[56];
  assign data_o[31352] = data_o[56];
  assign data_o[31416] = data_o[56];
  assign data_o[31480] = data_o[56];
  assign data_o[31544] = data_o[56];
  assign data_o[31608] = data_o[56];
  assign data_o[31672] = data_o[56];
  assign data_o[31736] = data_o[56];
  assign data_o[31800] = data_o[56];
  assign data_o[31864] = data_o[56];
  assign data_o[31928] = data_o[56];
  assign data_o[31992] = data_o[56];
  assign data_o[119] = data_o[55];
  assign data_o[183] = data_o[55];
  assign data_o[247] = data_o[55];
  assign data_o[311] = data_o[55];
  assign data_o[375] = data_o[55];
  assign data_o[439] = data_o[55];
  assign data_o[503] = data_o[55];
  assign data_o[567] = data_o[55];
  assign data_o[631] = data_o[55];
  assign data_o[695] = data_o[55];
  assign data_o[759] = data_o[55];
  assign data_o[823] = data_o[55];
  assign data_o[887] = data_o[55];
  assign data_o[951] = data_o[55];
  assign data_o[1015] = data_o[55];
  assign data_o[1079] = data_o[55];
  assign data_o[1143] = data_o[55];
  assign data_o[1207] = data_o[55];
  assign data_o[1271] = data_o[55];
  assign data_o[1335] = data_o[55];
  assign data_o[1399] = data_o[55];
  assign data_o[1463] = data_o[55];
  assign data_o[1527] = data_o[55];
  assign data_o[1591] = data_o[55];
  assign data_o[1655] = data_o[55];
  assign data_o[1719] = data_o[55];
  assign data_o[1783] = data_o[55];
  assign data_o[1847] = data_o[55];
  assign data_o[1911] = data_o[55];
  assign data_o[1975] = data_o[55];
  assign data_o[2039] = data_o[55];
  assign data_o[2103] = data_o[55];
  assign data_o[2167] = data_o[55];
  assign data_o[2231] = data_o[55];
  assign data_o[2295] = data_o[55];
  assign data_o[2359] = data_o[55];
  assign data_o[2423] = data_o[55];
  assign data_o[2487] = data_o[55];
  assign data_o[2551] = data_o[55];
  assign data_o[2615] = data_o[55];
  assign data_o[2679] = data_o[55];
  assign data_o[2743] = data_o[55];
  assign data_o[2807] = data_o[55];
  assign data_o[2871] = data_o[55];
  assign data_o[2935] = data_o[55];
  assign data_o[2999] = data_o[55];
  assign data_o[3063] = data_o[55];
  assign data_o[3127] = data_o[55];
  assign data_o[3191] = data_o[55];
  assign data_o[3255] = data_o[55];
  assign data_o[3319] = data_o[55];
  assign data_o[3383] = data_o[55];
  assign data_o[3447] = data_o[55];
  assign data_o[3511] = data_o[55];
  assign data_o[3575] = data_o[55];
  assign data_o[3639] = data_o[55];
  assign data_o[3703] = data_o[55];
  assign data_o[3767] = data_o[55];
  assign data_o[3831] = data_o[55];
  assign data_o[3895] = data_o[55];
  assign data_o[3959] = data_o[55];
  assign data_o[4023] = data_o[55];
  assign data_o[4087] = data_o[55];
  assign data_o[4151] = data_o[55];
  assign data_o[4215] = data_o[55];
  assign data_o[4279] = data_o[55];
  assign data_o[4343] = data_o[55];
  assign data_o[4407] = data_o[55];
  assign data_o[4471] = data_o[55];
  assign data_o[4535] = data_o[55];
  assign data_o[4599] = data_o[55];
  assign data_o[4663] = data_o[55];
  assign data_o[4727] = data_o[55];
  assign data_o[4791] = data_o[55];
  assign data_o[4855] = data_o[55];
  assign data_o[4919] = data_o[55];
  assign data_o[4983] = data_o[55];
  assign data_o[5047] = data_o[55];
  assign data_o[5111] = data_o[55];
  assign data_o[5175] = data_o[55];
  assign data_o[5239] = data_o[55];
  assign data_o[5303] = data_o[55];
  assign data_o[5367] = data_o[55];
  assign data_o[5431] = data_o[55];
  assign data_o[5495] = data_o[55];
  assign data_o[5559] = data_o[55];
  assign data_o[5623] = data_o[55];
  assign data_o[5687] = data_o[55];
  assign data_o[5751] = data_o[55];
  assign data_o[5815] = data_o[55];
  assign data_o[5879] = data_o[55];
  assign data_o[5943] = data_o[55];
  assign data_o[6007] = data_o[55];
  assign data_o[6071] = data_o[55];
  assign data_o[6135] = data_o[55];
  assign data_o[6199] = data_o[55];
  assign data_o[6263] = data_o[55];
  assign data_o[6327] = data_o[55];
  assign data_o[6391] = data_o[55];
  assign data_o[6455] = data_o[55];
  assign data_o[6519] = data_o[55];
  assign data_o[6583] = data_o[55];
  assign data_o[6647] = data_o[55];
  assign data_o[6711] = data_o[55];
  assign data_o[6775] = data_o[55];
  assign data_o[6839] = data_o[55];
  assign data_o[6903] = data_o[55];
  assign data_o[6967] = data_o[55];
  assign data_o[7031] = data_o[55];
  assign data_o[7095] = data_o[55];
  assign data_o[7159] = data_o[55];
  assign data_o[7223] = data_o[55];
  assign data_o[7287] = data_o[55];
  assign data_o[7351] = data_o[55];
  assign data_o[7415] = data_o[55];
  assign data_o[7479] = data_o[55];
  assign data_o[7543] = data_o[55];
  assign data_o[7607] = data_o[55];
  assign data_o[7671] = data_o[55];
  assign data_o[7735] = data_o[55];
  assign data_o[7799] = data_o[55];
  assign data_o[7863] = data_o[55];
  assign data_o[7927] = data_o[55];
  assign data_o[7991] = data_o[55];
  assign data_o[8055] = data_o[55];
  assign data_o[8119] = data_o[55];
  assign data_o[8183] = data_o[55];
  assign data_o[8247] = data_o[55];
  assign data_o[8311] = data_o[55];
  assign data_o[8375] = data_o[55];
  assign data_o[8439] = data_o[55];
  assign data_o[8503] = data_o[55];
  assign data_o[8567] = data_o[55];
  assign data_o[8631] = data_o[55];
  assign data_o[8695] = data_o[55];
  assign data_o[8759] = data_o[55];
  assign data_o[8823] = data_o[55];
  assign data_o[8887] = data_o[55];
  assign data_o[8951] = data_o[55];
  assign data_o[9015] = data_o[55];
  assign data_o[9079] = data_o[55];
  assign data_o[9143] = data_o[55];
  assign data_o[9207] = data_o[55];
  assign data_o[9271] = data_o[55];
  assign data_o[9335] = data_o[55];
  assign data_o[9399] = data_o[55];
  assign data_o[9463] = data_o[55];
  assign data_o[9527] = data_o[55];
  assign data_o[9591] = data_o[55];
  assign data_o[9655] = data_o[55];
  assign data_o[9719] = data_o[55];
  assign data_o[9783] = data_o[55];
  assign data_o[9847] = data_o[55];
  assign data_o[9911] = data_o[55];
  assign data_o[9975] = data_o[55];
  assign data_o[10039] = data_o[55];
  assign data_o[10103] = data_o[55];
  assign data_o[10167] = data_o[55];
  assign data_o[10231] = data_o[55];
  assign data_o[10295] = data_o[55];
  assign data_o[10359] = data_o[55];
  assign data_o[10423] = data_o[55];
  assign data_o[10487] = data_o[55];
  assign data_o[10551] = data_o[55];
  assign data_o[10615] = data_o[55];
  assign data_o[10679] = data_o[55];
  assign data_o[10743] = data_o[55];
  assign data_o[10807] = data_o[55];
  assign data_o[10871] = data_o[55];
  assign data_o[10935] = data_o[55];
  assign data_o[10999] = data_o[55];
  assign data_o[11063] = data_o[55];
  assign data_o[11127] = data_o[55];
  assign data_o[11191] = data_o[55];
  assign data_o[11255] = data_o[55];
  assign data_o[11319] = data_o[55];
  assign data_o[11383] = data_o[55];
  assign data_o[11447] = data_o[55];
  assign data_o[11511] = data_o[55];
  assign data_o[11575] = data_o[55];
  assign data_o[11639] = data_o[55];
  assign data_o[11703] = data_o[55];
  assign data_o[11767] = data_o[55];
  assign data_o[11831] = data_o[55];
  assign data_o[11895] = data_o[55];
  assign data_o[11959] = data_o[55];
  assign data_o[12023] = data_o[55];
  assign data_o[12087] = data_o[55];
  assign data_o[12151] = data_o[55];
  assign data_o[12215] = data_o[55];
  assign data_o[12279] = data_o[55];
  assign data_o[12343] = data_o[55];
  assign data_o[12407] = data_o[55];
  assign data_o[12471] = data_o[55];
  assign data_o[12535] = data_o[55];
  assign data_o[12599] = data_o[55];
  assign data_o[12663] = data_o[55];
  assign data_o[12727] = data_o[55];
  assign data_o[12791] = data_o[55];
  assign data_o[12855] = data_o[55];
  assign data_o[12919] = data_o[55];
  assign data_o[12983] = data_o[55];
  assign data_o[13047] = data_o[55];
  assign data_o[13111] = data_o[55];
  assign data_o[13175] = data_o[55];
  assign data_o[13239] = data_o[55];
  assign data_o[13303] = data_o[55];
  assign data_o[13367] = data_o[55];
  assign data_o[13431] = data_o[55];
  assign data_o[13495] = data_o[55];
  assign data_o[13559] = data_o[55];
  assign data_o[13623] = data_o[55];
  assign data_o[13687] = data_o[55];
  assign data_o[13751] = data_o[55];
  assign data_o[13815] = data_o[55];
  assign data_o[13879] = data_o[55];
  assign data_o[13943] = data_o[55];
  assign data_o[14007] = data_o[55];
  assign data_o[14071] = data_o[55];
  assign data_o[14135] = data_o[55];
  assign data_o[14199] = data_o[55];
  assign data_o[14263] = data_o[55];
  assign data_o[14327] = data_o[55];
  assign data_o[14391] = data_o[55];
  assign data_o[14455] = data_o[55];
  assign data_o[14519] = data_o[55];
  assign data_o[14583] = data_o[55];
  assign data_o[14647] = data_o[55];
  assign data_o[14711] = data_o[55];
  assign data_o[14775] = data_o[55];
  assign data_o[14839] = data_o[55];
  assign data_o[14903] = data_o[55];
  assign data_o[14967] = data_o[55];
  assign data_o[15031] = data_o[55];
  assign data_o[15095] = data_o[55];
  assign data_o[15159] = data_o[55];
  assign data_o[15223] = data_o[55];
  assign data_o[15287] = data_o[55];
  assign data_o[15351] = data_o[55];
  assign data_o[15415] = data_o[55];
  assign data_o[15479] = data_o[55];
  assign data_o[15543] = data_o[55];
  assign data_o[15607] = data_o[55];
  assign data_o[15671] = data_o[55];
  assign data_o[15735] = data_o[55];
  assign data_o[15799] = data_o[55];
  assign data_o[15863] = data_o[55];
  assign data_o[15927] = data_o[55];
  assign data_o[15991] = data_o[55];
  assign data_o[16055] = data_o[55];
  assign data_o[16119] = data_o[55];
  assign data_o[16183] = data_o[55];
  assign data_o[16247] = data_o[55];
  assign data_o[16311] = data_o[55];
  assign data_o[16375] = data_o[55];
  assign data_o[16439] = data_o[55];
  assign data_o[16503] = data_o[55];
  assign data_o[16567] = data_o[55];
  assign data_o[16631] = data_o[55];
  assign data_o[16695] = data_o[55];
  assign data_o[16759] = data_o[55];
  assign data_o[16823] = data_o[55];
  assign data_o[16887] = data_o[55];
  assign data_o[16951] = data_o[55];
  assign data_o[17015] = data_o[55];
  assign data_o[17079] = data_o[55];
  assign data_o[17143] = data_o[55];
  assign data_o[17207] = data_o[55];
  assign data_o[17271] = data_o[55];
  assign data_o[17335] = data_o[55];
  assign data_o[17399] = data_o[55];
  assign data_o[17463] = data_o[55];
  assign data_o[17527] = data_o[55];
  assign data_o[17591] = data_o[55];
  assign data_o[17655] = data_o[55];
  assign data_o[17719] = data_o[55];
  assign data_o[17783] = data_o[55];
  assign data_o[17847] = data_o[55];
  assign data_o[17911] = data_o[55];
  assign data_o[17975] = data_o[55];
  assign data_o[18039] = data_o[55];
  assign data_o[18103] = data_o[55];
  assign data_o[18167] = data_o[55];
  assign data_o[18231] = data_o[55];
  assign data_o[18295] = data_o[55];
  assign data_o[18359] = data_o[55];
  assign data_o[18423] = data_o[55];
  assign data_o[18487] = data_o[55];
  assign data_o[18551] = data_o[55];
  assign data_o[18615] = data_o[55];
  assign data_o[18679] = data_o[55];
  assign data_o[18743] = data_o[55];
  assign data_o[18807] = data_o[55];
  assign data_o[18871] = data_o[55];
  assign data_o[18935] = data_o[55];
  assign data_o[18999] = data_o[55];
  assign data_o[19063] = data_o[55];
  assign data_o[19127] = data_o[55];
  assign data_o[19191] = data_o[55];
  assign data_o[19255] = data_o[55];
  assign data_o[19319] = data_o[55];
  assign data_o[19383] = data_o[55];
  assign data_o[19447] = data_o[55];
  assign data_o[19511] = data_o[55];
  assign data_o[19575] = data_o[55];
  assign data_o[19639] = data_o[55];
  assign data_o[19703] = data_o[55];
  assign data_o[19767] = data_o[55];
  assign data_o[19831] = data_o[55];
  assign data_o[19895] = data_o[55];
  assign data_o[19959] = data_o[55];
  assign data_o[20023] = data_o[55];
  assign data_o[20087] = data_o[55];
  assign data_o[20151] = data_o[55];
  assign data_o[20215] = data_o[55];
  assign data_o[20279] = data_o[55];
  assign data_o[20343] = data_o[55];
  assign data_o[20407] = data_o[55];
  assign data_o[20471] = data_o[55];
  assign data_o[20535] = data_o[55];
  assign data_o[20599] = data_o[55];
  assign data_o[20663] = data_o[55];
  assign data_o[20727] = data_o[55];
  assign data_o[20791] = data_o[55];
  assign data_o[20855] = data_o[55];
  assign data_o[20919] = data_o[55];
  assign data_o[20983] = data_o[55];
  assign data_o[21047] = data_o[55];
  assign data_o[21111] = data_o[55];
  assign data_o[21175] = data_o[55];
  assign data_o[21239] = data_o[55];
  assign data_o[21303] = data_o[55];
  assign data_o[21367] = data_o[55];
  assign data_o[21431] = data_o[55];
  assign data_o[21495] = data_o[55];
  assign data_o[21559] = data_o[55];
  assign data_o[21623] = data_o[55];
  assign data_o[21687] = data_o[55];
  assign data_o[21751] = data_o[55];
  assign data_o[21815] = data_o[55];
  assign data_o[21879] = data_o[55];
  assign data_o[21943] = data_o[55];
  assign data_o[22007] = data_o[55];
  assign data_o[22071] = data_o[55];
  assign data_o[22135] = data_o[55];
  assign data_o[22199] = data_o[55];
  assign data_o[22263] = data_o[55];
  assign data_o[22327] = data_o[55];
  assign data_o[22391] = data_o[55];
  assign data_o[22455] = data_o[55];
  assign data_o[22519] = data_o[55];
  assign data_o[22583] = data_o[55];
  assign data_o[22647] = data_o[55];
  assign data_o[22711] = data_o[55];
  assign data_o[22775] = data_o[55];
  assign data_o[22839] = data_o[55];
  assign data_o[22903] = data_o[55];
  assign data_o[22967] = data_o[55];
  assign data_o[23031] = data_o[55];
  assign data_o[23095] = data_o[55];
  assign data_o[23159] = data_o[55];
  assign data_o[23223] = data_o[55];
  assign data_o[23287] = data_o[55];
  assign data_o[23351] = data_o[55];
  assign data_o[23415] = data_o[55];
  assign data_o[23479] = data_o[55];
  assign data_o[23543] = data_o[55];
  assign data_o[23607] = data_o[55];
  assign data_o[23671] = data_o[55];
  assign data_o[23735] = data_o[55];
  assign data_o[23799] = data_o[55];
  assign data_o[23863] = data_o[55];
  assign data_o[23927] = data_o[55];
  assign data_o[23991] = data_o[55];
  assign data_o[24055] = data_o[55];
  assign data_o[24119] = data_o[55];
  assign data_o[24183] = data_o[55];
  assign data_o[24247] = data_o[55];
  assign data_o[24311] = data_o[55];
  assign data_o[24375] = data_o[55];
  assign data_o[24439] = data_o[55];
  assign data_o[24503] = data_o[55];
  assign data_o[24567] = data_o[55];
  assign data_o[24631] = data_o[55];
  assign data_o[24695] = data_o[55];
  assign data_o[24759] = data_o[55];
  assign data_o[24823] = data_o[55];
  assign data_o[24887] = data_o[55];
  assign data_o[24951] = data_o[55];
  assign data_o[25015] = data_o[55];
  assign data_o[25079] = data_o[55];
  assign data_o[25143] = data_o[55];
  assign data_o[25207] = data_o[55];
  assign data_o[25271] = data_o[55];
  assign data_o[25335] = data_o[55];
  assign data_o[25399] = data_o[55];
  assign data_o[25463] = data_o[55];
  assign data_o[25527] = data_o[55];
  assign data_o[25591] = data_o[55];
  assign data_o[25655] = data_o[55];
  assign data_o[25719] = data_o[55];
  assign data_o[25783] = data_o[55];
  assign data_o[25847] = data_o[55];
  assign data_o[25911] = data_o[55];
  assign data_o[25975] = data_o[55];
  assign data_o[26039] = data_o[55];
  assign data_o[26103] = data_o[55];
  assign data_o[26167] = data_o[55];
  assign data_o[26231] = data_o[55];
  assign data_o[26295] = data_o[55];
  assign data_o[26359] = data_o[55];
  assign data_o[26423] = data_o[55];
  assign data_o[26487] = data_o[55];
  assign data_o[26551] = data_o[55];
  assign data_o[26615] = data_o[55];
  assign data_o[26679] = data_o[55];
  assign data_o[26743] = data_o[55];
  assign data_o[26807] = data_o[55];
  assign data_o[26871] = data_o[55];
  assign data_o[26935] = data_o[55];
  assign data_o[26999] = data_o[55];
  assign data_o[27063] = data_o[55];
  assign data_o[27127] = data_o[55];
  assign data_o[27191] = data_o[55];
  assign data_o[27255] = data_o[55];
  assign data_o[27319] = data_o[55];
  assign data_o[27383] = data_o[55];
  assign data_o[27447] = data_o[55];
  assign data_o[27511] = data_o[55];
  assign data_o[27575] = data_o[55];
  assign data_o[27639] = data_o[55];
  assign data_o[27703] = data_o[55];
  assign data_o[27767] = data_o[55];
  assign data_o[27831] = data_o[55];
  assign data_o[27895] = data_o[55];
  assign data_o[27959] = data_o[55];
  assign data_o[28023] = data_o[55];
  assign data_o[28087] = data_o[55];
  assign data_o[28151] = data_o[55];
  assign data_o[28215] = data_o[55];
  assign data_o[28279] = data_o[55];
  assign data_o[28343] = data_o[55];
  assign data_o[28407] = data_o[55];
  assign data_o[28471] = data_o[55];
  assign data_o[28535] = data_o[55];
  assign data_o[28599] = data_o[55];
  assign data_o[28663] = data_o[55];
  assign data_o[28727] = data_o[55];
  assign data_o[28791] = data_o[55];
  assign data_o[28855] = data_o[55];
  assign data_o[28919] = data_o[55];
  assign data_o[28983] = data_o[55];
  assign data_o[29047] = data_o[55];
  assign data_o[29111] = data_o[55];
  assign data_o[29175] = data_o[55];
  assign data_o[29239] = data_o[55];
  assign data_o[29303] = data_o[55];
  assign data_o[29367] = data_o[55];
  assign data_o[29431] = data_o[55];
  assign data_o[29495] = data_o[55];
  assign data_o[29559] = data_o[55];
  assign data_o[29623] = data_o[55];
  assign data_o[29687] = data_o[55];
  assign data_o[29751] = data_o[55];
  assign data_o[29815] = data_o[55];
  assign data_o[29879] = data_o[55];
  assign data_o[29943] = data_o[55];
  assign data_o[30007] = data_o[55];
  assign data_o[30071] = data_o[55];
  assign data_o[30135] = data_o[55];
  assign data_o[30199] = data_o[55];
  assign data_o[30263] = data_o[55];
  assign data_o[30327] = data_o[55];
  assign data_o[30391] = data_o[55];
  assign data_o[30455] = data_o[55];
  assign data_o[30519] = data_o[55];
  assign data_o[30583] = data_o[55];
  assign data_o[30647] = data_o[55];
  assign data_o[30711] = data_o[55];
  assign data_o[30775] = data_o[55];
  assign data_o[30839] = data_o[55];
  assign data_o[30903] = data_o[55];
  assign data_o[30967] = data_o[55];
  assign data_o[31031] = data_o[55];
  assign data_o[31095] = data_o[55];
  assign data_o[31159] = data_o[55];
  assign data_o[31223] = data_o[55];
  assign data_o[31287] = data_o[55];
  assign data_o[31351] = data_o[55];
  assign data_o[31415] = data_o[55];
  assign data_o[31479] = data_o[55];
  assign data_o[31543] = data_o[55];
  assign data_o[31607] = data_o[55];
  assign data_o[31671] = data_o[55];
  assign data_o[31735] = data_o[55];
  assign data_o[31799] = data_o[55];
  assign data_o[31863] = data_o[55];
  assign data_o[31927] = data_o[55];
  assign data_o[31991] = data_o[55];
  assign data_o[118] = data_o[54];
  assign data_o[182] = data_o[54];
  assign data_o[246] = data_o[54];
  assign data_o[310] = data_o[54];
  assign data_o[374] = data_o[54];
  assign data_o[438] = data_o[54];
  assign data_o[502] = data_o[54];
  assign data_o[566] = data_o[54];
  assign data_o[630] = data_o[54];
  assign data_o[694] = data_o[54];
  assign data_o[758] = data_o[54];
  assign data_o[822] = data_o[54];
  assign data_o[886] = data_o[54];
  assign data_o[950] = data_o[54];
  assign data_o[1014] = data_o[54];
  assign data_o[1078] = data_o[54];
  assign data_o[1142] = data_o[54];
  assign data_o[1206] = data_o[54];
  assign data_o[1270] = data_o[54];
  assign data_o[1334] = data_o[54];
  assign data_o[1398] = data_o[54];
  assign data_o[1462] = data_o[54];
  assign data_o[1526] = data_o[54];
  assign data_o[1590] = data_o[54];
  assign data_o[1654] = data_o[54];
  assign data_o[1718] = data_o[54];
  assign data_o[1782] = data_o[54];
  assign data_o[1846] = data_o[54];
  assign data_o[1910] = data_o[54];
  assign data_o[1974] = data_o[54];
  assign data_o[2038] = data_o[54];
  assign data_o[2102] = data_o[54];
  assign data_o[2166] = data_o[54];
  assign data_o[2230] = data_o[54];
  assign data_o[2294] = data_o[54];
  assign data_o[2358] = data_o[54];
  assign data_o[2422] = data_o[54];
  assign data_o[2486] = data_o[54];
  assign data_o[2550] = data_o[54];
  assign data_o[2614] = data_o[54];
  assign data_o[2678] = data_o[54];
  assign data_o[2742] = data_o[54];
  assign data_o[2806] = data_o[54];
  assign data_o[2870] = data_o[54];
  assign data_o[2934] = data_o[54];
  assign data_o[2998] = data_o[54];
  assign data_o[3062] = data_o[54];
  assign data_o[3126] = data_o[54];
  assign data_o[3190] = data_o[54];
  assign data_o[3254] = data_o[54];
  assign data_o[3318] = data_o[54];
  assign data_o[3382] = data_o[54];
  assign data_o[3446] = data_o[54];
  assign data_o[3510] = data_o[54];
  assign data_o[3574] = data_o[54];
  assign data_o[3638] = data_o[54];
  assign data_o[3702] = data_o[54];
  assign data_o[3766] = data_o[54];
  assign data_o[3830] = data_o[54];
  assign data_o[3894] = data_o[54];
  assign data_o[3958] = data_o[54];
  assign data_o[4022] = data_o[54];
  assign data_o[4086] = data_o[54];
  assign data_o[4150] = data_o[54];
  assign data_o[4214] = data_o[54];
  assign data_o[4278] = data_o[54];
  assign data_o[4342] = data_o[54];
  assign data_o[4406] = data_o[54];
  assign data_o[4470] = data_o[54];
  assign data_o[4534] = data_o[54];
  assign data_o[4598] = data_o[54];
  assign data_o[4662] = data_o[54];
  assign data_o[4726] = data_o[54];
  assign data_o[4790] = data_o[54];
  assign data_o[4854] = data_o[54];
  assign data_o[4918] = data_o[54];
  assign data_o[4982] = data_o[54];
  assign data_o[5046] = data_o[54];
  assign data_o[5110] = data_o[54];
  assign data_o[5174] = data_o[54];
  assign data_o[5238] = data_o[54];
  assign data_o[5302] = data_o[54];
  assign data_o[5366] = data_o[54];
  assign data_o[5430] = data_o[54];
  assign data_o[5494] = data_o[54];
  assign data_o[5558] = data_o[54];
  assign data_o[5622] = data_o[54];
  assign data_o[5686] = data_o[54];
  assign data_o[5750] = data_o[54];
  assign data_o[5814] = data_o[54];
  assign data_o[5878] = data_o[54];
  assign data_o[5942] = data_o[54];
  assign data_o[6006] = data_o[54];
  assign data_o[6070] = data_o[54];
  assign data_o[6134] = data_o[54];
  assign data_o[6198] = data_o[54];
  assign data_o[6262] = data_o[54];
  assign data_o[6326] = data_o[54];
  assign data_o[6390] = data_o[54];
  assign data_o[6454] = data_o[54];
  assign data_o[6518] = data_o[54];
  assign data_o[6582] = data_o[54];
  assign data_o[6646] = data_o[54];
  assign data_o[6710] = data_o[54];
  assign data_o[6774] = data_o[54];
  assign data_o[6838] = data_o[54];
  assign data_o[6902] = data_o[54];
  assign data_o[6966] = data_o[54];
  assign data_o[7030] = data_o[54];
  assign data_o[7094] = data_o[54];
  assign data_o[7158] = data_o[54];
  assign data_o[7222] = data_o[54];
  assign data_o[7286] = data_o[54];
  assign data_o[7350] = data_o[54];
  assign data_o[7414] = data_o[54];
  assign data_o[7478] = data_o[54];
  assign data_o[7542] = data_o[54];
  assign data_o[7606] = data_o[54];
  assign data_o[7670] = data_o[54];
  assign data_o[7734] = data_o[54];
  assign data_o[7798] = data_o[54];
  assign data_o[7862] = data_o[54];
  assign data_o[7926] = data_o[54];
  assign data_o[7990] = data_o[54];
  assign data_o[8054] = data_o[54];
  assign data_o[8118] = data_o[54];
  assign data_o[8182] = data_o[54];
  assign data_o[8246] = data_o[54];
  assign data_o[8310] = data_o[54];
  assign data_o[8374] = data_o[54];
  assign data_o[8438] = data_o[54];
  assign data_o[8502] = data_o[54];
  assign data_o[8566] = data_o[54];
  assign data_o[8630] = data_o[54];
  assign data_o[8694] = data_o[54];
  assign data_o[8758] = data_o[54];
  assign data_o[8822] = data_o[54];
  assign data_o[8886] = data_o[54];
  assign data_o[8950] = data_o[54];
  assign data_o[9014] = data_o[54];
  assign data_o[9078] = data_o[54];
  assign data_o[9142] = data_o[54];
  assign data_o[9206] = data_o[54];
  assign data_o[9270] = data_o[54];
  assign data_o[9334] = data_o[54];
  assign data_o[9398] = data_o[54];
  assign data_o[9462] = data_o[54];
  assign data_o[9526] = data_o[54];
  assign data_o[9590] = data_o[54];
  assign data_o[9654] = data_o[54];
  assign data_o[9718] = data_o[54];
  assign data_o[9782] = data_o[54];
  assign data_o[9846] = data_o[54];
  assign data_o[9910] = data_o[54];
  assign data_o[9974] = data_o[54];
  assign data_o[10038] = data_o[54];
  assign data_o[10102] = data_o[54];
  assign data_o[10166] = data_o[54];
  assign data_o[10230] = data_o[54];
  assign data_o[10294] = data_o[54];
  assign data_o[10358] = data_o[54];
  assign data_o[10422] = data_o[54];
  assign data_o[10486] = data_o[54];
  assign data_o[10550] = data_o[54];
  assign data_o[10614] = data_o[54];
  assign data_o[10678] = data_o[54];
  assign data_o[10742] = data_o[54];
  assign data_o[10806] = data_o[54];
  assign data_o[10870] = data_o[54];
  assign data_o[10934] = data_o[54];
  assign data_o[10998] = data_o[54];
  assign data_o[11062] = data_o[54];
  assign data_o[11126] = data_o[54];
  assign data_o[11190] = data_o[54];
  assign data_o[11254] = data_o[54];
  assign data_o[11318] = data_o[54];
  assign data_o[11382] = data_o[54];
  assign data_o[11446] = data_o[54];
  assign data_o[11510] = data_o[54];
  assign data_o[11574] = data_o[54];
  assign data_o[11638] = data_o[54];
  assign data_o[11702] = data_o[54];
  assign data_o[11766] = data_o[54];
  assign data_o[11830] = data_o[54];
  assign data_o[11894] = data_o[54];
  assign data_o[11958] = data_o[54];
  assign data_o[12022] = data_o[54];
  assign data_o[12086] = data_o[54];
  assign data_o[12150] = data_o[54];
  assign data_o[12214] = data_o[54];
  assign data_o[12278] = data_o[54];
  assign data_o[12342] = data_o[54];
  assign data_o[12406] = data_o[54];
  assign data_o[12470] = data_o[54];
  assign data_o[12534] = data_o[54];
  assign data_o[12598] = data_o[54];
  assign data_o[12662] = data_o[54];
  assign data_o[12726] = data_o[54];
  assign data_o[12790] = data_o[54];
  assign data_o[12854] = data_o[54];
  assign data_o[12918] = data_o[54];
  assign data_o[12982] = data_o[54];
  assign data_o[13046] = data_o[54];
  assign data_o[13110] = data_o[54];
  assign data_o[13174] = data_o[54];
  assign data_o[13238] = data_o[54];
  assign data_o[13302] = data_o[54];
  assign data_o[13366] = data_o[54];
  assign data_o[13430] = data_o[54];
  assign data_o[13494] = data_o[54];
  assign data_o[13558] = data_o[54];
  assign data_o[13622] = data_o[54];
  assign data_o[13686] = data_o[54];
  assign data_o[13750] = data_o[54];
  assign data_o[13814] = data_o[54];
  assign data_o[13878] = data_o[54];
  assign data_o[13942] = data_o[54];
  assign data_o[14006] = data_o[54];
  assign data_o[14070] = data_o[54];
  assign data_o[14134] = data_o[54];
  assign data_o[14198] = data_o[54];
  assign data_o[14262] = data_o[54];
  assign data_o[14326] = data_o[54];
  assign data_o[14390] = data_o[54];
  assign data_o[14454] = data_o[54];
  assign data_o[14518] = data_o[54];
  assign data_o[14582] = data_o[54];
  assign data_o[14646] = data_o[54];
  assign data_o[14710] = data_o[54];
  assign data_o[14774] = data_o[54];
  assign data_o[14838] = data_o[54];
  assign data_o[14902] = data_o[54];
  assign data_o[14966] = data_o[54];
  assign data_o[15030] = data_o[54];
  assign data_o[15094] = data_o[54];
  assign data_o[15158] = data_o[54];
  assign data_o[15222] = data_o[54];
  assign data_o[15286] = data_o[54];
  assign data_o[15350] = data_o[54];
  assign data_o[15414] = data_o[54];
  assign data_o[15478] = data_o[54];
  assign data_o[15542] = data_o[54];
  assign data_o[15606] = data_o[54];
  assign data_o[15670] = data_o[54];
  assign data_o[15734] = data_o[54];
  assign data_o[15798] = data_o[54];
  assign data_o[15862] = data_o[54];
  assign data_o[15926] = data_o[54];
  assign data_o[15990] = data_o[54];
  assign data_o[16054] = data_o[54];
  assign data_o[16118] = data_o[54];
  assign data_o[16182] = data_o[54];
  assign data_o[16246] = data_o[54];
  assign data_o[16310] = data_o[54];
  assign data_o[16374] = data_o[54];
  assign data_o[16438] = data_o[54];
  assign data_o[16502] = data_o[54];
  assign data_o[16566] = data_o[54];
  assign data_o[16630] = data_o[54];
  assign data_o[16694] = data_o[54];
  assign data_o[16758] = data_o[54];
  assign data_o[16822] = data_o[54];
  assign data_o[16886] = data_o[54];
  assign data_o[16950] = data_o[54];
  assign data_o[17014] = data_o[54];
  assign data_o[17078] = data_o[54];
  assign data_o[17142] = data_o[54];
  assign data_o[17206] = data_o[54];
  assign data_o[17270] = data_o[54];
  assign data_o[17334] = data_o[54];
  assign data_o[17398] = data_o[54];
  assign data_o[17462] = data_o[54];
  assign data_o[17526] = data_o[54];
  assign data_o[17590] = data_o[54];
  assign data_o[17654] = data_o[54];
  assign data_o[17718] = data_o[54];
  assign data_o[17782] = data_o[54];
  assign data_o[17846] = data_o[54];
  assign data_o[17910] = data_o[54];
  assign data_o[17974] = data_o[54];
  assign data_o[18038] = data_o[54];
  assign data_o[18102] = data_o[54];
  assign data_o[18166] = data_o[54];
  assign data_o[18230] = data_o[54];
  assign data_o[18294] = data_o[54];
  assign data_o[18358] = data_o[54];
  assign data_o[18422] = data_o[54];
  assign data_o[18486] = data_o[54];
  assign data_o[18550] = data_o[54];
  assign data_o[18614] = data_o[54];
  assign data_o[18678] = data_o[54];
  assign data_o[18742] = data_o[54];
  assign data_o[18806] = data_o[54];
  assign data_o[18870] = data_o[54];
  assign data_o[18934] = data_o[54];
  assign data_o[18998] = data_o[54];
  assign data_o[19062] = data_o[54];
  assign data_o[19126] = data_o[54];
  assign data_o[19190] = data_o[54];
  assign data_o[19254] = data_o[54];
  assign data_o[19318] = data_o[54];
  assign data_o[19382] = data_o[54];
  assign data_o[19446] = data_o[54];
  assign data_o[19510] = data_o[54];
  assign data_o[19574] = data_o[54];
  assign data_o[19638] = data_o[54];
  assign data_o[19702] = data_o[54];
  assign data_o[19766] = data_o[54];
  assign data_o[19830] = data_o[54];
  assign data_o[19894] = data_o[54];
  assign data_o[19958] = data_o[54];
  assign data_o[20022] = data_o[54];
  assign data_o[20086] = data_o[54];
  assign data_o[20150] = data_o[54];
  assign data_o[20214] = data_o[54];
  assign data_o[20278] = data_o[54];
  assign data_o[20342] = data_o[54];
  assign data_o[20406] = data_o[54];
  assign data_o[20470] = data_o[54];
  assign data_o[20534] = data_o[54];
  assign data_o[20598] = data_o[54];
  assign data_o[20662] = data_o[54];
  assign data_o[20726] = data_o[54];
  assign data_o[20790] = data_o[54];
  assign data_o[20854] = data_o[54];
  assign data_o[20918] = data_o[54];
  assign data_o[20982] = data_o[54];
  assign data_o[21046] = data_o[54];
  assign data_o[21110] = data_o[54];
  assign data_o[21174] = data_o[54];
  assign data_o[21238] = data_o[54];
  assign data_o[21302] = data_o[54];
  assign data_o[21366] = data_o[54];
  assign data_o[21430] = data_o[54];
  assign data_o[21494] = data_o[54];
  assign data_o[21558] = data_o[54];
  assign data_o[21622] = data_o[54];
  assign data_o[21686] = data_o[54];
  assign data_o[21750] = data_o[54];
  assign data_o[21814] = data_o[54];
  assign data_o[21878] = data_o[54];
  assign data_o[21942] = data_o[54];
  assign data_o[22006] = data_o[54];
  assign data_o[22070] = data_o[54];
  assign data_o[22134] = data_o[54];
  assign data_o[22198] = data_o[54];
  assign data_o[22262] = data_o[54];
  assign data_o[22326] = data_o[54];
  assign data_o[22390] = data_o[54];
  assign data_o[22454] = data_o[54];
  assign data_o[22518] = data_o[54];
  assign data_o[22582] = data_o[54];
  assign data_o[22646] = data_o[54];
  assign data_o[22710] = data_o[54];
  assign data_o[22774] = data_o[54];
  assign data_o[22838] = data_o[54];
  assign data_o[22902] = data_o[54];
  assign data_o[22966] = data_o[54];
  assign data_o[23030] = data_o[54];
  assign data_o[23094] = data_o[54];
  assign data_o[23158] = data_o[54];
  assign data_o[23222] = data_o[54];
  assign data_o[23286] = data_o[54];
  assign data_o[23350] = data_o[54];
  assign data_o[23414] = data_o[54];
  assign data_o[23478] = data_o[54];
  assign data_o[23542] = data_o[54];
  assign data_o[23606] = data_o[54];
  assign data_o[23670] = data_o[54];
  assign data_o[23734] = data_o[54];
  assign data_o[23798] = data_o[54];
  assign data_o[23862] = data_o[54];
  assign data_o[23926] = data_o[54];
  assign data_o[23990] = data_o[54];
  assign data_o[24054] = data_o[54];
  assign data_o[24118] = data_o[54];
  assign data_o[24182] = data_o[54];
  assign data_o[24246] = data_o[54];
  assign data_o[24310] = data_o[54];
  assign data_o[24374] = data_o[54];
  assign data_o[24438] = data_o[54];
  assign data_o[24502] = data_o[54];
  assign data_o[24566] = data_o[54];
  assign data_o[24630] = data_o[54];
  assign data_o[24694] = data_o[54];
  assign data_o[24758] = data_o[54];
  assign data_o[24822] = data_o[54];
  assign data_o[24886] = data_o[54];
  assign data_o[24950] = data_o[54];
  assign data_o[25014] = data_o[54];
  assign data_o[25078] = data_o[54];
  assign data_o[25142] = data_o[54];
  assign data_o[25206] = data_o[54];
  assign data_o[25270] = data_o[54];
  assign data_o[25334] = data_o[54];
  assign data_o[25398] = data_o[54];
  assign data_o[25462] = data_o[54];
  assign data_o[25526] = data_o[54];
  assign data_o[25590] = data_o[54];
  assign data_o[25654] = data_o[54];
  assign data_o[25718] = data_o[54];
  assign data_o[25782] = data_o[54];
  assign data_o[25846] = data_o[54];
  assign data_o[25910] = data_o[54];
  assign data_o[25974] = data_o[54];
  assign data_o[26038] = data_o[54];
  assign data_o[26102] = data_o[54];
  assign data_o[26166] = data_o[54];
  assign data_o[26230] = data_o[54];
  assign data_o[26294] = data_o[54];
  assign data_o[26358] = data_o[54];
  assign data_o[26422] = data_o[54];
  assign data_o[26486] = data_o[54];
  assign data_o[26550] = data_o[54];
  assign data_o[26614] = data_o[54];
  assign data_o[26678] = data_o[54];
  assign data_o[26742] = data_o[54];
  assign data_o[26806] = data_o[54];
  assign data_o[26870] = data_o[54];
  assign data_o[26934] = data_o[54];
  assign data_o[26998] = data_o[54];
  assign data_o[27062] = data_o[54];
  assign data_o[27126] = data_o[54];
  assign data_o[27190] = data_o[54];
  assign data_o[27254] = data_o[54];
  assign data_o[27318] = data_o[54];
  assign data_o[27382] = data_o[54];
  assign data_o[27446] = data_o[54];
  assign data_o[27510] = data_o[54];
  assign data_o[27574] = data_o[54];
  assign data_o[27638] = data_o[54];
  assign data_o[27702] = data_o[54];
  assign data_o[27766] = data_o[54];
  assign data_o[27830] = data_o[54];
  assign data_o[27894] = data_o[54];
  assign data_o[27958] = data_o[54];
  assign data_o[28022] = data_o[54];
  assign data_o[28086] = data_o[54];
  assign data_o[28150] = data_o[54];
  assign data_o[28214] = data_o[54];
  assign data_o[28278] = data_o[54];
  assign data_o[28342] = data_o[54];
  assign data_o[28406] = data_o[54];
  assign data_o[28470] = data_o[54];
  assign data_o[28534] = data_o[54];
  assign data_o[28598] = data_o[54];
  assign data_o[28662] = data_o[54];
  assign data_o[28726] = data_o[54];
  assign data_o[28790] = data_o[54];
  assign data_o[28854] = data_o[54];
  assign data_o[28918] = data_o[54];
  assign data_o[28982] = data_o[54];
  assign data_o[29046] = data_o[54];
  assign data_o[29110] = data_o[54];
  assign data_o[29174] = data_o[54];
  assign data_o[29238] = data_o[54];
  assign data_o[29302] = data_o[54];
  assign data_o[29366] = data_o[54];
  assign data_o[29430] = data_o[54];
  assign data_o[29494] = data_o[54];
  assign data_o[29558] = data_o[54];
  assign data_o[29622] = data_o[54];
  assign data_o[29686] = data_o[54];
  assign data_o[29750] = data_o[54];
  assign data_o[29814] = data_o[54];
  assign data_o[29878] = data_o[54];
  assign data_o[29942] = data_o[54];
  assign data_o[30006] = data_o[54];
  assign data_o[30070] = data_o[54];
  assign data_o[30134] = data_o[54];
  assign data_o[30198] = data_o[54];
  assign data_o[30262] = data_o[54];
  assign data_o[30326] = data_o[54];
  assign data_o[30390] = data_o[54];
  assign data_o[30454] = data_o[54];
  assign data_o[30518] = data_o[54];
  assign data_o[30582] = data_o[54];
  assign data_o[30646] = data_o[54];
  assign data_o[30710] = data_o[54];
  assign data_o[30774] = data_o[54];
  assign data_o[30838] = data_o[54];
  assign data_o[30902] = data_o[54];
  assign data_o[30966] = data_o[54];
  assign data_o[31030] = data_o[54];
  assign data_o[31094] = data_o[54];
  assign data_o[31158] = data_o[54];
  assign data_o[31222] = data_o[54];
  assign data_o[31286] = data_o[54];
  assign data_o[31350] = data_o[54];
  assign data_o[31414] = data_o[54];
  assign data_o[31478] = data_o[54];
  assign data_o[31542] = data_o[54];
  assign data_o[31606] = data_o[54];
  assign data_o[31670] = data_o[54];
  assign data_o[31734] = data_o[54];
  assign data_o[31798] = data_o[54];
  assign data_o[31862] = data_o[54];
  assign data_o[31926] = data_o[54];
  assign data_o[31990] = data_o[54];
  assign data_o[117] = data_o[53];
  assign data_o[181] = data_o[53];
  assign data_o[245] = data_o[53];
  assign data_o[309] = data_o[53];
  assign data_o[373] = data_o[53];
  assign data_o[437] = data_o[53];
  assign data_o[501] = data_o[53];
  assign data_o[565] = data_o[53];
  assign data_o[629] = data_o[53];
  assign data_o[693] = data_o[53];
  assign data_o[757] = data_o[53];
  assign data_o[821] = data_o[53];
  assign data_o[885] = data_o[53];
  assign data_o[949] = data_o[53];
  assign data_o[1013] = data_o[53];
  assign data_o[1077] = data_o[53];
  assign data_o[1141] = data_o[53];
  assign data_o[1205] = data_o[53];
  assign data_o[1269] = data_o[53];
  assign data_o[1333] = data_o[53];
  assign data_o[1397] = data_o[53];
  assign data_o[1461] = data_o[53];
  assign data_o[1525] = data_o[53];
  assign data_o[1589] = data_o[53];
  assign data_o[1653] = data_o[53];
  assign data_o[1717] = data_o[53];
  assign data_o[1781] = data_o[53];
  assign data_o[1845] = data_o[53];
  assign data_o[1909] = data_o[53];
  assign data_o[1973] = data_o[53];
  assign data_o[2037] = data_o[53];
  assign data_o[2101] = data_o[53];
  assign data_o[2165] = data_o[53];
  assign data_o[2229] = data_o[53];
  assign data_o[2293] = data_o[53];
  assign data_o[2357] = data_o[53];
  assign data_o[2421] = data_o[53];
  assign data_o[2485] = data_o[53];
  assign data_o[2549] = data_o[53];
  assign data_o[2613] = data_o[53];
  assign data_o[2677] = data_o[53];
  assign data_o[2741] = data_o[53];
  assign data_o[2805] = data_o[53];
  assign data_o[2869] = data_o[53];
  assign data_o[2933] = data_o[53];
  assign data_o[2997] = data_o[53];
  assign data_o[3061] = data_o[53];
  assign data_o[3125] = data_o[53];
  assign data_o[3189] = data_o[53];
  assign data_o[3253] = data_o[53];
  assign data_o[3317] = data_o[53];
  assign data_o[3381] = data_o[53];
  assign data_o[3445] = data_o[53];
  assign data_o[3509] = data_o[53];
  assign data_o[3573] = data_o[53];
  assign data_o[3637] = data_o[53];
  assign data_o[3701] = data_o[53];
  assign data_o[3765] = data_o[53];
  assign data_o[3829] = data_o[53];
  assign data_o[3893] = data_o[53];
  assign data_o[3957] = data_o[53];
  assign data_o[4021] = data_o[53];
  assign data_o[4085] = data_o[53];
  assign data_o[4149] = data_o[53];
  assign data_o[4213] = data_o[53];
  assign data_o[4277] = data_o[53];
  assign data_o[4341] = data_o[53];
  assign data_o[4405] = data_o[53];
  assign data_o[4469] = data_o[53];
  assign data_o[4533] = data_o[53];
  assign data_o[4597] = data_o[53];
  assign data_o[4661] = data_o[53];
  assign data_o[4725] = data_o[53];
  assign data_o[4789] = data_o[53];
  assign data_o[4853] = data_o[53];
  assign data_o[4917] = data_o[53];
  assign data_o[4981] = data_o[53];
  assign data_o[5045] = data_o[53];
  assign data_o[5109] = data_o[53];
  assign data_o[5173] = data_o[53];
  assign data_o[5237] = data_o[53];
  assign data_o[5301] = data_o[53];
  assign data_o[5365] = data_o[53];
  assign data_o[5429] = data_o[53];
  assign data_o[5493] = data_o[53];
  assign data_o[5557] = data_o[53];
  assign data_o[5621] = data_o[53];
  assign data_o[5685] = data_o[53];
  assign data_o[5749] = data_o[53];
  assign data_o[5813] = data_o[53];
  assign data_o[5877] = data_o[53];
  assign data_o[5941] = data_o[53];
  assign data_o[6005] = data_o[53];
  assign data_o[6069] = data_o[53];
  assign data_o[6133] = data_o[53];
  assign data_o[6197] = data_o[53];
  assign data_o[6261] = data_o[53];
  assign data_o[6325] = data_o[53];
  assign data_o[6389] = data_o[53];
  assign data_o[6453] = data_o[53];
  assign data_o[6517] = data_o[53];
  assign data_o[6581] = data_o[53];
  assign data_o[6645] = data_o[53];
  assign data_o[6709] = data_o[53];
  assign data_o[6773] = data_o[53];
  assign data_o[6837] = data_o[53];
  assign data_o[6901] = data_o[53];
  assign data_o[6965] = data_o[53];
  assign data_o[7029] = data_o[53];
  assign data_o[7093] = data_o[53];
  assign data_o[7157] = data_o[53];
  assign data_o[7221] = data_o[53];
  assign data_o[7285] = data_o[53];
  assign data_o[7349] = data_o[53];
  assign data_o[7413] = data_o[53];
  assign data_o[7477] = data_o[53];
  assign data_o[7541] = data_o[53];
  assign data_o[7605] = data_o[53];
  assign data_o[7669] = data_o[53];
  assign data_o[7733] = data_o[53];
  assign data_o[7797] = data_o[53];
  assign data_o[7861] = data_o[53];
  assign data_o[7925] = data_o[53];
  assign data_o[7989] = data_o[53];
  assign data_o[8053] = data_o[53];
  assign data_o[8117] = data_o[53];
  assign data_o[8181] = data_o[53];
  assign data_o[8245] = data_o[53];
  assign data_o[8309] = data_o[53];
  assign data_o[8373] = data_o[53];
  assign data_o[8437] = data_o[53];
  assign data_o[8501] = data_o[53];
  assign data_o[8565] = data_o[53];
  assign data_o[8629] = data_o[53];
  assign data_o[8693] = data_o[53];
  assign data_o[8757] = data_o[53];
  assign data_o[8821] = data_o[53];
  assign data_o[8885] = data_o[53];
  assign data_o[8949] = data_o[53];
  assign data_o[9013] = data_o[53];
  assign data_o[9077] = data_o[53];
  assign data_o[9141] = data_o[53];
  assign data_o[9205] = data_o[53];
  assign data_o[9269] = data_o[53];
  assign data_o[9333] = data_o[53];
  assign data_o[9397] = data_o[53];
  assign data_o[9461] = data_o[53];
  assign data_o[9525] = data_o[53];
  assign data_o[9589] = data_o[53];
  assign data_o[9653] = data_o[53];
  assign data_o[9717] = data_o[53];
  assign data_o[9781] = data_o[53];
  assign data_o[9845] = data_o[53];
  assign data_o[9909] = data_o[53];
  assign data_o[9973] = data_o[53];
  assign data_o[10037] = data_o[53];
  assign data_o[10101] = data_o[53];
  assign data_o[10165] = data_o[53];
  assign data_o[10229] = data_o[53];
  assign data_o[10293] = data_o[53];
  assign data_o[10357] = data_o[53];
  assign data_o[10421] = data_o[53];
  assign data_o[10485] = data_o[53];
  assign data_o[10549] = data_o[53];
  assign data_o[10613] = data_o[53];
  assign data_o[10677] = data_o[53];
  assign data_o[10741] = data_o[53];
  assign data_o[10805] = data_o[53];
  assign data_o[10869] = data_o[53];
  assign data_o[10933] = data_o[53];
  assign data_o[10997] = data_o[53];
  assign data_o[11061] = data_o[53];
  assign data_o[11125] = data_o[53];
  assign data_o[11189] = data_o[53];
  assign data_o[11253] = data_o[53];
  assign data_o[11317] = data_o[53];
  assign data_o[11381] = data_o[53];
  assign data_o[11445] = data_o[53];
  assign data_o[11509] = data_o[53];
  assign data_o[11573] = data_o[53];
  assign data_o[11637] = data_o[53];
  assign data_o[11701] = data_o[53];
  assign data_o[11765] = data_o[53];
  assign data_o[11829] = data_o[53];
  assign data_o[11893] = data_o[53];
  assign data_o[11957] = data_o[53];
  assign data_o[12021] = data_o[53];
  assign data_o[12085] = data_o[53];
  assign data_o[12149] = data_o[53];
  assign data_o[12213] = data_o[53];
  assign data_o[12277] = data_o[53];
  assign data_o[12341] = data_o[53];
  assign data_o[12405] = data_o[53];
  assign data_o[12469] = data_o[53];
  assign data_o[12533] = data_o[53];
  assign data_o[12597] = data_o[53];
  assign data_o[12661] = data_o[53];
  assign data_o[12725] = data_o[53];
  assign data_o[12789] = data_o[53];
  assign data_o[12853] = data_o[53];
  assign data_o[12917] = data_o[53];
  assign data_o[12981] = data_o[53];
  assign data_o[13045] = data_o[53];
  assign data_o[13109] = data_o[53];
  assign data_o[13173] = data_o[53];
  assign data_o[13237] = data_o[53];
  assign data_o[13301] = data_o[53];
  assign data_o[13365] = data_o[53];
  assign data_o[13429] = data_o[53];
  assign data_o[13493] = data_o[53];
  assign data_o[13557] = data_o[53];
  assign data_o[13621] = data_o[53];
  assign data_o[13685] = data_o[53];
  assign data_o[13749] = data_o[53];
  assign data_o[13813] = data_o[53];
  assign data_o[13877] = data_o[53];
  assign data_o[13941] = data_o[53];
  assign data_o[14005] = data_o[53];
  assign data_o[14069] = data_o[53];
  assign data_o[14133] = data_o[53];
  assign data_o[14197] = data_o[53];
  assign data_o[14261] = data_o[53];
  assign data_o[14325] = data_o[53];
  assign data_o[14389] = data_o[53];
  assign data_o[14453] = data_o[53];
  assign data_o[14517] = data_o[53];
  assign data_o[14581] = data_o[53];
  assign data_o[14645] = data_o[53];
  assign data_o[14709] = data_o[53];
  assign data_o[14773] = data_o[53];
  assign data_o[14837] = data_o[53];
  assign data_o[14901] = data_o[53];
  assign data_o[14965] = data_o[53];
  assign data_o[15029] = data_o[53];
  assign data_o[15093] = data_o[53];
  assign data_o[15157] = data_o[53];
  assign data_o[15221] = data_o[53];
  assign data_o[15285] = data_o[53];
  assign data_o[15349] = data_o[53];
  assign data_o[15413] = data_o[53];
  assign data_o[15477] = data_o[53];
  assign data_o[15541] = data_o[53];
  assign data_o[15605] = data_o[53];
  assign data_o[15669] = data_o[53];
  assign data_o[15733] = data_o[53];
  assign data_o[15797] = data_o[53];
  assign data_o[15861] = data_o[53];
  assign data_o[15925] = data_o[53];
  assign data_o[15989] = data_o[53];
  assign data_o[16053] = data_o[53];
  assign data_o[16117] = data_o[53];
  assign data_o[16181] = data_o[53];
  assign data_o[16245] = data_o[53];
  assign data_o[16309] = data_o[53];
  assign data_o[16373] = data_o[53];
  assign data_o[16437] = data_o[53];
  assign data_o[16501] = data_o[53];
  assign data_o[16565] = data_o[53];
  assign data_o[16629] = data_o[53];
  assign data_o[16693] = data_o[53];
  assign data_o[16757] = data_o[53];
  assign data_o[16821] = data_o[53];
  assign data_o[16885] = data_o[53];
  assign data_o[16949] = data_o[53];
  assign data_o[17013] = data_o[53];
  assign data_o[17077] = data_o[53];
  assign data_o[17141] = data_o[53];
  assign data_o[17205] = data_o[53];
  assign data_o[17269] = data_o[53];
  assign data_o[17333] = data_o[53];
  assign data_o[17397] = data_o[53];
  assign data_o[17461] = data_o[53];
  assign data_o[17525] = data_o[53];
  assign data_o[17589] = data_o[53];
  assign data_o[17653] = data_o[53];
  assign data_o[17717] = data_o[53];
  assign data_o[17781] = data_o[53];
  assign data_o[17845] = data_o[53];
  assign data_o[17909] = data_o[53];
  assign data_o[17973] = data_o[53];
  assign data_o[18037] = data_o[53];
  assign data_o[18101] = data_o[53];
  assign data_o[18165] = data_o[53];
  assign data_o[18229] = data_o[53];
  assign data_o[18293] = data_o[53];
  assign data_o[18357] = data_o[53];
  assign data_o[18421] = data_o[53];
  assign data_o[18485] = data_o[53];
  assign data_o[18549] = data_o[53];
  assign data_o[18613] = data_o[53];
  assign data_o[18677] = data_o[53];
  assign data_o[18741] = data_o[53];
  assign data_o[18805] = data_o[53];
  assign data_o[18869] = data_o[53];
  assign data_o[18933] = data_o[53];
  assign data_o[18997] = data_o[53];
  assign data_o[19061] = data_o[53];
  assign data_o[19125] = data_o[53];
  assign data_o[19189] = data_o[53];
  assign data_o[19253] = data_o[53];
  assign data_o[19317] = data_o[53];
  assign data_o[19381] = data_o[53];
  assign data_o[19445] = data_o[53];
  assign data_o[19509] = data_o[53];
  assign data_o[19573] = data_o[53];
  assign data_o[19637] = data_o[53];
  assign data_o[19701] = data_o[53];
  assign data_o[19765] = data_o[53];
  assign data_o[19829] = data_o[53];
  assign data_o[19893] = data_o[53];
  assign data_o[19957] = data_o[53];
  assign data_o[20021] = data_o[53];
  assign data_o[20085] = data_o[53];
  assign data_o[20149] = data_o[53];
  assign data_o[20213] = data_o[53];
  assign data_o[20277] = data_o[53];
  assign data_o[20341] = data_o[53];
  assign data_o[20405] = data_o[53];
  assign data_o[20469] = data_o[53];
  assign data_o[20533] = data_o[53];
  assign data_o[20597] = data_o[53];
  assign data_o[20661] = data_o[53];
  assign data_o[20725] = data_o[53];
  assign data_o[20789] = data_o[53];
  assign data_o[20853] = data_o[53];
  assign data_o[20917] = data_o[53];
  assign data_o[20981] = data_o[53];
  assign data_o[21045] = data_o[53];
  assign data_o[21109] = data_o[53];
  assign data_o[21173] = data_o[53];
  assign data_o[21237] = data_o[53];
  assign data_o[21301] = data_o[53];
  assign data_o[21365] = data_o[53];
  assign data_o[21429] = data_o[53];
  assign data_o[21493] = data_o[53];
  assign data_o[21557] = data_o[53];
  assign data_o[21621] = data_o[53];
  assign data_o[21685] = data_o[53];
  assign data_o[21749] = data_o[53];
  assign data_o[21813] = data_o[53];
  assign data_o[21877] = data_o[53];
  assign data_o[21941] = data_o[53];
  assign data_o[22005] = data_o[53];
  assign data_o[22069] = data_o[53];
  assign data_o[22133] = data_o[53];
  assign data_o[22197] = data_o[53];
  assign data_o[22261] = data_o[53];
  assign data_o[22325] = data_o[53];
  assign data_o[22389] = data_o[53];
  assign data_o[22453] = data_o[53];
  assign data_o[22517] = data_o[53];
  assign data_o[22581] = data_o[53];
  assign data_o[22645] = data_o[53];
  assign data_o[22709] = data_o[53];
  assign data_o[22773] = data_o[53];
  assign data_o[22837] = data_o[53];
  assign data_o[22901] = data_o[53];
  assign data_o[22965] = data_o[53];
  assign data_o[23029] = data_o[53];
  assign data_o[23093] = data_o[53];
  assign data_o[23157] = data_o[53];
  assign data_o[23221] = data_o[53];
  assign data_o[23285] = data_o[53];
  assign data_o[23349] = data_o[53];
  assign data_o[23413] = data_o[53];
  assign data_o[23477] = data_o[53];
  assign data_o[23541] = data_o[53];
  assign data_o[23605] = data_o[53];
  assign data_o[23669] = data_o[53];
  assign data_o[23733] = data_o[53];
  assign data_o[23797] = data_o[53];
  assign data_o[23861] = data_o[53];
  assign data_o[23925] = data_o[53];
  assign data_o[23989] = data_o[53];
  assign data_o[24053] = data_o[53];
  assign data_o[24117] = data_o[53];
  assign data_o[24181] = data_o[53];
  assign data_o[24245] = data_o[53];
  assign data_o[24309] = data_o[53];
  assign data_o[24373] = data_o[53];
  assign data_o[24437] = data_o[53];
  assign data_o[24501] = data_o[53];
  assign data_o[24565] = data_o[53];
  assign data_o[24629] = data_o[53];
  assign data_o[24693] = data_o[53];
  assign data_o[24757] = data_o[53];
  assign data_o[24821] = data_o[53];
  assign data_o[24885] = data_o[53];
  assign data_o[24949] = data_o[53];
  assign data_o[25013] = data_o[53];
  assign data_o[25077] = data_o[53];
  assign data_o[25141] = data_o[53];
  assign data_o[25205] = data_o[53];
  assign data_o[25269] = data_o[53];
  assign data_o[25333] = data_o[53];
  assign data_o[25397] = data_o[53];
  assign data_o[25461] = data_o[53];
  assign data_o[25525] = data_o[53];
  assign data_o[25589] = data_o[53];
  assign data_o[25653] = data_o[53];
  assign data_o[25717] = data_o[53];
  assign data_o[25781] = data_o[53];
  assign data_o[25845] = data_o[53];
  assign data_o[25909] = data_o[53];
  assign data_o[25973] = data_o[53];
  assign data_o[26037] = data_o[53];
  assign data_o[26101] = data_o[53];
  assign data_o[26165] = data_o[53];
  assign data_o[26229] = data_o[53];
  assign data_o[26293] = data_o[53];
  assign data_o[26357] = data_o[53];
  assign data_o[26421] = data_o[53];
  assign data_o[26485] = data_o[53];
  assign data_o[26549] = data_o[53];
  assign data_o[26613] = data_o[53];
  assign data_o[26677] = data_o[53];
  assign data_o[26741] = data_o[53];
  assign data_o[26805] = data_o[53];
  assign data_o[26869] = data_o[53];
  assign data_o[26933] = data_o[53];
  assign data_o[26997] = data_o[53];
  assign data_o[27061] = data_o[53];
  assign data_o[27125] = data_o[53];
  assign data_o[27189] = data_o[53];
  assign data_o[27253] = data_o[53];
  assign data_o[27317] = data_o[53];
  assign data_o[27381] = data_o[53];
  assign data_o[27445] = data_o[53];
  assign data_o[27509] = data_o[53];
  assign data_o[27573] = data_o[53];
  assign data_o[27637] = data_o[53];
  assign data_o[27701] = data_o[53];
  assign data_o[27765] = data_o[53];
  assign data_o[27829] = data_o[53];
  assign data_o[27893] = data_o[53];
  assign data_o[27957] = data_o[53];
  assign data_o[28021] = data_o[53];
  assign data_o[28085] = data_o[53];
  assign data_o[28149] = data_o[53];
  assign data_o[28213] = data_o[53];
  assign data_o[28277] = data_o[53];
  assign data_o[28341] = data_o[53];
  assign data_o[28405] = data_o[53];
  assign data_o[28469] = data_o[53];
  assign data_o[28533] = data_o[53];
  assign data_o[28597] = data_o[53];
  assign data_o[28661] = data_o[53];
  assign data_o[28725] = data_o[53];
  assign data_o[28789] = data_o[53];
  assign data_o[28853] = data_o[53];
  assign data_o[28917] = data_o[53];
  assign data_o[28981] = data_o[53];
  assign data_o[29045] = data_o[53];
  assign data_o[29109] = data_o[53];
  assign data_o[29173] = data_o[53];
  assign data_o[29237] = data_o[53];
  assign data_o[29301] = data_o[53];
  assign data_o[29365] = data_o[53];
  assign data_o[29429] = data_o[53];
  assign data_o[29493] = data_o[53];
  assign data_o[29557] = data_o[53];
  assign data_o[29621] = data_o[53];
  assign data_o[29685] = data_o[53];
  assign data_o[29749] = data_o[53];
  assign data_o[29813] = data_o[53];
  assign data_o[29877] = data_o[53];
  assign data_o[29941] = data_o[53];
  assign data_o[30005] = data_o[53];
  assign data_o[30069] = data_o[53];
  assign data_o[30133] = data_o[53];
  assign data_o[30197] = data_o[53];
  assign data_o[30261] = data_o[53];
  assign data_o[30325] = data_o[53];
  assign data_o[30389] = data_o[53];
  assign data_o[30453] = data_o[53];
  assign data_o[30517] = data_o[53];
  assign data_o[30581] = data_o[53];
  assign data_o[30645] = data_o[53];
  assign data_o[30709] = data_o[53];
  assign data_o[30773] = data_o[53];
  assign data_o[30837] = data_o[53];
  assign data_o[30901] = data_o[53];
  assign data_o[30965] = data_o[53];
  assign data_o[31029] = data_o[53];
  assign data_o[31093] = data_o[53];
  assign data_o[31157] = data_o[53];
  assign data_o[31221] = data_o[53];
  assign data_o[31285] = data_o[53];
  assign data_o[31349] = data_o[53];
  assign data_o[31413] = data_o[53];
  assign data_o[31477] = data_o[53];
  assign data_o[31541] = data_o[53];
  assign data_o[31605] = data_o[53];
  assign data_o[31669] = data_o[53];
  assign data_o[31733] = data_o[53];
  assign data_o[31797] = data_o[53];
  assign data_o[31861] = data_o[53];
  assign data_o[31925] = data_o[53];
  assign data_o[31989] = data_o[53];
  assign data_o[116] = data_o[52];
  assign data_o[180] = data_o[52];
  assign data_o[244] = data_o[52];
  assign data_o[308] = data_o[52];
  assign data_o[372] = data_o[52];
  assign data_o[436] = data_o[52];
  assign data_o[500] = data_o[52];
  assign data_o[564] = data_o[52];
  assign data_o[628] = data_o[52];
  assign data_o[692] = data_o[52];
  assign data_o[756] = data_o[52];
  assign data_o[820] = data_o[52];
  assign data_o[884] = data_o[52];
  assign data_o[948] = data_o[52];
  assign data_o[1012] = data_o[52];
  assign data_o[1076] = data_o[52];
  assign data_o[1140] = data_o[52];
  assign data_o[1204] = data_o[52];
  assign data_o[1268] = data_o[52];
  assign data_o[1332] = data_o[52];
  assign data_o[1396] = data_o[52];
  assign data_o[1460] = data_o[52];
  assign data_o[1524] = data_o[52];
  assign data_o[1588] = data_o[52];
  assign data_o[1652] = data_o[52];
  assign data_o[1716] = data_o[52];
  assign data_o[1780] = data_o[52];
  assign data_o[1844] = data_o[52];
  assign data_o[1908] = data_o[52];
  assign data_o[1972] = data_o[52];
  assign data_o[2036] = data_o[52];
  assign data_o[2100] = data_o[52];
  assign data_o[2164] = data_o[52];
  assign data_o[2228] = data_o[52];
  assign data_o[2292] = data_o[52];
  assign data_o[2356] = data_o[52];
  assign data_o[2420] = data_o[52];
  assign data_o[2484] = data_o[52];
  assign data_o[2548] = data_o[52];
  assign data_o[2612] = data_o[52];
  assign data_o[2676] = data_o[52];
  assign data_o[2740] = data_o[52];
  assign data_o[2804] = data_o[52];
  assign data_o[2868] = data_o[52];
  assign data_o[2932] = data_o[52];
  assign data_o[2996] = data_o[52];
  assign data_o[3060] = data_o[52];
  assign data_o[3124] = data_o[52];
  assign data_o[3188] = data_o[52];
  assign data_o[3252] = data_o[52];
  assign data_o[3316] = data_o[52];
  assign data_o[3380] = data_o[52];
  assign data_o[3444] = data_o[52];
  assign data_o[3508] = data_o[52];
  assign data_o[3572] = data_o[52];
  assign data_o[3636] = data_o[52];
  assign data_o[3700] = data_o[52];
  assign data_o[3764] = data_o[52];
  assign data_o[3828] = data_o[52];
  assign data_o[3892] = data_o[52];
  assign data_o[3956] = data_o[52];
  assign data_o[4020] = data_o[52];
  assign data_o[4084] = data_o[52];
  assign data_o[4148] = data_o[52];
  assign data_o[4212] = data_o[52];
  assign data_o[4276] = data_o[52];
  assign data_o[4340] = data_o[52];
  assign data_o[4404] = data_o[52];
  assign data_o[4468] = data_o[52];
  assign data_o[4532] = data_o[52];
  assign data_o[4596] = data_o[52];
  assign data_o[4660] = data_o[52];
  assign data_o[4724] = data_o[52];
  assign data_o[4788] = data_o[52];
  assign data_o[4852] = data_o[52];
  assign data_o[4916] = data_o[52];
  assign data_o[4980] = data_o[52];
  assign data_o[5044] = data_o[52];
  assign data_o[5108] = data_o[52];
  assign data_o[5172] = data_o[52];
  assign data_o[5236] = data_o[52];
  assign data_o[5300] = data_o[52];
  assign data_o[5364] = data_o[52];
  assign data_o[5428] = data_o[52];
  assign data_o[5492] = data_o[52];
  assign data_o[5556] = data_o[52];
  assign data_o[5620] = data_o[52];
  assign data_o[5684] = data_o[52];
  assign data_o[5748] = data_o[52];
  assign data_o[5812] = data_o[52];
  assign data_o[5876] = data_o[52];
  assign data_o[5940] = data_o[52];
  assign data_o[6004] = data_o[52];
  assign data_o[6068] = data_o[52];
  assign data_o[6132] = data_o[52];
  assign data_o[6196] = data_o[52];
  assign data_o[6260] = data_o[52];
  assign data_o[6324] = data_o[52];
  assign data_o[6388] = data_o[52];
  assign data_o[6452] = data_o[52];
  assign data_o[6516] = data_o[52];
  assign data_o[6580] = data_o[52];
  assign data_o[6644] = data_o[52];
  assign data_o[6708] = data_o[52];
  assign data_o[6772] = data_o[52];
  assign data_o[6836] = data_o[52];
  assign data_o[6900] = data_o[52];
  assign data_o[6964] = data_o[52];
  assign data_o[7028] = data_o[52];
  assign data_o[7092] = data_o[52];
  assign data_o[7156] = data_o[52];
  assign data_o[7220] = data_o[52];
  assign data_o[7284] = data_o[52];
  assign data_o[7348] = data_o[52];
  assign data_o[7412] = data_o[52];
  assign data_o[7476] = data_o[52];
  assign data_o[7540] = data_o[52];
  assign data_o[7604] = data_o[52];
  assign data_o[7668] = data_o[52];
  assign data_o[7732] = data_o[52];
  assign data_o[7796] = data_o[52];
  assign data_o[7860] = data_o[52];
  assign data_o[7924] = data_o[52];
  assign data_o[7988] = data_o[52];
  assign data_o[8052] = data_o[52];
  assign data_o[8116] = data_o[52];
  assign data_o[8180] = data_o[52];
  assign data_o[8244] = data_o[52];
  assign data_o[8308] = data_o[52];
  assign data_o[8372] = data_o[52];
  assign data_o[8436] = data_o[52];
  assign data_o[8500] = data_o[52];
  assign data_o[8564] = data_o[52];
  assign data_o[8628] = data_o[52];
  assign data_o[8692] = data_o[52];
  assign data_o[8756] = data_o[52];
  assign data_o[8820] = data_o[52];
  assign data_o[8884] = data_o[52];
  assign data_o[8948] = data_o[52];
  assign data_o[9012] = data_o[52];
  assign data_o[9076] = data_o[52];
  assign data_o[9140] = data_o[52];
  assign data_o[9204] = data_o[52];
  assign data_o[9268] = data_o[52];
  assign data_o[9332] = data_o[52];
  assign data_o[9396] = data_o[52];
  assign data_o[9460] = data_o[52];
  assign data_o[9524] = data_o[52];
  assign data_o[9588] = data_o[52];
  assign data_o[9652] = data_o[52];
  assign data_o[9716] = data_o[52];
  assign data_o[9780] = data_o[52];
  assign data_o[9844] = data_o[52];
  assign data_o[9908] = data_o[52];
  assign data_o[9972] = data_o[52];
  assign data_o[10036] = data_o[52];
  assign data_o[10100] = data_o[52];
  assign data_o[10164] = data_o[52];
  assign data_o[10228] = data_o[52];
  assign data_o[10292] = data_o[52];
  assign data_o[10356] = data_o[52];
  assign data_o[10420] = data_o[52];
  assign data_o[10484] = data_o[52];
  assign data_o[10548] = data_o[52];
  assign data_o[10612] = data_o[52];
  assign data_o[10676] = data_o[52];
  assign data_o[10740] = data_o[52];
  assign data_o[10804] = data_o[52];
  assign data_o[10868] = data_o[52];
  assign data_o[10932] = data_o[52];
  assign data_o[10996] = data_o[52];
  assign data_o[11060] = data_o[52];
  assign data_o[11124] = data_o[52];
  assign data_o[11188] = data_o[52];
  assign data_o[11252] = data_o[52];
  assign data_o[11316] = data_o[52];
  assign data_o[11380] = data_o[52];
  assign data_o[11444] = data_o[52];
  assign data_o[11508] = data_o[52];
  assign data_o[11572] = data_o[52];
  assign data_o[11636] = data_o[52];
  assign data_o[11700] = data_o[52];
  assign data_o[11764] = data_o[52];
  assign data_o[11828] = data_o[52];
  assign data_o[11892] = data_o[52];
  assign data_o[11956] = data_o[52];
  assign data_o[12020] = data_o[52];
  assign data_o[12084] = data_o[52];
  assign data_o[12148] = data_o[52];
  assign data_o[12212] = data_o[52];
  assign data_o[12276] = data_o[52];
  assign data_o[12340] = data_o[52];
  assign data_o[12404] = data_o[52];
  assign data_o[12468] = data_o[52];
  assign data_o[12532] = data_o[52];
  assign data_o[12596] = data_o[52];
  assign data_o[12660] = data_o[52];
  assign data_o[12724] = data_o[52];
  assign data_o[12788] = data_o[52];
  assign data_o[12852] = data_o[52];
  assign data_o[12916] = data_o[52];
  assign data_o[12980] = data_o[52];
  assign data_o[13044] = data_o[52];
  assign data_o[13108] = data_o[52];
  assign data_o[13172] = data_o[52];
  assign data_o[13236] = data_o[52];
  assign data_o[13300] = data_o[52];
  assign data_o[13364] = data_o[52];
  assign data_o[13428] = data_o[52];
  assign data_o[13492] = data_o[52];
  assign data_o[13556] = data_o[52];
  assign data_o[13620] = data_o[52];
  assign data_o[13684] = data_o[52];
  assign data_o[13748] = data_o[52];
  assign data_o[13812] = data_o[52];
  assign data_o[13876] = data_o[52];
  assign data_o[13940] = data_o[52];
  assign data_o[14004] = data_o[52];
  assign data_o[14068] = data_o[52];
  assign data_o[14132] = data_o[52];
  assign data_o[14196] = data_o[52];
  assign data_o[14260] = data_o[52];
  assign data_o[14324] = data_o[52];
  assign data_o[14388] = data_o[52];
  assign data_o[14452] = data_o[52];
  assign data_o[14516] = data_o[52];
  assign data_o[14580] = data_o[52];
  assign data_o[14644] = data_o[52];
  assign data_o[14708] = data_o[52];
  assign data_o[14772] = data_o[52];
  assign data_o[14836] = data_o[52];
  assign data_o[14900] = data_o[52];
  assign data_o[14964] = data_o[52];
  assign data_o[15028] = data_o[52];
  assign data_o[15092] = data_o[52];
  assign data_o[15156] = data_o[52];
  assign data_o[15220] = data_o[52];
  assign data_o[15284] = data_o[52];
  assign data_o[15348] = data_o[52];
  assign data_o[15412] = data_o[52];
  assign data_o[15476] = data_o[52];
  assign data_o[15540] = data_o[52];
  assign data_o[15604] = data_o[52];
  assign data_o[15668] = data_o[52];
  assign data_o[15732] = data_o[52];
  assign data_o[15796] = data_o[52];
  assign data_o[15860] = data_o[52];
  assign data_o[15924] = data_o[52];
  assign data_o[15988] = data_o[52];
  assign data_o[16052] = data_o[52];
  assign data_o[16116] = data_o[52];
  assign data_o[16180] = data_o[52];
  assign data_o[16244] = data_o[52];
  assign data_o[16308] = data_o[52];
  assign data_o[16372] = data_o[52];
  assign data_o[16436] = data_o[52];
  assign data_o[16500] = data_o[52];
  assign data_o[16564] = data_o[52];
  assign data_o[16628] = data_o[52];
  assign data_o[16692] = data_o[52];
  assign data_o[16756] = data_o[52];
  assign data_o[16820] = data_o[52];
  assign data_o[16884] = data_o[52];
  assign data_o[16948] = data_o[52];
  assign data_o[17012] = data_o[52];
  assign data_o[17076] = data_o[52];
  assign data_o[17140] = data_o[52];
  assign data_o[17204] = data_o[52];
  assign data_o[17268] = data_o[52];
  assign data_o[17332] = data_o[52];
  assign data_o[17396] = data_o[52];
  assign data_o[17460] = data_o[52];
  assign data_o[17524] = data_o[52];
  assign data_o[17588] = data_o[52];
  assign data_o[17652] = data_o[52];
  assign data_o[17716] = data_o[52];
  assign data_o[17780] = data_o[52];
  assign data_o[17844] = data_o[52];
  assign data_o[17908] = data_o[52];
  assign data_o[17972] = data_o[52];
  assign data_o[18036] = data_o[52];
  assign data_o[18100] = data_o[52];
  assign data_o[18164] = data_o[52];
  assign data_o[18228] = data_o[52];
  assign data_o[18292] = data_o[52];
  assign data_o[18356] = data_o[52];
  assign data_o[18420] = data_o[52];
  assign data_o[18484] = data_o[52];
  assign data_o[18548] = data_o[52];
  assign data_o[18612] = data_o[52];
  assign data_o[18676] = data_o[52];
  assign data_o[18740] = data_o[52];
  assign data_o[18804] = data_o[52];
  assign data_o[18868] = data_o[52];
  assign data_o[18932] = data_o[52];
  assign data_o[18996] = data_o[52];
  assign data_o[19060] = data_o[52];
  assign data_o[19124] = data_o[52];
  assign data_o[19188] = data_o[52];
  assign data_o[19252] = data_o[52];
  assign data_o[19316] = data_o[52];
  assign data_o[19380] = data_o[52];
  assign data_o[19444] = data_o[52];
  assign data_o[19508] = data_o[52];
  assign data_o[19572] = data_o[52];
  assign data_o[19636] = data_o[52];
  assign data_o[19700] = data_o[52];
  assign data_o[19764] = data_o[52];
  assign data_o[19828] = data_o[52];
  assign data_o[19892] = data_o[52];
  assign data_o[19956] = data_o[52];
  assign data_o[20020] = data_o[52];
  assign data_o[20084] = data_o[52];
  assign data_o[20148] = data_o[52];
  assign data_o[20212] = data_o[52];
  assign data_o[20276] = data_o[52];
  assign data_o[20340] = data_o[52];
  assign data_o[20404] = data_o[52];
  assign data_o[20468] = data_o[52];
  assign data_o[20532] = data_o[52];
  assign data_o[20596] = data_o[52];
  assign data_o[20660] = data_o[52];
  assign data_o[20724] = data_o[52];
  assign data_o[20788] = data_o[52];
  assign data_o[20852] = data_o[52];
  assign data_o[20916] = data_o[52];
  assign data_o[20980] = data_o[52];
  assign data_o[21044] = data_o[52];
  assign data_o[21108] = data_o[52];
  assign data_o[21172] = data_o[52];
  assign data_o[21236] = data_o[52];
  assign data_o[21300] = data_o[52];
  assign data_o[21364] = data_o[52];
  assign data_o[21428] = data_o[52];
  assign data_o[21492] = data_o[52];
  assign data_o[21556] = data_o[52];
  assign data_o[21620] = data_o[52];
  assign data_o[21684] = data_o[52];
  assign data_o[21748] = data_o[52];
  assign data_o[21812] = data_o[52];
  assign data_o[21876] = data_o[52];
  assign data_o[21940] = data_o[52];
  assign data_o[22004] = data_o[52];
  assign data_o[22068] = data_o[52];
  assign data_o[22132] = data_o[52];
  assign data_o[22196] = data_o[52];
  assign data_o[22260] = data_o[52];
  assign data_o[22324] = data_o[52];
  assign data_o[22388] = data_o[52];
  assign data_o[22452] = data_o[52];
  assign data_o[22516] = data_o[52];
  assign data_o[22580] = data_o[52];
  assign data_o[22644] = data_o[52];
  assign data_o[22708] = data_o[52];
  assign data_o[22772] = data_o[52];
  assign data_o[22836] = data_o[52];
  assign data_o[22900] = data_o[52];
  assign data_o[22964] = data_o[52];
  assign data_o[23028] = data_o[52];
  assign data_o[23092] = data_o[52];
  assign data_o[23156] = data_o[52];
  assign data_o[23220] = data_o[52];
  assign data_o[23284] = data_o[52];
  assign data_o[23348] = data_o[52];
  assign data_o[23412] = data_o[52];
  assign data_o[23476] = data_o[52];
  assign data_o[23540] = data_o[52];
  assign data_o[23604] = data_o[52];
  assign data_o[23668] = data_o[52];
  assign data_o[23732] = data_o[52];
  assign data_o[23796] = data_o[52];
  assign data_o[23860] = data_o[52];
  assign data_o[23924] = data_o[52];
  assign data_o[23988] = data_o[52];
  assign data_o[24052] = data_o[52];
  assign data_o[24116] = data_o[52];
  assign data_o[24180] = data_o[52];
  assign data_o[24244] = data_o[52];
  assign data_o[24308] = data_o[52];
  assign data_o[24372] = data_o[52];
  assign data_o[24436] = data_o[52];
  assign data_o[24500] = data_o[52];
  assign data_o[24564] = data_o[52];
  assign data_o[24628] = data_o[52];
  assign data_o[24692] = data_o[52];
  assign data_o[24756] = data_o[52];
  assign data_o[24820] = data_o[52];
  assign data_o[24884] = data_o[52];
  assign data_o[24948] = data_o[52];
  assign data_o[25012] = data_o[52];
  assign data_o[25076] = data_o[52];
  assign data_o[25140] = data_o[52];
  assign data_o[25204] = data_o[52];
  assign data_o[25268] = data_o[52];
  assign data_o[25332] = data_o[52];
  assign data_o[25396] = data_o[52];
  assign data_o[25460] = data_o[52];
  assign data_o[25524] = data_o[52];
  assign data_o[25588] = data_o[52];
  assign data_o[25652] = data_o[52];
  assign data_o[25716] = data_o[52];
  assign data_o[25780] = data_o[52];
  assign data_o[25844] = data_o[52];
  assign data_o[25908] = data_o[52];
  assign data_o[25972] = data_o[52];
  assign data_o[26036] = data_o[52];
  assign data_o[26100] = data_o[52];
  assign data_o[26164] = data_o[52];
  assign data_o[26228] = data_o[52];
  assign data_o[26292] = data_o[52];
  assign data_o[26356] = data_o[52];
  assign data_o[26420] = data_o[52];
  assign data_o[26484] = data_o[52];
  assign data_o[26548] = data_o[52];
  assign data_o[26612] = data_o[52];
  assign data_o[26676] = data_o[52];
  assign data_o[26740] = data_o[52];
  assign data_o[26804] = data_o[52];
  assign data_o[26868] = data_o[52];
  assign data_o[26932] = data_o[52];
  assign data_o[26996] = data_o[52];
  assign data_o[27060] = data_o[52];
  assign data_o[27124] = data_o[52];
  assign data_o[27188] = data_o[52];
  assign data_o[27252] = data_o[52];
  assign data_o[27316] = data_o[52];
  assign data_o[27380] = data_o[52];
  assign data_o[27444] = data_o[52];
  assign data_o[27508] = data_o[52];
  assign data_o[27572] = data_o[52];
  assign data_o[27636] = data_o[52];
  assign data_o[27700] = data_o[52];
  assign data_o[27764] = data_o[52];
  assign data_o[27828] = data_o[52];
  assign data_o[27892] = data_o[52];
  assign data_o[27956] = data_o[52];
  assign data_o[28020] = data_o[52];
  assign data_o[28084] = data_o[52];
  assign data_o[28148] = data_o[52];
  assign data_o[28212] = data_o[52];
  assign data_o[28276] = data_o[52];
  assign data_o[28340] = data_o[52];
  assign data_o[28404] = data_o[52];
  assign data_o[28468] = data_o[52];
  assign data_o[28532] = data_o[52];
  assign data_o[28596] = data_o[52];
  assign data_o[28660] = data_o[52];
  assign data_o[28724] = data_o[52];
  assign data_o[28788] = data_o[52];
  assign data_o[28852] = data_o[52];
  assign data_o[28916] = data_o[52];
  assign data_o[28980] = data_o[52];
  assign data_o[29044] = data_o[52];
  assign data_o[29108] = data_o[52];
  assign data_o[29172] = data_o[52];
  assign data_o[29236] = data_o[52];
  assign data_o[29300] = data_o[52];
  assign data_o[29364] = data_o[52];
  assign data_o[29428] = data_o[52];
  assign data_o[29492] = data_o[52];
  assign data_o[29556] = data_o[52];
  assign data_o[29620] = data_o[52];
  assign data_o[29684] = data_o[52];
  assign data_o[29748] = data_o[52];
  assign data_o[29812] = data_o[52];
  assign data_o[29876] = data_o[52];
  assign data_o[29940] = data_o[52];
  assign data_o[30004] = data_o[52];
  assign data_o[30068] = data_o[52];
  assign data_o[30132] = data_o[52];
  assign data_o[30196] = data_o[52];
  assign data_o[30260] = data_o[52];
  assign data_o[30324] = data_o[52];
  assign data_o[30388] = data_o[52];
  assign data_o[30452] = data_o[52];
  assign data_o[30516] = data_o[52];
  assign data_o[30580] = data_o[52];
  assign data_o[30644] = data_o[52];
  assign data_o[30708] = data_o[52];
  assign data_o[30772] = data_o[52];
  assign data_o[30836] = data_o[52];
  assign data_o[30900] = data_o[52];
  assign data_o[30964] = data_o[52];
  assign data_o[31028] = data_o[52];
  assign data_o[31092] = data_o[52];
  assign data_o[31156] = data_o[52];
  assign data_o[31220] = data_o[52];
  assign data_o[31284] = data_o[52];
  assign data_o[31348] = data_o[52];
  assign data_o[31412] = data_o[52];
  assign data_o[31476] = data_o[52];
  assign data_o[31540] = data_o[52];
  assign data_o[31604] = data_o[52];
  assign data_o[31668] = data_o[52];
  assign data_o[31732] = data_o[52];
  assign data_o[31796] = data_o[52];
  assign data_o[31860] = data_o[52];
  assign data_o[31924] = data_o[52];
  assign data_o[31988] = data_o[52];
  assign data_o[115] = data_o[51];
  assign data_o[179] = data_o[51];
  assign data_o[243] = data_o[51];
  assign data_o[307] = data_o[51];
  assign data_o[371] = data_o[51];
  assign data_o[435] = data_o[51];
  assign data_o[499] = data_o[51];
  assign data_o[563] = data_o[51];
  assign data_o[627] = data_o[51];
  assign data_o[691] = data_o[51];
  assign data_o[755] = data_o[51];
  assign data_o[819] = data_o[51];
  assign data_o[883] = data_o[51];
  assign data_o[947] = data_o[51];
  assign data_o[1011] = data_o[51];
  assign data_o[1075] = data_o[51];
  assign data_o[1139] = data_o[51];
  assign data_o[1203] = data_o[51];
  assign data_o[1267] = data_o[51];
  assign data_o[1331] = data_o[51];
  assign data_o[1395] = data_o[51];
  assign data_o[1459] = data_o[51];
  assign data_o[1523] = data_o[51];
  assign data_o[1587] = data_o[51];
  assign data_o[1651] = data_o[51];
  assign data_o[1715] = data_o[51];
  assign data_o[1779] = data_o[51];
  assign data_o[1843] = data_o[51];
  assign data_o[1907] = data_o[51];
  assign data_o[1971] = data_o[51];
  assign data_o[2035] = data_o[51];
  assign data_o[2099] = data_o[51];
  assign data_o[2163] = data_o[51];
  assign data_o[2227] = data_o[51];
  assign data_o[2291] = data_o[51];
  assign data_o[2355] = data_o[51];
  assign data_o[2419] = data_o[51];
  assign data_o[2483] = data_o[51];
  assign data_o[2547] = data_o[51];
  assign data_o[2611] = data_o[51];
  assign data_o[2675] = data_o[51];
  assign data_o[2739] = data_o[51];
  assign data_o[2803] = data_o[51];
  assign data_o[2867] = data_o[51];
  assign data_o[2931] = data_o[51];
  assign data_o[2995] = data_o[51];
  assign data_o[3059] = data_o[51];
  assign data_o[3123] = data_o[51];
  assign data_o[3187] = data_o[51];
  assign data_o[3251] = data_o[51];
  assign data_o[3315] = data_o[51];
  assign data_o[3379] = data_o[51];
  assign data_o[3443] = data_o[51];
  assign data_o[3507] = data_o[51];
  assign data_o[3571] = data_o[51];
  assign data_o[3635] = data_o[51];
  assign data_o[3699] = data_o[51];
  assign data_o[3763] = data_o[51];
  assign data_o[3827] = data_o[51];
  assign data_o[3891] = data_o[51];
  assign data_o[3955] = data_o[51];
  assign data_o[4019] = data_o[51];
  assign data_o[4083] = data_o[51];
  assign data_o[4147] = data_o[51];
  assign data_o[4211] = data_o[51];
  assign data_o[4275] = data_o[51];
  assign data_o[4339] = data_o[51];
  assign data_o[4403] = data_o[51];
  assign data_o[4467] = data_o[51];
  assign data_o[4531] = data_o[51];
  assign data_o[4595] = data_o[51];
  assign data_o[4659] = data_o[51];
  assign data_o[4723] = data_o[51];
  assign data_o[4787] = data_o[51];
  assign data_o[4851] = data_o[51];
  assign data_o[4915] = data_o[51];
  assign data_o[4979] = data_o[51];
  assign data_o[5043] = data_o[51];
  assign data_o[5107] = data_o[51];
  assign data_o[5171] = data_o[51];
  assign data_o[5235] = data_o[51];
  assign data_o[5299] = data_o[51];
  assign data_o[5363] = data_o[51];
  assign data_o[5427] = data_o[51];
  assign data_o[5491] = data_o[51];
  assign data_o[5555] = data_o[51];
  assign data_o[5619] = data_o[51];
  assign data_o[5683] = data_o[51];
  assign data_o[5747] = data_o[51];
  assign data_o[5811] = data_o[51];
  assign data_o[5875] = data_o[51];
  assign data_o[5939] = data_o[51];
  assign data_o[6003] = data_o[51];
  assign data_o[6067] = data_o[51];
  assign data_o[6131] = data_o[51];
  assign data_o[6195] = data_o[51];
  assign data_o[6259] = data_o[51];
  assign data_o[6323] = data_o[51];
  assign data_o[6387] = data_o[51];
  assign data_o[6451] = data_o[51];
  assign data_o[6515] = data_o[51];
  assign data_o[6579] = data_o[51];
  assign data_o[6643] = data_o[51];
  assign data_o[6707] = data_o[51];
  assign data_o[6771] = data_o[51];
  assign data_o[6835] = data_o[51];
  assign data_o[6899] = data_o[51];
  assign data_o[6963] = data_o[51];
  assign data_o[7027] = data_o[51];
  assign data_o[7091] = data_o[51];
  assign data_o[7155] = data_o[51];
  assign data_o[7219] = data_o[51];
  assign data_o[7283] = data_o[51];
  assign data_o[7347] = data_o[51];
  assign data_o[7411] = data_o[51];
  assign data_o[7475] = data_o[51];
  assign data_o[7539] = data_o[51];
  assign data_o[7603] = data_o[51];
  assign data_o[7667] = data_o[51];
  assign data_o[7731] = data_o[51];
  assign data_o[7795] = data_o[51];
  assign data_o[7859] = data_o[51];
  assign data_o[7923] = data_o[51];
  assign data_o[7987] = data_o[51];
  assign data_o[8051] = data_o[51];
  assign data_o[8115] = data_o[51];
  assign data_o[8179] = data_o[51];
  assign data_o[8243] = data_o[51];
  assign data_o[8307] = data_o[51];
  assign data_o[8371] = data_o[51];
  assign data_o[8435] = data_o[51];
  assign data_o[8499] = data_o[51];
  assign data_o[8563] = data_o[51];
  assign data_o[8627] = data_o[51];
  assign data_o[8691] = data_o[51];
  assign data_o[8755] = data_o[51];
  assign data_o[8819] = data_o[51];
  assign data_o[8883] = data_o[51];
  assign data_o[8947] = data_o[51];
  assign data_o[9011] = data_o[51];
  assign data_o[9075] = data_o[51];
  assign data_o[9139] = data_o[51];
  assign data_o[9203] = data_o[51];
  assign data_o[9267] = data_o[51];
  assign data_o[9331] = data_o[51];
  assign data_o[9395] = data_o[51];
  assign data_o[9459] = data_o[51];
  assign data_o[9523] = data_o[51];
  assign data_o[9587] = data_o[51];
  assign data_o[9651] = data_o[51];
  assign data_o[9715] = data_o[51];
  assign data_o[9779] = data_o[51];
  assign data_o[9843] = data_o[51];
  assign data_o[9907] = data_o[51];
  assign data_o[9971] = data_o[51];
  assign data_o[10035] = data_o[51];
  assign data_o[10099] = data_o[51];
  assign data_o[10163] = data_o[51];
  assign data_o[10227] = data_o[51];
  assign data_o[10291] = data_o[51];
  assign data_o[10355] = data_o[51];
  assign data_o[10419] = data_o[51];
  assign data_o[10483] = data_o[51];
  assign data_o[10547] = data_o[51];
  assign data_o[10611] = data_o[51];
  assign data_o[10675] = data_o[51];
  assign data_o[10739] = data_o[51];
  assign data_o[10803] = data_o[51];
  assign data_o[10867] = data_o[51];
  assign data_o[10931] = data_o[51];
  assign data_o[10995] = data_o[51];
  assign data_o[11059] = data_o[51];
  assign data_o[11123] = data_o[51];
  assign data_o[11187] = data_o[51];
  assign data_o[11251] = data_o[51];
  assign data_o[11315] = data_o[51];
  assign data_o[11379] = data_o[51];
  assign data_o[11443] = data_o[51];
  assign data_o[11507] = data_o[51];
  assign data_o[11571] = data_o[51];
  assign data_o[11635] = data_o[51];
  assign data_o[11699] = data_o[51];
  assign data_o[11763] = data_o[51];
  assign data_o[11827] = data_o[51];
  assign data_o[11891] = data_o[51];
  assign data_o[11955] = data_o[51];
  assign data_o[12019] = data_o[51];
  assign data_o[12083] = data_o[51];
  assign data_o[12147] = data_o[51];
  assign data_o[12211] = data_o[51];
  assign data_o[12275] = data_o[51];
  assign data_o[12339] = data_o[51];
  assign data_o[12403] = data_o[51];
  assign data_o[12467] = data_o[51];
  assign data_o[12531] = data_o[51];
  assign data_o[12595] = data_o[51];
  assign data_o[12659] = data_o[51];
  assign data_o[12723] = data_o[51];
  assign data_o[12787] = data_o[51];
  assign data_o[12851] = data_o[51];
  assign data_o[12915] = data_o[51];
  assign data_o[12979] = data_o[51];
  assign data_o[13043] = data_o[51];
  assign data_o[13107] = data_o[51];
  assign data_o[13171] = data_o[51];
  assign data_o[13235] = data_o[51];
  assign data_o[13299] = data_o[51];
  assign data_o[13363] = data_o[51];
  assign data_o[13427] = data_o[51];
  assign data_o[13491] = data_o[51];
  assign data_o[13555] = data_o[51];
  assign data_o[13619] = data_o[51];
  assign data_o[13683] = data_o[51];
  assign data_o[13747] = data_o[51];
  assign data_o[13811] = data_o[51];
  assign data_o[13875] = data_o[51];
  assign data_o[13939] = data_o[51];
  assign data_o[14003] = data_o[51];
  assign data_o[14067] = data_o[51];
  assign data_o[14131] = data_o[51];
  assign data_o[14195] = data_o[51];
  assign data_o[14259] = data_o[51];
  assign data_o[14323] = data_o[51];
  assign data_o[14387] = data_o[51];
  assign data_o[14451] = data_o[51];
  assign data_o[14515] = data_o[51];
  assign data_o[14579] = data_o[51];
  assign data_o[14643] = data_o[51];
  assign data_o[14707] = data_o[51];
  assign data_o[14771] = data_o[51];
  assign data_o[14835] = data_o[51];
  assign data_o[14899] = data_o[51];
  assign data_o[14963] = data_o[51];
  assign data_o[15027] = data_o[51];
  assign data_o[15091] = data_o[51];
  assign data_o[15155] = data_o[51];
  assign data_o[15219] = data_o[51];
  assign data_o[15283] = data_o[51];
  assign data_o[15347] = data_o[51];
  assign data_o[15411] = data_o[51];
  assign data_o[15475] = data_o[51];
  assign data_o[15539] = data_o[51];
  assign data_o[15603] = data_o[51];
  assign data_o[15667] = data_o[51];
  assign data_o[15731] = data_o[51];
  assign data_o[15795] = data_o[51];
  assign data_o[15859] = data_o[51];
  assign data_o[15923] = data_o[51];
  assign data_o[15987] = data_o[51];
  assign data_o[16051] = data_o[51];
  assign data_o[16115] = data_o[51];
  assign data_o[16179] = data_o[51];
  assign data_o[16243] = data_o[51];
  assign data_o[16307] = data_o[51];
  assign data_o[16371] = data_o[51];
  assign data_o[16435] = data_o[51];
  assign data_o[16499] = data_o[51];
  assign data_o[16563] = data_o[51];
  assign data_o[16627] = data_o[51];
  assign data_o[16691] = data_o[51];
  assign data_o[16755] = data_o[51];
  assign data_o[16819] = data_o[51];
  assign data_o[16883] = data_o[51];
  assign data_o[16947] = data_o[51];
  assign data_o[17011] = data_o[51];
  assign data_o[17075] = data_o[51];
  assign data_o[17139] = data_o[51];
  assign data_o[17203] = data_o[51];
  assign data_o[17267] = data_o[51];
  assign data_o[17331] = data_o[51];
  assign data_o[17395] = data_o[51];
  assign data_o[17459] = data_o[51];
  assign data_o[17523] = data_o[51];
  assign data_o[17587] = data_o[51];
  assign data_o[17651] = data_o[51];
  assign data_o[17715] = data_o[51];
  assign data_o[17779] = data_o[51];
  assign data_o[17843] = data_o[51];
  assign data_o[17907] = data_o[51];
  assign data_o[17971] = data_o[51];
  assign data_o[18035] = data_o[51];
  assign data_o[18099] = data_o[51];
  assign data_o[18163] = data_o[51];
  assign data_o[18227] = data_o[51];
  assign data_o[18291] = data_o[51];
  assign data_o[18355] = data_o[51];
  assign data_o[18419] = data_o[51];
  assign data_o[18483] = data_o[51];
  assign data_o[18547] = data_o[51];
  assign data_o[18611] = data_o[51];
  assign data_o[18675] = data_o[51];
  assign data_o[18739] = data_o[51];
  assign data_o[18803] = data_o[51];
  assign data_o[18867] = data_o[51];
  assign data_o[18931] = data_o[51];
  assign data_o[18995] = data_o[51];
  assign data_o[19059] = data_o[51];
  assign data_o[19123] = data_o[51];
  assign data_o[19187] = data_o[51];
  assign data_o[19251] = data_o[51];
  assign data_o[19315] = data_o[51];
  assign data_o[19379] = data_o[51];
  assign data_o[19443] = data_o[51];
  assign data_o[19507] = data_o[51];
  assign data_o[19571] = data_o[51];
  assign data_o[19635] = data_o[51];
  assign data_o[19699] = data_o[51];
  assign data_o[19763] = data_o[51];
  assign data_o[19827] = data_o[51];
  assign data_o[19891] = data_o[51];
  assign data_o[19955] = data_o[51];
  assign data_o[20019] = data_o[51];
  assign data_o[20083] = data_o[51];
  assign data_o[20147] = data_o[51];
  assign data_o[20211] = data_o[51];
  assign data_o[20275] = data_o[51];
  assign data_o[20339] = data_o[51];
  assign data_o[20403] = data_o[51];
  assign data_o[20467] = data_o[51];
  assign data_o[20531] = data_o[51];
  assign data_o[20595] = data_o[51];
  assign data_o[20659] = data_o[51];
  assign data_o[20723] = data_o[51];
  assign data_o[20787] = data_o[51];
  assign data_o[20851] = data_o[51];
  assign data_o[20915] = data_o[51];
  assign data_o[20979] = data_o[51];
  assign data_o[21043] = data_o[51];
  assign data_o[21107] = data_o[51];
  assign data_o[21171] = data_o[51];
  assign data_o[21235] = data_o[51];
  assign data_o[21299] = data_o[51];
  assign data_o[21363] = data_o[51];
  assign data_o[21427] = data_o[51];
  assign data_o[21491] = data_o[51];
  assign data_o[21555] = data_o[51];
  assign data_o[21619] = data_o[51];
  assign data_o[21683] = data_o[51];
  assign data_o[21747] = data_o[51];
  assign data_o[21811] = data_o[51];
  assign data_o[21875] = data_o[51];
  assign data_o[21939] = data_o[51];
  assign data_o[22003] = data_o[51];
  assign data_o[22067] = data_o[51];
  assign data_o[22131] = data_o[51];
  assign data_o[22195] = data_o[51];
  assign data_o[22259] = data_o[51];
  assign data_o[22323] = data_o[51];
  assign data_o[22387] = data_o[51];
  assign data_o[22451] = data_o[51];
  assign data_o[22515] = data_o[51];
  assign data_o[22579] = data_o[51];
  assign data_o[22643] = data_o[51];
  assign data_o[22707] = data_o[51];
  assign data_o[22771] = data_o[51];
  assign data_o[22835] = data_o[51];
  assign data_o[22899] = data_o[51];
  assign data_o[22963] = data_o[51];
  assign data_o[23027] = data_o[51];
  assign data_o[23091] = data_o[51];
  assign data_o[23155] = data_o[51];
  assign data_o[23219] = data_o[51];
  assign data_o[23283] = data_o[51];
  assign data_o[23347] = data_o[51];
  assign data_o[23411] = data_o[51];
  assign data_o[23475] = data_o[51];
  assign data_o[23539] = data_o[51];
  assign data_o[23603] = data_o[51];
  assign data_o[23667] = data_o[51];
  assign data_o[23731] = data_o[51];
  assign data_o[23795] = data_o[51];
  assign data_o[23859] = data_o[51];
  assign data_o[23923] = data_o[51];
  assign data_o[23987] = data_o[51];
  assign data_o[24051] = data_o[51];
  assign data_o[24115] = data_o[51];
  assign data_o[24179] = data_o[51];
  assign data_o[24243] = data_o[51];
  assign data_o[24307] = data_o[51];
  assign data_o[24371] = data_o[51];
  assign data_o[24435] = data_o[51];
  assign data_o[24499] = data_o[51];
  assign data_o[24563] = data_o[51];
  assign data_o[24627] = data_o[51];
  assign data_o[24691] = data_o[51];
  assign data_o[24755] = data_o[51];
  assign data_o[24819] = data_o[51];
  assign data_o[24883] = data_o[51];
  assign data_o[24947] = data_o[51];
  assign data_o[25011] = data_o[51];
  assign data_o[25075] = data_o[51];
  assign data_o[25139] = data_o[51];
  assign data_o[25203] = data_o[51];
  assign data_o[25267] = data_o[51];
  assign data_o[25331] = data_o[51];
  assign data_o[25395] = data_o[51];
  assign data_o[25459] = data_o[51];
  assign data_o[25523] = data_o[51];
  assign data_o[25587] = data_o[51];
  assign data_o[25651] = data_o[51];
  assign data_o[25715] = data_o[51];
  assign data_o[25779] = data_o[51];
  assign data_o[25843] = data_o[51];
  assign data_o[25907] = data_o[51];
  assign data_o[25971] = data_o[51];
  assign data_o[26035] = data_o[51];
  assign data_o[26099] = data_o[51];
  assign data_o[26163] = data_o[51];
  assign data_o[26227] = data_o[51];
  assign data_o[26291] = data_o[51];
  assign data_o[26355] = data_o[51];
  assign data_o[26419] = data_o[51];
  assign data_o[26483] = data_o[51];
  assign data_o[26547] = data_o[51];
  assign data_o[26611] = data_o[51];
  assign data_o[26675] = data_o[51];
  assign data_o[26739] = data_o[51];
  assign data_o[26803] = data_o[51];
  assign data_o[26867] = data_o[51];
  assign data_o[26931] = data_o[51];
  assign data_o[26995] = data_o[51];
  assign data_o[27059] = data_o[51];
  assign data_o[27123] = data_o[51];
  assign data_o[27187] = data_o[51];
  assign data_o[27251] = data_o[51];
  assign data_o[27315] = data_o[51];
  assign data_o[27379] = data_o[51];
  assign data_o[27443] = data_o[51];
  assign data_o[27507] = data_o[51];
  assign data_o[27571] = data_o[51];
  assign data_o[27635] = data_o[51];
  assign data_o[27699] = data_o[51];
  assign data_o[27763] = data_o[51];
  assign data_o[27827] = data_o[51];
  assign data_o[27891] = data_o[51];
  assign data_o[27955] = data_o[51];
  assign data_o[28019] = data_o[51];
  assign data_o[28083] = data_o[51];
  assign data_o[28147] = data_o[51];
  assign data_o[28211] = data_o[51];
  assign data_o[28275] = data_o[51];
  assign data_o[28339] = data_o[51];
  assign data_o[28403] = data_o[51];
  assign data_o[28467] = data_o[51];
  assign data_o[28531] = data_o[51];
  assign data_o[28595] = data_o[51];
  assign data_o[28659] = data_o[51];
  assign data_o[28723] = data_o[51];
  assign data_o[28787] = data_o[51];
  assign data_o[28851] = data_o[51];
  assign data_o[28915] = data_o[51];
  assign data_o[28979] = data_o[51];
  assign data_o[29043] = data_o[51];
  assign data_o[29107] = data_o[51];
  assign data_o[29171] = data_o[51];
  assign data_o[29235] = data_o[51];
  assign data_o[29299] = data_o[51];
  assign data_o[29363] = data_o[51];
  assign data_o[29427] = data_o[51];
  assign data_o[29491] = data_o[51];
  assign data_o[29555] = data_o[51];
  assign data_o[29619] = data_o[51];
  assign data_o[29683] = data_o[51];
  assign data_o[29747] = data_o[51];
  assign data_o[29811] = data_o[51];
  assign data_o[29875] = data_o[51];
  assign data_o[29939] = data_o[51];
  assign data_o[30003] = data_o[51];
  assign data_o[30067] = data_o[51];
  assign data_o[30131] = data_o[51];
  assign data_o[30195] = data_o[51];
  assign data_o[30259] = data_o[51];
  assign data_o[30323] = data_o[51];
  assign data_o[30387] = data_o[51];
  assign data_o[30451] = data_o[51];
  assign data_o[30515] = data_o[51];
  assign data_o[30579] = data_o[51];
  assign data_o[30643] = data_o[51];
  assign data_o[30707] = data_o[51];
  assign data_o[30771] = data_o[51];
  assign data_o[30835] = data_o[51];
  assign data_o[30899] = data_o[51];
  assign data_o[30963] = data_o[51];
  assign data_o[31027] = data_o[51];
  assign data_o[31091] = data_o[51];
  assign data_o[31155] = data_o[51];
  assign data_o[31219] = data_o[51];
  assign data_o[31283] = data_o[51];
  assign data_o[31347] = data_o[51];
  assign data_o[31411] = data_o[51];
  assign data_o[31475] = data_o[51];
  assign data_o[31539] = data_o[51];
  assign data_o[31603] = data_o[51];
  assign data_o[31667] = data_o[51];
  assign data_o[31731] = data_o[51];
  assign data_o[31795] = data_o[51];
  assign data_o[31859] = data_o[51];
  assign data_o[31923] = data_o[51];
  assign data_o[31987] = data_o[51];
  assign data_o[114] = data_o[50];
  assign data_o[178] = data_o[50];
  assign data_o[242] = data_o[50];
  assign data_o[306] = data_o[50];
  assign data_o[370] = data_o[50];
  assign data_o[434] = data_o[50];
  assign data_o[498] = data_o[50];
  assign data_o[562] = data_o[50];
  assign data_o[626] = data_o[50];
  assign data_o[690] = data_o[50];
  assign data_o[754] = data_o[50];
  assign data_o[818] = data_o[50];
  assign data_o[882] = data_o[50];
  assign data_o[946] = data_o[50];
  assign data_o[1010] = data_o[50];
  assign data_o[1074] = data_o[50];
  assign data_o[1138] = data_o[50];
  assign data_o[1202] = data_o[50];
  assign data_o[1266] = data_o[50];
  assign data_o[1330] = data_o[50];
  assign data_o[1394] = data_o[50];
  assign data_o[1458] = data_o[50];
  assign data_o[1522] = data_o[50];
  assign data_o[1586] = data_o[50];
  assign data_o[1650] = data_o[50];
  assign data_o[1714] = data_o[50];
  assign data_o[1778] = data_o[50];
  assign data_o[1842] = data_o[50];
  assign data_o[1906] = data_o[50];
  assign data_o[1970] = data_o[50];
  assign data_o[2034] = data_o[50];
  assign data_o[2098] = data_o[50];
  assign data_o[2162] = data_o[50];
  assign data_o[2226] = data_o[50];
  assign data_o[2290] = data_o[50];
  assign data_o[2354] = data_o[50];
  assign data_o[2418] = data_o[50];
  assign data_o[2482] = data_o[50];
  assign data_o[2546] = data_o[50];
  assign data_o[2610] = data_o[50];
  assign data_o[2674] = data_o[50];
  assign data_o[2738] = data_o[50];
  assign data_o[2802] = data_o[50];
  assign data_o[2866] = data_o[50];
  assign data_o[2930] = data_o[50];
  assign data_o[2994] = data_o[50];
  assign data_o[3058] = data_o[50];
  assign data_o[3122] = data_o[50];
  assign data_o[3186] = data_o[50];
  assign data_o[3250] = data_o[50];
  assign data_o[3314] = data_o[50];
  assign data_o[3378] = data_o[50];
  assign data_o[3442] = data_o[50];
  assign data_o[3506] = data_o[50];
  assign data_o[3570] = data_o[50];
  assign data_o[3634] = data_o[50];
  assign data_o[3698] = data_o[50];
  assign data_o[3762] = data_o[50];
  assign data_o[3826] = data_o[50];
  assign data_o[3890] = data_o[50];
  assign data_o[3954] = data_o[50];
  assign data_o[4018] = data_o[50];
  assign data_o[4082] = data_o[50];
  assign data_o[4146] = data_o[50];
  assign data_o[4210] = data_o[50];
  assign data_o[4274] = data_o[50];
  assign data_o[4338] = data_o[50];
  assign data_o[4402] = data_o[50];
  assign data_o[4466] = data_o[50];
  assign data_o[4530] = data_o[50];
  assign data_o[4594] = data_o[50];
  assign data_o[4658] = data_o[50];
  assign data_o[4722] = data_o[50];
  assign data_o[4786] = data_o[50];
  assign data_o[4850] = data_o[50];
  assign data_o[4914] = data_o[50];
  assign data_o[4978] = data_o[50];
  assign data_o[5042] = data_o[50];
  assign data_o[5106] = data_o[50];
  assign data_o[5170] = data_o[50];
  assign data_o[5234] = data_o[50];
  assign data_o[5298] = data_o[50];
  assign data_o[5362] = data_o[50];
  assign data_o[5426] = data_o[50];
  assign data_o[5490] = data_o[50];
  assign data_o[5554] = data_o[50];
  assign data_o[5618] = data_o[50];
  assign data_o[5682] = data_o[50];
  assign data_o[5746] = data_o[50];
  assign data_o[5810] = data_o[50];
  assign data_o[5874] = data_o[50];
  assign data_o[5938] = data_o[50];
  assign data_o[6002] = data_o[50];
  assign data_o[6066] = data_o[50];
  assign data_o[6130] = data_o[50];
  assign data_o[6194] = data_o[50];
  assign data_o[6258] = data_o[50];
  assign data_o[6322] = data_o[50];
  assign data_o[6386] = data_o[50];
  assign data_o[6450] = data_o[50];
  assign data_o[6514] = data_o[50];
  assign data_o[6578] = data_o[50];
  assign data_o[6642] = data_o[50];
  assign data_o[6706] = data_o[50];
  assign data_o[6770] = data_o[50];
  assign data_o[6834] = data_o[50];
  assign data_o[6898] = data_o[50];
  assign data_o[6962] = data_o[50];
  assign data_o[7026] = data_o[50];
  assign data_o[7090] = data_o[50];
  assign data_o[7154] = data_o[50];
  assign data_o[7218] = data_o[50];
  assign data_o[7282] = data_o[50];
  assign data_o[7346] = data_o[50];
  assign data_o[7410] = data_o[50];
  assign data_o[7474] = data_o[50];
  assign data_o[7538] = data_o[50];
  assign data_o[7602] = data_o[50];
  assign data_o[7666] = data_o[50];
  assign data_o[7730] = data_o[50];
  assign data_o[7794] = data_o[50];
  assign data_o[7858] = data_o[50];
  assign data_o[7922] = data_o[50];
  assign data_o[7986] = data_o[50];
  assign data_o[8050] = data_o[50];
  assign data_o[8114] = data_o[50];
  assign data_o[8178] = data_o[50];
  assign data_o[8242] = data_o[50];
  assign data_o[8306] = data_o[50];
  assign data_o[8370] = data_o[50];
  assign data_o[8434] = data_o[50];
  assign data_o[8498] = data_o[50];
  assign data_o[8562] = data_o[50];
  assign data_o[8626] = data_o[50];
  assign data_o[8690] = data_o[50];
  assign data_o[8754] = data_o[50];
  assign data_o[8818] = data_o[50];
  assign data_o[8882] = data_o[50];
  assign data_o[8946] = data_o[50];
  assign data_o[9010] = data_o[50];
  assign data_o[9074] = data_o[50];
  assign data_o[9138] = data_o[50];
  assign data_o[9202] = data_o[50];
  assign data_o[9266] = data_o[50];
  assign data_o[9330] = data_o[50];
  assign data_o[9394] = data_o[50];
  assign data_o[9458] = data_o[50];
  assign data_o[9522] = data_o[50];
  assign data_o[9586] = data_o[50];
  assign data_o[9650] = data_o[50];
  assign data_o[9714] = data_o[50];
  assign data_o[9778] = data_o[50];
  assign data_o[9842] = data_o[50];
  assign data_o[9906] = data_o[50];
  assign data_o[9970] = data_o[50];
  assign data_o[10034] = data_o[50];
  assign data_o[10098] = data_o[50];
  assign data_o[10162] = data_o[50];
  assign data_o[10226] = data_o[50];
  assign data_o[10290] = data_o[50];
  assign data_o[10354] = data_o[50];
  assign data_o[10418] = data_o[50];
  assign data_o[10482] = data_o[50];
  assign data_o[10546] = data_o[50];
  assign data_o[10610] = data_o[50];
  assign data_o[10674] = data_o[50];
  assign data_o[10738] = data_o[50];
  assign data_o[10802] = data_o[50];
  assign data_o[10866] = data_o[50];
  assign data_o[10930] = data_o[50];
  assign data_o[10994] = data_o[50];
  assign data_o[11058] = data_o[50];
  assign data_o[11122] = data_o[50];
  assign data_o[11186] = data_o[50];
  assign data_o[11250] = data_o[50];
  assign data_o[11314] = data_o[50];
  assign data_o[11378] = data_o[50];
  assign data_o[11442] = data_o[50];
  assign data_o[11506] = data_o[50];
  assign data_o[11570] = data_o[50];
  assign data_o[11634] = data_o[50];
  assign data_o[11698] = data_o[50];
  assign data_o[11762] = data_o[50];
  assign data_o[11826] = data_o[50];
  assign data_o[11890] = data_o[50];
  assign data_o[11954] = data_o[50];
  assign data_o[12018] = data_o[50];
  assign data_o[12082] = data_o[50];
  assign data_o[12146] = data_o[50];
  assign data_o[12210] = data_o[50];
  assign data_o[12274] = data_o[50];
  assign data_o[12338] = data_o[50];
  assign data_o[12402] = data_o[50];
  assign data_o[12466] = data_o[50];
  assign data_o[12530] = data_o[50];
  assign data_o[12594] = data_o[50];
  assign data_o[12658] = data_o[50];
  assign data_o[12722] = data_o[50];
  assign data_o[12786] = data_o[50];
  assign data_o[12850] = data_o[50];
  assign data_o[12914] = data_o[50];
  assign data_o[12978] = data_o[50];
  assign data_o[13042] = data_o[50];
  assign data_o[13106] = data_o[50];
  assign data_o[13170] = data_o[50];
  assign data_o[13234] = data_o[50];
  assign data_o[13298] = data_o[50];
  assign data_o[13362] = data_o[50];
  assign data_o[13426] = data_o[50];
  assign data_o[13490] = data_o[50];
  assign data_o[13554] = data_o[50];
  assign data_o[13618] = data_o[50];
  assign data_o[13682] = data_o[50];
  assign data_o[13746] = data_o[50];
  assign data_o[13810] = data_o[50];
  assign data_o[13874] = data_o[50];
  assign data_o[13938] = data_o[50];
  assign data_o[14002] = data_o[50];
  assign data_o[14066] = data_o[50];
  assign data_o[14130] = data_o[50];
  assign data_o[14194] = data_o[50];
  assign data_o[14258] = data_o[50];
  assign data_o[14322] = data_o[50];
  assign data_o[14386] = data_o[50];
  assign data_o[14450] = data_o[50];
  assign data_o[14514] = data_o[50];
  assign data_o[14578] = data_o[50];
  assign data_o[14642] = data_o[50];
  assign data_o[14706] = data_o[50];
  assign data_o[14770] = data_o[50];
  assign data_o[14834] = data_o[50];
  assign data_o[14898] = data_o[50];
  assign data_o[14962] = data_o[50];
  assign data_o[15026] = data_o[50];
  assign data_o[15090] = data_o[50];
  assign data_o[15154] = data_o[50];
  assign data_o[15218] = data_o[50];
  assign data_o[15282] = data_o[50];
  assign data_o[15346] = data_o[50];
  assign data_o[15410] = data_o[50];
  assign data_o[15474] = data_o[50];
  assign data_o[15538] = data_o[50];
  assign data_o[15602] = data_o[50];
  assign data_o[15666] = data_o[50];
  assign data_o[15730] = data_o[50];
  assign data_o[15794] = data_o[50];
  assign data_o[15858] = data_o[50];
  assign data_o[15922] = data_o[50];
  assign data_o[15986] = data_o[50];
  assign data_o[16050] = data_o[50];
  assign data_o[16114] = data_o[50];
  assign data_o[16178] = data_o[50];
  assign data_o[16242] = data_o[50];
  assign data_o[16306] = data_o[50];
  assign data_o[16370] = data_o[50];
  assign data_o[16434] = data_o[50];
  assign data_o[16498] = data_o[50];
  assign data_o[16562] = data_o[50];
  assign data_o[16626] = data_o[50];
  assign data_o[16690] = data_o[50];
  assign data_o[16754] = data_o[50];
  assign data_o[16818] = data_o[50];
  assign data_o[16882] = data_o[50];
  assign data_o[16946] = data_o[50];
  assign data_o[17010] = data_o[50];
  assign data_o[17074] = data_o[50];
  assign data_o[17138] = data_o[50];
  assign data_o[17202] = data_o[50];
  assign data_o[17266] = data_o[50];
  assign data_o[17330] = data_o[50];
  assign data_o[17394] = data_o[50];
  assign data_o[17458] = data_o[50];
  assign data_o[17522] = data_o[50];
  assign data_o[17586] = data_o[50];
  assign data_o[17650] = data_o[50];
  assign data_o[17714] = data_o[50];
  assign data_o[17778] = data_o[50];
  assign data_o[17842] = data_o[50];
  assign data_o[17906] = data_o[50];
  assign data_o[17970] = data_o[50];
  assign data_o[18034] = data_o[50];
  assign data_o[18098] = data_o[50];
  assign data_o[18162] = data_o[50];
  assign data_o[18226] = data_o[50];
  assign data_o[18290] = data_o[50];
  assign data_o[18354] = data_o[50];
  assign data_o[18418] = data_o[50];
  assign data_o[18482] = data_o[50];
  assign data_o[18546] = data_o[50];
  assign data_o[18610] = data_o[50];
  assign data_o[18674] = data_o[50];
  assign data_o[18738] = data_o[50];
  assign data_o[18802] = data_o[50];
  assign data_o[18866] = data_o[50];
  assign data_o[18930] = data_o[50];
  assign data_o[18994] = data_o[50];
  assign data_o[19058] = data_o[50];
  assign data_o[19122] = data_o[50];
  assign data_o[19186] = data_o[50];
  assign data_o[19250] = data_o[50];
  assign data_o[19314] = data_o[50];
  assign data_o[19378] = data_o[50];
  assign data_o[19442] = data_o[50];
  assign data_o[19506] = data_o[50];
  assign data_o[19570] = data_o[50];
  assign data_o[19634] = data_o[50];
  assign data_o[19698] = data_o[50];
  assign data_o[19762] = data_o[50];
  assign data_o[19826] = data_o[50];
  assign data_o[19890] = data_o[50];
  assign data_o[19954] = data_o[50];
  assign data_o[20018] = data_o[50];
  assign data_o[20082] = data_o[50];
  assign data_o[20146] = data_o[50];
  assign data_o[20210] = data_o[50];
  assign data_o[20274] = data_o[50];
  assign data_o[20338] = data_o[50];
  assign data_o[20402] = data_o[50];
  assign data_o[20466] = data_o[50];
  assign data_o[20530] = data_o[50];
  assign data_o[20594] = data_o[50];
  assign data_o[20658] = data_o[50];
  assign data_o[20722] = data_o[50];
  assign data_o[20786] = data_o[50];
  assign data_o[20850] = data_o[50];
  assign data_o[20914] = data_o[50];
  assign data_o[20978] = data_o[50];
  assign data_o[21042] = data_o[50];
  assign data_o[21106] = data_o[50];
  assign data_o[21170] = data_o[50];
  assign data_o[21234] = data_o[50];
  assign data_o[21298] = data_o[50];
  assign data_o[21362] = data_o[50];
  assign data_o[21426] = data_o[50];
  assign data_o[21490] = data_o[50];
  assign data_o[21554] = data_o[50];
  assign data_o[21618] = data_o[50];
  assign data_o[21682] = data_o[50];
  assign data_o[21746] = data_o[50];
  assign data_o[21810] = data_o[50];
  assign data_o[21874] = data_o[50];
  assign data_o[21938] = data_o[50];
  assign data_o[22002] = data_o[50];
  assign data_o[22066] = data_o[50];
  assign data_o[22130] = data_o[50];
  assign data_o[22194] = data_o[50];
  assign data_o[22258] = data_o[50];
  assign data_o[22322] = data_o[50];
  assign data_o[22386] = data_o[50];
  assign data_o[22450] = data_o[50];
  assign data_o[22514] = data_o[50];
  assign data_o[22578] = data_o[50];
  assign data_o[22642] = data_o[50];
  assign data_o[22706] = data_o[50];
  assign data_o[22770] = data_o[50];
  assign data_o[22834] = data_o[50];
  assign data_o[22898] = data_o[50];
  assign data_o[22962] = data_o[50];
  assign data_o[23026] = data_o[50];
  assign data_o[23090] = data_o[50];
  assign data_o[23154] = data_o[50];
  assign data_o[23218] = data_o[50];
  assign data_o[23282] = data_o[50];
  assign data_o[23346] = data_o[50];
  assign data_o[23410] = data_o[50];
  assign data_o[23474] = data_o[50];
  assign data_o[23538] = data_o[50];
  assign data_o[23602] = data_o[50];
  assign data_o[23666] = data_o[50];
  assign data_o[23730] = data_o[50];
  assign data_o[23794] = data_o[50];
  assign data_o[23858] = data_o[50];
  assign data_o[23922] = data_o[50];
  assign data_o[23986] = data_o[50];
  assign data_o[24050] = data_o[50];
  assign data_o[24114] = data_o[50];
  assign data_o[24178] = data_o[50];
  assign data_o[24242] = data_o[50];
  assign data_o[24306] = data_o[50];
  assign data_o[24370] = data_o[50];
  assign data_o[24434] = data_o[50];
  assign data_o[24498] = data_o[50];
  assign data_o[24562] = data_o[50];
  assign data_o[24626] = data_o[50];
  assign data_o[24690] = data_o[50];
  assign data_o[24754] = data_o[50];
  assign data_o[24818] = data_o[50];
  assign data_o[24882] = data_o[50];
  assign data_o[24946] = data_o[50];
  assign data_o[25010] = data_o[50];
  assign data_o[25074] = data_o[50];
  assign data_o[25138] = data_o[50];
  assign data_o[25202] = data_o[50];
  assign data_o[25266] = data_o[50];
  assign data_o[25330] = data_o[50];
  assign data_o[25394] = data_o[50];
  assign data_o[25458] = data_o[50];
  assign data_o[25522] = data_o[50];
  assign data_o[25586] = data_o[50];
  assign data_o[25650] = data_o[50];
  assign data_o[25714] = data_o[50];
  assign data_o[25778] = data_o[50];
  assign data_o[25842] = data_o[50];
  assign data_o[25906] = data_o[50];
  assign data_o[25970] = data_o[50];
  assign data_o[26034] = data_o[50];
  assign data_o[26098] = data_o[50];
  assign data_o[26162] = data_o[50];
  assign data_o[26226] = data_o[50];
  assign data_o[26290] = data_o[50];
  assign data_o[26354] = data_o[50];
  assign data_o[26418] = data_o[50];
  assign data_o[26482] = data_o[50];
  assign data_o[26546] = data_o[50];
  assign data_o[26610] = data_o[50];
  assign data_o[26674] = data_o[50];
  assign data_o[26738] = data_o[50];
  assign data_o[26802] = data_o[50];
  assign data_o[26866] = data_o[50];
  assign data_o[26930] = data_o[50];
  assign data_o[26994] = data_o[50];
  assign data_o[27058] = data_o[50];
  assign data_o[27122] = data_o[50];
  assign data_o[27186] = data_o[50];
  assign data_o[27250] = data_o[50];
  assign data_o[27314] = data_o[50];
  assign data_o[27378] = data_o[50];
  assign data_o[27442] = data_o[50];
  assign data_o[27506] = data_o[50];
  assign data_o[27570] = data_o[50];
  assign data_o[27634] = data_o[50];
  assign data_o[27698] = data_o[50];
  assign data_o[27762] = data_o[50];
  assign data_o[27826] = data_o[50];
  assign data_o[27890] = data_o[50];
  assign data_o[27954] = data_o[50];
  assign data_o[28018] = data_o[50];
  assign data_o[28082] = data_o[50];
  assign data_o[28146] = data_o[50];
  assign data_o[28210] = data_o[50];
  assign data_o[28274] = data_o[50];
  assign data_o[28338] = data_o[50];
  assign data_o[28402] = data_o[50];
  assign data_o[28466] = data_o[50];
  assign data_o[28530] = data_o[50];
  assign data_o[28594] = data_o[50];
  assign data_o[28658] = data_o[50];
  assign data_o[28722] = data_o[50];
  assign data_o[28786] = data_o[50];
  assign data_o[28850] = data_o[50];
  assign data_o[28914] = data_o[50];
  assign data_o[28978] = data_o[50];
  assign data_o[29042] = data_o[50];
  assign data_o[29106] = data_o[50];
  assign data_o[29170] = data_o[50];
  assign data_o[29234] = data_o[50];
  assign data_o[29298] = data_o[50];
  assign data_o[29362] = data_o[50];
  assign data_o[29426] = data_o[50];
  assign data_o[29490] = data_o[50];
  assign data_o[29554] = data_o[50];
  assign data_o[29618] = data_o[50];
  assign data_o[29682] = data_o[50];
  assign data_o[29746] = data_o[50];
  assign data_o[29810] = data_o[50];
  assign data_o[29874] = data_o[50];
  assign data_o[29938] = data_o[50];
  assign data_o[30002] = data_o[50];
  assign data_o[30066] = data_o[50];
  assign data_o[30130] = data_o[50];
  assign data_o[30194] = data_o[50];
  assign data_o[30258] = data_o[50];
  assign data_o[30322] = data_o[50];
  assign data_o[30386] = data_o[50];
  assign data_o[30450] = data_o[50];
  assign data_o[30514] = data_o[50];
  assign data_o[30578] = data_o[50];
  assign data_o[30642] = data_o[50];
  assign data_o[30706] = data_o[50];
  assign data_o[30770] = data_o[50];
  assign data_o[30834] = data_o[50];
  assign data_o[30898] = data_o[50];
  assign data_o[30962] = data_o[50];
  assign data_o[31026] = data_o[50];
  assign data_o[31090] = data_o[50];
  assign data_o[31154] = data_o[50];
  assign data_o[31218] = data_o[50];
  assign data_o[31282] = data_o[50];
  assign data_o[31346] = data_o[50];
  assign data_o[31410] = data_o[50];
  assign data_o[31474] = data_o[50];
  assign data_o[31538] = data_o[50];
  assign data_o[31602] = data_o[50];
  assign data_o[31666] = data_o[50];
  assign data_o[31730] = data_o[50];
  assign data_o[31794] = data_o[50];
  assign data_o[31858] = data_o[50];
  assign data_o[31922] = data_o[50];
  assign data_o[31986] = data_o[50];
  assign data_o[113] = data_o[49];
  assign data_o[177] = data_o[49];
  assign data_o[241] = data_o[49];
  assign data_o[305] = data_o[49];
  assign data_o[369] = data_o[49];
  assign data_o[433] = data_o[49];
  assign data_o[497] = data_o[49];
  assign data_o[561] = data_o[49];
  assign data_o[625] = data_o[49];
  assign data_o[689] = data_o[49];
  assign data_o[753] = data_o[49];
  assign data_o[817] = data_o[49];
  assign data_o[881] = data_o[49];
  assign data_o[945] = data_o[49];
  assign data_o[1009] = data_o[49];
  assign data_o[1073] = data_o[49];
  assign data_o[1137] = data_o[49];
  assign data_o[1201] = data_o[49];
  assign data_o[1265] = data_o[49];
  assign data_o[1329] = data_o[49];
  assign data_o[1393] = data_o[49];
  assign data_o[1457] = data_o[49];
  assign data_o[1521] = data_o[49];
  assign data_o[1585] = data_o[49];
  assign data_o[1649] = data_o[49];
  assign data_o[1713] = data_o[49];
  assign data_o[1777] = data_o[49];
  assign data_o[1841] = data_o[49];
  assign data_o[1905] = data_o[49];
  assign data_o[1969] = data_o[49];
  assign data_o[2033] = data_o[49];
  assign data_o[2097] = data_o[49];
  assign data_o[2161] = data_o[49];
  assign data_o[2225] = data_o[49];
  assign data_o[2289] = data_o[49];
  assign data_o[2353] = data_o[49];
  assign data_o[2417] = data_o[49];
  assign data_o[2481] = data_o[49];
  assign data_o[2545] = data_o[49];
  assign data_o[2609] = data_o[49];
  assign data_o[2673] = data_o[49];
  assign data_o[2737] = data_o[49];
  assign data_o[2801] = data_o[49];
  assign data_o[2865] = data_o[49];
  assign data_o[2929] = data_o[49];
  assign data_o[2993] = data_o[49];
  assign data_o[3057] = data_o[49];
  assign data_o[3121] = data_o[49];
  assign data_o[3185] = data_o[49];
  assign data_o[3249] = data_o[49];
  assign data_o[3313] = data_o[49];
  assign data_o[3377] = data_o[49];
  assign data_o[3441] = data_o[49];
  assign data_o[3505] = data_o[49];
  assign data_o[3569] = data_o[49];
  assign data_o[3633] = data_o[49];
  assign data_o[3697] = data_o[49];
  assign data_o[3761] = data_o[49];
  assign data_o[3825] = data_o[49];
  assign data_o[3889] = data_o[49];
  assign data_o[3953] = data_o[49];
  assign data_o[4017] = data_o[49];
  assign data_o[4081] = data_o[49];
  assign data_o[4145] = data_o[49];
  assign data_o[4209] = data_o[49];
  assign data_o[4273] = data_o[49];
  assign data_o[4337] = data_o[49];
  assign data_o[4401] = data_o[49];
  assign data_o[4465] = data_o[49];
  assign data_o[4529] = data_o[49];
  assign data_o[4593] = data_o[49];
  assign data_o[4657] = data_o[49];
  assign data_o[4721] = data_o[49];
  assign data_o[4785] = data_o[49];
  assign data_o[4849] = data_o[49];
  assign data_o[4913] = data_o[49];
  assign data_o[4977] = data_o[49];
  assign data_o[5041] = data_o[49];
  assign data_o[5105] = data_o[49];
  assign data_o[5169] = data_o[49];
  assign data_o[5233] = data_o[49];
  assign data_o[5297] = data_o[49];
  assign data_o[5361] = data_o[49];
  assign data_o[5425] = data_o[49];
  assign data_o[5489] = data_o[49];
  assign data_o[5553] = data_o[49];
  assign data_o[5617] = data_o[49];
  assign data_o[5681] = data_o[49];
  assign data_o[5745] = data_o[49];
  assign data_o[5809] = data_o[49];
  assign data_o[5873] = data_o[49];
  assign data_o[5937] = data_o[49];
  assign data_o[6001] = data_o[49];
  assign data_o[6065] = data_o[49];
  assign data_o[6129] = data_o[49];
  assign data_o[6193] = data_o[49];
  assign data_o[6257] = data_o[49];
  assign data_o[6321] = data_o[49];
  assign data_o[6385] = data_o[49];
  assign data_o[6449] = data_o[49];
  assign data_o[6513] = data_o[49];
  assign data_o[6577] = data_o[49];
  assign data_o[6641] = data_o[49];
  assign data_o[6705] = data_o[49];
  assign data_o[6769] = data_o[49];
  assign data_o[6833] = data_o[49];
  assign data_o[6897] = data_o[49];
  assign data_o[6961] = data_o[49];
  assign data_o[7025] = data_o[49];
  assign data_o[7089] = data_o[49];
  assign data_o[7153] = data_o[49];
  assign data_o[7217] = data_o[49];
  assign data_o[7281] = data_o[49];
  assign data_o[7345] = data_o[49];
  assign data_o[7409] = data_o[49];
  assign data_o[7473] = data_o[49];
  assign data_o[7537] = data_o[49];
  assign data_o[7601] = data_o[49];
  assign data_o[7665] = data_o[49];
  assign data_o[7729] = data_o[49];
  assign data_o[7793] = data_o[49];
  assign data_o[7857] = data_o[49];
  assign data_o[7921] = data_o[49];
  assign data_o[7985] = data_o[49];
  assign data_o[8049] = data_o[49];
  assign data_o[8113] = data_o[49];
  assign data_o[8177] = data_o[49];
  assign data_o[8241] = data_o[49];
  assign data_o[8305] = data_o[49];
  assign data_o[8369] = data_o[49];
  assign data_o[8433] = data_o[49];
  assign data_o[8497] = data_o[49];
  assign data_o[8561] = data_o[49];
  assign data_o[8625] = data_o[49];
  assign data_o[8689] = data_o[49];
  assign data_o[8753] = data_o[49];
  assign data_o[8817] = data_o[49];
  assign data_o[8881] = data_o[49];
  assign data_o[8945] = data_o[49];
  assign data_o[9009] = data_o[49];
  assign data_o[9073] = data_o[49];
  assign data_o[9137] = data_o[49];
  assign data_o[9201] = data_o[49];
  assign data_o[9265] = data_o[49];
  assign data_o[9329] = data_o[49];
  assign data_o[9393] = data_o[49];
  assign data_o[9457] = data_o[49];
  assign data_o[9521] = data_o[49];
  assign data_o[9585] = data_o[49];
  assign data_o[9649] = data_o[49];
  assign data_o[9713] = data_o[49];
  assign data_o[9777] = data_o[49];
  assign data_o[9841] = data_o[49];
  assign data_o[9905] = data_o[49];
  assign data_o[9969] = data_o[49];
  assign data_o[10033] = data_o[49];
  assign data_o[10097] = data_o[49];
  assign data_o[10161] = data_o[49];
  assign data_o[10225] = data_o[49];
  assign data_o[10289] = data_o[49];
  assign data_o[10353] = data_o[49];
  assign data_o[10417] = data_o[49];
  assign data_o[10481] = data_o[49];
  assign data_o[10545] = data_o[49];
  assign data_o[10609] = data_o[49];
  assign data_o[10673] = data_o[49];
  assign data_o[10737] = data_o[49];
  assign data_o[10801] = data_o[49];
  assign data_o[10865] = data_o[49];
  assign data_o[10929] = data_o[49];
  assign data_o[10993] = data_o[49];
  assign data_o[11057] = data_o[49];
  assign data_o[11121] = data_o[49];
  assign data_o[11185] = data_o[49];
  assign data_o[11249] = data_o[49];
  assign data_o[11313] = data_o[49];
  assign data_o[11377] = data_o[49];
  assign data_o[11441] = data_o[49];
  assign data_o[11505] = data_o[49];
  assign data_o[11569] = data_o[49];
  assign data_o[11633] = data_o[49];
  assign data_o[11697] = data_o[49];
  assign data_o[11761] = data_o[49];
  assign data_o[11825] = data_o[49];
  assign data_o[11889] = data_o[49];
  assign data_o[11953] = data_o[49];
  assign data_o[12017] = data_o[49];
  assign data_o[12081] = data_o[49];
  assign data_o[12145] = data_o[49];
  assign data_o[12209] = data_o[49];
  assign data_o[12273] = data_o[49];
  assign data_o[12337] = data_o[49];
  assign data_o[12401] = data_o[49];
  assign data_o[12465] = data_o[49];
  assign data_o[12529] = data_o[49];
  assign data_o[12593] = data_o[49];
  assign data_o[12657] = data_o[49];
  assign data_o[12721] = data_o[49];
  assign data_o[12785] = data_o[49];
  assign data_o[12849] = data_o[49];
  assign data_o[12913] = data_o[49];
  assign data_o[12977] = data_o[49];
  assign data_o[13041] = data_o[49];
  assign data_o[13105] = data_o[49];
  assign data_o[13169] = data_o[49];
  assign data_o[13233] = data_o[49];
  assign data_o[13297] = data_o[49];
  assign data_o[13361] = data_o[49];
  assign data_o[13425] = data_o[49];
  assign data_o[13489] = data_o[49];
  assign data_o[13553] = data_o[49];
  assign data_o[13617] = data_o[49];
  assign data_o[13681] = data_o[49];
  assign data_o[13745] = data_o[49];
  assign data_o[13809] = data_o[49];
  assign data_o[13873] = data_o[49];
  assign data_o[13937] = data_o[49];
  assign data_o[14001] = data_o[49];
  assign data_o[14065] = data_o[49];
  assign data_o[14129] = data_o[49];
  assign data_o[14193] = data_o[49];
  assign data_o[14257] = data_o[49];
  assign data_o[14321] = data_o[49];
  assign data_o[14385] = data_o[49];
  assign data_o[14449] = data_o[49];
  assign data_o[14513] = data_o[49];
  assign data_o[14577] = data_o[49];
  assign data_o[14641] = data_o[49];
  assign data_o[14705] = data_o[49];
  assign data_o[14769] = data_o[49];
  assign data_o[14833] = data_o[49];
  assign data_o[14897] = data_o[49];
  assign data_o[14961] = data_o[49];
  assign data_o[15025] = data_o[49];
  assign data_o[15089] = data_o[49];
  assign data_o[15153] = data_o[49];
  assign data_o[15217] = data_o[49];
  assign data_o[15281] = data_o[49];
  assign data_o[15345] = data_o[49];
  assign data_o[15409] = data_o[49];
  assign data_o[15473] = data_o[49];
  assign data_o[15537] = data_o[49];
  assign data_o[15601] = data_o[49];
  assign data_o[15665] = data_o[49];
  assign data_o[15729] = data_o[49];
  assign data_o[15793] = data_o[49];
  assign data_o[15857] = data_o[49];
  assign data_o[15921] = data_o[49];
  assign data_o[15985] = data_o[49];
  assign data_o[16049] = data_o[49];
  assign data_o[16113] = data_o[49];
  assign data_o[16177] = data_o[49];
  assign data_o[16241] = data_o[49];
  assign data_o[16305] = data_o[49];
  assign data_o[16369] = data_o[49];
  assign data_o[16433] = data_o[49];
  assign data_o[16497] = data_o[49];
  assign data_o[16561] = data_o[49];
  assign data_o[16625] = data_o[49];
  assign data_o[16689] = data_o[49];
  assign data_o[16753] = data_o[49];
  assign data_o[16817] = data_o[49];
  assign data_o[16881] = data_o[49];
  assign data_o[16945] = data_o[49];
  assign data_o[17009] = data_o[49];
  assign data_o[17073] = data_o[49];
  assign data_o[17137] = data_o[49];
  assign data_o[17201] = data_o[49];
  assign data_o[17265] = data_o[49];
  assign data_o[17329] = data_o[49];
  assign data_o[17393] = data_o[49];
  assign data_o[17457] = data_o[49];
  assign data_o[17521] = data_o[49];
  assign data_o[17585] = data_o[49];
  assign data_o[17649] = data_o[49];
  assign data_o[17713] = data_o[49];
  assign data_o[17777] = data_o[49];
  assign data_o[17841] = data_o[49];
  assign data_o[17905] = data_o[49];
  assign data_o[17969] = data_o[49];
  assign data_o[18033] = data_o[49];
  assign data_o[18097] = data_o[49];
  assign data_o[18161] = data_o[49];
  assign data_o[18225] = data_o[49];
  assign data_o[18289] = data_o[49];
  assign data_o[18353] = data_o[49];
  assign data_o[18417] = data_o[49];
  assign data_o[18481] = data_o[49];
  assign data_o[18545] = data_o[49];
  assign data_o[18609] = data_o[49];
  assign data_o[18673] = data_o[49];
  assign data_o[18737] = data_o[49];
  assign data_o[18801] = data_o[49];
  assign data_o[18865] = data_o[49];
  assign data_o[18929] = data_o[49];
  assign data_o[18993] = data_o[49];
  assign data_o[19057] = data_o[49];
  assign data_o[19121] = data_o[49];
  assign data_o[19185] = data_o[49];
  assign data_o[19249] = data_o[49];
  assign data_o[19313] = data_o[49];
  assign data_o[19377] = data_o[49];
  assign data_o[19441] = data_o[49];
  assign data_o[19505] = data_o[49];
  assign data_o[19569] = data_o[49];
  assign data_o[19633] = data_o[49];
  assign data_o[19697] = data_o[49];
  assign data_o[19761] = data_o[49];
  assign data_o[19825] = data_o[49];
  assign data_o[19889] = data_o[49];
  assign data_o[19953] = data_o[49];
  assign data_o[20017] = data_o[49];
  assign data_o[20081] = data_o[49];
  assign data_o[20145] = data_o[49];
  assign data_o[20209] = data_o[49];
  assign data_o[20273] = data_o[49];
  assign data_o[20337] = data_o[49];
  assign data_o[20401] = data_o[49];
  assign data_o[20465] = data_o[49];
  assign data_o[20529] = data_o[49];
  assign data_o[20593] = data_o[49];
  assign data_o[20657] = data_o[49];
  assign data_o[20721] = data_o[49];
  assign data_o[20785] = data_o[49];
  assign data_o[20849] = data_o[49];
  assign data_o[20913] = data_o[49];
  assign data_o[20977] = data_o[49];
  assign data_o[21041] = data_o[49];
  assign data_o[21105] = data_o[49];
  assign data_o[21169] = data_o[49];
  assign data_o[21233] = data_o[49];
  assign data_o[21297] = data_o[49];
  assign data_o[21361] = data_o[49];
  assign data_o[21425] = data_o[49];
  assign data_o[21489] = data_o[49];
  assign data_o[21553] = data_o[49];
  assign data_o[21617] = data_o[49];
  assign data_o[21681] = data_o[49];
  assign data_o[21745] = data_o[49];
  assign data_o[21809] = data_o[49];
  assign data_o[21873] = data_o[49];
  assign data_o[21937] = data_o[49];
  assign data_o[22001] = data_o[49];
  assign data_o[22065] = data_o[49];
  assign data_o[22129] = data_o[49];
  assign data_o[22193] = data_o[49];
  assign data_o[22257] = data_o[49];
  assign data_o[22321] = data_o[49];
  assign data_o[22385] = data_o[49];
  assign data_o[22449] = data_o[49];
  assign data_o[22513] = data_o[49];
  assign data_o[22577] = data_o[49];
  assign data_o[22641] = data_o[49];
  assign data_o[22705] = data_o[49];
  assign data_o[22769] = data_o[49];
  assign data_o[22833] = data_o[49];
  assign data_o[22897] = data_o[49];
  assign data_o[22961] = data_o[49];
  assign data_o[23025] = data_o[49];
  assign data_o[23089] = data_o[49];
  assign data_o[23153] = data_o[49];
  assign data_o[23217] = data_o[49];
  assign data_o[23281] = data_o[49];
  assign data_o[23345] = data_o[49];
  assign data_o[23409] = data_o[49];
  assign data_o[23473] = data_o[49];
  assign data_o[23537] = data_o[49];
  assign data_o[23601] = data_o[49];
  assign data_o[23665] = data_o[49];
  assign data_o[23729] = data_o[49];
  assign data_o[23793] = data_o[49];
  assign data_o[23857] = data_o[49];
  assign data_o[23921] = data_o[49];
  assign data_o[23985] = data_o[49];
  assign data_o[24049] = data_o[49];
  assign data_o[24113] = data_o[49];
  assign data_o[24177] = data_o[49];
  assign data_o[24241] = data_o[49];
  assign data_o[24305] = data_o[49];
  assign data_o[24369] = data_o[49];
  assign data_o[24433] = data_o[49];
  assign data_o[24497] = data_o[49];
  assign data_o[24561] = data_o[49];
  assign data_o[24625] = data_o[49];
  assign data_o[24689] = data_o[49];
  assign data_o[24753] = data_o[49];
  assign data_o[24817] = data_o[49];
  assign data_o[24881] = data_o[49];
  assign data_o[24945] = data_o[49];
  assign data_o[25009] = data_o[49];
  assign data_o[25073] = data_o[49];
  assign data_o[25137] = data_o[49];
  assign data_o[25201] = data_o[49];
  assign data_o[25265] = data_o[49];
  assign data_o[25329] = data_o[49];
  assign data_o[25393] = data_o[49];
  assign data_o[25457] = data_o[49];
  assign data_o[25521] = data_o[49];
  assign data_o[25585] = data_o[49];
  assign data_o[25649] = data_o[49];
  assign data_o[25713] = data_o[49];
  assign data_o[25777] = data_o[49];
  assign data_o[25841] = data_o[49];
  assign data_o[25905] = data_o[49];
  assign data_o[25969] = data_o[49];
  assign data_o[26033] = data_o[49];
  assign data_o[26097] = data_o[49];
  assign data_o[26161] = data_o[49];
  assign data_o[26225] = data_o[49];
  assign data_o[26289] = data_o[49];
  assign data_o[26353] = data_o[49];
  assign data_o[26417] = data_o[49];
  assign data_o[26481] = data_o[49];
  assign data_o[26545] = data_o[49];
  assign data_o[26609] = data_o[49];
  assign data_o[26673] = data_o[49];
  assign data_o[26737] = data_o[49];
  assign data_o[26801] = data_o[49];
  assign data_o[26865] = data_o[49];
  assign data_o[26929] = data_o[49];
  assign data_o[26993] = data_o[49];
  assign data_o[27057] = data_o[49];
  assign data_o[27121] = data_o[49];
  assign data_o[27185] = data_o[49];
  assign data_o[27249] = data_o[49];
  assign data_o[27313] = data_o[49];
  assign data_o[27377] = data_o[49];
  assign data_o[27441] = data_o[49];
  assign data_o[27505] = data_o[49];
  assign data_o[27569] = data_o[49];
  assign data_o[27633] = data_o[49];
  assign data_o[27697] = data_o[49];
  assign data_o[27761] = data_o[49];
  assign data_o[27825] = data_o[49];
  assign data_o[27889] = data_o[49];
  assign data_o[27953] = data_o[49];
  assign data_o[28017] = data_o[49];
  assign data_o[28081] = data_o[49];
  assign data_o[28145] = data_o[49];
  assign data_o[28209] = data_o[49];
  assign data_o[28273] = data_o[49];
  assign data_o[28337] = data_o[49];
  assign data_o[28401] = data_o[49];
  assign data_o[28465] = data_o[49];
  assign data_o[28529] = data_o[49];
  assign data_o[28593] = data_o[49];
  assign data_o[28657] = data_o[49];
  assign data_o[28721] = data_o[49];
  assign data_o[28785] = data_o[49];
  assign data_o[28849] = data_o[49];
  assign data_o[28913] = data_o[49];
  assign data_o[28977] = data_o[49];
  assign data_o[29041] = data_o[49];
  assign data_o[29105] = data_o[49];
  assign data_o[29169] = data_o[49];
  assign data_o[29233] = data_o[49];
  assign data_o[29297] = data_o[49];
  assign data_o[29361] = data_o[49];
  assign data_o[29425] = data_o[49];
  assign data_o[29489] = data_o[49];
  assign data_o[29553] = data_o[49];
  assign data_o[29617] = data_o[49];
  assign data_o[29681] = data_o[49];
  assign data_o[29745] = data_o[49];
  assign data_o[29809] = data_o[49];
  assign data_o[29873] = data_o[49];
  assign data_o[29937] = data_o[49];
  assign data_o[30001] = data_o[49];
  assign data_o[30065] = data_o[49];
  assign data_o[30129] = data_o[49];
  assign data_o[30193] = data_o[49];
  assign data_o[30257] = data_o[49];
  assign data_o[30321] = data_o[49];
  assign data_o[30385] = data_o[49];
  assign data_o[30449] = data_o[49];
  assign data_o[30513] = data_o[49];
  assign data_o[30577] = data_o[49];
  assign data_o[30641] = data_o[49];
  assign data_o[30705] = data_o[49];
  assign data_o[30769] = data_o[49];
  assign data_o[30833] = data_o[49];
  assign data_o[30897] = data_o[49];
  assign data_o[30961] = data_o[49];
  assign data_o[31025] = data_o[49];
  assign data_o[31089] = data_o[49];
  assign data_o[31153] = data_o[49];
  assign data_o[31217] = data_o[49];
  assign data_o[31281] = data_o[49];
  assign data_o[31345] = data_o[49];
  assign data_o[31409] = data_o[49];
  assign data_o[31473] = data_o[49];
  assign data_o[31537] = data_o[49];
  assign data_o[31601] = data_o[49];
  assign data_o[31665] = data_o[49];
  assign data_o[31729] = data_o[49];
  assign data_o[31793] = data_o[49];
  assign data_o[31857] = data_o[49];
  assign data_o[31921] = data_o[49];
  assign data_o[31985] = data_o[49];
  assign data_o[112] = data_o[48];
  assign data_o[176] = data_o[48];
  assign data_o[240] = data_o[48];
  assign data_o[304] = data_o[48];
  assign data_o[368] = data_o[48];
  assign data_o[432] = data_o[48];
  assign data_o[496] = data_o[48];
  assign data_o[560] = data_o[48];
  assign data_o[624] = data_o[48];
  assign data_o[688] = data_o[48];
  assign data_o[752] = data_o[48];
  assign data_o[816] = data_o[48];
  assign data_o[880] = data_o[48];
  assign data_o[944] = data_o[48];
  assign data_o[1008] = data_o[48];
  assign data_o[1072] = data_o[48];
  assign data_o[1136] = data_o[48];
  assign data_o[1200] = data_o[48];
  assign data_o[1264] = data_o[48];
  assign data_o[1328] = data_o[48];
  assign data_o[1392] = data_o[48];
  assign data_o[1456] = data_o[48];
  assign data_o[1520] = data_o[48];
  assign data_o[1584] = data_o[48];
  assign data_o[1648] = data_o[48];
  assign data_o[1712] = data_o[48];
  assign data_o[1776] = data_o[48];
  assign data_o[1840] = data_o[48];
  assign data_o[1904] = data_o[48];
  assign data_o[1968] = data_o[48];
  assign data_o[2032] = data_o[48];
  assign data_o[2096] = data_o[48];
  assign data_o[2160] = data_o[48];
  assign data_o[2224] = data_o[48];
  assign data_o[2288] = data_o[48];
  assign data_o[2352] = data_o[48];
  assign data_o[2416] = data_o[48];
  assign data_o[2480] = data_o[48];
  assign data_o[2544] = data_o[48];
  assign data_o[2608] = data_o[48];
  assign data_o[2672] = data_o[48];
  assign data_o[2736] = data_o[48];
  assign data_o[2800] = data_o[48];
  assign data_o[2864] = data_o[48];
  assign data_o[2928] = data_o[48];
  assign data_o[2992] = data_o[48];
  assign data_o[3056] = data_o[48];
  assign data_o[3120] = data_o[48];
  assign data_o[3184] = data_o[48];
  assign data_o[3248] = data_o[48];
  assign data_o[3312] = data_o[48];
  assign data_o[3376] = data_o[48];
  assign data_o[3440] = data_o[48];
  assign data_o[3504] = data_o[48];
  assign data_o[3568] = data_o[48];
  assign data_o[3632] = data_o[48];
  assign data_o[3696] = data_o[48];
  assign data_o[3760] = data_o[48];
  assign data_o[3824] = data_o[48];
  assign data_o[3888] = data_o[48];
  assign data_o[3952] = data_o[48];
  assign data_o[4016] = data_o[48];
  assign data_o[4080] = data_o[48];
  assign data_o[4144] = data_o[48];
  assign data_o[4208] = data_o[48];
  assign data_o[4272] = data_o[48];
  assign data_o[4336] = data_o[48];
  assign data_o[4400] = data_o[48];
  assign data_o[4464] = data_o[48];
  assign data_o[4528] = data_o[48];
  assign data_o[4592] = data_o[48];
  assign data_o[4656] = data_o[48];
  assign data_o[4720] = data_o[48];
  assign data_o[4784] = data_o[48];
  assign data_o[4848] = data_o[48];
  assign data_o[4912] = data_o[48];
  assign data_o[4976] = data_o[48];
  assign data_o[5040] = data_o[48];
  assign data_o[5104] = data_o[48];
  assign data_o[5168] = data_o[48];
  assign data_o[5232] = data_o[48];
  assign data_o[5296] = data_o[48];
  assign data_o[5360] = data_o[48];
  assign data_o[5424] = data_o[48];
  assign data_o[5488] = data_o[48];
  assign data_o[5552] = data_o[48];
  assign data_o[5616] = data_o[48];
  assign data_o[5680] = data_o[48];
  assign data_o[5744] = data_o[48];
  assign data_o[5808] = data_o[48];
  assign data_o[5872] = data_o[48];
  assign data_o[5936] = data_o[48];
  assign data_o[6000] = data_o[48];
  assign data_o[6064] = data_o[48];
  assign data_o[6128] = data_o[48];
  assign data_o[6192] = data_o[48];
  assign data_o[6256] = data_o[48];
  assign data_o[6320] = data_o[48];
  assign data_o[6384] = data_o[48];
  assign data_o[6448] = data_o[48];
  assign data_o[6512] = data_o[48];
  assign data_o[6576] = data_o[48];
  assign data_o[6640] = data_o[48];
  assign data_o[6704] = data_o[48];
  assign data_o[6768] = data_o[48];
  assign data_o[6832] = data_o[48];
  assign data_o[6896] = data_o[48];
  assign data_o[6960] = data_o[48];
  assign data_o[7024] = data_o[48];
  assign data_o[7088] = data_o[48];
  assign data_o[7152] = data_o[48];
  assign data_o[7216] = data_o[48];
  assign data_o[7280] = data_o[48];
  assign data_o[7344] = data_o[48];
  assign data_o[7408] = data_o[48];
  assign data_o[7472] = data_o[48];
  assign data_o[7536] = data_o[48];
  assign data_o[7600] = data_o[48];
  assign data_o[7664] = data_o[48];
  assign data_o[7728] = data_o[48];
  assign data_o[7792] = data_o[48];
  assign data_o[7856] = data_o[48];
  assign data_o[7920] = data_o[48];
  assign data_o[7984] = data_o[48];
  assign data_o[8048] = data_o[48];
  assign data_o[8112] = data_o[48];
  assign data_o[8176] = data_o[48];
  assign data_o[8240] = data_o[48];
  assign data_o[8304] = data_o[48];
  assign data_o[8368] = data_o[48];
  assign data_o[8432] = data_o[48];
  assign data_o[8496] = data_o[48];
  assign data_o[8560] = data_o[48];
  assign data_o[8624] = data_o[48];
  assign data_o[8688] = data_o[48];
  assign data_o[8752] = data_o[48];
  assign data_o[8816] = data_o[48];
  assign data_o[8880] = data_o[48];
  assign data_o[8944] = data_o[48];
  assign data_o[9008] = data_o[48];
  assign data_o[9072] = data_o[48];
  assign data_o[9136] = data_o[48];
  assign data_o[9200] = data_o[48];
  assign data_o[9264] = data_o[48];
  assign data_o[9328] = data_o[48];
  assign data_o[9392] = data_o[48];
  assign data_o[9456] = data_o[48];
  assign data_o[9520] = data_o[48];
  assign data_o[9584] = data_o[48];
  assign data_o[9648] = data_o[48];
  assign data_o[9712] = data_o[48];
  assign data_o[9776] = data_o[48];
  assign data_o[9840] = data_o[48];
  assign data_o[9904] = data_o[48];
  assign data_o[9968] = data_o[48];
  assign data_o[10032] = data_o[48];
  assign data_o[10096] = data_o[48];
  assign data_o[10160] = data_o[48];
  assign data_o[10224] = data_o[48];
  assign data_o[10288] = data_o[48];
  assign data_o[10352] = data_o[48];
  assign data_o[10416] = data_o[48];
  assign data_o[10480] = data_o[48];
  assign data_o[10544] = data_o[48];
  assign data_o[10608] = data_o[48];
  assign data_o[10672] = data_o[48];
  assign data_o[10736] = data_o[48];
  assign data_o[10800] = data_o[48];
  assign data_o[10864] = data_o[48];
  assign data_o[10928] = data_o[48];
  assign data_o[10992] = data_o[48];
  assign data_o[11056] = data_o[48];
  assign data_o[11120] = data_o[48];
  assign data_o[11184] = data_o[48];
  assign data_o[11248] = data_o[48];
  assign data_o[11312] = data_o[48];
  assign data_o[11376] = data_o[48];
  assign data_o[11440] = data_o[48];
  assign data_o[11504] = data_o[48];
  assign data_o[11568] = data_o[48];
  assign data_o[11632] = data_o[48];
  assign data_o[11696] = data_o[48];
  assign data_o[11760] = data_o[48];
  assign data_o[11824] = data_o[48];
  assign data_o[11888] = data_o[48];
  assign data_o[11952] = data_o[48];
  assign data_o[12016] = data_o[48];
  assign data_o[12080] = data_o[48];
  assign data_o[12144] = data_o[48];
  assign data_o[12208] = data_o[48];
  assign data_o[12272] = data_o[48];
  assign data_o[12336] = data_o[48];
  assign data_o[12400] = data_o[48];
  assign data_o[12464] = data_o[48];
  assign data_o[12528] = data_o[48];
  assign data_o[12592] = data_o[48];
  assign data_o[12656] = data_o[48];
  assign data_o[12720] = data_o[48];
  assign data_o[12784] = data_o[48];
  assign data_o[12848] = data_o[48];
  assign data_o[12912] = data_o[48];
  assign data_o[12976] = data_o[48];
  assign data_o[13040] = data_o[48];
  assign data_o[13104] = data_o[48];
  assign data_o[13168] = data_o[48];
  assign data_o[13232] = data_o[48];
  assign data_o[13296] = data_o[48];
  assign data_o[13360] = data_o[48];
  assign data_o[13424] = data_o[48];
  assign data_o[13488] = data_o[48];
  assign data_o[13552] = data_o[48];
  assign data_o[13616] = data_o[48];
  assign data_o[13680] = data_o[48];
  assign data_o[13744] = data_o[48];
  assign data_o[13808] = data_o[48];
  assign data_o[13872] = data_o[48];
  assign data_o[13936] = data_o[48];
  assign data_o[14000] = data_o[48];
  assign data_o[14064] = data_o[48];
  assign data_o[14128] = data_o[48];
  assign data_o[14192] = data_o[48];
  assign data_o[14256] = data_o[48];
  assign data_o[14320] = data_o[48];
  assign data_o[14384] = data_o[48];
  assign data_o[14448] = data_o[48];
  assign data_o[14512] = data_o[48];
  assign data_o[14576] = data_o[48];
  assign data_o[14640] = data_o[48];
  assign data_o[14704] = data_o[48];
  assign data_o[14768] = data_o[48];
  assign data_o[14832] = data_o[48];
  assign data_o[14896] = data_o[48];
  assign data_o[14960] = data_o[48];
  assign data_o[15024] = data_o[48];
  assign data_o[15088] = data_o[48];
  assign data_o[15152] = data_o[48];
  assign data_o[15216] = data_o[48];
  assign data_o[15280] = data_o[48];
  assign data_o[15344] = data_o[48];
  assign data_o[15408] = data_o[48];
  assign data_o[15472] = data_o[48];
  assign data_o[15536] = data_o[48];
  assign data_o[15600] = data_o[48];
  assign data_o[15664] = data_o[48];
  assign data_o[15728] = data_o[48];
  assign data_o[15792] = data_o[48];
  assign data_o[15856] = data_o[48];
  assign data_o[15920] = data_o[48];
  assign data_o[15984] = data_o[48];
  assign data_o[16048] = data_o[48];
  assign data_o[16112] = data_o[48];
  assign data_o[16176] = data_o[48];
  assign data_o[16240] = data_o[48];
  assign data_o[16304] = data_o[48];
  assign data_o[16368] = data_o[48];
  assign data_o[16432] = data_o[48];
  assign data_o[16496] = data_o[48];
  assign data_o[16560] = data_o[48];
  assign data_o[16624] = data_o[48];
  assign data_o[16688] = data_o[48];
  assign data_o[16752] = data_o[48];
  assign data_o[16816] = data_o[48];
  assign data_o[16880] = data_o[48];
  assign data_o[16944] = data_o[48];
  assign data_o[17008] = data_o[48];
  assign data_o[17072] = data_o[48];
  assign data_o[17136] = data_o[48];
  assign data_o[17200] = data_o[48];
  assign data_o[17264] = data_o[48];
  assign data_o[17328] = data_o[48];
  assign data_o[17392] = data_o[48];
  assign data_o[17456] = data_o[48];
  assign data_o[17520] = data_o[48];
  assign data_o[17584] = data_o[48];
  assign data_o[17648] = data_o[48];
  assign data_o[17712] = data_o[48];
  assign data_o[17776] = data_o[48];
  assign data_o[17840] = data_o[48];
  assign data_o[17904] = data_o[48];
  assign data_o[17968] = data_o[48];
  assign data_o[18032] = data_o[48];
  assign data_o[18096] = data_o[48];
  assign data_o[18160] = data_o[48];
  assign data_o[18224] = data_o[48];
  assign data_o[18288] = data_o[48];
  assign data_o[18352] = data_o[48];
  assign data_o[18416] = data_o[48];
  assign data_o[18480] = data_o[48];
  assign data_o[18544] = data_o[48];
  assign data_o[18608] = data_o[48];
  assign data_o[18672] = data_o[48];
  assign data_o[18736] = data_o[48];
  assign data_o[18800] = data_o[48];
  assign data_o[18864] = data_o[48];
  assign data_o[18928] = data_o[48];
  assign data_o[18992] = data_o[48];
  assign data_o[19056] = data_o[48];
  assign data_o[19120] = data_o[48];
  assign data_o[19184] = data_o[48];
  assign data_o[19248] = data_o[48];
  assign data_o[19312] = data_o[48];
  assign data_o[19376] = data_o[48];
  assign data_o[19440] = data_o[48];
  assign data_o[19504] = data_o[48];
  assign data_o[19568] = data_o[48];
  assign data_o[19632] = data_o[48];
  assign data_o[19696] = data_o[48];
  assign data_o[19760] = data_o[48];
  assign data_o[19824] = data_o[48];
  assign data_o[19888] = data_o[48];
  assign data_o[19952] = data_o[48];
  assign data_o[20016] = data_o[48];
  assign data_o[20080] = data_o[48];
  assign data_o[20144] = data_o[48];
  assign data_o[20208] = data_o[48];
  assign data_o[20272] = data_o[48];
  assign data_o[20336] = data_o[48];
  assign data_o[20400] = data_o[48];
  assign data_o[20464] = data_o[48];
  assign data_o[20528] = data_o[48];
  assign data_o[20592] = data_o[48];
  assign data_o[20656] = data_o[48];
  assign data_o[20720] = data_o[48];
  assign data_o[20784] = data_o[48];
  assign data_o[20848] = data_o[48];
  assign data_o[20912] = data_o[48];
  assign data_o[20976] = data_o[48];
  assign data_o[21040] = data_o[48];
  assign data_o[21104] = data_o[48];
  assign data_o[21168] = data_o[48];
  assign data_o[21232] = data_o[48];
  assign data_o[21296] = data_o[48];
  assign data_o[21360] = data_o[48];
  assign data_o[21424] = data_o[48];
  assign data_o[21488] = data_o[48];
  assign data_o[21552] = data_o[48];
  assign data_o[21616] = data_o[48];
  assign data_o[21680] = data_o[48];
  assign data_o[21744] = data_o[48];
  assign data_o[21808] = data_o[48];
  assign data_o[21872] = data_o[48];
  assign data_o[21936] = data_o[48];
  assign data_o[22000] = data_o[48];
  assign data_o[22064] = data_o[48];
  assign data_o[22128] = data_o[48];
  assign data_o[22192] = data_o[48];
  assign data_o[22256] = data_o[48];
  assign data_o[22320] = data_o[48];
  assign data_o[22384] = data_o[48];
  assign data_o[22448] = data_o[48];
  assign data_o[22512] = data_o[48];
  assign data_o[22576] = data_o[48];
  assign data_o[22640] = data_o[48];
  assign data_o[22704] = data_o[48];
  assign data_o[22768] = data_o[48];
  assign data_o[22832] = data_o[48];
  assign data_o[22896] = data_o[48];
  assign data_o[22960] = data_o[48];
  assign data_o[23024] = data_o[48];
  assign data_o[23088] = data_o[48];
  assign data_o[23152] = data_o[48];
  assign data_o[23216] = data_o[48];
  assign data_o[23280] = data_o[48];
  assign data_o[23344] = data_o[48];
  assign data_o[23408] = data_o[48];
  assign data_o[23472] = data_o[48];
  assign data_o[23536] = data_o[48];
  assign data_o[23600] = data_o[48];
  assign data_o[23664] = data_o[48];
  assign data_o[23728] = data_o[48];
  assign data_o[23792] = data_o[48];
  assign data_o[23856] = data_o[48];
  assign data_o[23920] = data_o[48];
  assign data_o[23984] = data_o[48];
  assign data_o[24048] = data_o[48];
  assign data_o[24112] = data_o[48];
  assign data_o[24176] = data_o[48];
  assign data_o[24240] = data_o[48];
  assign data_o[24304] = data_o[48];
  assign data_o[24368] = data_o[48];
  assign data_o[24432] = data_o[48];
  assign data_o[24496] = data_o[48];
  assign data_o[24560] = data_o[48];
  assign data_o[24624] = data_o[48];
  assign data_o[24688] = data_o[48];
  assign data_o[24752] = data_o[48];
  assign data_o[24816] = data_o[48];
  assign data_o[24880] = data_o[48];
  assign data_o[24944] = data_o[48];
  assign data_o[25008] = data_o[48];
  assign data_o[25072] = data_o[48];
  assign data_o[25136] = data_o[48];
  assign data_o[25200] = data_o[48];
  assign data_o[25264] = data_o[48];
  assign data_o[25328] = data_o[48];
  assign data_o[25392] = data_o[48];
  assign data_o[25456] = data_o[48];
  assign data_o[25520] = data_o[48];
  assign data_o[25584] = data_o[48];
  assign data_o[25648] = data_o[48];
  assign data_o[25712] = data_o[48];
  assign data_o[25776] = data_o[48];
  assign data_o[25840] = data_o[48];
  assign data_o[25904] = data_o[48];
  assign data_o[25968] = data_o[48];
  assign data_o[26032] = data_o[48];
  assign data_o[26096] = data_o[48];
  assign data_o[26160] = data_o[48];
  assign data_o[26224] = data_o[48];
  assign data_o[26288] = data_o[48];
  assign data_o[26352] = data_o[48];
  assign data_o[26416] = data_o[48];
  assign data_o[26480] = data_o[48];
  assign data_o[26544] = data_o[48];
  assign data_o[26608] = data_o[48];
  assign data_o[26672] = data_o[48];
  assign data_o[26736] = data_o[48];
  assign data_o[26800] = data_o[48];
  assign data_o[26864] = data_o[48];
  assign data_o[26928] = data_o[48];
  assign data_o[26992] = data_o[48];
  assign data_o[27056] = data_o[48];
  assign data_o[27120] = data_o[48];
  assign data_o[27184] = data_o[48];
  assign data_o[27248] = data_o[48];
  assign data_o[27312] = data_o[48];
  assign data_o[27376] = data_o[48];
  assign data_o[27440] = data_o[48];
  assign data_o[27504] = data_o[48];
  assign data_o[27568] = data_o[48];
  assign data_o[27632] = data_o[48];
  assign data_o[27696] = data_o[48];
  assign data_o[27760] = data_o[48];
  assign data_o[27824] = data_o[48];
  assign data_o[27888] = data_o[48];
  assign data_o[27952] = data_o[48];
  assign data_o[28016] = data_o[48];
  assign data_o[28080] = data_o[48];
  assign data_o[28144] = data_o[48];
  assign data_o[28208] = data_o[48];
  assign data_o[28272] = data_o[48];
  assign data_o[28336] = data_o[48];
  assign data_o[28400] = data_o[48];
  assign data_o[28464] = data_o[48];
  assign data_o[28528] = data_o[48];
  assign data_o[28592] = data_o[48];
  assign data_o[28656] = data_o[48];
  assign data_o[28720] = data_o[48];
  assign data_o[28784] = data_o[48];
  assign data_o[28848] = data_o[48];
  assign data_o[28912] = data_o[48];
  assign data_o[28976] = data_o[48];
  assign data_o[29040] = data_o[48];
  assign data_o[29104] = data_o[48];
  assign data_o[29168] = data_o[48];
  assign data_o[29232] = data_o[48];
  assign data_o[29296] = data_o[48];
  assign data_o[29360] = data_o[48];
  assign data_o[29424] = data_o[48];
  assign data_o[29488] = data_o[48];
  assign data_o[29552] = data_o[48];
  assign data_o[29616] = data_o[48];
  assign data_o[29680] = data_o[48];
  assign data_o[29744] = data_o[48];
  assign data_o[29808] = data_o[48];
  assign data_o[29872] = data_o[48];
  assign data_o[29936] = data_o[48];
  assign data_o[30000] = data_o[48];
  assign data_o[30064] = data_o[48];
  assign data_o[30128] = data_o[48];
  assign data_o[30192] = data_o[48];
  assign data_o[30256] = data_o[48];
  assign data_o[30320] = data_o[48];
  assign data_o[30384] = data_o[48];
  assign data_o[30448] = data_o[48];
  assign data_o[30512] = data_o[48];
  assign data_o[30576] = data_o[48];
  assign data_o[30640] = data_o[48];
  assign data_o[30704] = data_o[48];
  assign data_o[30768] = data_o[48];
  assign data_o[30832] = data_o[48];
  assign data_o[30896] = data_o[48];
  assign data_o[30960] = data_o[48];
  assign data_o[31024] = data_o[48];
  assign data_o[31088] = data_o[48];
  assign data_o[31152] = data_o[48];
  assign data_o[31216] = data_o[48];
  assign data_o[31280] = data_o[48];
  assign data_o[31344] = data_o[48];
  assign data_o[31408] = data_o[48];
  assign data_o[31472] = data_o[48];
  assign data_o[31536] = data_o[48];
  assign data_o[31600] = data_o[48];
  assign data_o[31664] = data_o[48];
  assign data_o[31728] = data_o[48];
  assign data_o[31792] = data_o[48];
  assign data_o[31856] = data_o[48];
  assign data_o[31920] = data_o[48];
  assign data_o[31984] = data_o[48];
  assign data_o[111] = data_o[47];
  assign data_o[175] = data_o[47];
  assign data_o[239] = data_o[47];
  assign data_o[303] = data_o[47];
  assign data_o[367] = data_o[47];
  assign data_o[431] = data_o[47];
  assign data_o[495] = data_o[47];
  assign data_o[559] = data_o[47];
  assign data_o[623] = data_o[47];
  assign data_o[687] = data_o[47];
  assign data_o[751] = data_o[47];
  assign data_o[815] = data_o[47];
  assign data_o[879] = data_o[47];
  assign data_o[943] = data_o[47];
  assign data_o[1007] = data_o[47];
  assign data_o[1071] = data_o[47];
  assign data_o[1135] = data_o[47];
  assign data_o[1199] = data_o[47];
  assign data_o[1263] = data_o[47];
  assign data_o[1327] = data_o[47];
  assign data_o[1391] = data_o[47];
  assign data_o[1455] = data_o[47];
  assign data_o[1519] = data_o[47];
  assign data_o[1583] = data_o[47];
  assign data_o[1647] = data_o[47];
  assign data_o[1711] = data_o[47];
  assign data_o[1775] = data_o[47];
  assign data_o[1839] = data_o[47];
  assign data_o[1903] = data_o[47];
  assign data_o[1967] = data_o[47];
  assign data_o[2031] = data_o[47];
  assign data_o[2095] = data_o[47];
  assign data_o[2159] = data_o[47];
  assign data_o[2223] = data_o[47];
  assign data_o[2287] = data_o[47];
  assign data_o[2351] = data_o[47];
  assign data_o[2415] = data_o[47];
  assign data_o[2479] = data_o[47];
  assign data_o[2543] = data_o[47];
  assign data_o[2607] = data_o[47];
  assign data_o[2671] = data_o[47];
  assign data_o[2735] = data_o[47];
  assign data_o[2799] = data_o[47];
  assign data_o[2863] = data_o[47];
  assign data_o[2927] = data_o[47];
  assign data_o[2991] = data_o[47];
  assign data_o[3055] = data_o[47];
  assign data_o[3119] = data_o[47];
  assign data_o[3183] = data_o[47];
  assign data_o[3247] = data_o[47];
  assign data_o[3311] = data_o[47];
  assign data_o[3375] = data_o[47];
  assign data_o[3439] = data_o[47];
  assign data_o[3503] = data_o[47];
  assign data_o[3567] = data_o[47];
  assign data_o[3631] = data_o[47];
  assign data_o[3695] = data_o[47];
  assign data_o[3759] = data_o[47];
  assign data_o[3823] = data_o[47];
  assign data_o[3887] = data_o[47];
  assign data_o[3951] = data_o[47];
  assign data_o[4015] = data_o[47];
  assign data_o[4079] = data_o[47];
  assign data_o[4143] = data_o[47];
  assign data_o[4207] = data_o[47];
  assign data_o[4271] = data_o[47];
  assign data_o[4335] = data_o[47];
  assign data_o[4399] = data_o[47];
  assign data_o[4463] = data_o[47];
  assign data_o[4527] = data_o[47];
  assign data_o[4591] = data_o[47];
  assign data_o[4655] = data_o[47];
  assign data_o[4719] = data_o[47];
  assign data_o[4783] = data_o[47];
  assign data_o[4847] = data_o[47];
  assign data_o[4911] = data_o[47];
  assign data_o[4975] = data_o[47];
  assign data_o[5039] = data_o[47];
  assign data_o[5103] = data_o[47];
  assign data_o[5167] = data_o[47];
  assign data_o[5231] = data_o[47];
  assign data_o[5295] = data_o[47];
  assign data_o[5359] = data_o[47];
  assign data_o[5423] = data_o[47];
  assign data_o[5487] = data_o[47];
  assign data_o[5551] = data_o[47];
  assign data_o[5615] = data_o[47];
  assign data_o[5679] = data_o[47];
  assign data_o[5743] = data_o[47];
  assign data_o[5807] = data_o[47];
  assign data_o[5871] = data_o[47];
  assign data_o[5935] = data_o[47];
  assign data_o[5999] = data_o[47];
  assign data_o[6063] = data_o[47];
  assign data_o[6127] = data_o[47];
  assign data_o[6191] = data_o[47];
  assign data_o[6255] = data_o[47];
  assign data_o[6319] = data_o[47];
  assign data_o[6383] = data_o[47];
  assign data_o[6447] = data_o[47];
  assign data_o[6511] = data_o[47];
  assign data_o[6575] = data_o[47];
  assign data_o[6639] = data_o[47];
  assign data_o[6703] = data_o[47];
  assign data_o[6767] = data_o[47];
  assign data_o[6831] = data_o[47];
  assign data_o[6895] = data_o[47];
  assign data_o[6959] = data_o[47];
  assign data_o[7023] = data_o[47];
  assign data_o[7087] = data_o[47];
  assign data_o[7151] = data_o[47];
  assign data_o[7215] = data_o[47];
  assign data_o[7279] = data_o[47];
  assign data_o[7343] = data_o[47];
  assign data_o[7407] = data_o[47];
  assign data_o[7471] = data_o[47];
  assign data_o[7535] = data_o[47];
  assign data_o[7599] = data_o[47];
  assign data_o[7663] = data_o[47];
  assign data_o[7727] = data_o[47];
  assign data_o[7791] = data_o[47];
  assign data_o[7855] = data_o[47];
  assign data_o[7919] = data_o[47];
  assign data_o[7983] = data_o[47];
  assign data_o[8047] = data_o[47];
  assign data_o[8111] = data_o[47];
  assign data_o[8175] = data_o[47];
  assign data_o[8239] = data_o[47];
  assign data_o[8303] = data_o[47];
  assign data_o[8367] = data_o[47];
  assign data_o[8431] = data_o[47];
  assign data_o[8495] = data_o[47];
  assign data_o[8559] = data_o[47];
  assign data_o[8623] = data_o[47];
  assign data_o[8687] = data_o[47];
  assign data_o[8751] = data_o[47];
  assign data_o[8815] = data_o[47];
  assign data_o[8879] = data_o[47];
  assign data_o[8943] = data_o[47];
  assign data_o[9007] = data_o[47];
  assign data_o[9071] = data_o[47];
  assign data_o[9135] = data_o[47];
  assign data_o[9199] = data_o[47];
  assign data_o[9263] = data_o[47];
  assign data_o[9327] = data_o[47];
  assign data_o[9391] = data_o[47];
  assign data_o[9455] = data_o[47];
  assign data_o[9519] = data_o[47];
  assign data_o[9583] = data_o[47];
  assign data_o[9647] = data_o[47];
  assign data_o[9711] = data_o[47];
  assign data_o[9775] = data_o[47];
  assign data_o[9839] = data_o[47];
  assign data_o[9903] = data_o[47];
  assign data_o[9967] = data_o[47];
  assign data_o[10031] = data_o[47];
  assign data_o[10095] = data_o[47];
  assign data_o[10159] = data_o[47];
  assign data_o[10223] = data_o[47];
  assign data_o[10287] = data_o[47];
  assign data_o[10351] = data_o[47];
  assign data_o[10415] = data_o[47];
  assign data_o[10479] = data_o[47];
  assign data_o[10543] = data_o[47];
  assign data_o[10607] = data_o[47];
  assign data_o[10671] = data_o[47];
  assign data_o[10735] = data_o[47];
  assign data_o[10799] = data_o[47];
  assign data_o[10863] = data_o[47];
  assign data_o[10927] = data_o[47];
  assign data_o[10991] = data_o[47];
  assign data_o[11055] = data_o[47];
  assign data_o[11119] = data_o[47];
  assign data_o[11183] = data_o[47];
  assign data_o[11247] = data_o[47];
  assign data_o[11311] = data_o[47];
  assign data_o[11375] = data_o[47];
  assign data_o[11439] = data_o[47];
  assign data_o[11503] = data_o[47];
  assign data_o[11567] = data_o[47];
  assign data_o[11631] = data_o[47];
  assign data_o[11695] = data_o[47];
  assign data_o[11759] = data_o[47];
  assign data_o[11823] = data_o[47];
  assign data_o[11887] = data_o[47];
  assign data_o[11951] = data_o[47];
  assign data_o[12015] = data_o[47];
  assign data_o[12079] = data_o[47];
  assign data_o[12143] = data_o[47];
  assign data_o[12207] = data_o[47];
  assign data_o[12271] = data_o[47];
  assign data_o[12335] = data_o[47];
  assign data_o[12399] = data_o[47];
  assign data_o[12463] = data_o[47];
  assign data_o[12527] = data_o[47];
  assign data_o[12591] = data_o[47];
  assign data_o[12655] = data_o[47];
  assign data_o[12719] = data_o[47];
  assign data_o[12783] = data_o[47];
  assign data_o[12847] = data_o[47];
  assign data_o[12911] = data_o[47];
  assign data_o[12975] = data_o[47];
  assign data_o[13039] = data_o[47];
  assign data_o[13103] = data_o[47];
  assign data_o[13167] = data_o[47];
  assign data_o[13231] = data_o[47];
  assign data_o[13295] = data_o[47];
  assign data_o[13359] = data_o[47];
  assign data_o[13423] = data_o[47];
  assign data_o[13487] = data_o[47];
  assign data_o[13551] = data_o[47];
  assign data_o[13615] = data_o[47];
  assign data_o[13679] = data_o[47];
  assign data_o[13743] = data_o[47];
  assign data_o[13807] = data_o[47];
  assign data_o[13871] = data_o[47];
  assign data_o[13935] = data_o[47];
  assign data_o[13999] = data_o[47];
  assign data_o[14063] = data_o[47];
  assign data_o[14127] = data_o[47];
  assign data_o[14191] = data_o[47];
  assign data_o[14255] = data_o[47];
  assign data_o[14319] = data_o[47];
  assign data_o[14383] = data_o[47];
  assign data_o[14447] = data_o[47];
  assign data_o[14511] = data_o[47];
  assign data_o[14575] = data_o[47];
  assign data_o[14639] = data_o[47];
  assign data_o[14703] = data_o[47];
  assign data_o[14767] = data_o[47];
  assign data_o[14831] = data_o[47];
  assign data_o[14895] = data_o[47];
  assign data_o[14959] = data_o[47];
  assign data_o[15023] = data_o[47];
  assign data_o[15087] = data_o[47];
  assign data_o[15151] = data_o[47];
  assign data_o[15215] = data_o[47];
  assign data_o[15279] = data_o[47];
  assign data_o[15343] = data_o[47];
  assign data_o[15407] = data_o[47];
  assign data_o[15471] = data_o[47];
  assign data_o[15535] = data_o[47];
  assign data_o[15599] = data_o[47];
  assign data_o[15663] = data_o[47];
  assign data_o[15727] = data_o[47];
  assign data_o[15791] = data_o[47];
  assign data_o[15855] = data_o[47];
  assign data_o[15919] = data_o[47];
  assign data_o[15983] = data_o[47];
  assign data_o[16047] = data_o[47];
  assign data_o[16111] = data_o[47];
  assign data_o[16175] = data_o[47];
  assign data_o[16239] = data_o[47];
  assign data_o[16303] = data_o[47];
  assign data_o[16367] = data_o[47];
  assign data_o[16431] = data_o[47];
  assign data_o[16495] = data_o[47];
  assign data_o[16559] = data_o[47];
  assign data_o[16623] = data_o[47];
  assign data_o[16687] = data_o[47];
  assign data_o[16751] = data_o[47];
  assign data_o[16815] = data_o[47];
  assign data_o[16879] = data_o[47];
  assign data_o[16943] = data_o[47];
  assign data_o[17007] = data_o[47];
  assign data_o[17071] = data_o[47];
  assign data_o[17135] = data_o[47];
  assign data_o[17199] = data_o[47];
  assign data_o[17263] = data_o[47];
  assign data_o[17327] = data_o[47];
  assign data_o[17391] = data_o[47];
  assign data_o[17455] = data_o[47];
  assign data_o[17519] = data_o[47];
  assign data_o[17583] = data_o[47];
  assign data_o[17647] = data_o[47];
  assign data_o[17711] = data_o[47];
  assign data_o[17775] = data_o[47];
  assign data_o[17839] = data_o[47];
  assign data_o[17903] = data_o[47];
  assign data_o[17967] = data_o[47];
  assign data_o[18031] = data_o[47];
  assign data_o[18095] = data_o[47];
  assign data_o[18159] = data_o[47];
  assign data_o[18223] = data_o[47];
  assign data_o[18287] = data_o[47];
  assign data_o[18351] = data_o[47];
  assign data_o[18415] = data_o[47];
  assign data_o[18479] = data_o[47];
  assign data_o[18543] = data_o[47];
  assign data_o[18607] = data_o[47];
  assign data_o[18671] = data_o[47];
  assign data_o[18735] = data_o[47];
  assign data_o[18799] = data_o[47];
  assign data_o[18863] = data_o[47];
  assign data_o[18927] = data_o[47];
  assign data_o[18991] = data_o[47];
  assign data_o[19055] = data_o[47];
  assign data_o[19119] = data_o[47];
  assign data_o[19183] = data_o[47];
  assign data_o[19247] = data_o[47];
  assign data_o[19311] = data_o[47];
  assign data_o[19375] = data_o[47];
  assign data_o[19439] = data_o[47];
  assign data_o[19503] = data_o[47];
  assign data_o[19567] = data_o[47];
  assign data_o[19631] = data_o[47];
  assign data_o[19695] = data_o[47];
  assign data_o[19759] = data_o[47];
  assign data_o[19823] = data_o[47];
  assign data_o[19887] = data_o[47];
  assign data_o[19951] = data_o[47];
  assign data_o[20015] = data_o[47];
  assign data_o[20079] = data_o[47];
  assign data_o[20143] = data_o[47];
  assign data_o[20207] = data_o[47];
  assign data_o[20271] = data_o[47];
  assign data_o[20335] = data_o[47];
  assign data_o[20399] = data_o[47];
  assign data_o[20463] = data_o[47];
  assign data_o[20527] = data_o[47];
  assign data_o[20591] = data_o[47];
  assign data_o[20655] = data_o[47];
  assign data_o[20719] = data_o[47];
  assign data_o[20783] = data_o[47];
  assign data_o[20847] = data_o[47];
  assign data_o[20911] = data_o[47];
  assign data_o[20975] = data_o[47];
  assign data_o[21039] = data_o[47];
  assign data_o[21103] = data_o[47];
  assign data_o[21167] = data_o[47];
  assign data_o[21231] = data_o[47];
  assign data_o[21295] = data_o[47];
  assign data_o[21359] = data_o[47];
  assign data_o[21423] = data_o[47];
  assign data_o[21487] = data_o[47];
  assign data_o[21551] = data_o[47];
  assign data_o[21615] = data_o[47];
  assign data_o[21679] = data_o[47];
  assign data_o[21743] = data_o[47];
  assign data_o[21807] = data_o[47];
  assign data_o[21871] = data_o[47];
  assign data_o[21935] = data_o[47];
  assign data_o[21999] = data_o[47];
  assign data_o[22063] = data_o[47];
  assign data_o[22127] = data_o[47];
  assign data_o[22191] = data_o[47];
  assign data_o[22255] = data_o[47];
  assign data_o[22319] = data_o[47];
  assign data_o[22383] = data_o[47];
  assign data_o[22447] = data_o[47];
  assign data_o[22511] = data_o[47];
  assign data_o[22575] = data_o[47];
  assign data_o[22639] = data_o[47];
  assign data_o[22703] = data_o[47];
  assign data_o[22767] = data_o[47];
  assign data_o[22831] = data_o[47];
  assign data_o[22895] = data_o[47];
  assign data_o[22959] = data_o[47];
  assign data_o[23023] = data_o[47];
  assign data_o[23087] = data_o[47];
  assign data_o[23151] = data_o[47];
  assign data_o[23215] = data_o[47];
  assign data_o[23279] = data_o[47];
  assign data_o[23343] = data_o[47];
  assign data_o[23407] = data_o[47];
  assign data_o[23471] = data_o[47];
  assign data_o[23535] = data_o[47];
  assign data_o[23599] = data_o[47];
  assign data_o[23663] = data_o[47];
  assign data_o[23727] = data_o[47];
  assign data_o[23791] = data_o[47];
  assign data_o[23855] = data_o[47];
  assign data_o[23919] = data_o[47];
  assign data_o[23983] = data_o[47];
  assign data_o[24047] = data_o[47];
  assign data_o[24111] = data_o[47];
  assign data_o[24175] = data_o[47];
  assign data_o[24239] = data_o[47];
  assign data_o[24303] = data_o[47];
  assign data_o[24367] = data_o[47];
  assign data_o[24431] = data_o[47];
  assign data_o[24495] = data_o[47];
  assign data_o[24559] = data_o[47];
  assign data_o[24623] = data_o[47];
  assign data_o[24687] = data_o[47];
  assign data_o[24751] = data_o[47];
  assign data_o[24815] = data_o[47];
  assign data_o[24879] = data_o[47];
  assign data_o[24943] = data_o[47];
  assign data_o[25007] = data_o[47];
  assign data_o[25071] = data_o[47];
  assign data_o[25135] = data_o[47];
  assign data_o[25199] = data_o[47];
  assign data_o[25263] = data_o[47];
  assign data_o[25327] = data_o[47];
  assign data_o[25391] = data_o[47];
  assign data_o[25455] = data_o[47];
  assign data_o[25519] = data_o[47];
  assign data_o[25583] = data_o[47];
  assign data_o[25647] = data_o[47];
  assign data_o[25711] = data_o[47];
  assign data_o[25775] = data_o[47];
  assign data_o[25839] = data_o[47];
  assign data_o[25903] = data_o[47];
  assign data_o[25967] = data_o[47];
  assign data_o[26031] = data_o[47];
  assign data_o[26095] = data_o[47];
  assign data_o[26159] = data_o[47];
  assign data_o[26223] = data_o[47];
  assign data_o[26287] = data_o[47];
  assign data_o[26351] = data_o[47];
  assign data_o[26415] = data_o[47];
  assign data_o[26479] = data_o[47];
  assign data_o[26543] = data_o[47];
  assign data_o[26607] = data_o[47];
  assign data_o[26671] = data_o[47];
  assign data_o[26735] = data_o[47];
  assign data_o[26799] = data_o[47];
  assign data_o[26863] = data_o[47];
  assign data_o[26927] = data_o[47];
  assign data_o[26991] = data_o[47];
  assign data_o[27055] = data_o[47];
  assign data_o[27119] = data_o[47];
  assign data_o[27183] = data_o[47];
  assign data_o[27247] = data_o[47];
  assign data_o[27311] = data_o[47];
  assign data_o[27375] = data_o[47];
  assign data_o[27439] = data_o[47];
  assign data_o[27503] = data_o[47];
  assign data_o[27567] = data_o[47];
  assign data_o[27631] = data_o[47];
  assign data_o[27695] = data_o[47];
  assign data_o[27759] = data_o[47];
  assign data_o[27823] = data_o[47];
  assign data_o[27887] = data_o[47];
  assign data_o[27951] = data_o[47];
  assign data_o[28015] = data_o[47];
  assign data_o[28079] = data_o[47];
  assign data_o[28143] = data_o[47];
  assign data_o[28207] = data_o[47];
  assign data_o[28271] = data_o[47];
  assign data_o[28335] = data_o[47];
  assign data_o[28399] = data_o[47];
  assign data_o[28463] = data_o[47];
  assign data_o[28527] = data_o[47];
  assign data_o[28591] = data_o[47];
  assign data_o[28655] = data_o[47];
  assign data_o[28719] = data_o[47];
  assign data_o[28783] = data_o[47];
  assign data_o[28847] = data_o[47];
  assign data_o[28911] = data_o[47];
  assign data_o[28975] = data_o[47];
  assign data_o[29039] = data_o[47];
  assign data_o[29103] = data_o[47];
  assign data_o[29167] = data_o[47];
  assign data_o[29231] = data_o[47];
  assign data_o[29295] = data_o[47];
  assign data_o[29359] = data_o[47];
  assign data_o[29423] = data_o[47];
  assign data_o[29487] = data_o[47];
  assign data_o[29551] = data_o[47];
  assign data_o[29615] = data_o[47];
  assign data_o[29679] = data_o[47];
  assign data_o[29743] = data_o[47];
  assign data_o[29807] = data_o[47];
  assign data_o[29871] = data_o[47];
  assign data_o[29935] = data_o[47];
  assign data_o[29999] = data_o[47];
  assign data_o[30063] = data_o[47];
  assign data_o[30127] = data_o[47];
  assign data_o[30191] = data_o[47];
  assign data_o[30255] = data_o[47];
  assign data_o[30319] = data_o[47];
  assign data_o[30383] = data_o[47];
  assign data_o[30447] = data_o[47];
  assign data_o[30511] = data_o[47];
  assign data_o[30575] = data_o[47];
  assign data_o[30639] = data_o[47];
  assign data_o[30703] = data_o[47];
  assign data_o[30767] = data_o[47];
  assign data_o[30831] = data_o[47];
  assign data_o[30895] = data_o[47];
  assign data_o[30959] = data_o[47];
  assign data_o[31023] = data_o[47];
  assign data_o[31087] = data_o[47];
  assign data_o[31151] = data_o[47];
  assign data_o[31215] = data_o[47];
  assign data_o[31279] = data_o[47];
  assign data_o[31343] = data_o[47];
  assign data_o[31407] = data_o[47];
  assign data_o[31471] = data_o[47];
  assign data_o[31535] = data_o[47];
  assign data_o[31599] = data_o[47];
  assign data_o[31663] = data_o[47];
  assign data_o[31727] = data_o[47];
  assign data_o[31791] = data_o[47];
  assign data_o[31855] = data_o[47];
  assign data_o[31919] = data_o[47];
  assign data_o[31983] = data_o[47];
  assign data_o[110] = data_o[46];
  assign data_o[174] = data_o[46];
  assign data_o[238] = data_o[46];
  assign data_o[302] = data_o[46];
  assign data_o[366] = data_o[46];
  assign data_o[430] = data_o[46];
  assign data_o[494] = data_o[46];
  assign data_o[558] = data_o[46];
  assign data_o[622] = data_o[46];
  assign data_o[686] = data_o[46];
  assign data_o[750] = data_o[46];
  assign data_o[814] = data_o[46];
  assign data_o[878] = data_o[46];
  assign data_o[942] = data_o[46];
  assign data_o[1006] = data_o[46];
  assign data_o[1070] = data_o[46];
  assign data_o[1134] = data_o[46];
  assign data_o[1198] = data_o[46];
  assign data_o[1262] = data_o[46];
  assign data_o[1326] = data_o[46];
  assign data_o[1390] = data_o[46];
  assign data_o[1454] = data_o[46];
  assign data_o[1518] = data_o[46];
  assign data_o[1582] = data_o[46];
  assign data_o[1646] = data_o[46];
  assign data_o[1710] = data_o[46];
  assign data_o[1774] = data_o[46];
  assign data_o[1838] = data_o[46];
  assign data_o[1902] = data_o[46];
  assign data_o[1966] = data_o[46];
  assign data_o[2030] = data_o[46];
  assign data_o[2094] = data_o[46];
  assign data_o[2158] = data_o[46];
  assign data_o[2222] = data_o[46];
  assign data_o[2286] = data_o[46];
  assign data_o[2350] = data_o[46];
  assign data_o[2414] = data_o[46];
  assign data_o[2478] = data_o[46];
  assign data_o[2542] = data_o[46];
  assign data_o[2606] = data_o[46];
  assign data_o[2670] = data_o[46];
  assign data_o[2734] = data_o[46];
  assign data_o[2798] = data_o[46];
  assign data_o[2862] = data_o[46];
  assign data_o[2926] = data_o[46];
  assign data_o[2990] = data_o[46];
  assign data_o[3054] = data_o[46];
  assign data_o[3118] = data_o[46];
  assign data_o[3182] = data_o[46];
  assign data_o[3246] = data_o[46];
  assign data_o[3310] = data_o[46];
  assign data_o[3374] = data_o[46];
  assign data_o[3438] = data_o[46];
  assign data_o[3502] = data_o[46];
  assign data_o[3566] = data_o[46];
  assign data_o[3630] = data_o[46];
  assign data_o[3694] = data_o[46];
  assign data_o[3758] = data_o[46];
  assign data_o[3822] = data_o[46];
  assign data_o[3886] = data_o[46];
  assign data_o[3950] = data_o[46];
  assign data_o[4014] = data_o[46];
  assign data_o[4078] = data_o[46];
  assign data_o[4142] = data_o[46];
  assign data_o[4206] = data_o[46];
  assign data_o[4270] = data_o[46];
  assign data_o[4334] = data_o[46];
  assign data_o[4398] = data_o[46];
  assign data_o[4462] = data_o[46];
  assign data_o[4526] = data_o[46];
  assign data_o[4590] = data_o[46];
  assign data_o[4654] = data_o[46];
  assign data_o[4718] = data_o[46];
  assign data_o[4782] = data_o[46];
  assign data_o[4846] = data_o[46];
  assign data_o[4910] = data_o[46];
  assign data_o[4974] = data_o[46];
  assign data_o[5038] = data_o[46];
  assign data_o[5102] = data_o[46];
  assign data_o[5166] = data_o[46];
  assign data_o[5230] = data_o[46];
  assign data_o[5294] = data_o[46];
  assign data_o[5358] = data_o[46];
  assign data_o[5422] = data_o[46];
  assign data_o[5486] = data_o[46];
  assign data_o[5550] = data_o[46];
  assign data_o[5614] = data_o[46];
  assign data_o[5678] = data_o[46];
  assign data_o[5742] = data_o[46];
  assign data_o[5806] = data_o[46];
  assign data_o[5870] = data_o[46];
  assign data_o[5934] = data_o[46];
  assign data_o[5998] = data_o[46];
  assign data_o[6062] = data_o[46];
  assign data_o[6126] = data_o[46];
  assign data_o[6190] = data_o[46];
  assign data_o[6254] = data_o[46];
  assign data_o[6318] = data_o[46];
  assign data_o[6382] = data_o[46];
  assign data_o[6446] = data_o[46];
  assign data_o[6510] = data_o[46];
  assign data_o[6574] = data_o[46];
  assign data_o[6638] = data_o[46];
  assign data_o[6702] = data_o[46];
  assign data_o[6766] = data_o[46];
  assign data_o[6830] = data_o[46];
  assign data_o[6894] = data_o[46];
  assign data_o[6958] = data_o[46];
  assign data_o[7022] = data_o[46];
  assign data_o[7086] = data_o[46];
  assign data_o[7150] = data_o[46];
  assign data_o[7214] = data_o[46];
  assign data_o[7278] = data_o[46];
  assign data_o[7342] = data_o[46];
  assign data_o[7406] = data_o[46];
  assign data_o[7470] = data_o[46];
  assign data_o[7534] = data_o[46];
  assign data_o[7598] = data_o[46];
  assign data_o[7662] = data_o[46];
  assign data_o[7726] = data_o[46];
  assign data_o[7790] = data_o[46];
  assign data_o[7854] = data_o[46];
  assign data_o[7918] = data_o[46];
  assign data_o[7982] = data_o[46];
  assign data_o[8046] = data_o[46];
  assign data_o[8110] = data_o[46];
  assign data_o[8174] = data_o[46];
  assign data_o[8238] = data_o[46];
  assign data_o[8302] = data_o[46];
  assign data_o[8366] = data_o[46];
  assign data_o[8430] = data_o[46];
  assign data_o[8494] = data_o[46];
  assign data_o[8558] = data_o[46];
  assign data_o[8622] = data_o[46];
  assign data_o[8686] = data_o[46];
  assign data_o[8750] = data_o[46];
  assign data_o[8814] = data_o[46];
  assign data_o[8878] = data_o[46];
  assign data_o[8942] = data_o[46];
  assign data_o[9006] = data_o[46];
  assign data_o[9070] = data_o[46];
  assign data_o[9134] = data_o[46];
  assign data_o[9198] = data_o[46];
  assign data_o[9262] = data_o[46];
  assign data_o[9326] = data_o[46];
  assign data_o[9390] = data_o[46];
  assign data_o[9454] = data_o[46];
  assign data_o[9518] = data_o[46];
  assign data_o[9582] = data_o[46];
  assign data_o[9646] = data_o[46];
  assign data_o[9710] = data_o[46];
  assign data_o[9774] = data_o[46];
  assign data_o[9838] = data_o[46];
  assign data_o[9902] = data_o[46];
  assign data_o[9966] = data_o[46];
  assign data_o[10030] = data_o[46];
  assign data_o[10094] = data_o[46];
  assign data_o[10158] = data_o[46];
  assign data_o[10222] = data_o[46];
  assign data_o[10286] = data_o[46];
  assign data_o[10350] = data_o[46];
  assign data_o[10414] = data_o[46];
  assign data_o[10478] = data_o[46];
  assign data_o[10542] = data_o[46];
  assign data_o[10606] = data_o[46];
  assign data_o[10670] = data_o[46];
  assign data_o[10734] = data_o[46];
  assign data_o[10798] = data_o[46];
  assign data_o[10862] = data_o[46];
  assign data_o[10926] = data_o[46];
  assign data_o[10990] = data_o[46];
  assign data_o[11054] = data_o[46];
  assign data_o[11118] = data_o[46];
  assign data_o[11182] = data_o[46];
  assign data_o[11246] = data_o[46];
  assign data_o[11310] = data_o[46];
  assign data_o[11374] = data_o[46];
  assign data_o[11438] = data_o[46];
  assign data_o[11502] = data_o[46];
  assign data_o[11566] = data_o[46];
  assign data_o[11630] = data_o[46];
  assign data_o[11694] = data_o[46];
  assign data_o[11758] = data_o[46];
  assign data_o[11822] = data_o[46];
  assign data_o[11886] = data_o[46];
  assign data_o[11950] = data_o[46];
  assign data_o[12014] = data_o[46];
  assign data_o[12078] = data_o[46];
  assign data_o[12142] = data_o[46];
  assign data_o[12206] = data_o[46];
  assign data_o[12270] = data_o[46];
  assign data_o[12334] = data_o[46];
  assign data_o[12398] = data_o[46];
  assign data_o[12462] = data_o[46];
  assign data_o[12526] = data_o[46];
  assign data_o[12590] = data_o[46];
  assign data_o[12654] = data_o[46];
  assign data_o[12718] = data_o[46];
  assign data_o[12782] = data_o[46];
  assign data_o[12846] = data_o[46];
  assign data_o[12910] = data_o[46];
  assign data_o[12974] = data_o[46];
  assign data_o[13038] = data_o[46];
  assign data_o[13102] = data_o[46];
  assign data_o[13166] = data_o[46];
  assign data_o[13230] = data_o[46];
  assign data_o[13294] = data_o[46];
  assign data_o[13358] = data_o[46];
  assign data_o[13422] = data_o[46];
  assign data_o[13486] = data_o[46];
  assign data_o[13550] = data_o[46];
  assign data_o[13614] = data_o[46];
  assign data_o[13678] = data_o[46];
  assign data_o[13742] = data_o[46];
  assign data_o[13806] = data_o[46];
  assign data_o[13870] = data_o[46];
  assign data_o[13934] = data_o[46];
  assign data_o[13998] = data_o[46];
  assign data_o[14062] = data_o[46];
  assign data_o[14126] = data_o[46];
  assign data_o[14190] = data_o[46];
  assign data_o[14254] = data_o[46];
  assign data_o[14318] = data_o[46];
  assign data_o[14382] = data_o[46];
  assign data_o[14446] = data_o[46];
  assign data_o[14510] = data_o[46];
  assign data_o[14574] = data_o[46];
  assign data_o[14638] = data_o[46];
  assign data_o[14702] = data_o[46];
  assign data_o[14766] = data_o[46];
  assign data_o[14830] = data_o[46];
  assign data_o[14894] = data_o[46];
  assign data_o[14958] = data_o[46];
  assign data_o[15022] = data_o[46];
  assign data_o[15086] = data_o[46];
  assign data_o[15150] = data_o[46];
  assign data_o[15214] = data_o[46];
  assign data_o[15278] = data_o[46];
  assign data_o[15342] = data_o[46];
  assign data_o[15406] = data_o[46];
  assign data_o[15470] = data_o[46];
  assign data_o[15534] = data_o[46];
  assign data_o[15598] = data_o[46];
  assign data_o[15662] = data_o[46];
  assign data_o[15726] = data_o[46];
  assign data_o[15790] = data_o[46];
  assign data_o[15854] = data_o[46];
  assign data_o[15918] = data_o[46];
  assign data_o[15982] = data_o[46];
  assign data_o[16046] = data_o[46];
  assign data_o[16110] = data_o[46];
  assign data_o[16174] = data_o[46];
  assign data_o[16238] = data_o[46];
  assign data_o[16302] = data_o[46];
  assign data_o[16366] = data_o[46];
  assign data_o[16430] = data_o[46];
  assign data_o[16494] = data_o[46];
  assign data_o[16558] = data_o[46];
  assign data_o[16622] = data_o[46];
  assign data_o[16686] = data_o[46];
  assign data_o[16750] = data_o[46];
  assign data_o[16814] = data_o[46];
  assign data_o[16878] = data_o[46];
  assign data_o[16942] = data_o[46];
  assign data_o[17006] = data_o[46];
  assign data_o[17070] = data_o[46];
  assign data_o[17134] = data_o[46];
  assign data_o[17198] = data_o[46];
  assign data_o[17262] = data_o[46];
  assign data_o[17326] = data_o[46];
  assign data_o[17390] = data_o[46];
  assign data_o[17454] = data_o[46];
  assign data_o[17518] = data_o[46];
  assign data_o[17582] = data_o[46];
  assign data_o[17646] = data_o[46];
  assign data_o[17710] = data_o[46];
  assign data_o[17774] = data_o[46];
  assign data_o[17838] = data_o[46];
  assign data_o[17902] = data_o[46];
  assign data_o[17966] = data_o[46];
  assign data_o[18030] = data_o[46];
  assign data_o[18094] = data_o[46];
  assign data_o[18158] = data_o[46];
  assign data_o[18222] = data_o[46];
  assign data_o[18286] = data_o[46];
  assign data_o[18350] = data_o[46];
  assign data_o[18414] = data_o[46];
  assign data_o[18478] = data_o[46];
  assign data_o[18542] = data_o[46];
  assign data_o[18606] = data_o[46];
  assign data_o[18670] = data_o[46];
  assign data_o[18734] = data_o[46];
  assign data_o[18798] = data_o[46];
  assign data_o[18862] = data_o[46];
  assign data_o[18926] = data_o[46];
  assign data_o[18990] = data_o[46];
  assign data_o[19054] = data_o[46];
  assign data_o[19118] = data_o[46];
  assign data_o[19182] = data_o[46];
  assign data_o[19246] = data_o[46];
  assign data_o[19310] = data_o[46];
  assign data_o[19374] = data_o[46];
  assign data_o[19438] = data_o[46];
  assign data_o[19502] = data_o[46];
  assign data_o[19566] = data_o[46];
  assign data_o[19630] = data_o[46];
  assign data_o[19694] = data_o[46];
  assign data_o[19758] = data_o[46];
  assign data_o[19822] = data_o[46];
  assign data_o[19886] = data_o[46];
  assign data_o[19950] = data_o[46];
  assign data_o[20014] = data_o[46];
  assign data_o[20078] = data_o[46];
  assign data_o[20142] = data_o[46];
  assign data_o[20206] = data_o[46];
  assign data_o[20270] = data_o[46];
  assign data_o[20334] = data_o[46];
  assign data_o[20398] = data_o[46];
  assign data_o[20462] = data_o[46];
  assign data_o[20526] = data_o[46];
  assign data_o[20590] = data_o[46];
  assign data_o[20654] = data_o[46];
  assign data_o[20718] = data_o[46];
  assign data_o[20782] = data_o[46];
  assign data_o[20846] = data_o[46];
  assign data_o[20910] = data_o[46];
  assign data_o[20974] = data_o[46];
  assign data_o[21038] = data_o[46];
  assign data_o[21102] = data_o[46];
  assign data_o[21166] = data_o[46];
  assign data_o[21230] = data_o[46];
  assign data_o[21294] = data_o[46];
  assign data_o[21358] = data_o[46];
  assign data_o[21422] = data_o[46];
  assign data_o[21486] = data_o[46];
  assign data_o[21550] = data_o[46];
  assign data_o[21614] = data_o[46];
  assign data_o[21678] = data_o[46];
  assign data_o[21742] = data_o[46];
  assign data_o[21806] = data_o[46];
  assign data_o[21870] = data_o[46];
  assign data_o[21934] = data_o[46];
  assign data_o[21998] = data_o[46];
  assign data_o[22062] = data_o[46];
  assign data_o[22126] = data_o[46];
  assign data_o[22190] = data_o[46];
  assign data_o[22254] = data_o[46];
  assign data_o[22318] = data_o[46];
  assign data_o[22382] = data_o[46];
  assign data_o[22446] = data_o[46];
  assign data_o[22510] = data_o[46];
  assign data_o[22574] = data_o[46];
  assign data_o[22638] = data_o[46];
  assign data_o[22702] = data_o[46];
  assign data_o[22766] = data_o[46];
  assign data_o[22830] = data_o[46];
  assign data_o[22894] = data_o[46];
  assign data_o[22958] = data_o[46];
  assign data_o[23022] = data_o[46];
  assign data_o[23086] = data_o[46];
  assign data_o[23150] = data_o[46];
  assign data_o[23214] = data_o[46];
  assign data_o[23278] = data_o[46];
  assign data_o[23342] = data_o[46];
  assign data_o[23406] = data_o[46];
  assign data_o[23470] = data_o[46];
  assign data_o[23534] = data_o[46];
  assign data_o[23598] = data_o[46];
  assign data_o[23662] = data_o[46];
  assign data_o[23726] = data_o[46];
  assign data_o[23790] = data_o[46];
  assign data_o[23854] = data_o[46];
  assign data_o[23918] = data_o[46];
  assign data_o[23982] = data_o[46];
  assign data_o[24046] = data_o[46];
  assign data_o[24110] = data_o[46];
  assign data_o[24174] = data_o[46];
  assign data_o[24238] = data_o[46];
  assign data_o[24302] = data_o[46];
  assign data_o[24366] = data_o[46];
  assign data_o[24430] = data_o[46];
  assign data_o[24494] = data_o[46];
  assign data_o[24558] = data_o[46];
  assign data_o[24622] = data_o[46];
  assign data_o[24686] = data_o[46];
  assign data_o[24750] = data_o[46];
  assign data_o[24814] = data_o[46];
  assign data_o[24878] = data_o[46];
  assign data_o[24942] = data_o[46];
  assign data_o[25006] = data_o[46];
  assign data_o[25070] = data_o[46];
  assign data_o[25134] = data_o[46];
  assign data_o[25198] = data_o[46];
  assign data_o[25262] = data_o[46];
  assign data_o[25326] = data_o[46];
  assign data_o[25390] = data_o[46];
  assign data_o[25454] = data_o[46];
  assign data_o[25518] = data_o[46];
  assign data_o[25582] = data_o[46];
  assign data_o[25646] = data_o[46];
  assign data_o[25710] = data_o[46];
  assign data_o[25774] = data_o[46];
  assign data_o[25838] = data_o[46];
  assign data_o[25902] = data_o[46];
  assign data_o[25966] = data_o[46];
  assign data_o[26030] = data_o[46];
  assign data_o[26094] = data_o[46];
  assign data_o[26158] = data_o[46];
  assign data_o[26222] = data_o[46];
  assign data_o[26286] = data_o[46];
  assign data_o[26350] = data_o[46];
  assign data_o[26414] = data_o[46];
  assign data_o[26478] = data_o[46];
  assign data_o[26542] = data_o[46];
  assign data_o[26606] = data_o[46];
  assign data_o[26670] = data_o[46];
  assign data_o[26734] = data_o[46];
  assign data_o[26798] = data_o[46];
  assign data_o[26862] = data_o[46];
  assign data_o[26926] = data_o[46];
  assign data_o[26990] = data_o[46];
  assign data_o[27054] = data_o[46];
  assign data_o[27118] = data_o[46];
  assign data_o[27182] = data_o[46];
  assign data_o[27246] = data_o[46];
  assign data_o[27310] = data_o[46];
  assign data_o[27374] = data_o[46];
  assign data_o[27438] = data_o[46];
  assign data_o[27502] = data_o[46];
  assign data_o[27566] = data_o[46];
  assign data_o[27630] = data_o[46];
  assign data_o[27694] = data_o[46];
  assign data_o[27758] = data_o[46];
  assign data_o[27822] = data_o[46];
  assign data_o[27886] = data_o[46];
  assign data_o[27950] = data_o[46];
  assign data_o[28014] = data_o[46];
  assign data_o[28078] = data_o[46];
  assign data_o[28142] = data_o[46];
  assign data_o[28206] = data_o[46];
  assign data_o[28270] = data_o[46];
  assign data_o[28334] = data_o[46];
  assign data_o[28398] = data_o[46];
  assign data_o[28462] = data_o[46];
  assign data_o[28526] = data_o[46];
  assign data_o[28590] = data_o[46];
  assign data_o[28654] = data_o[46];
  assign data_o[28718] = data_o[46];
  assign data_o[28782] = data_o[46];
  assign data_o[28846] = data_o[46];
  assign data_o[28910] = data_o[46];
  assign data_o[28974] = data_o[46];
  assign data_o[29038] = data_o[46];
  assign data_o[29102] = data_o[46];
  assign data_o[29166] = data_o[46];
  assign data_o[29230] = data_o[46];
  assign data_o[29294] = data_o[46];
  assign data_o[29358] = data_o[46];
  assign data_o[29422] = data_o[46];
  assign data_o[29486] = data_o[46];
  assign data_o[29550] = data_o[46];
  assign data_o[29614] = data_o[46];
  assign data_o[29678] = data_o[46];
  assign data_o[29742] = data_o[46];
  assign data_o[29806] = data_o[46];
  assign data_o[29870] = data_o[46];
  assign data_o[29934] = data_o[46];
  assign data_o[29998] = data_o[46];
  assign data_o[30062] = data_o[46];
  assign data_o[30126] = data_o[46];
  assign data_o[30190] = data_o[46];
  assign data_o[30254] = data_o[46];
  assign data_o[30318] = data_o[46];
  assign data_o[30382] = data_o[46];
  assign data_o[30446] = data_o[46];
  assign data_o[30510] = data_o[46];
  assign data_o[30574] = data_o[46];
  assign data_o[30638] = data_o[46];
  assign data_o[30702] = data_o[46];
  assign data_o[30766] = data_o[46];
  assign data_o[30830] = data_o[46];
  assign data_o[30894] = data_o[46];
  assign data_o[30958] = data_o[46];
  assign data_o[31022] = data_o[46];
  assign data_o[31086] = data_o[46];
  assign data_o[31150] = data_o[46];
  assign data_o[31214] = data_o[46];
  assign data_o[31278] = data_o[46];
  assign data_o[31342] = data_o[46];
  assign data_o[31406] = data_o[46];
  assign data_o[31470] = data_o[46];
  assign data_o[31534] = data_o[46];
  assign data_o[31598] = data_o[46];
  assign data_o[31662] = data_o[46];
  assign data_o[31726] = data_o[46];
  assign data_o[31790] = data_o[46];
  assign data_o[31854] = data_o[46];
  assign data_o[31918] = data_o[46];
  assign data_o[31982] = data_o[46];
  assign data_o[109] = data_o[45];
  assign data_o[173] = data_o[45];
  assign data_o[237] = data_o[45];
  assign data_o[301] = data_o[45];
  assign data_o[365] = data_o[45];
  assign data_o[429] = data_o[45];
  assign data_o[493] = data_o[45];
  assign data_o[557] = data_o[45];
  assign data_o[621] = data_o[45];
  assign data_o[685] = data_o[45];
  assign data_o[749] = data_o[45];
  assign data_o[813] = data_o[45];
  assign data_o[877] = data_o[45];
  assign data_o[941] = data_o[45];
  assign data_o[1005] = data_o[45];
  assign data_o[1069] = data_o[45];
  assign data_o[1133] = data_o[45];
  assign data_o[1197] = data_o[45];
  assign data_o[1261] = data_o[45];
  assign data_o[1325] = data_o[45];
  assign data_o[1389] = data_o[45];
  assign data_o[1453] = data_o[45];
  assign data_o[1517] = data_o[45];
  assign data_o[1581] = data_o[45];
  assign data_o[1645] = data_o[45];
  assign data_o[1709] = data_o[45];
  assign data_o[1773] = data_o[45];
  assign data_o[1837] = data_o[45];
  assign data_o[1901] = data_o[45];
  assign data_o[1965] = data_o[45];
  assign data_o[2029] = data_o[45];
  assign data_o[2093] = data_o[45];
  assign data_o[2157] = data_o[45];
  assign data_o[2221] = data_o[45];
  assign data_o[2285] = data_o[45];
  assign data_o[2349] = data_o[45];
  assign data_o[2413] = data_o[45];
  assign data_o[2477] = data_o[45];
  assign data_o[2541] = data_o[45];
  assign data_o[2605] = data_o[45];
  assign data_o[2669] = data_o[45];
  assign data_o[2733] = data_o[45];
  assign data_o[2797] = data_o[45];
  assign data_o[2861] = data_o[45];
  assign data_o[2925] = data_o[45];
  assign data_o[2989] = data_o[45];
  assign data_o[3053] = data_o[45];
  assign data_o[3117] = data_o[45];
  assign data_o[3181] = data_o[45];
  assign data_o[3245] = data_o[45];
  assign data_o[3309] = data_o[45];
  assign data_o[3373] = data_o[45];
  assign data_o[3437] = data_o[45];
  assign data_o[3501] = data_o[45];
  assign data_o[3565] = data_o[45];
  assign data_o[3629] = data_o[45];
  assign data_o[3693] = data_o[45];
  assign data_o[3757] = data_o[45];
  assign data_o[3821] = data_o[45];
  assign data_o[3885] = data_o[45];
  assign data_o[3949] = data_o[45];
  assign data_o[4013] = data_o[45];
  assign data_o[4077] = data_o[45];
  assign data_o[4141] = data_o[45];
  assign data_o[4205] = data_o[45];
  assign data_o[4269] = data_o[45];
  assign data_o[4333] = data_o[45];
  assign data_o[4397] = data_o[45];
  assign data_o[4461] = data_o[45];
  assign data_o[4525] = data_o[45];
  assign data_o[4589] = data_o[45];
  assign data_o[4653] = data_o[45];
  assign data_o[4717] = data_o[45];
  assign data_o[4781] = data_o[45];
  assign data_o[4845] = data_o[45];
  assign data_o[4909] = data_o[45];
  assign data_o[4973] = data_o[45];
  assign data_o[5037] = data_o[45];
  assign data_o[5101] = data_o[45];
  assign data_o[5165] = data_o[45];
  assign data_o[5229] = data_o[45];
  assign data_o[5293] = data_o[45];
  assign data_o[5357] = data_o[45];
  assign data_o[5421] = data_o[45];
  assign data_o[5485] = data_o[45];
  assign data_o[5549] = data_o[45];
  assign data_o[5613] = data_o[45];
  assign data_o[5677] = data_o[45];
  assign data_o[5741] = data_o[45];
  assign data_o[5805] = data_o[45];
  assign data_o[5869] = data_o[45];
  assign data_o[5933] = data_o[45];
  assign data_o[5997] = data_o[45];
  assign data_o[6061] = data_o[45];
  assign data_o[6125] = data_o[45];
  assign data_o[6189] = data_o[45];
  assign data_o[6253] = data_o[45];
  assign data_o[6317] = data_o[45];
  assign data_o[6381] = data_o[45];
  assign data_o[6445] = data_o[45];
  assign data_o[6509] = data_o[45];
  assign data_o[6573] = data_o[45];
  assign data_o[6637] = data_o[45];
  assign data_o[6701] = data_o[45];
  assign data_o[6765] = data_o[45];
  assign data_o[6829] = data_o[45];
  assign data_o[6893] = data_o[45];
  assign data_o[6957] = data_o[45];
  assign data_o[7021] = data_o[45];
  assign data_o[7085] = data_o[45];
  assign data_o[7149] = data_o[45];
  assign data_o[7213] = data_o[45];
  assign data_o[7277] = data_o[45];
  assign data_o[7341] = data_o[45];
  assign data_o[7405] = data_o[45];
  assign data_o[7469] = data_o[45];
  assign data_o[7533] = data_o[45];
  assign data_o[7597] = data_o[45];
  assign data_o[7661] = data_o[45];
  assign data_o[7725] = data_o[45];
  assign data_o[7789] = data_o[45];
  assign data_o[7853] = data_o[45];
  assign data_o[7917] = data_o[45];
  assign data_o[7981] = data_o[45];
  assign data_o[8045] = data_o[45];
  assign data_o[8109] = data_o[45];
  assign data_o[8173] = data_o[45];
  assign data_o[8237] = data_o[45];
  assign data_o[8301] = data_o[45];
  assign data_o[8365] = data_o[45];
  assign data_o[8429] = data_o[45];
  assign data_o[8493] = data_o[45];
  assign data_o[8557] = data_o[45];
  assign data_o[8621] = data_o[45];
  assign data_o[8685] = data_o[45];
  assign data_o[8749] = data_o[45];
  assign data_o[8813] = data_o[45];
  assign data_o[8877] = data_o[45];
  assign data_o[8941] = data_o[45];
  assign data_o[9005] = data_o[45];
  assign data_o[9069] = data_o[45];
  assign data_o[9133] = data_o[45];
  assign data_o[9197] = data_o[45];
  assign data_o[9261] = data_o[45];
  assign data_o[9325] = data_o[45];
  assign data_o[9389] = data_o[45];
  assign data_o[9453] = data_o[45];
  assign data_o[9517] = data_o[45];
  assign data_o[9581] = data_o[45];
  assign data_o[9645] = data_o[45];
  assign data_o[9709] = data_o[45];
  assign data_o[9773] = data_o[45];
  assign data_o[9837] = data_o[45];
  assign data_o[9901] = data_o[45];
  assign data_o[9965] = data_o[45];
  assign data_o[10029] = data_o[45];
  assign data_o[10093] = data_o[45];
  assign data_o[10157] = data_o[45];
  assign data_o[10221] = data_o[45];
  assign data_o[10285] = data_o[45];
  assign data_o[10349] = data_o[45];
  assign data_o[10413] = data_o[45];
  assign data_o[10477] = data_o[45];
  assign data_o[10541] = data_o[45];
  assign data_o[10605] = data_o[45];
  assign data_o[10669] = data_o[45];
  assign data_o[10733] = data_o[45];
  assign data_o[10797] = data_o[45];
  assign data_o[10861] = data_o[45];
  assign data_o[10925] = data_o[45];
  assign data_o[10989] = data_o[45];
  assign data_o[11053] = data_o[45];
  assign data_o[11117] = data_o[45];
  assign data_o[11181] = data_o[45];
  assign data_o[11245] = data_o[45];
  assign data_o[11309] = data_o[45];
  assign data_o[11373] = data_o[45];
  assign data_o[11437] = data_o[45];
  assign data_o[11501] = data_o[45];
  assign data_o[11565] = data_o[45];
  assign data_o[11629] = data_o[45];
  assign data_o[11693] = data_o[45];
  assign data_o[11757] = data_o[45];
  assign data_o[11821] = data_o[45];
  assign data_o[11885] = data_o[45];
  assign data_o[11949] = data_o[45];
  assign data_o[12013] = data_o[45];
  assign data_o[12077] = data_o[45];
  assign data_o[12141] = data_o[45];
  assign data_o[12205] = data_o[45];
  assign data_o[12269] = data_o[45];
  assign data_o[12333] = data_o[45];
  assign data_o[12397] = data_o[45];
  assign data_o[12461] = data_o[45];
  assign data_o[12525] = data_o[45];
  assign data_o[12589] = data_o[45];
  assign data_o[12653] = data_o[45];
  assign data_o[12717] = data_o[45];
  assign data_o[12781] = data_o[45];
  assign data_o[12845] = data_o[45];
  assign data_o[12909] = data_o[45];
  assign data_o[12973] = data_o[45];
  assign data_o[13037] = data_o[45];
  assign data_o[13101] = data_o[45];
  assign data_o[13165] = data_o[45];
  assign data_o[13229] = data_o[45];
  assign data_o[13293] = data_o[45];
  assign data_o[13357] = data_o[45];
  assign data_o[13421] = data_o[45];
  assign data_o[13485] = data_o[45];
  assign data_o[13549] = data_o[45];
  assign data_o[13613] = data_o[45];
  assign data_o[13677] = data_o[45];
  assign data_o[13741] = data_o[45];
  assign data_o[13805] = data_o[45];
  assign data_o[13869] = data_o[45];
  assign data_o[13933] = data_o[45];
  assign data_o[13997] = data_o[45];
  assign data_o[14061] = data_o[45];
  assign data_o[14125] = data_o[45];
  assign data_o[14189] = data_o[45];
  assign data_o[14253] = data_o[45];
  assign data_o[14317] = data_o[45];
  assign data_o[14381] = data_o[45];
  assign data_o[14445] = data_o[45];
  assign data_o[14509] = data_o[45];
  assign data_o[14573] = data_o[45];
  assign data_o[14637] = data_o[45];
  assign data_o[14701] = data_o[45];
  assign data_o[14765] = data_o[45];
  assign data_o[14829] = data_o[45];
  assign data_o[14893] = data_o[45];
  assign data_o[14957] = data_o[45];
  assign data_o[15021] = data_o[45];
  assign data_o[15085] = data_o[45];
  assign data_o[15149] = data_o[45];
  assign data_o[15213] = data_o[45];
  assign data_o[15277] = data_o[45];
  assign data_o[15341] = data_o[45];
  assign data_o[15405] = data_o[45];
  assign data_o[15469] = data_o[45];
  assign data_o[15533] = data_o[45];
  assign data_o[15597] = data_o[45];
  assign data_o[15661] = data_o[45];
  assign data_o[15725] = data_o[45];
  assign data_o[15789] = data_o[45];
  assign data_o[15853] = data_o[45];
  assign data_o[15917] = data_o[45];
  assign data_o[15981] = data_o[45];
  assign data_o[16045] = data_o[45];
  assign data_o[16109] = data_o[45];
  assign data_o[16173] = data_o[45];
  assign data_o[16237] = data_o[45];
  assign data_o[16301] = data_o[45];
  assign data_o[16365] = data_o[45];
  assign data_o[16429] = data_o[45];
  assign data_o[16493] = data_o[45];
  assign data_o[16557] = data_o[45];
  assign data_o[16621] = data_o[45];
  assign data_o[16685] = data_o[45];
  assign data_o[16749] = data_o[45];
  assign data_o[16813] = data_o[45];
  assign data_o[16877] = data_o[45];
  assign data_o[16941] = data_o[45];
  assign data_o[17005] = data_o[45];
  assign data_o[17069] = data_o[45];
  assign data_o[17133] = data_o[45];
  assign data_o[17197] = data_o[45];
  assign data_o[17261] = data_o[45];
  assign data_o[17325] = data_o[45];
  assign data_o[17389] = data_o[45];
  assign data_o[17453] = data_o[45];
  assign data_o[17517] = data_o[45];
  assign data_o[17581] = data_o[45];
  assign data_o[17645] = data_o[45];
  assign data_o[17709] = data_o[45];
  assign data_o[17773] = data_o[45];
  assign data_o[17837] = data_o[45];
  assign data_o[17901] = data_o[45];
  assign data_o[17965] = data_o[45];
  assign data_o[18029] = data_o[45];
  assign data_o[18093] = data_o[45];
  assign data_o[18157] = data_o[45];
  assign data_o[18221] = data_o[45];
  assign data_o[18285] = data_o[45];
  assign data_o[18349] = data_o[45];
  assign data_o[18413] = data_o[45];
  assign data_o[18477] = data_o[45];
  assign data_o[18541] = data_o[45];
  assign data_o[18605] = data_o[45];
  assign data_o[18669] = data_o[45];
  assign data_o[18733] = data_o[45];
  assign data_o[18797] = data_o[45];
  assign data_o[18861] = data_o[45];
  assign data_o[18925] = data_o[45];
  assign data_o[18989] = data_o[45];
  assign data_o[19053] = data_o[45];
  assign data_o[19117] = data_o[45];
  assign data_o[19181] = data_o[45];
  assign data_o[19245] = data_o[45];
  assign data_o[19309] = data_o[45];
  assign data_o[19373] = data_o[45];
  assign data_o[19437] = data_o[45];
  assign data_o[19501] = data_o[45];
  assign data_o[19565] = data_o[45];
  assign data_o[19629] = data_o[45];
  assign data_o[19693] = data_o[45];
  assign data_o[19757] = data_o[45];
  assign data_o[19821] = data_o[45];
  assign data_o[19885] = data_o[45];
  assign data_o[19949] = data_o[45];
  assign data_o[20013] = data_o[45];
  assign data_o[20077] = data_o[45];
  assign data_o[20141] = data_o[45];
  assign data_o[20205] = data_o[45];
  assign data_o[20269] = data_o[45];
  assign data_o[20333] = data_o[45];
  assign data_o[20397] = data_o[45];
  assign data_o[20461] = data_o[45];
  assign data_o[20525] = data_o[45];
  assign data_o[20589] = data_o[45];
  assign data_o[20653] = data_o[45];
  assign data_o[20717] = data_o[45];
  assign data_o[20781] = data_o[45];
  assign data_o[20845] = data_o[45];
  assign data_o[20909] = data_o[45];
  assign data_o[20973] = data_o[45];
  assign data_o[21037] = data_o[45];
  assign data_o[21101] = data_o[45];
  assign data_o[21165] = data_o[45];
  assign data_o[21229] = data_o[45];
  assign data_o[21293] = data_o[45];
  assign data_o[21357] = data_o[45];
  assign data_o[21421] = data_o[45];
  assign data_o[21485] = data_o[45];
  assign data_o[21549] = data_o[45];
  assign data_o[21613] = data_o[45];
  assign data_o[21677] = data_o[45];
  assign data_o[21741] = data_o[45];
  assign data_o[21805] = data_o[45];
  assign data_o[21869] = data_o[45];
  assign data_o[21933] = data_o[45];
  assign data_o[21997] = data_o[45];
  assign data_o[22061] = data_o[45];
  assign data_o[22125] = data_o[45];
  assign data_o[22189] = data_o[45];
  assign data_o[22253] = data_o[45];
  assign data_o[22317] = data_o[45];
  assign data_o[22381] = data_o[45];
  assign data_o[22445] = data_o[45];
  assign data_o[22509] = data_o[45];
  assign data_o[22573] = data_o[45];
  assign data_o[22637] = data_o[45];
  assign data_o[22701] = data_o[45];
  assign data_o[22765] = data_o[45];
  assign data_o[22829] = data_o[45];
  assign data_o[22893] = data_o[45];
  assign data_o[22957] = data_o[45];
  assign data_o[23021] = data_o[45];
  assign data_o[23085] = data_o[45];
  assign data_o[23149] = data_o[45];
  assign data_o[23213] = data_o[45];
  assign data_o[23277] = data_o[45];
  assign data_o[23341] = data_o[45];
  assign data_o[23405] = data_o[45];
  assign data_o[23469] = data_o[45];
  assign data_o[23533] = data_o[45];
  assign data_o[23597] = data_o[45];
  assign data_o[23661] = data_o[45];
  assign data_o[23725] = data_o[45];
  assign data_o[23789] = data_o[45];
  assign data_o[23853] = data_o[45];
  assign data_o[23917] = data_o[45];
  assign data_o[23981] = data_o[45];
  assign data_o[24045] = data_o[45];
  assign data_o[24109] = data_o[45];
  assign data_o[24173] = data_o[45];
  assign data_o[24237] = data_o[45];
  assign data_o[24301] = data_o[45];
  assign data_o[24365] = data_o[45];
  assign data_o[24429] = data_o[45];
  assign data_o[24493] = data_o[45];
  assign data_o[24557] = data_o[45];
  assign data_o[24621] = data_o[45];
  assign data_o[24685] = data_o[45];
  assign data_o[24749] = data_o[45];
  assign data_o[24813] = data_o[45];
  assign data_o[24877] = data_o[45];
  assign data_o[24941] = data_o[45];
  assign data_o[25005] = data_o[45];
  assign data_o[25069] = data_o[45];
  assign data_o[25133] = data_o[45];
  assign data_o[25197] = data_o[45];
  assign data_o[25261] = data_o[45];
  assign data_o[25325] = data_o[45];
  assign data_o[25389] = data_o[45];
  assign data_o[25453] = data_o[45];
  assign data_o[25517] = data_o[45];
  assign data_o[25581] = data_o[45];
  assign data_o[25645] = data_o[45];
  assign data_o[25709] = data_o[45];
  assign data_o[25773] = data_o[45];
  assign data_o[25837] = data_o[45];
  assign data_o[25901] = data_o[45];
  assign data_o[25965] = data_o[45];
  assign data_o[26029] = data_o[45];
  assign data_o[26093] = data_o[45];
  assign data_o[26157] = data_o[45];
  assign data_o[26221] = data_o[45];
  assign data_o[26285] = data_o[45];
  assign data_o[26349] = data_o[45];
  assign data_o[26413] = data_o[45];
  assign data_o[26477] = data_o[45];
  assign data_o[26541] = data_o[45];
  assign data_o[26605] = data_o[45];
  assign data_o[26669] = data_o[45];
  assign data_o[26733] = data_o[45];
  assign data_o[26797] = data_o[45];
  assign data_o[26861] = data_o[45];
  assign data_o[26925] = data_o[45];
  assign data_o[26989] = data_o[45];
  assign data_o[27053] = data_o[45];
  assign data_o[27117] = data_o[45];
  assign data_o[27181] = data_o[45];
  assign data_o[27245] = data_o[45];
  assign data_o[27309] = data_o[45];
  assign data_o[27373] = data_o[45];
  assign data_o[27437] = data_o[45];
  assign data_o[27501] = data_o[45];
  assign data_o[27565] = data_o[45];
  assign data_o[27629] = data_o[45];
  assign data_o[27693] = data_o[45];
  assign data_o[27757] = data_o[45];
  assign data_o[27821] = data_o[45];
  assign data_o[27885] = data_o[45];
  assign data_o[27949] = data_o[45];
  assign data_o[28013] = data_o[45];
  assign data_o[28077] = data_o[45];
  assign data_o[28141] = data_o[45];
  assign data_o[28205] = data_o[45];
  assign data_o[28269] = data_o[45];
  assign data_o[28333] = data_o[45];
  assign data_o[28397] = data_o[45];
  assign data_o[28461] = data_o[45];
  assign data_o[28525] = data_o[45];
  assign data_o[28589] = data_o[45];
  assign data_o[28653] = data_o[45];
  assign data_o[28717] = data_o[45];
  assign data_o[28781] = data_o[45];
  assign data_o[28845] = data_o[45];
  assign data_o[28909] = data_o[45];
  assign data_o[28973] = data_o[45];
  assign data_o[29037] = data_o[45];
  assign data_o[29101] = data_o[45];
  assign data_o[29165] = data_o[45];
  assign data_o[29229] = data_o[45];
  assign data_o[29293] = data_o[45];
  assign data_o[29357] = data_o[45];
  assign data_o[29421] = data_o[45];
  assign data_o[29485] = data_o[45];
  assign data_o[29549] = data_o[45];
  assign data_o[29613] = data_o[45];
  assign data_o[29677] = data_o[45];
  assign data_o[29741] = data_o[45];
  assign data_o[29805] = data_o[45];
  assign data_o[29869] = data_o[45];
  assign data_o[29933] = data_o[45];
  assign data_o[29997] = data_o[45];
  assign data_o[30061] = data_o[45];
  assign data_o[30125] = data_o[45];
  assign data_o[30189] = data_o[45];
  assign data_o[30253] = data_o[45];
  assign data_o[30317] = data_o[45];
  assign data_o[30381] = data_o[45];
  assign data_o[30445] = data_o[45];
  assign data_o[30509] = data_o[45];
  assign data_o[30573] = data_o[45];
  assign data_o[30637] = data_o[45];
  assign data_o[30701] = data_o[45];
  assign data_o[30765] = data_o[45];
  assign data_o[30829] = data_o[45];
  assign data_o[30893] = data_o[45];
  assign data_o[30957] = data_o[45];
  assign data_o[31021] = data_o[45];
  assign data_o[31085] = data_o[45];
  assign data_o[31149] = data_o[45];
  assign data_o[31213] = data_o[45];
  assign data_o[31277] = data_o[45];
  assign data_o[31341] = data_o[45];
  assign data_o[31405] = data_o[45];
  assign data_o[31469] = data_o[45];
  assign data_o[31533] = data_o[45];
  assign data_o[31597] = data_o[45];
  assign data_o[31661] = data_o[45];
  assign data_o[31725] = data_o[45];
  assign data_o[31789] = data_o[45];
  assign data_o[31853] = data_o[45];
  assign data_o[31917] = data_o[45];
  assign data_o[31981] = data_o[45];
  assign data_o[108] = data_o[44];
  assign data_o[172] = data_o[44];
  assign data_o[236] = data_o[44];
  assign data_o[300] = data_o[44];
  assign data_o[364] = data_o[44];
  assign data_o[428] = data_o[44];
  assign data_o[492] = data_o[44];
  assign data_o[556] = data_o[44];
  assign data_o[620] = data_o[44];
  assign data_o[684] = data_o[44];
  assign data_o[748] = data_o[44];
  assign data_o[812] = data_o[44];
  assign data_o[876] = data_o[44];
  assign data_o[940] = data_o[44];
  assign data_o[1004] = data_o[44];
  assign data_o[1068] = data_o[44];
  assign data_o[1132] = data_o[44];
  assign data_o[1196] = data_o[44];
  assign data_o[1260] = data_o[44];
  assign data_o[1324] = data_o[44];
  assign data_o[1388] = data_o[44];
  assign data_o[1452] = data_o[44];
  assign data_o[1516] = data_o[44];
  assign data_o[1580] = data_o[44];
  assign data_o[1644] = data_o[44];
  assign data_o[1708] = data_o[44];
  assign data_o[1772] = data_o[44];
  assign data_o[1836] = data_o[44];
  assign data_o[1900] = data_o[44];
  assign data_o[1964] = data_o[44];
  assign data_o[2028] = data_o[44];
  assign data_o[2092] = data_o[44];
  assign data_o[2156] = data_o[44];
  assign data_o[2220] = data_o[44];
  assign data_o[2284] = data_o[44];
  assign data_o[2348] = data_o[44];
  assign data_o[2412] = data_o[44];
  assign data_o[2476] = data_o[44];
  assign data_o[2540] = data_o[44];
  assign data_o[2604] = data_o[44];
  assign data_o[2668] = data_o[44];
  assign data_o[2732] = data_o[44];
  assign data_o[2796] = data_o[44];
  assign data_o[2860] = data_o[44];
  assign data_o[2924] = data_o[44];
  assign data_o[2988] = data_o[44];
  assign data_o[3052] = data_o[44];
  assign data_o[3116] = data_o[44];
  assign data_o[3180] = data_o[44];
  assign data_o[3244] = data_o[44];
  assign data_o[3308] = data_o[44];
  assign data_o[3372] = data_o[44];
  assign data_o[3436] = data_o[44];
  assign data_o[3500] = data_o[44];
  assign data_o[3564] = data_o[44];
  assign data_o[3628] = data_o[44];
  assign data_o[3692] = data_o[44];
  assign data_o[3756] = data_o[44];
  assign data_o[3820] = data_o[44];
  assign data_o[3884] = data_o[44];
  assign data_o[3948] = data_o[44];
  assign data_o[4012] = data_o[44];
  assign data_o[4076] = data_o[44];
  assign data_o[4140] = data_o[44];
  assign data_o[4204] = data_o[44];
  assign data_o[4268] = data_o[44];
  assign data_o[4332] = data_o[44];
  assign data_o[4396] = data_o[44];
  assign data_o[4460] = data_o[44];
  assign data_o[4524] = data_o[44];
  assign data_o[4588] = data_o[44];
  assign data_o[4652] = data_o[44];
  assign data_o[4716] = data_o[44];
  assign data_o[4780] = data_o[44];
  assign data_o[4844] = data_o[44];
  assign data_o[4908] = data_o[44];
  assign data_o[4972] = data_o[44];
  assign data_o[5036] = data_o[44];
  assign data_o[5100] = data_o[44];
  assign data_o[5164] = data_o[44];
  assign data_o[5228] = data_o[44];
  assign data_o[5292] = data_o[44];
  assign data_o[5356] = data_o[44];
  assign data_o[5420] = data_o[44];
  assign data_o[5484] = data_o[44];
  assign data_o[5548] = data_o[44];
  assign data_o[5612] = data_o[44];
  assign data_o[5676] = data_o[44];
  assign data_o[5740] = data_o[44];
  assign data_o[5804] = data_o[44];
  assign data_o[5868] = data_o[44];
  assign data_o[5932] = data_o[44];
  assign data_o[5996] = data_o[44];
  assign data_o[6060] = data_o[44];
  assign data_o[6124] = data_o[44];
  assign data_o[6188] = data_o[44];
  assign data_o[6252] = data_o[44];
  assign data_o[6316] = data_o[44];
  assign data_o[6380] = data_o[44];
  assign data_o[6444] = data_o[44];
  assign data_o[6508] = data_o[44];
  assign data_o[6572] = data_o[44];
  assign data_o[6636] = data_o[44];
  assign data_o[6700] = data_o[44];
  assign data_o[6764] = data_o[44];
  assign data_o[6828] = data_o[44];
  assign data_o[6892] = data_o[44];
  assign data_o[6956] = data_o[44];
  assign data_o[7020] = data_o[44];
  assign data_o[7084] = data_o[44];
  assign data_o[7148] = data_o[44];
  assign data_o[7212] = data_o[44];
  assign data_o[7276] = data_o[44];
  assign data_o[7340] = data_o[44];
  assign data_o[7404] = data_o[44];
  assign data_o[7468] = data_o[44];
  assign data_o[7532] = data_o[44];
  assign data_o[7596] = data_o[44];
  assign data_o[7660] = data_o[44];
  assign data_o[7724] = data_o[44];
  assign data_o[7788] = data_o[44];
  assign data_o[7852] = data_o[44];
  assign data_o[7916] = data_o[44];
  assign data_o[7980] = data_o[44];
  assign data_o[8044] = data_o[44];
  assign data_o[8108] = data_o[44];
  assign data_o[8172] = data_o[44];
  assign data_o[8236] = data_o[44];
  assign data_o[8300] = data_o[44];
  assign data_o[8364] = data_o[44];
  assign data_o[8428] = data_o[44];
  assign data_o[8492] = data_o[44];
  assign data_o[8556] = data_o[44];
  assign data_o[8620] = data_o[44];
  assign data_o[8684] = data_o[44];
  assign data_o[8748] = data_o[44];
  assign data_o[8812] = data_o[44];
  assign data_o[8876] = data_o[44];
  assign data_o[8940] = data_o[44];
  assign data_o[9004] = data_o[44];
  assign data_o[9068] = data_o[44];
  assign data_o[9132] = data_o[44];
  assign data_o[9196] = data_o[44];
  assign data_o[9260] = data_o[44];
  assign data_o[9324] = data_o[44];
  assign data_o[9388] = data_o[44];
  assign data_o[9452] = data_o[44];
  assign data_o[9516] = data_o[44];
  assign data_o[9580] = data_o[44];
  assign data_o[9644] = data_o[44];
  assign data_o[9708] = data_o[44];
  assign data_o[9772] = data_o[44];
  assign data_o[9836] = data_o[44];
  assign data_o[9900] = data_o[44];
  assign data_o[9964] = data_o[44];
  assign data_o[10028] = data_o[44];
  assign data_o[10092] = data_o[44];
  assign data_o[10156] = data_o[44];
  assign data_o[10220] = data_o[44];
  assign data_o[10284] = data_o[44];
  assign data_o[10348] = data_o[44];
  assign data_o[10412] = data_o[44];
  assign data_o[10476] = data_o[44];
  assign data_o[10540] = data_o[44];
  assign data_o[10604] = data_o[44];
  assign data_o[10668] = data_o[44];
  assign data_o[10732] = data_o[44];
  assign data_o[10796] = data_o[44];
  assign data_o[10860] = data_o[44];
  assign data_o[10924] = data_o[44];
  assign data_o[10988] = data_o[44];
  assign data_o[11052] = data_o[44];
  assign data_o[11116] = data_o[44];
  assign data_o[11180] = data_o[44];
  assign data_o[11244] = data_o[44];
  assign data_o[11308] = data_o[44];
  assign data_o[11372] = data_o[44];
  assign data_o[11436] = data_o[44];
  assign data_o[11500] = data_o[44];
  assign data_o[11564] = data_o[44];
  assign data_o[11628] = data_o[44];
  assign data_o[11692] = data_o[44];
  assign data_o[11756] = data_o[44];
  assign data_o[11820] = data_o[44];
  assign data_o[11884] = data_o[44];
  assign data_o[11948] = data_o[44];
  assign data_o[12012] = data_o[44];
  assign data_o[12076] = data_o[44];
  assign data_o[12140] = data_o[44];
  assign data_o[12204] = data_o[44];
  assign data_o[12268] = data_o[44];
  assign data_o[12332] = data_o[44];
  assign data_o[12396] = data_o[44];
  assign data_o[12460] = data_o[44];
  assign data_o[12524] = data_o[44];
  assign data_o[12588] = data_o[44];
  assign data_o[12652] = data_o[44];
  assign data_o[12716] = data_o[44];
  assign data_o[12780] = data_o[44];
  assign data_o[12844] = data_o[44];
  assign data_o[12908] = data_o[44];
  assign data_o[12972] = data_o[44];
  assign data_o[13036] = data_o[44];
  assign data_o[13100] = data_o[44];
  assign data_o[13164] = data_o[44];
  assign data_o[13228] = data_o[44];
  assign data_o[13292] = data_o[44];
  assign data_o[13356] = data_o[44];
  assign data_o[13420] = data_o[44];
  assign data_o[13484] = data_o[44];
  assign data_o[13548] = data_o[44];
  assign data_o[13612] = data_o[44];
  assign data_o[13676] = data_o[44];
  assign data_o[13740] = data_o[44];
  assign data_o[13804] = data_o[44];
  assign data_o[13868] = data_o[44];
  assign data_o[13932] = data_o[44];
  assign data_o[13996] = data_o[44];
  assign data_o[14060] = data_o[44];
  assign data_o[14124] = data_o[44];
  assign data_o[14188] = data_o[44];
  assign data_o[14252] = data_o[44];
  assign data_o[14316] = data_o[44];
  assign data_o[14380] = data_o[44];
  assign data_o[14444] = data_o[44];
  assign data_o[14508] = data_o[44];
  assign data_o[14572] = data_o[44];
  assign data_o[14636] = data_o[44];
  assign data_o[14700] = data_o[44];
  assign data_o[14764] = data_o[44];
  assign data_o[14828] = data_o[44];
  assign data_o[14892] = data_o[44];
  assign data_o[14956] = data_o[44];
  assign data_o[15020] = data_o[44];
  assign data_o[15084] = data_o[44];
  assign data_o[15148] = data_o[44];
  assign data_o[15212] = data_o[44];
  assign data_o[15276] = data_o[44];
  assign data_o[15340] = data_o[44];
  assign data_o[15404] = data_o[44];
  assign data_o[15468] = data_o[44];
  assign data_o[15532] = data_o[44];
  assign data_o[15596] = data_o[44];
  assign data_o[15660] = data_o[44];
  assign data_o[15724] = data_o[44];
  assign data_o[15788] = data_o[44];
  assign data_o[15852] = data_o[44];
  assign data_o[15916] = data_o[44];
  assign data_o[15980] = data_o[44];
  assign data_o[16044] = data_o[44];
  assign data_o[16108] = data_o[44];
  assign data_o[16172] = data_o[44];
  assign data_o[16236] = data_o[44];
  assign data_o[16300] = data_o[44];
  assign data_o[16364] = data_o[44];
  assign data_o[16428] = data_o[44];
  assign data_o[16492] = data_o[44];
  assign data_o[16556] = data_o[44];
  assign data_o[16620] = data_o[44];
  assign data_o[16684] = data_o[44];
  assign data_o[16748] = data_o[44];
  assign data_o[16812] = data_o[44];
  assign data_o[16876] = data_o[44];
  assign data_o[16940] = data_o[44];
  assign data_o[17004] = data_o[44];
  assign data_o[17068] = data_o[44];
  assign data_o[17132] = data_o[44];
  assign data_o[17196] = data_o[44];
  assign data_o[17260] = data_o[44];
  assign data_o[17324] = data_o[44];
  assign data_o[17388] = data_o[44];
  assign data_o[17452] = data_o[44];
  assign data_o[17516] = data_o[44];
  assign data_o[17580] = data_o[44];
  assign data_o[17644] = data_o[44];
  assign data_o[17708] = data_o[44];
  assign data_o[17772] = data_o[44];
  assign data_o[17836] = data_o[44];
  assign data_o[17900] = data_o[44];
  assign data_o[17964] = data_o[44];
  assign data_o[18028] = data_o[44];
  assign data_o[18092] = data_o[44];
  assign data_o[18156] = data_o[44];
  assign data_o[18220] = data_o[44];
  assign data_o[18284] = data_o[44];
  assign data_o[18348] = data_o[44];
  assign data_o[18412] = data_o[44];
  assign data_o[18476] = data_o[44];
  assign data_o[18540] = data_o[44];
  assign data_o[18604] = data_o[44];
  assign data_o[18668] = data_o[44];
  assign data_o[18732] = data_o[44];
  assign data_o[18796] = data_o[44];
  assign data_o[18860] = data_o[44];
  assign data_o[18924] = data_o[44];
  assign data_o[18988] = data_o[44];
  assign data_o[19052] = data_o[44];
  assign data_o[19116] = data_o[44];
  assign data_o[19180] = data_o[44];
  assign data_o[19244] = data_o[44];
  assign data_o[19308] = data_o[44];
  assign data_o[19372] = data_o[44];
  assign data_o[19436] = data_o[44];
  assign data_o[19500] = data_o[44];
  assign data_o[19564] = data_o[44];
  assign data_o[19628] = data_o[44];
  assign data_o[19692] = data_o[44];
  assign data_o[19756] = data_o[44];
  assign data_o[19820] = data_o[44];
  assign data_o[19884] = data_o[44];
  assign data_o[19948] = data_o[44];
  assign data_o[20012] = data_o[44];
  assign data_o[20076] = data_o[44];
  assign data_o[20140] = data_o[44];
  assign data_o[20204] = data_o[44];
  assign data_o[20268] = data_o[44];
  assign data_o[20332] = data_o[44];
  assign data_o[20396] = data_o[44];
  assign data_o[20460] = data_o[44];
  assign data_o[20524] = data_o[44];
  assign data_o[20588] = data_o[44];
  assign data_o[20652] = data_o[44];
  assign data_o[20716] = data_o[44];
  assign data_o[20780] = data_o[44];
  assign data_o[20844] = data_o[44];
  assign data_o[20908] = data_o[44];
  assign data_o[20972] = data_o[44];
  assign data_o[21036] = data_o[44];
  assign data_o[21100] = data_o[44];
  assign data_o[21164] = data_o[44];
  assign data_o[21228] = data_o[44];
  assign data_o[21292] = data_o[44];
  assign data_o[21356] = data_o[44];
  assign data_o[21420] = data_o[44];
  assign data_o[21484] = data_o[44];
  assign data_o[21548] = data_o[44];
  assign data_o[21612] = data_o[44];
  assign data_o[21676] = data_o[44];
  assign data_o[21740] = data_o[44];
  assign data_o[21804] = data_o[44];
  assign data_o[21868] = data_o[44];
  assign data_o[21932] = data_o[44];
  assign data_o[21996] = data_o[44];
  assign data_o[22060] = data_o[44];
  assign data_o[22124] = data_o[44];
  assign data_o[22188] = data_o[44];
  assign data_o[22252] = data_o[44];
  assign data_o[22316] = data_o[44];
  assign data_o[22380] = data_o[44];
  assign data_o[22444] = data_o[44];
  assign data_o[22508] = data_o[44];
  assign data_o[22572] = data_o[44];
  assign data_o[22636] = data_o[44];
  assign data_o[22700] = data_o[44];
  assign data_o[22764] = data_o[44];
  assign data_o[22828] = data_o[44];
  assign data_o[22892] = data_o[44];
  assign data_o[22956] = data_o[44];
  assign data_o[23020] = data_o[44];
  assign data_o[23084] = data_o[44];
  assign data_o[23148] = data_o[44];
  assign data_o[23212] = data_o[44];
  assign data_o[23276] = data_o[44];
  assign data_o[23340] = data_o[44];
  assign data_o[23404] = data_o[44];
  assign data_o[23468] = data_o[44];
  assign data_o[23532] = data_o[44];
  assign data_o[23596] = data_o[44];
  assign data_o[23660] = data_o[44];
  assign data_o[23724] = data_o[44];
  assign data_o[23788] = data_o[44];
  assign data_o[23852] = data_o[44];
  assign data_o[23916] = data_o[44];
  assign data_o[23980] = data_o[44];
  assign data_o[24044] = data_o[44];
  assign data_o[24108] = data_o[44];
  assign data_o[24172] = data_o[44];
  assign data_o[24236] = data_o[44];
  assign data_o[24300] = data_o[44];
  assign data_o[24364] = data_o[44];
  assign data_o[24428] = data_o[44];
  assign data_o[24492] = data_o[44];
  assign data_o[24556] = data_o[44];
  assign data_o[24620] = data_o[44];
  assign data_o[24684] = data_o[44];
  assign data_o[24748] = data_o[44];
  assign data_o[24812] = data_o[44];
  assign data_o[24876] = data_o[44];
  assign data_o[24940] = data_o[44];
  assign data_o[25004] = data_o[44];
  assign data_o[25068] = data_o[44];
  assign data_o[25132] = data_o[44];
  assign data_o[25196] = data_o[44];
  assign data_o[25260] = data_o[44];
  assign data_o[25324] = data_o[44];
  assign data_o[25388] = data_o[44];
  assign data_o[25452] = data_o[44];
  assign data_o[25516] = data_o[44];
  assign data_o[25580] = data_o[44];
  assign data_o[25644] = data_o[44];
  assign data_o[25708] = data_o[44];
  assign data_o[25772] = data_o[44];
  assign data_o[25836] = data_o[44];
  assign data_o[25900] = data_o[44];
  assign data_o[25964] = data_o[44];
  assign data_o[26028] = data_o[44];
  assign data_o[26092] = data_o[44];
  assign data_o[26156] = data_o[44];
  assign data_o[26220] = data_o[44];
  assign data_o[26284] = data_o[44];
  assign data_o[26348] = data_o[44];
  assign data_o[26412] = data_o[44];
  assign data_o[26476] = data_o[44];
  assign data_o[26540] = data_o[44];
  assign data_o[26604] = data_o[44];
  assign data_o[26668] = data_o[44];
  assign data_o[26732] = data_o[44];
  assign data_o[26796] = data_o[44];
  assign data_o[26860] = data_o[44];
  assign data_o[26924] = data_o[44];
  assign data_o[26988] = data_o[44];
  assign data_o[27052] = data_o[44];
  assign data_o[27116] = data_o[44];
  assign data_o[27180] = data_o[44];
  assign data_o[27244] = data_o[44];
  assign data_o[27308] = data_o[44];
  assign data_o[27372] = data_o[44];
  assign data_o[27436] = data_o[44];
  assign data_o[27500] = data_o[44];
  assign data_o[27564] = data_o[44];
  assign data_o[27628] = data_o[44];
  assign data_o[27692] = data_o[44];
  assign data_o[27756] = data_o[44];
  assign data_o[27820] = data_o[44];
  assign data_o[27884] = data_o[44];
  assign data_o[27948] = data_o[44];
  assign data_o[28012] = data_o[44];
  assign data_o[28076] = data_o[44];
  assign data_o[28140] = data_o[44];
  assign data_o[28204] = data_o[44];
  assign data_o[28268] = data_o[44];
  assign data_o[28332] = data_o[44];
  assign data_o[28396] = data_o[44];
  assign data_o[28460] = data_o[44];
  assign data_o[28524] = data_o[44];
  assign data_o[28588] = data_o[44];
  assign data_o[28652] = data_o[44];
  assign data_o[28716] = data_o[44];
  assign data_o[28780] = data_o[44];
  assign data_o[28844] = data_o[44];
  assign data_o[28908] = data_o[44];
  assign data_o[28972] = data_o[44];
  assign data_o[29036] = data_o[44];
  assign data_o[29100] = data_o[44];
  assign data_o[29164] = data_o[44];
  assign data_o[29228] = data_o[44];
  assign data_o[29292] = data_o[44];
  assign data_o[29356] = data_o[44];
  assign data_o[29420] = data_o[44];
  assign data_o[29484] = data_o[44];
  assign data_o[29548] = data_o[44];
  assign data_o[29612] = data_o[44];
  assign data_o[29676] = data_o[44];
  assign data_o[29740] = data_o[44];
  assign data_o[29804] = data_o[44];
  assign data_o[29868] = data_o[44];
  assign data_o[29932] = data_o[44];
  assign data_o[29996] = data_o[44];
  assign data_o[30060] = data_o[44];
  assign data_o[30124] = data_o[44];
  assign data_o[30188] = data_o[44];
  assign data_o[30252] = data_o[44];
  assign data_o[30316] = data_o[44];
  assign data_o[30380] = data_o[44];
  assign data_o[30444] = data_o[44];
  assign data_o[30508] = data_o[44];
  assign data_o[30572] = data_o[44];
  assign data_o[30636] = data_o[44];
  assign data_o[30700] = data_o[44];
  assign data_o[30764] = data_o[44];
  assign data_o[30828] = data_o[44];
  assign data_o[30892] = data_o[44];
  assign data_o[30956] = data_o[44];
  assign data_o[31020] = data_o[44];
  assign data_o[31084] = data_o[44];
  assign data_o[31148] = data_o[44];
  assign data_o[31212] = data_o[44];
  assign data_o[31276] = data_o[44];
  assign data_o[31340] = data_o[44];
  assign data_o[31404] = data_o[44];
  assign data_o[31468] = data_o[44];
  assign data_o[31532] = data_o[44];
  assign data_o[31596] = data_o[44];
  assign data_o[31660] = data_o[44];
  assign data_o[31724] = data_o[44];
  assign data_o[31788] = data_o[44];
  assign data_o[31852] = data_o[44];
  assign data_o[31916] = data_o[44];
  assign data_o[31980] = data_o[44];
  assign data_o[107] = data_o[43];
  assign data_o[171] = data_o[43];
  assign data_o[235] = data_o[43];
  assign data_o[299] = data_o[43];
  assign data_o[363] = data_o[43];
  assign data_o[427] = data_o[43];
  assign data_o[491] = data_o[43];
  assign data_o[555] = data_o[43];
  assign data_o[619] = data_o[43];
  assign data_o[683] = data_o[43];
  assign data_o[747] = data_o[43];
  assign data_o[811] = data_o[43];
  assign data_o[875] = data_o[43];
  assign data_o[939] = data_o[43];
  assign data_o[1003] = data_o[43];
  assign data_o[1067] = data_o[43];
  assign data_o[1131] = data_o[43];
  assign data_o[1195] = data_o[43];
  assign data_o[1259] = data_o[43];
  assign data_o[1323] = data_o[43];
  assign data_o[1387] = data_o[43];
  assign data_o[1451] = data_o[43];
  assign data_o[1515] = data_o[43];
  assign data_o[1579] = data_o[43];
  assign data_o[1643] = data_o[43];
  assign data_o[1707] = data_o[43];
  assign data_o[1771] = data_o[43];
  assign data_o[1835] = data_o[43];
  assign data_o[1899] = data_o[43];
  assign data_o[1963] = data_o[43];
  assign data_o[2027] = data_o[43];
  assign data_o[2091] = data_o[43];
  assign data_o[2155] = data_o[43];
  assign data_o[2219] = data_o[43];
  assign data_o[2283] = data_o[43];
  assign data_o[2347] = data_o[43];
  assign data_o[2411] = data_o[43];
  assign data_o[2475] = data_o[43];
  assign data_o[2539] = data_o[43];
  assign data_o[2603] = data_o[43];
  assign data_o[2667] = data_o[43];
  assign data_o[2731] = data_o[43];
  assign data_o[2795] = data_o[43];
  assign data_o[2859] = data_o[43];
  assign data_o[2923] = data_o[43];
  assign data_o[2987] = data_o[43];
  assign data_o[3051] = data_o[43];
  assign data_o[3115] = data_o[43];
  assign data_o[3179] = data_o[43];
  assign data_o[3243] = data_o[43];
  assign data_o[3307] = data_o[43];
  assign data_o[3371] = data_o[43];
  assign data_o[3435] = data_o[43];
  assign data_o[3499] = data_o[43];
  assign data_o[3563] = data_o[43];
  assign data_o[3627] = data_o[43];
  assign data_o[3691] = data_o[43];
  assign data_o[3755] = data_o[43];
  assign data_o[3819] = data_o[43];
  assign data_o[3883] = data_o[43];
  assign data_o[3947] = data_o[43];
  assign data_o[4011] = data_o[43];
  assign data_o[4075] = data_o[43];
  assign data_o[4139] = data_o[43];
  assign data_o[4203] = data_o[43];
  assign data_o[4267] = data_o[43];
  assign data_o[4331] = data_o[43];
  assign data_o[4395] = data_o[43];
  assign data_o[4459] = data_o[43];
  assign data_o[4523] = data_o[43];
  assign data_o[4587] = data_o[43];
  assign data_o[4651] = data_o[43];
  assign data_o[4715] = data_o[43];
  assign data_o[4779] = data_o[43];
  assign data_o[4843] = data_o[43];
  assign data_o[4907] = data_o[43];
  assign data_o[4971] = data_o[43];
  assign data_o[5035] = data_o[43];
  assign data_o[5099] = data_o[43];
  assign data_o[5163] = data_o[43];
  assign data_o[5227] = data_o[43];
  assign data_o[5291] = data_o[43];
  assign data_o[5355] = data_o[43];
  assign data_o[5419] = data_o[43];
  assign data_o[5483] = data_o[43];
  assign data_o[5547] = data_o[43];
  assign data_o[5611] = data_o[43];
  assign data_o[5675] = data_o[43];
  assign data_o[5739] = data_o[43];
  assign data_o[5803] = data_o[43];
  assign data_o[5867] = data_o[43];
  assign data_o[5931] = data_o[43];
  assign data_o[5995] = data_o[43];
  assign data_o[6059] = data_o[43];
  assign data_o[6123] = data_o[43];
  assign data_o[6187] = data_o[43];
  assign data_o[6251] = data_o[43];
  assign data_o[6315] = data_o[43];
  assign data_o[6379] = data_o[43];
  assign data_o[6443] = data_o[43];
  assign data_o[6507] = data_o[43];
  assign data_o[6571] = data_o[43];
  assign data_o[6635] = data_o[43];
  assign data_o[6699] = data_o[43];
  assign data_o[6763] = data_o[43];
  assign data_o[6827] = data_o[43];
  assign data_o[6891] = data_o[43];
  assign data_o[6955] = data_o[43];
  assign data_o[7019] = data_o[43];
  assign data_o[7083] = data_o[43];
  assign data_o[7147] = data_o[43];
  assign data_o[7211] = data_o[43];
  assign data_o[7275] = data_o[43];
  assign data_o[7339] = data_o[43];
  assign data_o[7403] = data_o[43];
  assign data_o[7467] = data_o[43];
  assign data_o[7531] = data_o[43];
  assign data_o[7595] = data_o[43];
  assign data_o[7659] = data_o[43];
  assign data_o[7723] = data_o[43];
  assign data_o[7787] = data_o[43];
  assign data_o[7851] = data_o[43];
  assign data_o[7915] = data_o[43];
  assign data_o[7979] = data_o[43];
  assign data_o[8043] = data_o[43];
  assign data_o[8107] = data_o[43];
  assign data_o[8171] = data_o[43];
  assign data_o[8235] = data_o[43];
  assign data_o[8299] = data_o[43];
  assign data_o[8363] = data_o[43];
  assign data_o[8427] = data_o[43];
  assign data_o[8491] = data_o[43];
  assign data_o[8555] = data_o[43];
  assign data_o[8619] = data_o[43];
  assign data_o[8683] = data_o[43];
  assign data_o[8747] = data_o[43];
  assign data_o[8811] = data_o[43];
  assign data_o[8875] = data_o[43];
  assign data_o[8939] = data_o[43];
  assign data_o[9003] = data_o[43];
  assign data_o[9067] = data_o[43];
  assign data_o[9131] = data_o[43];
  assign data_o[9195] = data_o[43];
  assign data_o[9259] = data_o[43];
  assign data_o[9323] = data_o[43];
  assign data_o[9387] = data_o[43];
  assign data_o[9451] = data_o[43];
  assign data_o[9515] = data_o[43];
  assign data_o[9579] = data_o[43];
  assign data_o[9643] = data_o[43];
  assign data_o[9707] = data_o[43];
  assign data_o[9771] = data_o[43];
  assign data_o[9835] = data_o[43];
  assign data_o[9899] = data_o[43];
  assign data_o[9963] = data_o[43];
  assign data_o[10027] = data_o[43];
  assign data_o[10091] = data_o[43];
  assign data_o[10155] = data_o[43];
  assign data_o[10219] = data_o[43];
  assign data_o[10283] = data_o[43];
  assign data_o[10347] = data_o[43];
  assign data_o[10411] = data_o[43];
  assign data_o[10475] = data_o[43];
  assign data_o[10539] = data_o[43];
  assign data_o[10603] = data_o[43];
  assign data_o[10667] = data_o[43];
  assign data_o[10731] = data_o[43];
  assign data_o[10795] = data_o[43];
  assign data_o[10859] = data_o[43];
  assign data_o[10923] = data_o[43];
  assign data_o[10987] = data_o[43];
  assign data_o[11051] = data_o[43];
  assign data_o[11115] = data_o[43];
  assign data_o[11179] = data_o[43];
  assign data_o[11243] = data_o[43];
  assign data_o[11307] = data_o[43];
  assign data_o[11371] = data_o[43];
  assign data_o[11435] = data_o[43];
  assign data_o[11499] = data_o[43];
  assign data_o[11563] = data_o[43];
  assign data_o[11627] = data_o[43];
  assign data_o[11691] = data_o[43];
  assign data_o[11755] = data_o[43];
  assign data_o[11819] = data_o[43];
  assign data_o[11883] = data_o[43];
  assign data_o[11947] = data_o[43];
  assign data_o[12011] = data_o[43];
  assign data_o[12075] = data_o[43];
  assign data_o[12139] = data_o[43];
  assign data_o[12203] = data_o[43];
  assign data_o[12267] = data_o[43];
  assign data_o[12331] = data_o[43];
  assign data_o[12395] = data_o[43];
  assign data_o[12459] = data_o[43];
  assign data_o[12523] = data_o[43];
  assign data_o[12587] = data_o[43];
  assign data_o[12651] = data_o[43];
  assign data_o[12715] = data_o[43];
  assign data_o[12779] = data_o[43];
  assign data_o[12843] = data_o[43];
  assign data_o[12907] = data_o[43];
  assign data_o[12971] = data_o[43];
  assign data_o[13035] = data_o[43];
  assign data_o[13099] = data_o[43];
  assign data_o[13163] = data_o[43];
  assign data_o[13227] = data_o[43];
  assign data_o[13291] = data_o[43];
  assign data_o[13355] = data_o[43];
  assign data_o[13419] = data_o[43];
  assign data_o[13483] = data_o[43];
  assign data_o[13547] = data_o[43];
  assign data_o[13611] = data_o[43];
  assign data_o[13675] = data_o[43];
  assign data_o[13739] = data_o[43];
  assign data_o[13803] = data_o[43];
  assign data_o[13867] = data_o[43];
  assign data_o[13931] = data_o[43];
  assign data_o[13995] = data_o[43];
  assign data_o[14059] = data_o[43];
  assign data_o[14123] = data_o[43];
  assign data_o[14187] = data_o[43];
  assign data_o[14251] = data_o[43];
  assign data_o[14315] = data_o[43];
  assign data_o[14379] = data_o[43];
  assign data_o[14443] = data_o[43];
  assign data_o[14507] = data_o[43];
  assign data_o[14571] = data_o[43];
  assign data_o[14635] = data_o[43];
  assign data_o[14699] = data_o[43];
  assign data_o[14763] = data_o[43];
  assign data_o[14827] = data_o[43];
  assign data_o[14891] = data_o[43];
  assign data_o[14955] = data_o[43];
  assign data_o[15019] = data_o[43];
  assign data_o[15083] = data_o[43];
  assign data_o[15147] = data_o[43];
  assign data_o[15211] = data_o[43];
  assign data_o[15275] = data_o[43];
  assign data_o[15339] = data_o[43];
  assign data_o[15403] = data_o[43];
  assign data_o[15467] = data_o[43];
  assign data_o[15531] = data_o[43];
  assign data_o[15595] = data_o[43];
  assign data_o[15659] = data_o[43];
  assign data_o[15723] = data_o[43];
  assign data_o[15787] = data_o[43];
  assign data_o[15851] = data_o[43];
  assign data_o[15915] = data_o[43];
  assign data_o[15979] = data_o[43];
  assign data_o[16043] = data_o[43];
  assign data_o[16107] = data_o[43];
  assign data_o[16171] = data_o[43];
  assign data_o[16235] = data_o[43];
  assign data_o[16299] = data_o[43];
  assign data_o[16363] = data_o[43];
  assign data_o[16427] = data_o[43];
  assign data_o[16491] = data_o[43];
  assign data_o[16555] = data_o[43];
  assign data_o[16619] = data_o[43];
  assign data_o[16683] = data_o[43];
  assign data_o[16747] = data_o[43];
  assign data_o[16811] = data_o[43];
  assign data_o[16875] = data_o[43];
  assign data_o[16939] = data_o[43];
  assign data_o[17003] = data_o[43];
  assign data_o[17067] = data_o[43];
  assign data_o[17131] = data_o[43];
  assign data_o[17195] = data_o[43];
  assign data_o[17259] = data_o[43];
  assign data_o[17323] = data_o[43];
  assign data_o[17387] = data_o[43];
  assign data_o[17451] = data_o[43];
  assign data_o[17515] = data_o[43];
  assign data_o[17579] = data_o[43];
  assign data_o[17643] = data_o[43];
  assign data_o[17707] = data_o[43];
  assign data_o[17771] = data_o[43];
  assign data_o[17835] = data_o[43];
  assign data_o[17899] = data_o[43];
  assign data_o[17963] = data_o[43];
  assign data_o[18027] = data_o[43];
  assign data_o[18091] = data_o[43];
  assign data_o[18155] = data_o[43];
  assign data_o[18219] = data_o[43];
  assign data_o[18283] = data_o[43];
  assign data_o[18347] = data_o[43];
  assign data_o[18411] = data_o[43];
  assign data_o[18475] = data_o[43];
  assign data_o[18539] = data_o[43];
  assign data_o[18603] = data_o[43];
  assign data_o[18667] = data_o[43];
  assign data_o[18731] = data_o[43];
  assign data_o[18795] = data_o[43];
  assign data_o[18859] = data_o[43];
  assign data_o[18923] = data_o[43];
  assign data_o[18987] = data_o[43];
  assign data_o[19051] = data_o[43];
  assign data_o[19115] = data_o[43];
  assign data_o[19179] = data_o[43];
  assign data_o[19243] = data_o[43];
  assign data_o[19307] = data_o[43];
  assign data_o[19371] = data_o[43];
  assign data_o[19435] = data_o[43];
  assign data_o[19499] = data_o[43];
  assign data_o[19563] = data_o[43];
  assign data_o[19627] = data_o[43];
  assign data_o[19691] = data_o[43];
  assign data_o[19755] = data_o[43];
  assign data_o[19819] = data_o[43];
  assign data_o[19883] = data_o[43];
  assign data_o[19947] = data_o[43];
  assign data_o[20011] = data_o[43];
  assign data_o[20075] = data_o[43];
  assign data_o[20139] = data_o[43];
  assign data_o[20203] = data_o[43];
  assign data_o[20267] = data_o[43];
  assign data_o[20331] = data_o[43];
  assign data_o[20395] = data_o[43];
  assign data_o[20459] = data_o[43];
  assign data_o[20523] = data_o[43];
  assign data_o[20587] = data_o[43];
  assign data_o[20651] = data_o[43];
  assign data_o[20715] = data_o[43];
  assign data_o[20779] = data_o[43];
  assign data_o[20843] = data_o[43];
  assign data_o[20907] = data_o[43];
  assign data_o[20971] = data_o[43];
  assign data_o[21035] = data_o[43];
  assign data_o[21099] = data_o[43];
  assign data_o[21163] = data_o[43];
  assign data_o[21227] = data_o[43];
  assign data_o[21291] = data_o[43];
  assign data_o[21355] = data_o[43];
  assign data_o[21419] = data_o[43];
  assign data_o[21483] = data_o[43];
  assign data_o[21547] = data_o[43];
  assign data_o[21611] = data_o[43];
  assign data_o[21675] = data_o[43];
  assign data_o[21739] = data_o[43];
  assign data_o[21803] = data_o[43];
  assign data_o[21867] = data_o[43];
  assign data_o[21931] = data_o[43];
  assign data_o[21995] = data_o[43];
  assign data_o[22059] = data_o[43];
  assign data_o[22123] = data_o[43];
  assign data_o[22187] = data_o[43];
  assign data_o[22251] = data_o[43];
  assign data_o[22315] = data_o[43];
  assign data_o[22379] = data_o[43];
  assign data_o[22443] = data_o[43];
  assign data_o[22507] = data_o[43];
  assign data_o[22571] = data_o[43];
  assign data_o[22635] = data_o[43];
  assign data_o[22699] = data_o[43];
  assign data_o[22763] = data_o[43];
  assign data_o[22827] = data_o[43];
  assign data_o[22891] = data_o[43];
  assign data_o[22955] = data_o[43];
  assign data_o[23019] = data_o[43];
  assign data_o[23083] = data_o[43];
  assign data_o[23147] = data_o[43];
  assign data_o[23211] = data_o[43];
  assign data_o[23275] = data_o[43];
  assign data_o[23339] = data_o[43];
  assign data_o[23403] = data_o[43];
  assign data_o[23467] = data_o[43];
  assign data_o[23531] = data_o[43];
  assign data_o[23595] = data_o[43];
  assign data_o[23659] = data_o[43];
  assign data_o[23723] = data_o[43];
  assign data_o[23787] = data_o[43];
  assign data_o[23851] = data_o[43];
  assign data_o[23915] = data_o[43];
  assign data_o[23979] = data_o[43];
  assign data_o[24043] = data_o[43];
  assign data_o[24107] = data_o[43];
  assign data_o[24171] = data_o[43];
  assign data_o[24235] = data_o[43];
  assign data_o[24299] = data_o[43];
  assign data_o[24363] = data_o[43];
  assign data_o[24427] = data_o[43];
  assign data_o[24491] = data_o[43];
  assign data_o[24555] = data_o[43];
  assign data_o[24619] = data_o[43];
  assign data_o[24683] = data_o[43];
  assign data_o[24747] = data_o[43];
  assign data_o[24811] = data_o[43];
  assign data_o[24875] = data_o[43];
  assign data_o[24939] = data_o[43];
  assign data_o[25003] = data_o[43];
  assign data_o[25067] = data_o[43];
  assign data_o[25131] = data_o[43];
  assign data_o[25195] = data_o[43];
  assign data_o[25259] = data_o[43];
  assign data_o[25323] = data_o[43];
  assign data_o[25387] = data_o[43];
  assign data_o[25451] = data_o[43];
  assign data_o[25515] = data_o[43];
  assign data_o[25579] = data_o[43];
  assign data_o[25643] = data_o[43];
  assign data_o[25707] = data_o[43];
  assign data_o[25771] = data_o[43];
  assign data_o[25835] = data_o[43];
  assign data_o[25899] = data_o[43];
  assign data_o[25963] = data_o[43];
  assign data_o[26027] = data_o[43];
  assign data_o[26091] = data_o[43];
  assign data_o[26155] = data_o[43];
  assign data_o[26219] = data_o[43];
  assign data_o[26283] = data_o[43];
  assign data_o[26347] = data_o[43];
  assign data_o[26411] = data_o[43];
  assign data_o[26475] = data_o[43];
  assign data_o[26539] = data_o[43];
  assign data_o[26603] = data_o[43];
  assign data_o[26667] = data_o[43];
  assign data_o[26731] = data_o[43];
  assign data_o[26795] = data_o[43];
  assign data_o[26859] = data_o[43];
  assign data_o[26923] = data_o[43];
  assign data_o[26987] = data_o[43];
  assign data_o[27051] = data_o[43];
  assign data_o[27115] = data_o[43];
  assign data_o[27179] = data_o[43];
  assign data_o[27243] = data_o[43];
  assign data_o[27307] = data_o[43];
  assign data_o[27371] = data_o[43];
  assign data_o[27435] = data_o[43];
  assign data_o[27499] = data_o[43];
  assign data_o[27563] = data_o[43];
  assign data_o[27627] = data_o[43];
  assign data_o[27691] = data_o[43];
  assign data_o[27755] = data_o[43];
  assign data_o[27819] = data_o[43];
  assign data_o[27883] = data_o[43];
  assign data_o[27947] = data_o[43];
  assign data_o[28011] = data_o[43];
  assign data_o[28075] = data_o[43];
  assign data_o[28139] = data_o[43];
  assign data_o[28203] = data_o[43];
  assign data_o[28267] = data_o[43];
  assign data_o[28331] = data_o[43];
  assign data_o[28395] = data_o[43];
  assign data_o[28459] = data_o[43];
  assign data_o[28523] = data_o[43];
  assign data_o[28587] = data_o[43];
  assign data_o[28651] = data_o[43];
  assign data_o[28715] = data_o[43];
  assign data_o[28779] = data_o[43];
  assign data_o[28843] = data_o[43];
  assign data_o[28907] = data_o[43];
  assign data_o[28971] = data_o[43];
  assign data_o[29035] = data_o[43];
  assign data_o[29099] = data_o[43];
  assign data_o[29163] = data_o[43];
  assign data_o[29227] = data_o[43];
  assign data_o[29291] = data_o[43];
  assign data_o[29355] = data_o[43];
  assign data_o[29419] = data_o[43];
  assign data_o[29483] = data_o[43];
  assign data_o[29547] = data_o[43];
  assign data_o[29611] = data_o[43];
  assign data_o[29675] = data_o[43];
  assign data_o[29739] = data_o[43];
  assign data_o[29803] = data_o[43];
  assign data_o[29867] = data_o[43];
  assign data_o[29931] = data_o[43];
  assign data_o[29995] = data_o[43];
  assign data_o[30059] = data_o[43];
  assign data_o[30123] = data_o[43];
  assign data_o[30187] = data_o[43];
  assign data_o[30251] = data_o[43];
  assign data_o[30315] = data_o[43];
  assign data_o[30379] = data_o[43];
  assign data_o[30443] = data_o[43];
  assign data_o[30507] = data_o[43];
  assign data_o[30571] = data_o[43];
  assign data_o[30635] = data_o[43];
  assign data_o[30699] = data_o[43];
  assign data_o[30763] = data_o[43];
  assign data_o[30827] = data_o[43];
  assign data_o[30891] = data_o[43];
  assign data_o[30955] = data_o[43];
  assign data_o[31019] = data_o[43];
  assign data_o[31083] = data_o[43];
  assign data_o[31147] = data_o[43];
  assign data_o[31211] = data_o[43];
  assign data_o[31275] = data_o[43];
  assign data_o[31339] = data_o[43];
  assign data_o[31403] = data_o[43];
  assign data_o[31467] = data_o[43];
  assign data_o[31531] = data_o[43];
  assign data_o[31595] = data_o[43];
  assign data_o[31659] = data_o[43];
  assign data_o[31723] = data_o[43];
  assign data_o[31787] = data_o[43];
  assign data_o[31851] = data_o[43];
  assign data_o[31915] = data_o[43];
  assign data_o[31979] = data_o[43];
  assign data_o[106] = data_o[42];
  assign data_o[170] = data_o[42];
  assign data_o[234] = data_o[42];
  assign data_o[298] = data_o[42];
  assign data_o[362] = data_o[42];
  assign data_o[426] = data_o[42];
  assign data_o[490] = data_o[42];
  assign data_o[554] = data_o[42];
  assign data_o[618] = data_o[42];
  assign data_o[682] = data_o[42];
  assign data_o[746] = data_o[42];
  assign data_o[810] = data_o[42];
  assign data_o[874] = data_o[42];
  assign data_o[938] = data_o[42];
  assign data_o[1002] = data_o[42];
  assign data_o[1066] = data_o[42];
  assign data_o[1130] = data_o[42];
  assign data_o[1194] = data_o[42];
  assign data_o[1258] = data_o[42];
  assign data_o[1322] = data_o[42];
  assign data_o[1386] = data_o[42];
  assign data_o[1450] = data_o[42];
  assign data_o[1514] = data_o[42];
  assign data_o[1578] = data_o[42];
  assign data_o[1642] = data_o[42];
  assign data_o[1706] = data_o[42];
  assign data_o[1770] = data_o[42];
  assign data_o[1834] = data_o[42];
  assign data_o[1898] = data_o[42];
  assign data_o[1962] = data_o[42];
  assign data_o[2026] = data_o[42];
  assign data_o[2090] = data_o[42];
  assign data_o[2154] = data_o[42];
  assign data_o[2218] = data_o[42];
  assign data_o[2282] = data_o[42];
  assign data_o[2346] = data_o[42];
  assign data_o[2410] = data_o[42];
  assign data_o[2474] = data_o[42];
  assign data_o[2538] = data_o[42];
  assign data_o[2602] = data_o[42];
  assign data_o[2666] = data_o[42];
  assign data_o[2730] = data_o[42];
  assign data_o[2794] = data_o[42];
  assign data_o[2858] = data_o[42];
  assign data_o[2922] = data_o[42];
  assign data_o[2986] = data_o[42];
  assign data_o[3050] = data_o[42];
  assign data_o[3114] = data_o[42];
  assign data_o[3178] = data_o[42];
  assign data_o[3242] = data_o[42];
  assign data_o[3306] = data_o[42];
  assign data_o[3370] = data_o[42];
  assign data_o[3434] = data_o[42];
  assign data_o[3498] = data_o[42];
  assign data_o[3562] = data_o[42];
  assign data_o[3626] = data_o[42];
  assign data_o[3690] = data_o[42];
  assign data_o[3754] = data_o[42];
  assign data_o[3818] = data_o[42];
  assign data_o[3882] = data_o[42];
  assign data_o[3946] = data_o[42];
  assign data_o[4010] = data_o[42];
  assign data_o[4074] = data_o[42];
  assign data_o[4138] = data_o[42];
  assign data_o[4202] = data_o[42];
  assign data_o[4266] = data_o[42];
  assign data_o[4330] = data_o[42];
  assign data_o[4394] = data_o[42];
  assign data_o[4458] = data_o[42];
  assign data_o[4522] = data_o[42];
  assign data_o[4586] = data_o[42];
  assign data_o[4650] = data_o[42];
  assign data_o[4714] = data_o[42];
  assign data_o[4778] = data_o[42];
  assign data_o[4842] = data_o[42];
  assign data_o[4906] = data_o[42];
  assign data_o[4970] = data_o[42];
  assign data_o[5034] = data_o[42];
  assign data_o[5098] = data_o[42];
  assign data_o[5162] = data_o[42];
  assign data_o[5226] = data_o[42];
  assign data_o[5290] = data_o[42];
  assign data_o[5354] = data_o[42];
  assign data_o[5418] = data_o[42];
  assign data_o[5482] = data_o[42];
  assign data_o[5546] = data_o[42];
  assign data_o[5610] = data_o[42];
  assign data_o[5674] = data_o[42];
  assign data_o[5738] = data_o[42];
  assign data_o[5802] = data_o[42];
  assign data_o[5866] = data_o[42];
  assign data_o[5930] = data_o[42];
  assign data_o[5994] = data_o[42];
  assign data_o[6058] = data_o[42];
  assign data_o[6122] = data_o[42];
  assign data_o[6186] = data_o[42];
  assign data_o[6250] = data_o[42];
  assign data_o[6314] = data_o[42];
  assign data_o[6378] = data_o[42];
  assign data_o[6442] = data_o[42];
  assign data_o[6506] = data_o[42];
  assign data_o[6570] = data_o[42];
  assign data_o[6634] = data_o[42];
  assign data_o[6698] = data_o[42];
  assign data_o[6762] = data_o[42];
  assign data_o[6826] = data_o[42];
  assign data_o[6890] = data_o[42];
  assign data_o[6954] = data_o[42];
  assign data_o[7018] = data_o[42];
  assign data_o[7082] = data_o[42];
  assign data_o[7146] = data_o[42];
  assign data_o[7210] = data_o[42];
  assign data_o[7274] = data_o[42];
  assign data_o[7338] = data_o[42];
  assign data_o[7402] = data_o[42];
  assign data_o[7466] = data_o[42];
  assign data_o[7530] = data_o[42];
  assign data_o[7594] = data_o[42];
  assign data_o[7658] = data_o[42];
  assign data_o[7722] = data_o[42];
  assign data_o[7786] = data_o[42];
  assign data_o[7850] = data_o[42];
  assign data_o[7914] = data_o[42];
  assign data_o[7978] = data_o[42];
  assign data_o[8042] = data_o[42];
  assign data_o[8106] = data_o[42];
  assign data_o[8170] = data_o[42];
  assign data_o[8234] = data_o[42];
  assign data_o[8298] = data_o[42];
  assign data_o[8362] = data_o[42];
  assign data_o[8426] = data_o[42];
  assign data_o[8490] = data_o[42];
  assign data_o[8554] = data_o[42];
  assign data_o[8618] = data_o[42];
  assign data_o[8682] = data_o[42];
  assign data_o[8746] = data_o[42];
  assign data_o[8810] = data_o[42];
  assign data_o[8874] = data_o[42];
  assign data_o[8938] = data_o[42];
  assign data_o[9002] = data_o[42];
  assign data_o[9066] = data_o[42];
  assign data_o[9130] = data_o[42];
  assign data_o[9194] = data_o[42];
  assign data_o[9258] = data_o[42];
  assign data_o[9322] = data_o[42];
  assign data_o[9386] = data_o[42];
  assign data_o[9450] = data_o[42];
  assign data_o[9514] = data_o[42];
  assign data_o[9578] = data_o[42];
  assign data_o[9642] = data_o[42];
  assign data_o[9706] = data_o[42];
  assign data_o[9770] = data_o[42];
  assign data_o[9834] = data_o[42];
  assign data_o[9898] = data_o[42];
  assign data_o[9962] = data_o[42];
  assign data_o[10026] = data_o[42];
  assign data_o[10090] = data_o[42];
  assign data_o[10154] = data_o[42];
  assign data_o[10218] = data_o[42];
  assign data_o[10282] = data_o[42];
  assign data_o[10346] = data_o[42];
  assign data_o[10410] = data_o[42];
  assign data_o[10474] = data_o[42];
  assign data_o[10538] = data_o[42];
  assign data_o[10602] = data_o[42];
  assign data_o[10666] = data_o[42];
  assign data_o[10730] = data_o[42];
  assign data_o[10794] = data_o[42];
  assign data_o[10858] = data_o[42];
  assign data_o[10922] = data_o[42];
  assign data_o[10986] = data_o[42];
  assign data_o[11050] = data_o[42];
  assign data_o[11114] = data_o[42];
  assign data_o[11178] = data_o[42];
  assign data_o[11242] = data_o[42];
  assign data_o[11306] = data_o[42];
  assign data_o[11370] = data_o[42];
  assign data_o[11434] = data_o[42];
  assign data_o[11498] = data_o[42];
  assign data_o[11562] = data_o[42];
  assign data_o[11626] = data_o[42];
  assign data_o[11690] = data_o[42];
  assign data_o[11754] = data_o[42];
  assign data_o[11818] = data_o[42];
  assign data_o[11882] = data_o[42];
  assign data_o[11946] = data_o[42];
  assign data_o[12010] = data_o[42];
  assign data_o[12074] = data_o[42];
  assign data_o[12138] = data_o[42];
  assign data_o[12202] = data_o[42];
  assign data_o[12266] = data_o[42];
  assign data_o[12330] = data_o[42];
  assign data_o[12394] = data_o[42];
  assign data_o[12458] = data_o[42];
  assign data_o[12522] = data_o[42];
  assign data_o[12586] = data_o[42];
  assign data_o[12650] = data_o[42];
  assign data_o[12714] = data_o[42];
  assign data_o[12778] = data_o[42];
  assign data_o[12842] = data_o[42];
  assign data_o[12906] = data_o[42];
  assign data_o[12970] = data_o[42];
  assign data_o[13034] = data_o[42];
  assign data_o[13098] = data_o[42];
  assign data_o[13162] = data_o[42];
  assign data_o[13226] = data_o[42];
  assign data_o[13290] = data_o[42];
  assign data_o[13354] = data_o[42];
  assign data_o[13418] = data_o[42];
  assign data_o[13482] = data_o[42];
  assign data_o[13546] = data_o[42];
  assign data_o[13610] = data_o[42];
  assign data_o[13674] = data_o[42];
  assign data_o[13738] = data_o[42];
  assign data_o[13802] = data_o[42];
  assign data_o[13866] = data_o[42];
  assign data_o[13930] = data_o[42];
  assign data_o[13994] = data_o[42];
  assign data_o[14058] = data_o[42];
  assign data_o[14122] = data_o[42];
  assign data_o[14186] = data_o[42];
  assign data_o[14250] = data_o[42];
  assign data_o[14314] = data_o[42];
  assign data_o[14378] = data_o[42];
  assign data_o[14442] = data_o[42];
  assign data_o[14506] = data_o[42];
  assign data_o[14570] = data_o[42];
  assign data_o[14634] = data_o[42];
  assign data_o[14698] = data_o[42];
  assign data_o[14762] = data_o[42];
  assign data_o[14826] = data_o[42];
  assign data_o[14890] = data_o[42];
  assign data_o[14954] = data_o[42];
  assign data_o[15018] = data_o[42];
  assign data_o[15082] = data_o[42];
  assign data_o[15146] = data_o[42];
  assign data_o[15210] = data_o[42];
  assign data_o[15274] = data_o[42];
  assign data_o[15338] = data_o[42];
  assign data_o[15402] = data_o[42];
  assign data_o[15466] = data_o[42];
  assign data_o[15530] = data_o[42];
  assign data_o[15594] = data_o[42];
  assign data_o[15658] = data_o[42];
  assign data_o[15722] = data_o[42];
  assign data_o[15786] = data_o[42];
  assign data_o[15850] = data_o[42];
  assign data_o[15914] = data_o[42];
  assign data_o[15978] = data_o[42];
  assign data_o[16042] = data_o[42];
  assign data_o[16106] = data_o[42];
  assign data_o[16170] = data_o[42];
  assign data_o[16234] = data_o[42];
  assign data_o[16298] = data_o[42];
  assign data_o[16362] = data_o[42];
  assign data_o[16426] = data_o[42];
  assign data_o[16490] = data_o[42];
  assign data_o[16554] = data_o[42];
  assign data_o[16618] = data_o[42];
  assign data_o[16682] = data_o[42];
  assign data_o[16746] = data_o[42];
  assign data_o[16810] = data_o[42];
  assign data_o[16874] = data_o[42];
  assign data_o[16938] = data_o[42];
  assign data_o[17002] = data_o[42];
  assign data_o[17066] = data_o[42];
  assign data_o[17130] = data_o[42];
  assign data_o[17194] = data_o[42];
  assign data_o[17258] = data_o[42];
  assign data_o[17322] = data_o[42];
  assign data_o[17386] = data_o[42];
  assign data_o[17450] = data_o[42];
  assign data_o[17514] = data_o[42];
  assign data_o[17578] = data_o[42];
  assign data_o[17642] = data_o[42];
  assign data_o[17706] = data_o[42];
  assign data_o[17770] = data_o[42];
  assign data_o[17834] = data_o[42];
  assign data_o[17898] = data_o[42];
  assign data_o[17962] = data_o[42];
  assign data_o[18026] = data_o[42];
  assign data_o[18090] = data_o[42];
  assign data_o[18154] = data_o[42];
  assign data_o[18218] = data_o[42];
  assign data_o[18282] = data_o[42];
  assign data_o[18346] = data_o[42];
  assign data_o[18410] = data_o[42];
  assign data_o[18474] = data_o[42];
  assign data_o[18538] = data_o[42];
  assign data_o[18602] = data_o[42];
  assign data_o[18666] = data_o[42];
  assign data_o[18730] = data_o[42];
  assign data_o[18794] = data_o[42];
  assign data_o[18858] = data_o[42];
  assign data_o[18922] = data_o[42];
  assign data_o[18986] = data_o[42];
  assign data_o[19050] = data_o[42];
  assign data_o[19114] = data_o[42];
  assign data_o[19178] = data_o[42];
  assign data_o[19242] = data_o[42];
  assign data_o[19306] = data_o[42];
  assign data_o[19370] = data_o[42];
  assign data_o[19434] = data_o[42];
  assign data_o[19498] = data_o[42];
  assign data_o[19562] = data_o[42];
  assign data_o[19626] = data_o[42];
  assign data_o[19690] = data_o[42];
  assign data_o[19754] = data_o[42];
  assign data_o[19818] = data_o[42];
  assign data_o[19882] = data_o[42];
  assign data_o[19946] = data_o[42];
  assign data_o[20010] = data_o[42];
  assign data_o[20074] = data_o[42];
  assign data_o[20138] = data_o[42];
  assign data_o[20202] = data_o[42];
  assign data_o[20266] = data_o[42];
  assign data_o[20330] = data_o[42];
  assign data_o[20394] = data_o[42];
  assign data_o[20458] = data_o[42];
  assign data_o[20522] = data_o[42];
  assign data_o[20586] = data_o[42];
  assign data_o[20650] = data_o[42];
  assign data_o[20714] = data_o[42];
  assign data_o[20778] = data_o[42];
  assign data_o[20842] = data_o[42];
  assign data_o[20906] = data_o[42];
  assign data_o[20970] = data_o[42];
  assign data_o[21034] = data_o[42];
  assign data_o[21098] = data_o[42];
  assign data_o[21162] = data_o[42];
  assign data_o[21226] = data_o[42];
  assign data_o[21290] = data_o[42];
  assign data_o[21354] = data_o[42];
  assign data_o[21418] = data_o[42];
  assign data_o[21482] = data_o[42];
  assign data_o[21546] = data_o[42];
  assign data_o[21610] = data_o[42];
  assign data_o[21674] = data_o[42];
  assign data_o[21738] = data_o[42];
  assign data_o[21802] = data_o[42];
  assign data_o[21866] = data_o[42];
  assign data_o[21930] = data_o[42];
  assign data_o[21994] = data_o[42];
  assign data_o[22058] = data_o[42];
  assign data_o[22122] = data_o[42];
  assign data_o[22186] = data_o[42];
  assign data_o[22250] = data_o[42];
  assign data_o[22314] = data_o[42];
  assign data_o[22378] = data_o[42];
  assign data_o[22442] = data_o[42];
  assign data_o[22506] = data_o[42];
  assign data_o[22570] = data_o[42];
  assign data_o[22634] = data_o[42];
  assign data_o[22698] = data_o[42];
  assign data_o[22762] = data_o[42];
  assign data_o[22826] = data_o[42];
  assign data_o[22890] = data_o[42];
  assign data_o[22954] = data_o[42];
  assign data_o[23018] = data_o[42];
  assign data_o[23082] = data_o[42];
  assign data_o[23146] = data_o[42];
  assign data_o[23210] = data_o[42];
  assign data_o[23274] = data_o[42];
  assign data_o[23338] = data_o[42];
  assign data_o[23402] = data_o[42];
  assign data_o[23466] = data_o[42];
  assign data_o[23530] = data_o[42];
  assign data_o[23594] = data_o[42];
  assign data_o[23658] = data_o[42];
  assign data_o[23722] = data_o[42];
  assign data_o[23786] = data_o[42];
  assign data_o[23850] = data_o[42];
  assign data_o[23914] = data_o[42];
  assign data_o[23978] = data_o[42];
  assign data_o[24042] = data_o[42];
  assign data_o[24106] = data_o[42];
  assign data_o[24170] = data_o[42];
  assign data_o[24234] = data_o[42];
  assign data_o[24298] = data_o[42];
  assign data_o[24362] = data_o[42];
  assign data_o[24426] = data_o[42];
  assign data_o[24490] = data_o[42];
  assign data_o[24554] = data_o[42];
  assign data_o[24618] = data_o[42];
  assign data_o[24682] = data_o[42];
  assign data_o[24746] = data_o[42];
  assign data_o[24810] = data_o[42];
  assign data_o[24874] = data_o[42];
  assign data_o[24938] = data_o[42];
  assign data_o[25002] = data_o[42];
  assign data_o[25066] = data_o[42];
  assign data_o[25130] = data_o[42];
  assign data_o[25194] = data_o[42];
  assign data_o[25258] = data_o[42];
  assign data_o[25322] = data_o[42];
  assign data_o[25386] = data_o[42];
  assign data_o[25450] = data_o[42];
  assign data_o[25514] = data_o[42];
  assign data_o[25578] = data_o[42];
  assign data_o[25642] = data_o[42];
  assign data_o[25706] = data_o[42];
  assign data_o[25770] = data_o[42];
  assign data_o[25834] = data_o[42];
  assign data_o[25898] = data_o[42];
  assign data_o[25962] = data_o[42];
  assign data_o[26026] = data_o[42];
  assign data_o[26090] = data_o[42];
  assign data_o[26154] = data_o[42];
  assign data_o[26218] = data_o[42];
  assign data_o[26282] = data_o[42];
  assign data_o[26346] = data_o[42];
  assign data_o[26410] = data_o[42];
  assign data_o[26474] = data_o[42];
  assign data_o[26538] = data_o[42];
  assign data_o[26602] = data_o[42];
  assign data_o[26666] = data_o[42];
  assign data_o[26730] = data_o[42];
  assign data_o[26794] = data_o[42];
  assign data_o[26858] = data_o[42];
  assign data_o[26922] = data_o[42];
  assign data_o[26986] = data_o[42];
  assign data_o[27050] = data_o[42];
  assign data_o[27114] = data_o[42];
  assign data_o[27178] = data_o[42];
  assign data_o[27242] = data_o[42];
  assign data_o[27306] = data_o[42];
  assign data_o[27370] = data_o[42];
  assign data_o[27434] = data_o[42];
  assign data_o[27498] = data_o[42];
  assign data_o[27562] = data_o[42];
  assign data_o[27626] = data_o[42];
  assign data_o[27690] = data_o[42];
  assign data_o[27754] = data_o[42];
  assign data_o[27818] = data_o[42];
  assign data_o[27882] = data_o[42];
  assign data_o[27946] = data_o[42];
  assign data_o[28010] = data_o[42];
  assign data_o[28074] = data_o[42];
  assign data_o[28138] = data_o[42];
  assign data_o[28202] = data_o[42];
  assign data_o[28266] = data_o[42];
  assign data_o[28330] = data_o[42];
  assign data_o[28394] = data_o[42];
  assign data_o[28458] = data_o[42];
  assign data_o[28522] = data_o[42];
  assign data_o[28586] = data_o[42];
  assign data_o[28650] = data_o[42];
  assign data_o[28714] = data_o[42];
  assign data_o[28778] = data_o[42];
  assign data_o[28842] = data_o[42];
  assign data_o[28906] = data_o[42];
  assign data_o[28970] = data_o[42];
  assign data_o[29034] = data_o[42];
  assign data_o[29098] = data_o[42];
  assign data_o[29162] = data_o[42];
  assign data_o[29226] = data_o[42];
  assign data_o[29290] = data_o[42];
  assign data_o[29354] = data_o[42];
  assign data_o[29418] = data_o[42];
  assign data_o[29482] = data_o[42];
  assign data_o[29546] = data_o[42];
  assign data_o[29610] = data_o[42];
  assign data_o[29674] = data_o[42];
  assign data_o[29738] = data_o[42];
  assign data_o[29802] = data_o[42];
  assign data_o[29866] = data_o[42];
  assign data_o[29930] = data_o[42];
  assign data_o[29994] = data_o[42];
  assign data_o[30058] = data_o[42];
  assign data_o[30122] = data_o[42];
  assign data_o[30186] = data_o[42];
  assign data_o[30250] = data_o[42];
  assign data_o[30314] = data_o[42];
  assign data_o[30378] = data_o[42];
  assign data_o[30442] = data_o[42];
  assign data_o[30506] = data_o[42];
  assign data_o[30570] = data_o[42];
  assign data_o[30634] = data_o[42];
  assign data_o[30698] = data_o[42];
  assign data_o[30762] = data_o[42];
  assign data_o[30826] = data_o[42];
  assign data_o[30890] = data_o[42];
  assign data_o[30954] = data_o[42];
  assign data_o[31018] = data_o[42];
  assign data_o[31082] = data_o[42];
  assign data_o[31146] = data_o[42];
  assign data_o[31210] = data_o[42];
  assign data_o[31274] = data_o[42];
  assign data_o[31338] = data_o[42];
  assign data_o[31402] = data_o[42];
  assign data_o[31466] = data_o[42];
  assign data_o[31530] = data_o[42];
  assign data_o[31594] = data_o[42];
  assign data_o[31658] = data_o[42];
  assign data_o[31722] = data_o[42];
  assign data_o[31786] = data_o[42];
  assign data_o[31850] = data_o[42];
  assign data_o[31914] = data_o[42];
  assign data_o[31978] = data_o[42];
  assign data_o[105] = data_o[41];
  assign data_o[169] = data_o[41];
  assign data_o[233] = data_o[41];
  assign data_o[297] = data_o[41];
  assign data_o[361] = data_o[41];
  assign data_o[425] = data_o[41];
  assign data_o[489] = data_o[41];
  assign data_o[553] = data_o[41];
  assign data_o[617] = data_o[41];
  assign data_o[681] = data_o[41];
  assign data_o[745] = data_o[41];
  assign data_o[809] = data_o[41];
  assign data_o[873] = data_o[41];
  assign data_o[937] = data_o[41];
  assign data_o[1001] = data_o[41];
  assign data_o[1065] = data_o[41];
  assign data_o[1129] = data_o[41];
  assign data_o[1193] = data_o[41];
  assign data_o[1257] = data_o[41];
  assign data_o[1321] = data_o[41];
  assign data_o[1385] = data_o[41];
  assign data_o[1449] = data_o[41];
  assign data_o[1513] = data_o[41];
  assign data_o[1577] = data_o[41];
  assign data_o[1641] = data_o[41];
  assign data_o[1705] = data_o[41];
  assign data_o[1769] = data_o[41];
  assign data_o[1833] = data_o[41];
  assign data_o[1897] = data_o[41];
  assign data_o[1961] = data_o[41];
  assign data_o[2025] = data_o[41];
  assign data_o[2089] = data_o[41];
  assign data_o[2153] = data_o[41];
  assign data_o[2217] = data_o[41];
  assign data_o[2281] = data_o[41];
  assign data_o[2345] = data_o[41];
  assign data_o[2409] = data_o[41];
  assign data_o[2473] = data_o[41];
  assign data_o[2537] = data_o[41];
  assign data_o[2601] = data_o[41];
  assign data_o[2665] = data_o[41];
  assign data_o[2729] = data_o[41];
  assign data_o[2793] = data_o[41];
  assign data_o[2857] = data_o[41];
  assign data_o[2921] = data_o[41];
  assign data_o[2985] = data_o[41];
  assign data_o[3049] = data_o[41];
  assign data_o[3113] = data_o[41];
  assign data_o[3177] = data_o[41];
  assign data_o[3241] = data_o[41];
  assign data_o[3305] = data_o[41];
  assign data_o[3369] = data_o[41];
  assign data_o[3433] = data_o[41];
  assign data_o[3497] = data_o[41];
  assign data_o[3561] = data_o[41];
  assign data_o[3625] = data_o[41];
  assign data_o[3689] = data_o[41];
  assign data_o[3753] = data_o[41];
  assign data_o[3817] = data_o[41];
  assign data_o[3881] = data_o[41];
  assign data_o[3945] = data_o[41];
  assign data_o[4009] = data_o[41];
  assign data_o[4073] = data_o[41];
  assign data_o[4137] = data_o[41];
  assign data_o[4201] = data_o[41];
  assign data_o[4265] = data_o[41];
  assign data_o[4329] = data_o[41];
  assign data_o[4393] = data_o[41];
  assign data_o[4457] = data_o[41];
  assign data_o[4521] = data_o[41];
  assign data_o[4585] = data_o[41];
  assign data_o[4649] = data_o[41];
  assign data_o[4713] = data_o[41];
  assign data_o[4777] = data_o[41];
  assign data_o[4841] = data_o[41];
  assign data_o[4905] = data_o[41];
  assign data_o[4969] = data_o[41];
  assign data_o[5033] = data_o[41];
  assign data_o[5097] = data_o[41];
  assign data_o[5161] = data_o[41];
  assign data_o[5225] = data_o[41];
  assign data_o[5289] = data_o[41];
  assign data_o[5353] = data_o[41];
  assign data_o[5417] = data_o[41];
  assign data_o[5481] = data_o[41];
  assign data_o[5545] = data_o[41];
  assign data_o[5609] = data_o[41];
  assign data_o[5673] = data_o[41];
  assign data_o[5737] = data_o[41];
  assign data_o[5801] = data_o[41];
  assign data_o[5865] = data_o[41];
  assign data_o[5929] = data_o[41];
  assign data_o[5993] = data_o[41];
  assign data_o[6057] = data_o[41];
  assign data_o[6121] = data_o[41];
  assign data_o[6185] = data_o[41];
  assign data_o[6249] = data_o[41];
  assign data_o[6313] = data_o[41];
  assign data_o[6377] = data_o[41];
  assign data_o[6441] = data_o[41];
  assign data_o[6505] = data_o[41];
  assign data_o[6569] = data_o[41];
  assign data_o[6633] = data_o[41];
  assign data_o[6697] = data_o[41];
  assign data_o[6761] = data_o[41];
  assign data_o[6825] = data_o[41];
  assign data_o[6889] = data_o[41];
  assign data_o[6953] = data_o[41];
  assign data_o[7017] = data_o[41];
  assign data_o[7081] = data_o[41];
  assign data_o[7145] = data_o[41];
  assign data_o[7209] = data_o[41];
  assign data_o[7273] = data_o[41];
  assign data_o[7337] = data_o[41];
  assign data_o[7401] = data_o[41];
  assign data_o[7465] = data_o[41];
  assign data_o[7529] = data_o[41];
  assign data_o[7593] = data_o[41];
  assign data_o[7657] = data_o[41];
  assign data_o[7721] = data_o[41];
  assign data_o[7785] = data_o[41];
  assign data_o[7849] = data_o[41];
  assign data_o[7913] = data_o[41];
  assign data_o[7977] = data_o[41];
  assign data_o[8041] = data_o[41];
  assign data_o[8105] = data_o[41];
  assign data_o[8169] = data_o[41];
  assign data_o[8233] = data_o[41];
  assign data_o[8297] = data_o[41];
  assign data_o[8361] = data_o[41];
  assign data_o[8425] = data_o[41];
  assign data_o[8489] = data_o[41];
  assign data_o[8553] = data_o[41];
  assign data_o[8617] = data_o[41];
  assign data_o[8681] = data_o[41];
  assign data_o[8745] = data_o[41];
  assign data_o[8809] = data_o[41];
  assign data_o[8873] = data_o[41];
  assign data_o[8937] = data_o[41];
  assign data_o[9001] = data_o[41];
  assign data_o[9065] = data_o[41];
  assign data_o[9129] = data_o[41];
  assign data_o[9193] = data_o[41];
  assign data_o[9257] = data_o[41];
  assign data_o[9321] = data_o[41];
  assign data_o[9385] = data_o[41];
  assign data_o[9449] = data_o[41];
  assign data_o[9513] = data_o[41];
  assign data_o[9577] = data_o[41];
  assign data_o[9641] = data_o[41];
  assign data_o[9705] = data_o[41];
  assign data_o[9769] = data_o[41];
  assign data_o[9833] = data_o[41];
  assign data_o[9897] = data_o[41];
  assign data_o[9961] = data_o[41];
  assign data_o[10025] = data_o[41];
  assign data_o[10089] = data_o[41];
  assign data_o[10153] = data_o[41];
  assign data_o[10217] = data_o[41];
  assign data_o[10281] = data_o[41];
  assign data_o[10345] = data_o[41];
  assign data_o[10409] = data_o[41];
  assign data_o[10473] = data_o[41];
  assign data_o[10537] = data_o[41];
  assign data_o[10601] = data_o[41];
  assign data_o[10665] = data_o[41];
  assign data_o[10729] = data_o[41];
  assign data_o[10793] = data_o[41];
  assign data_o[10857] = data_o[41];
  assign data_o[10921] = data_o[41];
  assign data_o[10985] = data_o[41];
  assign data_o[11049] = data_o[41];
  assign data_o[11113] = data_o[41];
  assign data_o[11177] = data_o[41];
  assign data_o[11241] = data_o[41];
  assign data_o[11305] = data_o[41];
  assign data_o[11369] = data_o[41];
  assign data_o[11433] = data_o[41];
  assign data_o[11497] = data_o[41];
  assign data_o[11561] = data_o[41];
  assign data_o[11625] = data_o[41];
  assign data_o[11689] = data_o[41];
  assign data_o[11753] = data_o[41];
  assign data_o[11817] = data_o[41];
  assign data_o[11881] = data_o[41];
  assign data_o[11945] = data_o[41];
  assign data_o[12009] = data_o[41];
  assign data_o[12073] = data_o[41];
  assign data_o[12137] = data_o[41];
  assign data_o[12201] = data_o[41];
  assign data_o[12265] = data_o[41];
  assign data_o[12329] = data_o[41];
  assign data_o[12393] = data_o[41];
  assign data_o[12457] = data_o[41];
  assign data_o[12521] = data_o[41];
  assign data_o[12585] = data_o[41];
  assign data_o[12649] = data_o[41];
  assign data_o[12713] = data_o[41];
  assign data_o[12777] = data_o[41];
  assign data_o[12841] = data_o[41];
  assign data_o[12905] = data_o[41];
  assign data_o[12969] = data_o[41];
  assign data_o[13033] = data_o[41];
  assign data_o[13097] = data_o[41];
  assign data_o[13161] = data_o[41];
  assign data_o[13225] = data_o[41];
  assign data_o[13289] = data_o[41];
  assign data_o[13353] = data_o[41];
  assign data_o[13417] = data_o[41];
  assign data_o[13481] = data_o[41];
  assign data_o[13545] = data_o[41];
  assign data_o[13609] = data_o[41];
  assign data_o[13673] = data_o[41];
  assign data_o[13737] = data_o[41];
  assign data_o[13801] = data_o[41];
  assign data_o[13865] = data_o[41];
  assign data_o[13929] = data_o[41];
  assign data_o[13993] = data_o[41];
  assign data_o[14057] = data_o[41];
  assign data_o[14121] = data_o[41];
  assign data_o[14185] = data_o[41];
  assign data_o[14249] = data_o[41];
  assign data_o[14313] = data_o[41];
  assign data_o[14377] = data_o[41];
  assign data_o[14441] = data_o[41];
  assign data_o[14505] = data_o[41];
  assign data_o[14569] = data_o[41];
  assign data_o[14633] = data_o[41];
  assign data_o[14697] = data_o[41];
  assign data_o[14761] = data_o[41];
  assign data_o[14825] = data_o[41];
  assign data_o[14889] = data_o[41];
  assign data_o[14953] = data_o[41];
  assign data_o[15017] = data_o[41];
  assign data_o[15081] = data_o[41];
  assign data_o[15145] = data_o[41];
  assign data_o[15209] = data_o[41];
  assign data_o[15273] = data_o[41];
  assign data_o[15337] = data_o[41];
  assign data_o[15401] = data_o[41];
  assign data_o[15465] = data_o[41];
  assign data_o[15529] = data_o[41];
  assign data_o[15593] = data_o[41];
  assign data_o[15657] = data_o[41];
  assign data_o[15721] = data_o[41];
  assign data_o[15785] = data_o[41];
  assign data_o[15849] = data_o[41];
  assign data_o[15913] = data_o[41];
  assign data_o[15977] = data_o[41];
  assign data_o[16041] = data_o[41];
  assign data_o[16105] = data_o[41];
  assign data_o[16169] = data_o[41];
  assign data_o[16233] = data_o[41];
  assign data_o[16297] = data_o[41];
  assign data_o[16361] = data_o[41];
  assign data_o[16425] = data_o[41];
  assign data_o[16489] = data_o[41];
  assign data_o[16553] = data_o[41];
  assign data_o[16617] = data_o[41];
  assign data_o[16681] = data_o[41];
  assign data_o[16745] = data_o[41];
  assign data_o[16809] = data_o[41];
  assign data_o[16873] = data_o[41];
  assign data_o[16937] = data_o[41];
  assign data_o[17001] = data_o[41];
  assign data_o[17065] = data_o[41];
  assign data_o[17129] = data_o[41];
  assign data_o[17193] = data_o[41];
  assign data_o[17257] = data_o[41];
  assign data_o[17321] = data_o[41];
  assign data_o[17385] = data_o[41];
  assign data_o[17449] = data_o[41];
  assign data_o[17513] = data_o[41];
  assign data_o[17577] = data_o[41];
  assign data_o[17641] = data_o[41];
  assign data_o[17705] = data_o[41];
  assign data_o[17769] = data_o[41];
  assign data_o[17833] = data_o[41];
  assign data_o[17897] = data_o[41];
  assign data_o[17961] = data_o[41];
  assign data_o[18025] = data_o[41];
  assign data_o[18089] = data_o[41];
  assign data_o[18153] = data_o[41];
  assign data_o[18217] = data_o[41];
  assign data_o[18281] = data_o[41];
  assign data_o[18345] = data_o[41];
  assign data_o[18409] = data_o[41];
  assign data_o[18473] = data_o[41];
  assign data_o[18537] = data_o[41];
  assign data_o[18601] = data_o[41];
  assign data_o[18665] = data_o[41];
  assign data_o[18729] = data_o[41];
  assign data_o[18793] = data_o[41];
  assign data_o[18857] = data_o[41];
  assign data_o[18921] = data_o[41];
  assign data_o[18985] = data_o[41];
  assign data_o[19049] = data_o[41];
  assign data_o[19113] = data_o[41];
  assign data_o[19177] = data_o[41];
  assign data_o[19241] = data_o[41];
  assign data_o[19305] = data_o[41];
  assign data_o[19369] = data_o[41];
  assign data_o[19433] = data_o[41];
  assign data_o[19497] = data_o[41];
  assign data_o[19561] = data_o[41];
  assign data_o[19625] = data_o[41];
  assign data_o[19689] = data_o[41];
  assign data_o[19753] = data_o[41];
  assign data_o[19817] = data_o[41];
  assign data_o[19881] = data_o[41];
  assign data_o[19945] = data_o[41];
  assign data_o[20009] = data_o[41];
  assign data_o[20073] = data_o[41];
  assign data_o[20137] = data_o[41];
  assign data_o[20201] = data_o[41];
  assign data_o[20265] = data_o[41];
  assign data_o[20329] = data_o[41];
  assign data_o[20393] = data_o[41];
  assign data_o[20457] = data_o[41];
  assign data_o[20521] = data_o[41];
  assign data_o[20585] = data_o[41];
  assign data_o[20649] = data_o[41];
  assign data_o[20713] = data_o[41];
  assign data_o[20777] = data_o[41];
  assign data_o[20841] = data_o[41];
  assign data_o[20905] = data_o[41];
  assign data_o[20969] = data_o[41];
  assign data_o[21033] = data_o[41];
  assign data_o[21097] = data_o[41];
  assign data_o[21161] = data_o[41];
  assign data_o[21225] = data_o[41];
  assign data_o[21289] = data_o[41];
  assign data_o[21353] = data_o[41];
  assign data_o[21417] = data_o[41];
  assign data_o[21481] = data_o[41];
  assign data_o[21545] = data_o[41];
  assign data_o[21609] = data_o[41];
  assign data_o[21673] = data_o[41];
  assign data_o[21737] = data_o[41];
  assign data_o[21801] = data_o[41];
  assign data_o[21865] = data_o[41];
  assign data_o[21929] = data_o[41];
  assign data_o[21993] = data_o[41];
  assign data_o[22057] = data_o[41];
  assign data_o[22121] = data_o[41];
  assign data_o[22185] = data_o[41];
  assign data_o[22249] = data_o[41];
  assign data_o[22313] = data_o[41];
  assign data_o[22377] = data_o[41];
  assign data_o[22441] = data_o[41];
  assign data_o[22505] = data_o[41];
  assign data_o[22569] = data_o[41];
  assign data_o[22633] = data_o[41];
  assign data_o[22697] = data_o[41];
  assign data_o[22761] = data_o[41];
  assign data_o[22825] = data_o[41];
  assign data_o[22889] = data_o[41];
  assign data_o[22953] = data_o[41];
  assign data_o[23017] = data_o[41];
  assign data_o[23081] = data_o[41];
  assign data_o[23145] = data_o[41];
  assign data_o[23209] = data_o[41];
  assign data_o[23273] = data_o[41];
  assign data_o[23337] = data_o[41];
  assign data_o[23401] = data_o[41];
  assign data_o[23465] = data_o[41];
  assign data_o[23529] = data_o[41];
  assign data_o[23593] = data_o[41];
  assign data_o[23657] = data_o[41];
  assign data_o[23721] = data_o[41];
  assign data_o[23785] = data_o[41];
  assign data_o[23849] = data_o[41];
  assign data_o[23913] = data_o[41];
  assign data_o[23977] = data_o[41];
  assign data_o[24041] = data_o[41];
  assign data_o[24105] = data_o[41];
  assign data_o[24169] = data_o[41];
  assign data_o[24233] = data_o[41];
  assign data_o[24297] = data_o[41];
  assign data_o[24361] = data_o[41];
  assign data_o[24425] = data_o[41];
  assign data_o[24489] = data_o[41];
  assign data_o[24553] = data_o[41];
  assign data_o[24617] = data_o[41];
  assign data_o[24681] = data_o[41];
  assign data_o[24745] = data_o[41];
  assign data_o[24809] = data_o[41];
  assign data_o[24873] = data_o[41];
  assign data_o[24937] = data_o[41];
  assign data_o[25001] = data_o[41];
  assign data_o[25065] = data_o[41];
  assign data_o[25129] = data_o[41];
  assign data_o[25193] = data_o[41];
  assign data_o[25257] = data_o[41];
  assign data_o[25321] = data_o[41];
  assign data_o[25385] = data_o[41];
  assign data_o[25449] = data_o[41];
  assign data_o[25513] = data_o[41];
  assign data_o[25577] = data_o[41];
  assign data_o[25641] = data_o[41];
  assign data_o[25705] = data_o[41];
  assign data_o[25769] = data_o[41];
  assign data_o[25833] = data_o[41];
  assign data_o[25897] = data_o[41];
  assign data_o[25961] = data_o[41];
  assign data_o[26025] = data_o[41];
  assign data_o[26089] = data_o[41];
  assign data_o[26153] = data_o[41];
  assign data_o[26217] = data_o[41];
  assign data_o[26281] = data_o[41];
  assign data_o[26345] = data_o[41];
  assign data_o[26409] = data_o[41];
  assign data_o[26473] = data_o[41];
  assign data_o[26537] = data_o[41];
  assign data_o[26601] = data_o[41];
  assign data_o[26665] = data_o[41];
  assign data_o[26729] = data_o[41];
  assign data_o[26793] = data_o[41];
  assign data_o[26857] = data_o[41];
  assign data_o[26921] = data_o[41];
  assign data_o[26985] = data_o[41];
  assign data_o[27049] = data_o[41];
  assign data_o[27113] = data_o[41];
  assign data_o[27177] = data_o[41];
  assign data_o[27241] = data_o[41];
  assign data_o[27305] = data_o[41];
  assign data_o[27369] = data_o[41];
  assign data_o[27433] = data_o[41];
  assign data_o[27497] = data_o[41];
  assign data_o[27561] = data_o[41];
  assign data_o[27625] = data_o[41];
  assign data_o[27689] = data_o[41];
  assign data_o[27753] = data_o[41];
  assign data_o[27817] = data_o[41];
  assign data_o[27881] = data_o[41];
  assign data_o[27945] = data_o[41];
  assign data_o[28009] = data_o[41];
  assign data_o[28073] = data_o[41];
  assign data_o[28137] = data_o[41];
  assign data_o[28201] = data_o[41];
  assign data_o[28265] = data_o[41];
  assign data_o[28329] = data_o[41];
  assign data_o[28393] = data_o[41];
  assign data_o[28457] = data_o[41];
  assign data_o[28521] = data_o[41];
  assign data_o[28585] = data_o[41];
  assign data_o[28649] = data_o[41];
  assign data_o[28713] = data_o[41];
  assign data_o[28777] = data_o[41];
  assign data_o[28841] = data_o[41];
  assign data_o[28905] = data_o[41];
  assign data_o[28969] = data_o[41];
  assign data_o[29033] = data_o[41];
  assign data_o[29097] = data_o[41];
  assign data_o[29161] = data_o[41];
  assign data_o[29225] = data_o[41];
  assign data_o[29289] = data_o[41];
  assign data_o[29353] = data_o[41];
  assign data_o[29417] = data_o[41];
  assign data_o[29481] = data_o[41];
  assign data_o[29545] = data_o[41];
  assign data_o[29609] = data_o[41];
  assign data_o[29673] = data_o[41];
  assign data_o[29737] = data_o[41];
  assign data_o[29801] = data_o[41];
  assign data_o[29865] = data_o[41];
  assign data_o[29929] = data_o[41];
  assign data_o[29993] = data_o[41];
  assign data_o[30057] = data_o[41];
  assign data_o[30121] = data_o[41];
  assign data_o[30185] = data_o[41];
  assign data_o[30249] = data_o[41];
  assign data_o[30313] = data_o[41];
  assign data_o[30377] = data_o[41];
  assign data_o[30441] = data_o[41];
  assign data_o[30505] = data_o[41];
  assign data_o[30569] = data_o[41];
  assign data_o[30633] = data_o[41];
  assign data_o[30697] = data_o[41];
  assign data_o[30761] = data_o[41];
  assign data_o[30825] = data_o[41];
  assign data_o[30889] = data_o[41];
  assign data_o[30953] = data_o[41];
  assign data_o[31017] = data_o[41];
  assign data_o[31081] = data_o[41];
  assign data_o[31145] = data_o[41];
  assign data_o[31209] = data_o[41];
  assign data_o[31273] = data_o[41];
  assign data_o[31337] = data_o[41];
  assign data_o[31401] = data_o[41];
  assign data_o[31465] = data_o[41];
  assign data_o[31529] = data_o[41];
  assign data_o[31593] = data_o[41];
  assign data_o[31657] = data_o[41];
  assign data_o[31721] = data_o[41];
  assign data_o[31785] = data_o[41];
  assign data_o[31849] = data_o[41];
  assign data_o[31913] = data_o[41];
  assign data_o[31977] = data_o[41];
  assign data_o[104] = data_o[40];
  assign data_o[168] = data_o[40];
  assign data_o[232] = data_o[40];
  assign data_o[296] = data_o[40];
  assign data_o[360] = data_o[40];
  assign data_o[424] = data_o[40];
  assign data_o[488] = data_o[40];
  assign data_o[552] = data_o[40];
  assign data_o[616] = data_o[40];
  assign data_o[680] = data_o[40];
  assign data_o[744] = data_o[40];
  assign data_o[808] = data_o[40];
  assign data_o[872] = data_o[40];
  assign data_o[936] = data_o[40];
  assign data_o[1000] = data_o[40];
  assign data_o[1064] = data_o[40];
  assign data_o[1128] = data_o[40];
  assign data_o[1192] = data_o[40];
  assign data_o[1256] = data_o[40];
  assign data_o[1320] = data_o[40];
  assign data_o[1384] = data_o[40];
  assign data_o[1448] = data_o[40];
  assign data_o[1512] = data_o[40];
  assign data_o[1576] = data_o[40];
  assign data_o[1640] = data_o[40];
  assign data_o[1704] = data_o[40];
  assign data_o[1768] = data_o[40];
  assign data_o[1832] = data_o[40];
  assign data_o[1896] = data_o[40];
  assign data_o[1960] = data_o[40];
  assign data_o[2024] = data_o[40];
  assign data_o[2088] = data_o[40];
  assign data_o[2152] = data_o[40];
  assign data_o[2216] = data_o[40];
  assign data_o[2280] = data_o[40];
  assign data_o[2344] = data_o[40];
  assign data_o[2408] = data_o[40];
  assign data_o[2472] = data_o[40];
  assign data_o[2536] = data_o[40];
  assign data_o[2600] = data_o[40];
  assign data_o[2664] = data_o[40];
  assign data_o[2728] = data_o[40];
  assign data_o[2792] = data_o[40];
  assign data_o[2856] = data_o[40];
  assign data_o[2920] = data_o[40];
  assign data_o[2984] = data_o[40];
  assign data_o[3048] = data_o[40];
  assign data_o[3112] = data_o[40];
  assign data_o[3176] = data_o[40];
  assign data_o[3240] = data_o[40];
  assign data_o[3304] = data_o[40];
  assign data_o[3368] = data_o[40];
  assign data_o[3432] = data_o[40];
  assign data_o[3496] = data_o[40];
  assign data_o[3560] = data_o[40];
  assign data_o[3624] = data_o[40];
  assign data_o[3688] = data_o[40];
  assign data_o[3752] = data_o[40];
  assign data_o[3816] = data_o[40];
  assign data_o[3880] = data_o[40];
  assign data_o[3944] = data_o[40];
  assign data_o[4008] = data_o[40];
  assign data_o[4072] = data_o[40];
  assign data_o[4136] = data_o[40];
  assign data_o[4200] = data_o[40];
  assign data_o[4264] = data_o[40];
  assign data_o[4328] = data_o[40];
  assign data_o[4392] = data_o[40];
  assign data_o[4456] = data_o[40];
  assign data_o[4520] = data_o[40];
  assign data_o[4584] = data_o[40];
  assign data_o[4648] = data_o[40];
  assign data_o[4712] = data_o[40];
  assign data_o[4776] = data_o[40];
  assign data_o[4840] = data_o[40];
  assign data_o[4904] = data_o[40];
  assign data_o[4968] = data_o[40];
  assign data_o[5032] = data_o[40];
  assign data_o[5096] = data_o[40];
  assign data_o[5160] = data_o[40];
  assign data_o[5224] = data_o[40];
  assign data_o[5288] = data_o[40];
  assign data_o[5352] = data_o[40];
  assign data_o[5416] = data_o[40];
  assign data_o[5480] = data_o[40];
  assign data_o[5544] = data_o[40];
  assign data_o[5608] = data_o[40];
  assign data_o[5672] = data_o[40];
  assign data_o[5736] = data_o[40];
  assign data_o[5800] = data_o[40];
  assign data_o[5864] = data_o[40];
  assign data_o[5928] = data_o[40];
  assign data_o[5992] = data_o[40];
  assign data_o[6056] = data_o[40];
  assign data_o[6120] = data_o[40];
  assign data_o[6184] = data_o[40];
  assign data_o[6248] = data_o[40];
  assign data_o[6312] = data_o[40];
  assign data_o[6376] = data_o[40];
  assign data_o[6440] = data_o[40];
  assign data_o[6504] = data_o[40];
  assign data_o[6568] = data_o[40];
  assign data_o[6632] = data_o[40];
  assign data_o[6696] = data_o[40];
  assign data_o[6760] = data_o[40];
  assign data_o[6824] = data_o[40];
  assign data_o[6888] = data_o[40];
  assign data_o[6952] = data_o[40];
  assign data_o[7016] = data_o[40];
  assign data_o[7080] = data_o[40];
  assign data_o[7144] = data_o[40];
  assign data_o[7208] = data_o[40];
  assign data_o[7272] = data_o[40];
  assign data_o[7336] = data_o[40];
  assign data_o[7400] = data_o[40];
  assign data_o[7464] = data_o[40];
  assign data_o[7528] = data_o[40];
  assign data_o[7592] = data_o[40];
  assign data_o[7656] = data_o[40];
  assign data_o[7720] = data_o[40];
  assign data_o[7784] = data_o[40];
  assign data_o[7848] = data_o[40];
  assign data_o[7912] = data_o[40];
  assign data_o[7976] = data_o[40];
  assign data_o[8040] = data_o[40];
  assign data_o[8104] = data_o[40];
  assign data_o[8168] = data_o[40];
  assign data_o[8232] = data_o[40];
  assign data_o[8296] = data_o[40];
  assign data_o[8360] = data_o[40];
  assign data_o[8424] = data_o[40];
  assign data_o[8488] = data_o[40];
  assign data_o[8552] = data_o[40];
  assign data_o[8616] = data_o[40];
  assign data_o[8680] = data_o[40];
  assign data_o[8744] = data_o[40];
  assign data_o[8808] = data_o[40];
  assign data_o[8872] = data_o[40];
  assign data_o[8936] = data_o[40];
  assign data_o[9000] = data_o[40];
  assign data_o[9064] = data_o[40];
  assign data_o[9128] = data_o[40];
  assign data_o[9192] = data_o[40];
  assign data_o[9256] = data_o[40];
  assign data_o[9320] = data_o[40];
  assign data_o[9384] = data_o[40];
  assign data_o[9448] = data_o[40];
  assign data_o[9512] = data_o[40];
  assign data_o[9576] = data_o[40];
  assign data_o[9640] = data_o[40];
  assign data_o[9704] = data_o[40];
  assign data_o[9768] = data_o[40];
  assign data_o[9832] = data_o[40];
  assign data_o[9896] = data_o[40];
  assign data_o[9960] = data_o[40];
  assign data_o[10024] = data_o[40];
  assign data_o[10088] = data_o[40];
  assign data_o[10152] = data_o[40];
  assign data_o[10216] = data_o[40];
  assign data_o[10280] = data_o[40];
  assign data_o[10344] = data_o[40];
  assign data_o[10408] = data_o[40];
  assign data_o[10472] = data_o[40];
  assign data_o[10536] = data_o[40];
  assign data_o[10600] = data_o[40];
  assign data_o[10664] = data_o[40];
  assign data_o[10728] = data_o[40];
  assign data_o[10792] = data_o[40];
  assign data_o[10856] = data_o[40];
  assign data_o[10920] = data_o[40];
  assign data_o[10984] = data_o[40];
  assign data_o[11048] = data_o[40];
  assign data_o[11112] = data_o[40];
  assign data_o[11176] = data_o[40];
  assign data_o[11240] = data_o[40];
  assign data_o[11304] = data_o[40];
  assign data_o[11368] = data_o[40];
  assign data_o[11432] = data_o[40];
  assign data_o[11496] = data_o[40];
  assign data_o[11560] = data_o[40];
  assign data_o[11624] = data_o[40];
  assign data_o[11688] = data_o[40];
  assign data_o[11752] = data_o[40];
  assign data_o[11816] = data_o[40];
  assign data_o[11880] = data_o[40];
  assign data_o[11944] = data_o[40];
  assign data_o[12008] = data_o[40];
  assign data_o[12072] = data_o[40];
  assign data_o[12136] = data_o[40];
  assign data_o[12200] = data_o[40];
  assign data_o[12264] = data_o[40];
  assign data_o[12328] = data_o[40];
  assign data_o[12392] = data_o[40];
  assign data_o[12456] = data_o[40];
  assign data_o[12520] = data_o[40];
  assign data_o[12584] = data_o[40];
  assign data_o[12648] = data_o[40];
  assign data_o[12712] = data_o[40];
  assign data_o[12776] = data_o[40];
  assign data_o[12840] = data_o[40];
  assign data_o[12904] = data_o[40];
  assign data_o[12968] = data_o[40];
  assign data_o[13032] = data_o[40];
  assign data_o[13096] = data_o[40];
  assign data_o[13160] = data_o[40];
  assign data_o[13224] = data_o[40];
  assign data_o[13288] = data_o[40];
  assign data_o[13352] = data_o[40];
  assign data_o[13416] = data_o[40];
  assign data_o[13480] = data_o[40];
  assign data_o[13544] = data_o[40];
  assign data_o[13608] = data_o[40];
  assign data_o[13672] = data_o[40];
  assign data_o[13736] = data_o[40];
  assign data_o[13800] = data_o[40];
  assign data_o[13864] = data_o[40];
  assign data_o[13928] = data_o[40];
  assign data_o[13992] = data_o[40];
  assign data_o[14056] = data_o[40];
  assign data_o[14120] = data_o[40];
  assign data_o[14184] = data_o[40];
  assign data_o[14248] = data_o[40];
  assign data_o[14312] = data_o[40];
  assign data_o[14376] = data_o[40];
  assign data_o[14440] = data_o[40];
  assign data_o[14504] = data_o[40];
  assign data_o[14568] = data_o[40];
  assign data_o[14632] = data_o[40];
  assign data_o[14696] = data_o[40];
  assign data_o[14760] = data_o[40];
  assign data_o[14824] = data_o[40];
  assign data_o[14888] = data_o[40];
  assign data_o[14952] = data_o[40];
  assign data_o[15016] = data_o[40];
  assign data_o[15080] = data_o[40];
  assign data_o[15144] = data_o[40];
  assign data_o[15208] = data_o[40];
  assign data_o[15272] = data_o[40];
  assign data_o[15336] = data_o[40];
  assign data_o[15400] = data_o[40];
  assign data_o[15464] = data_o[40];
  assign data_o[15528] = data_o[40];
  assign data_o[15592] = data_o[40];
  assign data_o[15656] = data_o[40];
  assign data_o[15720] = data_o[40];
  assign data_o[15784] = data_o[40];
  assign data_o[15848] = data_o[40];
  assign data_o[15912] = data_o[40];
  assign data_o[15976] = data_o[40];
  assign data_o[16040] = data_o[40];
  assign data_o[16104] = data_o[40];
  assign data_o[16168] = data_o[40];
  assign data_o[16232] = data_o[40];
  assign data_o[16296] = data_o[40];
  assign data_o[16360] = data_o[40];
  assign data_o[16424] = data_o[40];
  assign data_o[16488] = data_o[40];
  assign data_o[16552] = data_o[40];
  assign data_o[16616] = data_o[40];
  assign data_o[16680] = data_o[40];
  assign data_o[16744] = data_o[40];
  assign data_o[16808] = data_o[40];
  assign data_o[16872] = data_o[40];
  assign data_o[16936] = data_o[40];
  assign data_o[17000] = data_o[40];
  assign data_o[17064] = data_o[40];
  assign data_o[17128] = data_o[40];
  assign data_o[17192] = data_o[40];
  assign data_o[17256] = data_o[40];
  assign data_o[17320] = data_o[40];
  assign data_o[17384] = data_o[40];
  assign data_o[17448] = data_o[40];
  assign data_o[17512] = data_o[40];
  assign data_o[17576] = data_o[40];
  assign data_o[17640] = data_o[40];
  assign data_o[17704] = data_o[40];
  assign data_o[17768] = data_o[40];
  assign data_o[17832] = data_o[40];
  assign data_o[17896] = data_o[40];
  assign data_o[17960] = data_o[40];
  assign data_o[18024] = data_o[40];
  assign data_o[18088] = data_o[40];
  assign data_o[18152] = data_o[40];
  assign data_o[18216] = data_o[40];
  assign data_o[18280] = data_o[40];
  assign data_o[18344] = data_o[40];
  assign data_o[18408] = data_o[40];
  assign data_o[18472] = data_o[40];
  assign data_o[18536] = data_o[40];
  assign data_o[18600] = data_o[40];
  assign data_o[18664] = data_o[40];
  assign data_o[18728] = data_o[40];
  assign data_o[18792] = data_o[40];
  assign data_o[18856] = data_o[40];
  assign data_o[18920] = data_o[40];
  assign data_o[18984] = data_o[40];
  assign data_o[19048] = data_o[40];
  assign data_o[19112] = data_o[40];
  assign data_o[19176] = data_o[40];
  assign data_o[19240] = data_o[40];
  assign data_o[19304] = data_o[40];
  assign data_o[19368] = data_o[40];
  assign data_o[19432] = data_o[40];
  assign data_o[19496] = data_o[40];
  assign data_o[19560] = data_o[40];
  assign data_o[19624] = data_o[40];
  assign data_o[19688] = data_o[40];
  assign data_o[19752] = data_o[40];
  assign data_o[19816] = data_o[40];
  assign data_o[19880] = data_o[40];
  assign data_o[19944] = data_o[40];
  assign data_o[20008] = data_o[40];
  assign data_o[20072] = data_o[40];
  assign data_o[20136] = data_o[40];
  assign data_o[20200] = data_o[40];
  assign data_o[20264] = data_o[40];
  assign data_o[20328] = data_o[40];
  assign data_o[20392] = data_o[40];
  assign data_o[20456] = data_o[40];
  assign data_o[20520] = data_o[40];
  assign data_o[20584] = data_o[40];
  assign data_o[20648] = data_o[40];
  assign data_o[20712] = data_o[40];
  assign data_o[20776] = data_o[40];
  assign data_o[20840] = data_o[40];
  assign data_o[20904] = data_o[40];
  assign data_o[20968] = data_o[40];
  assign data_o[21032] = data_o[40];
  assign data_o[21096] = data_o[40];
  assign data_o[21160] = data_o[40];
  assign data_o[21224] = data_o[40];
  assign data_o[21288] = data_o[40];
  assign data_o[21352] = data_o[40];
  assign data_o[21416] = data_o[40];
  assign data_o[21480] = data_o[40];
  assign data_o[21544] = data_o[40];
  assign data_o[21608] = data_o[40];
  assign data_o[21672] = data_o[40];
  assign data_o[21736] = data_o[40];
  assign data_o[21800] = data_o[40];
  assign data_o[21864] = data_o[40];
  assign data_o[21928] = data_o[40];
  assign data_o[21992] = data_o[40];
  assign data_o[22056] = data_o[40];
  assign data_o[22120] = data_o[40];
  assign data_o[22184] = data_o[40];
  assign data_o[22248] = data_o[40];
  assign data_o[22312] = data_o[40];
  assign data_o[22376] = data_o[40];
  assign data_o[22440] = data_o[40];
  assign data_o[22504] = data_o[40];
  assign data_o[22568] = data_o[40];
  assign data_o[22632] = data_o[40];
  assign data_o[22696] = data_o[40];
  assign data_o[22760] = data_o[40];
  assign data_o[22824] = data_o[40];
  assign data_o[22888] = data_o[40];
  assign data_o[22952] = data_o[40];
  assign data_o[23016] = data_o[40];
  assign data_o[23080] = data_o[40];
  assign data_o[23144] = data_o[40];
  assign data_o[23208] = data_o[40];
  assign data_o[23272] = data_o[40];
  assign data_o[23336] = data_o[40];
  assign data_o[23400] = data_o[40];
  assign data_o[23464] = data_o[40];
  assign data_o[23528] = data_o[40];
  assign data_o[23592] = data_o[40];
  assign data_o[23656] = data_o[40];
  assign data_o[23720] = data_o[40];
  assign data_o[23784] = data_o[40];
  assign data_o[23848] = data_o[40];
  assign data_o[23912] = data_o[40];
  assign data_o[23976] = data_o[40];
  assign data_o[24040] = data_o[40];
  assign data_o[24104] = data_o[40];
  assign data_o[24168] = data_o[40];
  assign data_o[24232] = data_o[40];
  assign data_o[24296] = data_o[40];
  assign data_o[24360] = data_o[40];
  assign data_o[24424] = data_o[40];
  assign data_o[24488] = data_o[40];
  assign data_o[24552] = data_o[40];
  assign data_o[24616] = data_o[40];
  assign data_o[24680] = data_o[40];
  assign data_o[24744] = data_o[40];
  assign data_o[24808] = data_o[40];
  assign data_o[24872] = data_o[40];
  assign data_o[24936] = data_o[40];
  assign data_o[25000] = data_o[40];
  assign data_o[25064] = data_o[40];
  assign data_o[25128] = data_o[40];
  assign data_o[25192] = data_o[40];
  assign data_o[25256] = data_o[40];
  assign data_o[25320] = data_o[40];
  assign data_o[25384] = data_o[40];
  assign data_o[25448] = data_o[40];
  assign data_o[25512] = data_o[40];
  assign data_o[25576] = data_o[40];
  assign data_o[25640] = data_o[40];
  assign data_o[25704] = data_o[40];
  assign data_o[25768] = data_o[40];
  assign data_o[25832] = data_o[40];
  assign data_o[25896] = data_o[40];
  assign data_o[25960] = data_o[40];
  assign data_o[26024] = data_o[40];
  assign data_o[26088] = data_o[40];
  assign data_o[26152] = data_o[40];
  assign data_o[26216] = data_o[40];
  assign data_o[26280] = data_o[40];
  assign data_o[26344] = data_o[40];
  assign data_o[26408] = data_o[40];
  assign data_o[26472] = data_o[40];
  assign data_o[26536] = data_o[40];
  assign data_o[26600] = data_o[40];
  assign data_o[26664] = data_o[40];
  assign data_o[26728] = data_o[40];
  assign data_o[26792] = data_o[40];
  assign data_o[26856] = data_o[40];
  assign data_o[26920] = data_o[40];
  assign data_o[26984] = data_o[40];
  assign data_o[27048] = data_o[40];
  assign data_o[27112] = data_o[40];
  assign data_o[27176] = data_o[40];
  assign data_o[27240] = data_o[40];
  assign data_o[27304] = data_o[40];
  assign data_o[27368] = data_o[40];
  assign data_o[27432] = data_o[40];
  assign data_o[27496] = data_o[40];
  assign data_o[27560] = data_o[40];
  assign data_o[27624] = data_o[40];
  assign data_o[27688] = data_o[40];
  assign data_o[27752] = data_o[40];
  assign data_o[27816] = data_o[40];
  assign data_o[27880] = data_o[40];
  assign data_o[27944] = data_o[40];
  assign data_o[28008] = data_o[40];
  assign data_o[28072] = data_o[40];
  assign data_o[28136] = data_o[40];
  assign data_o[28200] = data_o[40];
  assign data_o[28264] = data_o[40];
  assign data_o[28328] = data_o[40];
  assign data_o[28392] = data_o[40];
  assign data_o[28456] = data_o[40];
  assign data_o[28520] = data_o[40];
  assign data_o[28584] = data_o[40];
  assign data_o[28648] = data_o[40];
  assign data_o[28712] = data_o[40];
  assign data_o[28776] = data_o[40];
  assign data_o[28840] = data_o[40];
  assign data_o[28904] = data_o[40];
  assign data_o[28968] = data_o[40];
  assign data_o[29032] = data_o[40];
  assign data_o[29096] = data_o[40];
  assign data_o[29160] = data_o[40];
  assign data_o[29224] = data_o[40];
  assign data_o[29288] = data_o[40];
  assign data_o[29352] = data_o[40];
  assign data_o[29416] = data_o[40];
  assign data_o[29480] = data_o[40];
  assign data_o[29544] = data_o[40];
  assign data_o[29608] = data_o[40];
  assign data_o[29672] = data_o[40];
  assign data_o[29736] = data_o[40];
  assign data_o[29800] = data_o[40];
  assign data_o[29864] = data_o[40];
  assign data_o[29928] = data_o[40];
  assign data_o[29992] = data_o[40];
  assign data_o[30056] = data_o[40];
  assign data_o[30120] = data_o[40];
  assign data_o[30184] = data_o[40];
  assign data_o[30248] = data_o[40];
  assign data_o[30312] = data_o[40];
  assign data_o[30376] = data_o[40];
  assign data_o[30440] = data_o[40];
  assign data_o[30504] = data_o[40];
  assign data_o[30568] = data_o[40];
  assign data_o[30632] = data_o[40];
  assign data_o[30696] = data_o[40];
  assign data_o[30760] = data_o[40];
  assign data_o[30824] = data_o[40];
  assign data_o[30888] = data_o[40];
  assign data_o[30952] = data_o[40];
  assign data_o[31016] = data_o[40];
  assign data_o[31080] = data_o[40];
  assign data_o[31144] = data_o[40];
  assign data_o[31208] = data_o[40];
  assign data_o[31272] = data_o[40];
  assign data_o[31336] = data_o[40];
  assign data_o[31400] = data_o[40];
  assign data_o[31464] = data_o[40];
  assign data_o[31528] = data_o[40];
  assign data_o[31592] = data_o[40];
  assign data_o[31656] = data_o[40];
  assign data_o[31720] = data_o[40];
  assign data_o[31784] = data_o[40];
  assign data_o[31848] = data_o[40];
  assign data_o[31912] = data_o[40];
  assign data_o[31976] = data_o[40];
  assign data_o[103] = data_o[39];
  assign data_o[167] = data_o[39];
  assign data_o[231] = data_o[39];
  assign data_o[295] = data_o[39];
  assign data_o[359] = data_o[39];
  assign data_o[423] = data_o[39];
  assign data_o[487] = data_o[39];
  assign data_o[551] = data_o[39];
  assign data_o[615] = data_o[39];
  assign data_o[679] = data_o[39];
  assign data_o[743] = data_o[39];
  assign data_o[807] = data_o[39];
  assign data_o[871] = data_o[39];
  assign data_o[935] = data_o[39];
  assign data_o[999] = data_o[39];
  assign data_o[1063] = data_o[39];
  assign data_o[1127] = data_o[39];
  assign data_o[1191] = data_o[39];
  assign data_o[1255] = data_o[39];
  assign data_o[1319] = data_o[39];
  assign data_o[1383] = data_o[39];
  assign data_o[1447] = data_o[39];
  assign data_o[1511] = data_o[39];
  assign data_o[1575] = data_o[39];
  assign data_o[1639] = data_o[39];
  assign data_o[1703] = data_o[39];
  assign data_o[1767] = data_o[39];
  assign data_o[1831] = data_o[39];
  assign data_o[1895] = data_o[39];
  assign data_o[1959] = data_o[39];
  assign data_o[2023] = data_o[39];
  assign data_o[2087] = data_o[39];
  assign data_o[2151] = data_o[39];
  assign data_o[2215] = data_o[39];
  assign data_o[2279] = data_o[39];
  assign data_o[2343] = data_o[39];
  assign data_o[2407] = data_o[39];
  assign data_o[2471] = data_o[39];
  assign data_o[2535] = data_o[39];
  assign data_o[2599] = data_o[39];
  assign data_o[2663] = data_o[39];
  assign data_o[2727] = data_o[39];
  assign data_o[2791] = data_o[39];
  assign data_o[2855] = data_o[39];
  assign data_o[2919] = data_o[39];
  assign data_o[2983] = data_o[39];
  assign data_o[3047] = data_o[39];
  assign data_o[3111] = data_o[39];
  assign data_o[3175] = data_o[39];
  assign data_o[3239] = data_o[39];
  assign data_o[3303] = data_o[39];
  assign data_o[3367] = data_o[39];
  assign data_o[3431] = data_o[39];
  assign data_o[3495] = data_o[39];
  assign data_o[3559] = data_o[39];
  assign data_o[3623] = data_o[39];
  assign data_o[3687] = data_o[39];
  assign data_o[3751] = data_o[39];
  assign data_o[3815] = data_o[39];
  assign data_o[3879] = data_o[39];
  assign data_o[3943] = data_o[39];
  assign data_o[4007] = data_o[39];
  assign data_o[4071] = data_o[39];
  assign data_o[4135] = data_o[39];
  assign data_o[4199] = data_o[39];
  assign data_o[4263] = data_o[39];
  assign data_o[4327] = data_o[39];
  assign data_o[4391] = data_o[39];
  assign data_o[4455] = data_o[39];
  assign data_o[4519] = data_o[39];
  assign data_o[4583] = data_o[39];
  assign data_o[4647] = data_o[39];
  assign data_o[4711] = data_o[39];
  assign data_o[4775] = data_o[39];
  assign data_o[4839] = data_o[39];
  assign data_o[4903] = data_o[39];
  assign data_o[4967] = data_o[39];
  assign data_o[5031] = data_o[39];
  assign data_o[5095] = data_o[39];
  assign data_o[5159] = data_o[39];
  assign data_o[5223] = data_o[39];
  assign data_o[5287] = data_o[39];
  assign data_o[5351] = data_o[39];
  assign data_o[5415] = data_o[39];
  assign data_o[5479] = data_o[39];
  assign data_o[5543] = data_o[39];
  assign data_o[5607] = data_o[39];
  assign data_o[5671] = data_o[39];
  assign data_o[5735] = data_o[39];
  assign data_o[5799] = data_o[39];
  assign data_o[5863] = data_o[39];
  assign data_o[5927] = data_o[39];
  assign data_o[5991] = data_o[39];
  assign data_o[6055] = data_o[39];
  assign data_o[6119] = data_o[39];
  assign data_o[6183] = data_o[39];
  assign data_o[6247] = data_o[39];
  assign data_o[6311] = data_o[39];
  assign data_o[6375] = data_o[39];
  assign data_o[6439] = data_o[39];
  assign data_o[6503] = data_o[39];
  assign data_o[6567] = data_o[39];
  assign data_o[6631] = data_o[39];
  assign data_o[6695] = data_o[39];
  assign data_o[6759] = data_o[39];
  assign data_o[6823] = data_o[39];
  assign data_o[6887] = data_o[39];
  assign data_o[6951] = data_o[39];
  assign data_o[7015] = data_o[39];
  assign data_o[7079] = data_o[39];
  assign data_o[7143] = data_o[39];
  assign data_o[7207] = data_o[39];
  assign data_o[7271] = data_o[39];
  assign data_o[7335] = data_o[39];
  assign data_o[7399] = data_o[39];
  assign data_o[7463] = data_o[39];
  assign data_o[7527] = data_o[39];
  assign data_o[7591] = data_o[39];
  assign data_o[7655] = data_o[39];
  assign data_o[7719] = data_o[39];
  assign data_o[7783] = data_o[39];
  assign data_o[7847] = data_o[39];
  assign data_o[7911] = data_o[39];
  assign data_o[7975] = data_o[39];
  assign data_o[8039] = data_o[39];
  assign data_o[8103] = data_o[39];
  assign data_o[8167] = data_o[39];
  assign data_o[8231] = data_o[39];
  assign data_o[8295] = data_o[39];
  assign data_o[8359] = data_o[39];
  assign data_o[8423] = data_o[39];
  assign data_o[8487] = data_o[39];
  assign data_o[8551] = data_o[39];
  assign data_o[8615] = data_o[39];
  assign data_o[8679] = data_o[39];
  assign data_o[8743] = data_o[39];
  assign data_o[8807] = data_o[39];
  assign data_o[8871] = data_o[39];
  assign data_o[8935] = data_o[39];
  assign data_o[8999] = data_o[39];
  assign data_o[9063] = data_o[39];
  assign data_o[9127] = data_o[39];
  assign data_o[9191] = data_o[39];
  assign data_o[9255] = data_o[39];
  assign data_o[9319] = data_o[39];
  assign data_o[9383] = data_o[39];
  assign data_o[9447] = data_o[39];
  assign data_o[9511] = data_o[39];
  assign data_o[9575] = data_o[39];
  assign data_o[9639] = data_o[39];
  assign data_o[9703] = data_o[39];
  assign data_o[9767] = data_o[39];
  assign data_o[9831] = data_o[39];
  assign data_o[9895] = data_o[39];
  assign data_o[9959] = data_o[39];
  assign data_o[10023] = data_o[39];
  assign data_o[10087] = data_o[39];
  assign data_o[10151] = data_o[39];
  assign data_o[10215] = data_o[39];
  assign data_o[10279] = data_o[39];
  assign data_o[10343] = data_o[39];
  assign data_o[10407] = data_o[39];
  assign data_o[10471] = data_o[39];
  assign data_o[10535] = data_o[39];
  assign data_o[10599] = data_o[39];
  assign data_o[10663] = data_o[39];
  assign data_o[10727] = data_o[39];
  assign data_o[10791] = data_o[39];
  assign data_o[10855] = data_o[39];
  assign data_o[10919] = data_o[39];
  assign data_o[10983] = data_o[39];
  assign data_o[11047] = data_o[39];
  assign data_o[11111] = data_o[39];
  assign data_o[11175] = data_o[39];
  assign data_o[11239] = data_o[39];
  assign data_o[11303] = data_o[39];
  assign data_o[11367] = data_o[39];
  assign data_o[11431] = data_o[39];
  assign data_o[11495] = data_o[39];
  assign data_o[11559] = data_o[39];
  assign data_o[11623] = data_o[39];
  assign data_o[11687] = data_o[39];
  assign data_o[11751] = data_o[39];
  assign data_o[11815] = data_o[39];
  assign data_o[11879] = data_o[39];
  assign data_o[11943] = data_o[39];
  assign data_o[12007] = data_o[39];
  assign data_o[12071] = data_o[39];
  assign data_o[12135] = data_o[39];
  assign data_o[12199] = data_o[39];
  assign data_o[12263] = data_o[39];
  assign data_o[12327] = data_o[39];
  assign data_o[12391] = data_o[39];
  assign data_o[12455] = data_o[39];
  assign data_o[12519] = data_o[39];
  assign data_o[12583] = data_o[39];
  assign data_o[12647] = data_o[39];
  assign data_o[12711] = data_o[39];
  assign data_o[12775] = data_o[39];
  assign data_o[12839] = data_o[39];
  assign data_o[12903] = data_o[39];
  assign data_o[12967] = data_o[39];
  assign data_o[13031] = data_o[39];
  assign data_o[13095] = data_o[39];
  assign data_o[13159] = data_o[39];
  assign data_o[13223] = data_o[39];
  assign data_o[13287] = data_o[39];
  assign data_o[13351] = data_o[39];
  assign data_o[13415] = data_o[39];
  assign data_o[13479] = data_o[39];
  assign data_o[13543] = data_o[39];
  assign data_o[13607] = data_o[39];
  assign data_o[13671] = data_o[39];
  assign data_o[13735] = data_o[39];
  assign data_o[13799] = data_o[39];
  assign data_o[13863] = data_o[39];
  assign data_o[13927] = data_o[39];
  assign data_o[13991] = data_o[39];
  assign data_o[14055] = data_o[39];
  assign data_o[14119] = data_o[39];
  assign data_o[14183] = data_o[39];
  assign data_o[14247] = data_o[39];
  assign data_o[14311] = data_o[39];
  assign data_o[14375] = data_o[39];
  assign data_o[14439] = data_o[39];
  assign data_o[14503] = data_o[39];
  assign data_o[14567] = data_o[39];
  assign data_o[14631] = data_o[39];
  assign data_o[14695] = data_o[39];
  assign data_o[14759] = data_o[39];
  assign data_o[14823] = data_o[39];
  assign data_o[14887] = data_o[39];
  assign data_o[14951] = data_o[39];
  assign data_o[15015] = data_o[39];
  assign data_o[15079] = data_o[39];
  assign data_o[15143] = data_o[39];
  assign data_o[15207] = data_o[39];
  assign data_o[15271] = data_o[39];
  assign data_o[15335] = data_o[39];
  assign data_o[15399] = data_o[39];
  assign data_o[15463] = data_o[39];
  assign data_o[15527] = data_o[39];
  assign data_o[15591] = data_o[39];
  assign data_o[15655] = data_o[39];
  assign data_o[15719] = data_o[39];
  assign data_o[15783] = data_o[39];
  assign data_o[15847] = data_o[39];
  assign data_o[15911] = data_o[39];
  assign data_o[15975] = data_o[39];
  assign data_o[16039] = data_o[39];
  assign data_o[16103] = data_o[39];
  assign data_o[16167] = data_o[39];
  assign data_o[16231] = data_o[39];
  assign data_o[16295] = data_o[39];
  assign data_o[16359] = data_o[39];
  assign data_o[16423] = data_o[39];
  assign data_o[16487] = data_o[39];
  assign data_o[16551] = data_o[39];
  assign data_o[16615] = data_o[39];
  assign data_o[16679] = data_o[39];
  assign data_o[16743] = data_o[39];
  assign data_o[16807] = data_o[39];
  assign data_o[16871] = data_o[39];
  assign data_o[16935] = data_o[39];
  assign data_o[16999] = data_o[39];
  assign data_o[17063] = data_o[39];
  assign data_o[17127] = data_o[39];
  assign data_o[17191] = data_o[39];
  assign data_o[17255] = data_o[39];
  assign data_o[17319] = data_o[39];
  assign data_o[17383] = data_o[39];
  assign data_o[17447] = data_o[39];
  assign data_o[17511] = data_o[39];
  assign data_o[17575] = data_o[39];
  assign data_o[17639] = data_o[39];
  assign data_o[17703] = data_o[39];
  assign data_o[17767] = data_o[39];
  assign data_o[17831] = data_o[39];
  assign data_o[17895] = data_o[39];
  assign data_o[17959] = data_o[39];
  assign data_o[18023] = data_o[39];
  assign data_o[18087] = data_o[39];
  assign data_o[18151] = data_o[39];
  assign data_o[18215] = data_o[39];
  assign data_o[18279] = data_o[39];
  assign data_o[18343] = data_o[39];
  assign data_o[18407] = data_o[39];
  assign data_o[18471] = data_o[39];
  assign data_o[18535] = data_o[39];
  assign data_o[18599] = data_o[39];
  assign data_o[18663] = data_o[39];
  assign data_o[18727] = data_o[39];
  assign data_o[18791] = data_o[39];
  assign data_o[18855] = data_o[39];
  assign data_o[18919] = data_o[39];
  assign data_o[18983] = data_o[39];
  assign data_o[19047] = data_o[39];
  assign data_o[19111] = data_o[39];
  assign data_o[19175] = data_o[39];
  assign data_o[19239] = data_o[39];
  assign data_o[19303] = data_o[39];
  assign data_o[19367] = data_o[39];
  assign data_o[19431] = data_o[39];
  assign data_o[19495] = data_o[39];
  assign data_o[19559] = data_o[39];
  assign data_o[19623] = data_o[39];
  assign data_o[19687] = data_o[39];
  assign data_o[19751] = data_o[39];
  assign data_o[19815] = data_o[39];
  assign data_o[19879] = data_o[39];
  assign data_o[19943] = data_o[39];
  assign data_o[20007] = data_o[39];
  assign data_o[20071] = data_o[39];
  assign data_o[20135] = data_o[39];
  assign data_o[20199] = data_o[39];
  assign data_o[20263] = data_o[39];
  assign data_o[20327] = data_o[39];
  assign data_o[20391] = data_o[39];
  assign data_o[20455] = data_o[39];
  assign data_o[20519] = data_o[39];
  assign data_o[20583] = data_o[39];
  assign data_o[20647] = data_o[39];
  assign data_o[20711] = data_o[39];
  assign data_o[20775] = data_o[39];
  assign data_o[20839] = data_o[39];
  assign data_o[20903] = data_o[39];
  assign data_o[20967] = data_o[39];
  assign data_o[21031] = data_o[39];
  assign data_o[21095] = data_o[39];
  assign data_o[21159] = data_o[39];
  assign data_o[21223] = data_o[39];
  assign data_o[21287] = data_o[39];
  assign data_o[21351] = data_o[39];
  assign data_o[21415] = data_o[39];
  assign data_o[21479] = data_o[39];
  assign data_o[21543] = data_o[39];
  assign data_o[21607] = data_o[39];
  assign data_o[21671] = data_o[39];
  assign data_o[21735] = data_o[39];
  assign data_o[21799] = data_o[39];
  assign data_o[21863] = data_o[39];
  assign data_o[21927] = data_o[39];
  assign data_o[21991] = data_o[39];
  assign data_o[22055] = data_o[39];
  assign data_o[22119] = data_o[39];
  assign data_o[22183] = data_o[39];
  assign data_o[22247] = data_o[39];
  assign data_o[22311] = data_o[39];
  assign data_o[22375] = data_o[39];
  assign data_o[22439] = data_o[39];
  assign data_o[22503] = data_o[39];
  assign data_o[22567] = data_o[39];
  assign data_o[22631] = data_o[39];
  assign data_o[22695] = data_o[39];
  assign data_o[22759] = data_o[39];
  assign data_o[22823] = data_o[39];
  assign data_o[22887] = data_o[39];
  assign data_o[22951] = data_o[39];
  assign data_o[23015] = data_o[39];
  assign data_o[23079] = data_o[39];
  assign data_o[23143] = data_o[39];
  assign data_o[23207] = data_o[39];
  assign data_o[23271] = data_o[39];
  assign data_o[23335] = data_o[39];
  assign data_o[23399] = data_o[39];
  assign data_o[23463] = data_o[39];
  assign data_o[23527] = data_o[39];
  assign data_o[23591] = data_o[39];
  assign data_o[23655] = data_o[39];
  assign data_o[23719] = data_o[39];
  assign data_o[23783] = data_o[39];
  assign data_o[23847] = data_o[39];
  assign data_o[23911] = data_o[39];
  assign data_o[23975] = data_o[39];
  assign data_o[24039] = data_o[39];
  assign data_o[24103] = data_o[39];
  assign data_o[24167] = data_o[39];
  assign data_o[24231] = data_o[39];
  assign data_o[24295] = data_o[39];
  assign data_o[24359] = data_o[39];
  assign data_o[24423] = data_o[39];
  assign data_o[24487] = data_o[39];
  assign data_o[24551] = data_o[39];
  assign data_o[24615] = data_o[39];
  assign data_o[24679] = data_o[39];
  assign data_o[24743] = data_o[39];
  assign data_o[24807] = data_o[39];
  assign data_o[24871] = data_o[39];
  assign data_o[24935] = data_o[39];
  assign data_o[24999] = data_o[39];
  assign data_o[25063] = data_o[39];
  assign data_o[25127] = data_o[39];
  assign data_o[25191] = data_o[39];
  assign data_o[25255] = data_o[39];
  assign data_o[25319] = data_o[39];
  assign data_o[25383] = data_o[39];
  assign data_o[25447] = data_o[39];
  assign data_o[25511] = data_o[39];
  assign data_o[25575] = data_o[39];
  assign data_o[25639] = data_o[39];
  assign data_o[25703] = data_o[39];
  assign data_o[25767] = data_o[39];
  assign data_o[25831] = data_o[39];
  assign data_o[25895] = data_o[39];
  assign data_o[25959] = data_o[39];
  assign data_o[26023] = data_o[39];
  assign data_o[26087] = data_o[39];
  assign data_o[26151] = data_o[39];
  assign data_o[26215] = data_o[39];
  assign data_o[26279] = data_o[39];
  assign data_o[26343] = data_o[39];
  assign data_o[26407] = data_o[39];
  assign data_o[26471] = data_o[39];
  assign data_o[26535] = data_o[39];
  assign data_o[26599] = data_o[39];
  assign data_o[26663] = data_o[39];
  assign data_o[26727] = data_o[39];
  assign data_o[26791] = data_o[39];
  assign data_o[26855] = data_o[39];
  assign data_o[26919] = data_o[39];
  assign data_o[26983] = data_o[39];
  assign data_o[27047] = data_o[39];
  assign data_o[27111] = data_o[39];
  assign data_o[27175] = data_o[39];
  assign data_o[27239] = data_o[39];
  assign data_o[27303] = data_o[39];
  assign data_o[27367] = data_o[39];
  assign data_o[27431] = data_o[39];
  assign data_o[27495] = data_o[39];
  assign data_o[27559] = data_o[39];
  assign data_o[27623] = data_o[39];
  assign data_o[27687] = data_o[39];
  assign data_o[27751] = data_o[39];
  assign data_o[27815] = data_o[39];
  assign data_o[27879] = data_o[39];
  assign data_o[27943] = data_o[39];
  assign data_o[28007] = data_o[39];
  assign data_o[28071] = data_o[39];
  assign data_o[28135] = data_o[39];
  assign data_o[28199] = data_o[39];
  assign data_o[28263] = data_o[39];
  assign data_o[28327] = data_o[39];
  assign data_o[28391] = data_o[39];
  assign data_o[28455] = data_o[39];
  assign data_o[28519] = data_o[39];
  assign data_o[28583] = data_o[39];
  assign data_o[28647] = data_o[39];
  assign data_o[28711] = data_o[39];
  assign data_o[28775] = data_o[39];
  assign data_o[28839] = data_o[39];
  assign data_o[28903] = data_o[39];
  assign data_o[28967] = data_o[39];
  assign data_o[29031] = data_o[39];
  assign data_o[29095] = data_o[39];
  assign data_o[29159] = data_o[39];
  assign data_o[29223] = data_o[39];
  assign data_o[29287] = data_o[39];
  assign data_o[29351] = data_o[39];
  assign data_o[29415] = data_o[39];
  assign data_o[29479] = data_o[39];
  assign data_o[29543] = data_o[39];
  assign data_o[29607] = data_o[39];
  assign data_o[29671] = data_o[39];
  assign data_o[29735] = data_o[39];
  assign data_o[29799] = data_o[39];
  assign data_o[29863] = data_o[39];
  assign data_o[29927] = data_o[39];
  assign data_o[29991] = data_o[39];
  assign data_o[30055] = data_o[39];
  assign data_o[30119] = data_o[39];
  assign data_o[30183] = data_o[39];
  assign data_o[30247] = data_o[39];
  assign data_o[30311] = data_o[39];
  assign data_o[30375] = data_o[39];
  assign data_o[30439] = data_o[39];
  assign data_o[30503] = data_o[39];
  assign data_o[30567] = data_o[39];
  assign data_o[30631] = data_o[39];
  assign data_o[30695] = data_o[39];
  assign data_o[30759] = data_o[39];
  assign data_o[30823] = data_o[39];
  assign data_o[30887] = data_o[39];
  assign data_o[30951] = data_o[39];
  assign data_o[31015] = data_o[39];
  assign data_o[31079] = data_o[39];
  assign data_o[31143] = data_o[39];
  assign data_o[31207] = data_o[39];
  assign data_o[31271] = data_o[39];
  assign data_o[31335] = data_o[39];
  assign data_o[31399] = data_o[39];
  assign data_o[31463] = data_o[39];
  assign data_o[31527] = data_o[39];
  assign data_o[31591] = data_o[39];
  assign data_o[31655] = data_o[39];
  assign data_o[31719] = data_o[39];
  assign data_o[31783] = data_o[39];
  assign data_o[31847] = data_o[39];
  assign data_o[31911] = data_o[39];
  assign data_o[31975] = data_o[39];
  assign data_o[102] = data_o[38];
  assign data_o[166] = data_o[38];
  assign data_o[230] = data_o[38];
  assign data_o[294] = data_o[38];
  assign data_o[358] = data_o[38];
  assign data_o[422] = data_o[38];
  assign data_o[486] = data_o[38];
  assign data_o[550] = data_o[38];
  assign data_o[614] = data_o[38];
  assign data_o[678] = data_o[38];
  assign data_o[742] = data_o[38];
  assign data_o[806] = data_o[38];
  assign data_o[870] = data_o[38];
  assign data_o[934] = data_o[38];
  assign data_o[998] = data_o[38];
  assign data_o[1062] = data_o[38];
  assign data_o[1126] = data_o[38];
  assign data_o[1190] = data_o[38];
  assign data_o[1254] = data_o[38];
  assign data_o[1318] = data_o[38];
  assign data_o[1382] = data_o[38];
  assign data_o[1446] = data_o[38];
  assign data_o[1510] = data_o[38];
  assign data_o[1574] = data_o[38];
  assign data_o[1638] = data_o[38];
  assign data_o[1702] = data_o[38];
  assign data_o[1766] = data_o[38];
  assign data_o[1830] = data_o[38];
  assign data_o[1894] = data_o[38];
  assign data_o[1958] = data_o[38];
  assign data_o[2022] = data_o[38];
  assign data_o[2086] = data_o[38];
  assign data_o[2150] = data_o[38];
  assign data_o[2214] = data_o[38];
  assign data_o[2278] = data_o[38];
  assign data_o[2342] = data_o[38];
  assign data_o[2406] = data_o[38];
  assign data_o[2470] = data_o[38];
  assign data_o[2534] = data_o[38];
  assign data_o[2598] = data_o[38];
  assign data_o[2662] = data_o[38];
  assign data_o[2726] = data_o[38];
  assign data_o[2790] = data_o[38];
  assign data_o[2854] = data_o[38];
  assign data_o[2918] = data_o[38];
  assign data_o[2982] = data_o[38];
  assign data_o[3046] = data_o[38];
  assign data_o[3110] = data_o[38];
  assign data_o[3174] = data_o[38];
  assign data_o[3238] = data_o[38];
  assign data_o[3302] = data_o[38];
  assign data_o[3366] = data_o[38];
  assign data_o[3430] = data_o[38];
  assign data_o[3494] = data_o[38];
  assign data_o[3558] = data_o[38];
  assign data_o[3622] = data_o[38];
  assign data_o[3686] = data_o[38];
  assign data_o[3750] = data_o[38];
  assign data_o[3814] = data_o[38];
  assign data_o[3878] = data_o[38];
  assign data_o[3942] = data_o[38];
  assign data_o[4006] = data_o[38];
  assign data_o[4070] = data_o[38];
  assign data_o[4134] = data_o[38];
  assign data_o[4198] = data_o[38];
  assign data_o[4262] = data_o[38];
  assign data_o[4326] = data_o[38];
  assign data_o[4390] = data_o[38];
  assign data_o[4454] = data_o[38];
  assign data_o[4518] = data_o[38];
  assign data_o[4582] = data_o[38];
  assign data_o[4646] = data_o[38];
  assign data_o[4710] = data_o[38];
  assign data_o[4774] = data_o[38];
  assign data_o[4838] = data_o[38];
  assign data_o[4902] = data_o[38];
  assign data_o[4966] = data_o[38];
  assign data_o[5030] = data_o[38];
  assign data_o[5094] = data_o[38];
  assign data_o[5158] = data_o[38];
  assign data_o[5222] = data_o[38];
  assign data_o[5286] = data_o[38];
  assign data_o[5350] = data_o[38];
  assign data_o[5414] = data_o[38];
  assign data_o[5478] = data_o[38];
  assign data_o[5542] = data_o[38];
  assign data_o[5606] = data_o[38];
  assign data_o[5670] = data_o[38];
  assign data_o[5734] = data_o[38];
  assign data_o[5798] = data_o[38];
  assign data_o[5862] = data_o[38];
  assign data_o[5926] = data_o[38];
  assign data_o[5990] = data_o[38];
  assign data_o[6054] = data_o[38];
  assign data_o[6118] = data_o[38];
  assign data_o[6182] = data_o[38];
  assign data_o[6246] = data_o[38];
  assign data_o[6310] = data_o[38];
  assign data_o[6374] = data_o[38];
  assign data_o[6438] = data_o[38];
  assign data_o[6502] = data_o[38];
  assign data_o[6566] = data_o[38];
  assign data_o[6630] = data_o[38];
  assign data_o[6694] = data_o[38];
  assign data_o[6758] = data_o[38];
  assign data_o[6822] = data_o[38];
  assign data_o[6886] = data_o[38];
  assign data_o[6950] = data_o[38];
  assign data_o[7014] = data_o[38];
  assign data_o[7078] = data_o[38];
  assign data_o[7142] = data_o[38];
  assign data_o[7206] = data_o[38];
  assign data_o[7270] = data_o[38];
  assign data_o[7334] = data_o[38];
  assign data_o[7398] = data_o[38];
  assign data_o[7462] = data_o[38];
  assign data_o[7526] = data_o[38];
  assign data_o[7590] = data_o[38];
  assign data_o[7654] = data_o[38];
  assign data_o[7718] = data_o[38];
  assign data_o[7782] = data_o[38];
  assign data_o[7846] = data_o[38];
  assign data_o[7910] = data_o[38];
  assign data_o[7974] = data_o[38];
  assign data_o[8038] = data_o[38];
  assign data_o[8102] = data_o[38];
  assign data_o[8166] = data_o[38];
  assign data_o[8230] = data_o[38];
  assign data_o[8294] = data_o[38];
  assign data_o[8358] = data_o[38];
  assign data_o[8422] = data_o[38];
  assign data_o[8486] = data_o[38];
  assign data_o[8550] = data_o[38];
  assign data_o[8614] = data_o[38];
  assign data_o[8678] = data_o[38];
  assign data_o[8742] = data_o[38];
  assign data_o[8806] = data_o[38];
  assign data_o[8870] = data_o[38];
  assign data_o[8934] = data_o[38];
  assign data_o[8998] = data_o[38];
  assign data_o[9062] = data_o[38];
  assign data_o[9126] = data_o[38];
  assign data_o[9190] = data_o[38];
  assign data_o[9254] = data_o[38];
  assign data_o[9318] = data_o[38];
  assign data_o[9382] = data_o[38];
  assign data_o[9446] = data_o[38];
  assign data_o[9510] = data_o[38];
  assign data_o[9574] = data_o[38];
  assign data_o[9638] = data_o[38];
  assign data_o[9702] = data_o[38];
  assign data_o[9766] = data_o[38];
  assign data_o[9830] = data_o[38];
  assign data_o[9894] = data_o[38];
  assign data_o[9958] = data_o[38];
  assign data_o[10022] = data_o[38];
  assign data_o[10086] = data_o[38];
  assign data_o[10150] = data_o[38];
  assign data_o[10214] = data_o[38];
  assign data_o[10278] = data_o[38];
  assign data_o[10342] = data_o[38];
  assign data_o[10406] = data_o[38];
  assign data_o[10470] = data_o[38];
  assign data_o[10534] = data_o[38];
  assign data_o[10598] = data_o[38];
  assign data_o[10662] = data_o[38];
  assign data_o[10726] = data_o[38];
  assign data_o[10790] = data_o[38];
  assign data_o[10854] = data_o[38];
  assign data_o[10918] = data_o[38];
  assign data_o[10982] = data_o[38];
  assign data_o[11046] = data_o[38];
  assign data_o[11110] = data_o[38];
  assign data_o[11174] = data_o[38];
  assign data_o[11238] = data_o[38];
  assign data_o[11302] = data_o[38];
  assign data_o[11366] = data_o[38];
  assign data_o[11430] = data_o[38];
  assign data_o[11494] = data_o[38];
  assign data_o[11558] = data_o[38];
  assign data_o[11622] = data_o[38];
  assign data_o[11686] = data_o[38];
  assign data_o[11750] = data_o[38];
  assign data_o[11814] = data_o[38];
  assign data_o[11878] = data_o[38];
  assign data_o[11942] = data_o[38];
  assign data_o[12006] = data_o[38];
  assign data_o[12070] = data_o[38];
  assign data_o[12134] = data_o[38];
  assign data_o[12198] = data_o[38];
  assign data_o[12262] = data_o[38];
  assign data_o[12326] = data_o[38];
  assign data_o[12390] = data_o[38];
  assign data_o[12454] = data_o[38];
  assign data_o[12518] = data_o[38];
  assign data_o[12582] = data_o[38];
  assign data_o[12646] = data_o[38];
  assign data_o[12710] = data_o[38];
  assign data_o[12774] = data_o[38];
  assign data_o[12838] = data_o[38];
  assign data_o[12902] = data_o[38];
  assign data_o[12966] = data_o[38];
  assign data_o[13030] = data_o[38];
  assign data_o[13094] = data_o[38];
  assign data_o[13158] = data_o[38];
  assign data_o[13222] = data_o[38];
  assign data_o[13286] = data_o[38];
  assign data_o[13350] = data_o[38];
  assign data_o[13414] = data_o[38];
  assign data_o[13478] = data_o[38];
  assign data_o[13542] = data_o[38];
  assign data_o[13606] = data_o[38];
  assign data_o[13670] = data_o[38];
  assign data_o[13734] = data_o[38];
  assign data_o[13798] = data_o[38];
  assign data_o[13862] = data_o[38];
  assign data_o[13926] = data_o[38];
  assign data_o[13990] = data_o[38];
  assign data_o[14054] = data_o[38];
  assign data_o[14118] = data_o[38];
  assign data_o[14182] = data_o[38];
  assign data_o[14246] = data_o[38];
  assign data_o[14310] = data_o[38];
  assign data_o[14374] = data_o[38];
  assign data_o[14438] = data_o[38];
  assign data_o[14502] = data_o[38];
  assign data_o[14566] = data_o[38];
  assign data_o[14630] = data_o[38];
  assign data_o[14694] = data_o[38];
  assign data_o[14758] = data_o[38];
  assign data_o[14822] = data_o[38];
  assign data_o[14886] = data_o[38];
  assign data_o[14950] = data_o[38];
  assign data_o[15014] = data_o[38];
  assign data_o[15078] = data_o[38];
  assign data_o[15142] = data_o[38];
  assign data_o[15206] = data_o[38];
  assign data_o[15270] = data_o[38];
  assign data_o[15334] = data_o[38];
  assign data_o[15398] = data_o[38];
  assign data_o[15462] = data_o[38];
  assign data_o[15526] = data_o[38];
  assign data_o[15590] = data_o[38];
  assign data_o[15654] = data_o[38];
  assign data_o[15718] = data_o[38];
  assign data_o[15782] = data_o[38];
  assign data_o[15846] = data_o[38];
  assign data_o[15910] = data_o[38];
  assign data_o[15974] = data_o[38];
  assign data_o[16038] = data_o[38];
  assign data_o[16102] = data_o[38];
  assign data_o[16166] = data_o[38];
  assign data_o[16230] = data_o[38];
  assign data_o[16294] = data_o[38];
  assign data_o[16358] = data_o[38];
  assign data_o[16422] = data_o[38];
  assign data_o[16486] = data_o[38];
  assign data_o[16550] = data_o[38];
  assign data_o[16614] = data_o[38];
  assign data_o[16678] = data_o[38];
  assign data_o[16742] = data_o[38];
  assign data_o[16806] = data_o[38];
  assign data_o[16870] = data_o[38];
  assign data_o[16934] = data_o[38];
  assign data_o[16998] = data_o[38];
  assign data_o[17062] = data_o[38];
  assign data_o[17126] = data_o[38];
  assign data_o[17190] = data_o[38];
  assign data_o[17254] = data_o[38];
  assign data_o[17318] = data_o[38];
  assign data_o[17382] = data_o[38];
  assign data_o[17446] = data_o[38];
  assign data_o[17510] = data_o[38];
  assign data_o[17574] = data_o[38];
  assign data_o[17638] = data_o[38];
  assign data_o[17702] = data_o[38];
  assign data_o[17766] = data_o[38];
  assign data_o[17830] = data_o[38];
  assign data_o[17894] = data_o[38];
  assign data_o[17958] = data_o[38];
  assign data_o[18022] = data_o[38];
  assign data_o[18086] = data_o[38];
  assign data_o[18150] = data_o[38];
  assign data_o[18214] = data_o[38];
  assign data_o[18278] = data_o[38];
  assign data_o[18342] = data_o[38];
  assign data_o[18406] = data_o[38];
  assign data_o[18470] = data_o[38];
  assign data_o[18534] = data_o[38];
  assign data_o[18598] = data_o[38];
  assign data_o[18662] = data_o[38];
  assign data_o[18726] = data_o[38];
  assign data_o[18790] = data_o[38];
  assign data_o[18854] = data_o[38];
  assign data_o[18918] = data_o[38];
  assign data_o[18982] = data_o[38];
  assign data_o[19046] = data_o[38];
  assign data_o[19110] = data_o[38];
  assign data_o[19174] = data_o[38];
  assign data_o[19238] = data_o[38];
  assign data_o[19302] = data_o[38];
  assign data_o[19366] = data_o[38];
  assign data_o[19430] = data_o[38];
  assign data_o[19494] = data_o[38];
  assign data_o[19558] = data_o[38];
  assign data_o[19622] = data_o[38];
  assign data_o[19686] = data_o[38];
  assign data_o[19750] = data_o[38];
  assign data_o[19814] = data_o[38];
  assign data_o[19878] = data_o[38];
  assign data_o[19942] = data_o[38];
  assign data_o[20006] = data_o[38];
  assign data_o[20070] = data_o[38];
  assign data_o[20134] = data_o[38];
  assign data_o[20198] = data_o[38];
  assign data_o[20262] = data_o[38];
  assign data_o[20326] = data_o[38];
  assign data_o[20390] = data_o[38];
  assign data_o[20454] = data_o[38];
  assign data_o[20518] = data_o[38];
  assign data_o[20582] = data_o[38];
  assign data_o[20646] = data_o[38];
  assign data_o[20710] = data_o[38];
  assign data_o[20774] = data_o[38];
  assign data_o[20838] = data_o[38];
  assign data_o[20902] = data_o[38];
  assign data_o[20966] = data_o[38];
  assign data_o[21030] = data_o[38];
  assign data_o[21094] = data_o[38];
  assign data_o[21158] = data_o[38];
  assign data_o[21222] = data_o[38];
  assign data_o[21286] = data_o[38];
  assign data_o[21350] = data_o[38];
  assign data_o[21414] = data_o[38];
  assign data_o[21478] = data_o[38];
  assign data_o[21542] = data_o[38];
  assign data_o[21606] = data_o[38];
  assign data_o[21670] = data_o[38];
  assign data_o[21734] = data_o[38];
  assign data_o[21798] = data_o[38];
  assign data_o[21862] = data_o[38];
  assign data_o[21926] = data_o[38];
  assign data_o[21990] = data_o[38];
  assign data_o[22054] = data_o[38];
  assign data_o[22118] = data_o[38];
  assign data_o[22182] = data_o[38];
  assign data_o[22246] = data_o[38];
  assign data_o[22310] = data_o[38];
  assign data_o[22374] = data_o[38];
  assign data_o[22438] = data_o[38];
  assign data_o[22502] = data_o[38];
  assign data_o[22566] = data_o[38];
  assign data_o[22630] = data_o[38];
  assign data_o[22694] = data_o[38];
  assign data_o[22758] = data_o[38];
  assign data_o[22822] = data_o[38];
  assign data_o[22886] = data_o[38];
  assign data_o[22950] = data_o[38];
  assign data_o[23014] = data_o[38];
  assign data_o[23078] = data_o[38];
  assign data_o[23142] = data_o[38];
  assign data_o[23206] = data_o[38];
  assign data_o[23270] = data_o[38];
  assign data_o[23334] = data_o[38];
  assign data_o[23398] = data_o[38];
  assign data_o[23462] = data_o[38];
  assign data_o[23526] = data_o[38];
  assign data_o[23590] = data_o[38];
  assign data_o[23654] = data_o[38];
  assign data_o[23718] = data_o[38];
  assign data_o[23782] = data_o[38];
  assign data_o[23846] = data_o[38];
  assign data_o[23910] = data_o[38];
  assign data_o[23974] = data_o[38];
  assign data_o[24038] = data_o[38];
  assign data_o[24102] = data_o[38];
  assign data_o[24166] = data_o[38];
  assign data_o[24230] = data_o[38];
  assign data_o[24294] = data_o[38];
  assign data_o[24358] = data_o[38];
  assign data_o[24422] = data_o[38];
  assign data_o[24486] = data_o[38];
  assign data_o[24550] = data_o[38];
  assign data_o[24614] = data_o[38];
  assign data_o[24678] = data_o[38];
  assign data_o[24742] = data_o[38];
  assign data_o[24806] = data_o[38];
  assign data_o[24870] = data_o[38];
  assign data_o[24934] = data_o[38];
  assign data_o[24998] = data_o[38];
  assign data_o[25062] = data_o[38];
  assign data_o[25126] = data_o[38];
  assign data_o[25190] = data_o[38];
  assign data_o[25254] = data_o[38];
  assign data_o[25318] = data_o[38];
  assign data_o[25382] = data_o[38];
  assign data_o[25446] = data_o[38];
  assign data_o[25510] = data_o[38];
  assign data_o[25574] = data_o[38];
  assign data_o[25638] = data_o[38];
  assign data_o[25702] = data_o[38];
  assign data_o[25766] = data_o[38];
  assign data_o[25830] = data_o[38];
  assign data_o[25894] = data_o[38];
  assign data_o[25958] = data_o[38];
  assign data_o[26022] = data_o[38];
  assign data_o[26086] = data_o[38];
  assign data_o[26150] = data_o[38];
  assign data_o[26214] = data_o[38];
  assign data_o[26278] = data_o[38];
  assign data_o[26342] = data_o[38];
  assign data_o[26406] = data_o[38];
  assign data_o[26470] = data_o[38];
  assign data_o[26534] = data_o[38];
  assign data_o[26598] = data_o[38];
  assign data_o[26662] = data_o[38];
  assign data_o[26726] = data_o[38];
  assign data_o[26790] = data_o[38];
  assign data_o[26854] = data_o[38];
  assign data_o[26918] = data_o[38];
  assign data_o[26982] = data_o[38];
  assign data_o[27046] = data_o[38];
  assign data_o[27110] = data_o[38];
  assign data_o[27174] = data_o[38];
  assign data_o[27238] = data_o[38];
  assign data_o[27302] = data_o[38];
  assign data_o[27366] = data_o[38];
  assign data_o[27430] = data_o[38];
  assign data_o[27494] = data_o[38];
  assign data_o[27558] = data_o[38];
  assign data_o[27622] = data_o[38];
  assign data_o[27686] = data_o[38];
  assign data_o[27750] = data_o[38];
  assign data_o[27814] = data_o[38];
  assign data_o[27878] = data_o[38];
  assign data_o[27942] = data_o[38];
  assign data_o[28006] = data_o[38];
  assign data_o[28070] = data_o[38];
  assign data_o[28134] = data_o[38];
  assign data_o[28198] = data_o[38];
  assign data_o[28262] = data_o[38];
  assign data_o[28326] = data_o[38];
  assign data_o[28390] = data_o[38];
  assign data_o[28454] = data_o[38];
  assign data_o[28518] = data_o[38];
  assign data_o[28582] = data_o[38];
  assign data_o[28646] = data_o[38];
  assign data_o[28710] = data_o[38];
  assign data_o[28774] = data_o[38];
  assign data_o[28838] = data_o[38];
  assign data_o[28902] = data_o[38];
  assign data_o[28966] = data_o[38];
  assign data_o[29030] = data_o[38];
  assign data_o[29094] = data_o[38];
  assign data_o[29158] = data_o[38];
  assign data_o[29222] = data_o[38];
  assign data_o[29286] = data_o[38];
  assign data_o[29350] = data_o[38];
  assign data_o[29414] = data_o[38];
  assign data_o[29478] = data_o[38];
  assign data_o[29542] = data_o[38];
  assign data_o[29606] = data_o[38];
  assign data_o[29670] = data_o[38];
  assign data_o[29734] = data_o[38];
  assign data_o[29798] = data_o[38];
  assign data_o[29862] = data_o[38];
  assign data_o[29926] = data_o[38];
  assign data_o[29990] = data_o[38];
  assign data_o[30054] = data_o[38];
  assign data_o[30118] = data_o[38];
  assign data_o[30182] = data_o[38];
  assign data_o[30246] = data_o[38];
  assign data_o[30310] = data_o[38];
  assign data_o[30374] = data_o[38];
  assign data_o[30438] = data_o[38];
  assign data_o[30502] = data_o[38];
  assign data_o[30566] = data_o[38];
  assign data_o[30630] = data_o[38];
  assign data_o[30694] = data_o[38];
  assign data_o[30758] = data_o[38];
  assign data_o[30822] = data_o[38];
  assign data_o[30886] = data_o[38];
  assign data_o[30950] = data_o[38];
  assign data_o[31014] = data_o[38];
  assign data_o[31078] = data_o[38];
  assign data_o[31142] = data_o[38];
  assign data_o[31206] = data_o[38];
  assign data_o[31270] = data_o[38];
  assign data_o[31334] = data_o[38];
  assign data_o[31398] = data_o[38];
  assign data_o[31462] = data_o[38];
  assign data_o[31526] = data_o[38];
  assign data_o[31590] = data_o[38];
  assign data_o[31654] = data_o[38];
  assign data_o[31718] = data_o[38];
  assign data_o[31782] = data_o[38];
  assign data_o[31846] = data_o[38];
  assign data_o[31910] = data_o[38];
  assign data_o[31974] = data_o[38];
  assign data_o[101] = data_o[37];
  assign data_o[165] = data_o[37];
  assign data_o[229] = data_o[37];
  assign data_o[293] = data_o[37];
  assign data_o[357] = data_o[37];
  assign data_o[421] = data_o[37];
  assign data_o[485] = data_o[37];
  assign data_o[549] = data_o[37];
  assign data_o[613] = data_o[37];
  assign data_o[677] = data_o[37];
  assign data_o[741] = data_o[37];
  assign data_o[805] = data_o[37];
  assign data_o[869] = data_o[37];
  assign data_o[933] = data_o[37];
  assign data_o[997] = data_o[37];
  assign data_o[1061] = data_o[37];
  assign data_o[1125] = data_o[37];
  assign data_o[1189] = data_o[37];
  assign data_o[1253] = data_o[37];
  assign data_o[1317] = data_o[37];
  assign data_o[1381] = data_o[37];
  assign data_o[1445] = data_o[37];
  assign data_o[1509] = data_o[37];
  assign data_o[1573] = data_o[37];
  assign data_o[1637] = data_o[37];
  assign data_o[1701] = data_o[37];
  assign data_o[1765] = data_o[37];
  assign data_o[1829] = data_o[37];
  assign data_o[1893] = data_o[37];
  assign data_o[1957] = data_o[37];
  assign data_o[2021] = data_o[37];
  assign data_o[2085] = data_o[37];
  assign data_o[2149] = data_o[37];
  assign data_o[2213] = data_o[37];
  assign data_o[2277] = data_o[37];
  assign data_o[2341] = data_o[37];
  assign data_o[2405] = data_o[37];
  assign data_o[2469] = data_o[37];
  assign data_o[2533] = data_o[37];
  assign data_o[2597] = data_o[37];
  assign data_o[2661] = data_o[37];
  assign data_o[2725] = data_o[37];
  assign data_o[2789] = data_o[37];
  assign data_o[2853] = data_o[37];
  assign data_o[2917] = data_o[37];
  assign data_o[2981] = data_o[37];
  assign data_o[3045] = data_o[37];
  assign data_o[3109] = data_o[37];
  assign data_o[3173] = data_o[37];
  assign data_o[3237] = data_o[37];
  assign data_o[3301] = data_o[37];
  assign data_o[3365] = data_o[37];
  assign data_o[3429] = data_o[37];
  assign data_o[3493] = data_o[37];
  assign data_o[3557] = data_o[37];
  assign data_o[3621] = data_o[37];
  assign data_o[3685] = data_o[37];
  assign data_o[3749] = data_o[37];
  assign data_o[3813] = data_o[37];
  assign data_o[3877] = data_o[37];
  assign data_o[3941] = data_o[37];
  assign data_o[4005] = data_o[37];
  assign data_o[4069] = data_o[37];
  assign data_o[4133] = data_o[37];
  assign data_o[4197] = data_o[37];
  assign data_o[4261] = data_o[37];
  assign data_o[4325] = data_o[37];
  assign data_o[4389] = data_o[37];
  assign data_o[4453] = data_o[37];
  assign data_o[4517] = data_o[37];
  assign data_o[4581] = data_o[37];
  assign data_o[4645] = data_o[37];
  assign data_o[4709] = data_o[37];
  assign data_o[4773] = data_o[37];
  assign data_o[4837] = data_o[37];
  assign data_o[4901] = data_o[37];
  assign data_o[4965] = data_o[37];
  assign data_o[5029] = data_o[37];
  assign data_o[5093] = data_o[37];
  assign data_o[5157] = data_o[37];
  assign data_o[5221] = data_o[37];
  assign data_o[5285] = data_o[37];
  assign data_o[5349] = data_o[37];
  assign data_o[5413] = data_o[37];
  assign data_o[5477] = data_o[37];
  assign data_o[5541] = data_o[37];
  assign data_o[5605] = data_o[37];
  assign data_o[5669] = data_o[37];
  assign data_o[5733] = data_o[37];
  assign data_o[5797] = data_o[37];
  assign data_o[5861] = data_o[37];
  assign data_o[5925] = data_o[37];
  assign data_o[5989] = data_o[37];
  assign data_o[6053] = data_o[37];
  assign data_o[6117] = data_o[37];
  assign data_o[6181] = data_o[37];
  assign data_o[6245] = data_o[37];
  assign data_o[6309] = data_o[37];
  assign data_o[6373] = data_o[37];
  assign data_o[6437] = data_o[37];
  assign data_o[6501] = data_o[37];
  assign data_o[6565] = data_o[37];
  assign data_o[6629] = data_o[37];
  assign data_o[6693] = data_o[37];
  assign data_o[6757] = data_o[37];
  assign data_o[6821] = data_o[37];
  assign data_o[6885] = data_o[37];
  assign data_o[6949] = data_o[37];
  assign data_o[7013] = data_o[37];
  assign data_o[7077] = data_o[37];
  assign data_o[7141] = data_o[37];
  assign data_o[7205] = data_o[37];
  assign data_o[7269] = data_o[37];
  assign data_o[7333] = data_o[37];
  assign data_o[7397] = data_o[37];
  assign data_o[7461] = data_o[37];
  assign data_o[7525] = data_o[37];
  assign data_o[7589] = data_o[37];
  assign data_o[7653] = data_o[37];
  assign data_o[7717] = data_o[37];
  assign data_o[7781] = data_o[37];
  assign data_o[7845] = data_o[37];
  assign data_o[7909] = data_o[37];
  assign data_o[7973] = data_o[37];
  assign data_o[8037] = data_o[37];
  assign data_o[8101] = data_o[37];
  assign data_o[8165] = data_o[37];
  assign data_o[8229] = data_o[37];
  assign data_o[8293] = data_o[37];
  assign data_o[8357] = data_o[37];
  assign data_o[8421] = data_o[37];
  assign data_o[8485] = data_o[37];
  assign data_o[8549] = data_o[37];
  assign data_o[8613] = data_o[37];
  assign data_o[8677] = data_o[37];
  assign data_o[8741] = data_o[37];
  assign data_o[8805] = data_o[37];
  assign data_o[8869] = data_o[37];
  assign data_o[8933] = data_o[37];
  assign data_o[8997] = data_o[37];
  assign data_o[9061] = data_o[37];
  assign data_o[9125] = data_o[37];
  assign data_o[9189] = data_o[37];
  assign data_o[9253] = data_o[37];
  assign data_o[9317] = data_o[37];
  assign data_o[9381] = data_o[37];
  assign data_o[9445] = data_o[37];
  assign data_o[9509] = data_o[37];
  assign data_o[9573] = data_o[37];
  assign data_o[9637] = data_o[37];
  assign data_o[9701] = data_o[37];
  assign data_o[9765] = data_o[37];
  assign data_o[9829] = data_o[37];
  assign data_o[9893] = data_o[37];
  assign data_o[9957] = data_o[37];
  assign data_o[10021] = data_o[37];
  assign data_o[10085] = data_o[37];
  assign data_o[10149] = data_o[37];
  assign data_o[10213] = data_o[37];
  assign data_o[10277] = data_o[37];
  assign data_o[10341] = data_o[37];
  assign data_o[10405] = data_o[37];
  assign data_o[10469] = data_o[37];
  assign data_o[10533] = data_o[37];
  assign data_o[10597] = data_o[37];
  assign data_o[10661] = data_o[37];
  assign data_o[10725] = data_o[37];
  assign data_o[10789] = data_o[37];
  assign data_o[10853] = data_o[37];
  assign data_o[10917] = data_o[37];
  assign data_o[10981] = data_o[37];
  assign data_o[11045] = data_o[37];
  assign data_o[11109] = data_o[37];
  assign data_o[11173] = data_o[37];
  assign data_o[11237] = data_o[37];
  assign data_o[11301] = data_o[37];
  assign data_o[11365] = data_o[37];
  assign data_o[11429] = data_o[37];
  assign data_o[11493] = data_o[37];
  assign data_o[11557] = data_o[37];
  assign data_o[11621] = data_o[37];
  assign data_o[11685] = data_o[37];
  assign data_o[11749] = data_o[37];
  assign data_o[11813] = data_o[37];
  assign data_o[11877] = data_o[37];
  assign data_o[11941] = data_o[37];
  assign data_o[12005] = data_o[37];
  assign data_o[12069] = data_o[37];
  assign data_o[12133] = data_o[37];
  assign data_o[12197] = data_o[37];
  assign data_o[12261] = data_o[37];
  assign data_o[12325] = data_o[37];
  assign data_o[12389] = data_o[37];
  assign data_o[12453] = data_o[37];
  assign data_o[12517] = data_o[37];
  assign data_o[12581] = data_o[37];
  assign data_o[12645] = data_o[37];
  assign data_o[12709] = data_o[37];
  assign data_o[12773] = data_o[37];
  assign data_o[12837] = data_o[37];
  assign data_o[12901] = data_o[37];
  assign data_o[12965] = data_o[37];
  assign data_o[13029] = data_o[37];
  assign data_o[13093] = data_o[37];
  assign data_o[13157] = data_o[37];
  assign data_o[13221] = data_o[37];
  assign data_o[13285] = data_o[37];
  assign data_o[13349] = data_o[37];
  assign data_o[13413] = data_o[37];
  assign data_o[13477] = data_o[37];
  assign data_o[13541] = data_o[37];
  assign data_o[13605] = data_o[37];
  assign data_o[13669] = data_o[37];
  assign data_o[13733] = data_o[37];
  assign data_o[13797] = data_o[37];
  assign data_o[13861] = data_o[37];
  assign data_o[13925] = data_o[37];
  assign data_o[13989] = data_o[37];
  assign data_o[14053] = data_o[37];
  assign data_o[14117] = data_o[37];
  assign data_o[14181] = data_o[37];
  assign data_o[14245] = data_o[37];
  assign data_o[14309] = data_o[37];
  assign data_o[14373] = data_o[37];
  assign data_o[14437] = data_o[37];
  assign data_o[14501] = data_o[37];
  assign data_o[14565] = data_o[37];
  assign data_o[14629] = data_o[37];
  assign data_o[14693] = data_o[37];
  assign data_o[14757] = data_o[37];
  assign data_o[14821] = data_o[37];
  assign data_o[14885] = data_o[37];
  assign data_o[14949] = data_o[37];
  assign data_o[15013] = data_o[37];
  assign data_o[15077] = data_o[37];
  assign data_o[15141] = data_o[37];
  assign data_o[15205] = data_o[37];
  assign data_o[15269] = data_o[37];
  assign data_o[15333] = data_o[37];
  assign data_o[15397] = data_o[37];
  assign data_o[15461] = data_o[37];
  assign data_o[15525] = data_o[37];
  assign data_o[15589] = data_o[37];
  assign data_o[15653] = data_o[37];
  assign data_o[15717] = data_o[37];
  assign data_o[15781] = data_o[37];
  assign data_o[15845] = data_o[37];
  assign data_o[15909] = data_o[37];
  assign data_o[15973] = data_o[37];
  assign data_o[16037] = data_o[37];
  assign data_o[16101] = data_o[37];
  assign data_o[16165] = data_o[37];
  assign data_o[16229] = data_o[37];
  assign data_o[16293] = data_o[37];
  assign data_o[16357] = data_o[37];
  assign data_o[16421] = data_o[37];
  assign data_o[16485] = data_o[37];
  assign data_o[16549] = data_o[37];
  assign data_o[16613] = data_o[37];
  assign data_o[16677] = data_o[37];
  assign data_o[16741] = data_o[37];
  assign data_o[16805] = data_o[37];
  assign data_o[16869] = data_o[37];
  assign data_o[16933] = data_o[37];
  assign data_o[16997] = data_o[37];
  assign data_o[17061] = data_o[37];
  assign data_o[17125] = data_o[37];
  assign data_o[17189] = data_o[37];
  assign data_o[17253] = data_o[37];
  assign data_o[17317] = data_o[37];
  assign data_o[17381] = data_o[37];
  assign data_o[17445] = data_o[37];
  assign data_o[17509] = data_o[37];
  assign data_o[17573] = data_o[37];
  assign data_o[17637] = data_o[37];
  assign data_o[17701] = data_o[37];
  assign data_o[17765] = data_o[37];
  assign data_o[17829] = data_o[37];
  assign data_o[17893] = data_o[37];
  assign data_o[17957] = data_o[37];
  assign data_o[18021] = data_o[37];
  assign data_o[18085] = data_o[37];
  assign data_o[18149] = data_o[37];
  assign data_o[18213] = data_o[37];
  assign data_o[18277] = data_o[37];
  assign data_o[18341] = data_o[37];
  assign data_o[18405] = data_o[37];
  assign data_o[18469] = data_o[37];
  assign data_o[18533] = data_o[37];
  assign data_o[18597] = data_o[37];
  assign data_o[18661] = data_o[37];
  assign data_o[18725] = data_o[37];
  assign data_o[18789] = data_o[37];
  assign data_o[18853] = data_o[37];
  assign data_o[18917] = data_o[37];
  assign data_o[18981] = data_o[37];
  assign data_o[19045] = data_o[37];
  assign data_o[19109] = data_o[37];
  assign data_o[19173] = data_o[37];
  assign data_o[19237] = data_o[37];
  assign data_o[19301] = data_o[37];
  assign data_o[19365] = data_o[37];
  assign data_o[19429] = data_o[37];
  assign data_o[19493] = data_o[37];
  assign data_o[19557] = data_o[37];
  assign data_o[19621] = data_o[37];
  assign data_o[19685] = data_o[37];
  assign data_o[19749] = data_o[37];
  assign data_o[19813] = data_o[37];
  assign data_o[19877] = data_o[37];
  assign data_o[19941] = data_o[37];
  assign data_o[20005] = data_o[37];
  assign data_o[20069] = data_o[37];
  assign data_o[20133] = data_o[37];
  assign data_o[20197] = data_o[37];
  assign data_o[20261] = data_o[37];
  assign data_o[20325] = data_o[37];
  assign data_o[20389] = data_o[37];
  assign data_o[20453] = data_o[37];
  assign data_o[20517] = data_o[37];
  assign data_o[20581] = data_o[37];
  assign data_o[20645] = data_o[37];
  assign data_o[20709] = data_o[37];
  assign data_o[20773] = data_o[37];
  assign data_o[20837] = data_o[37];
  assign data_o[20901] = data_o[37];
  assign data_o[20965] = data_o[37];
  assign data_o[21029] = data_o[37];
  assign data_o[21093] = data_o[37];
  assign data_o[21157] = data_o[37];
  assign data_o[21221] = data_o[37];
  assign data_o[21285] = data_o[37];
  assign data_o[21349] = data_o[37];
  assign data_o[21413] = data_o[37];
  assign data_o[21477] = data_o[37];
  assign data_o[21541] = data_o[37];
  assign data_o[21605] = data_o[37];
  assign data_o[21669] = data_o[37];
  assign data_o[21733] = data_o[37];
  assign data_o[21797] = data_o[37];
  assign data_o[21861] = data_o[37];
  assign data_o[21925] = data_o[37];
  assign data_o[21989] = data_o[37];
  assign data_o[22053] = data_o[37];
  assign data_o[22117] = data_o[37];
  assign data_o[22181] = data_o[37];
  assign data_o[22245] = data_o[37];
  assign data_o[22309] = data_o[37];
  assign data_o[22373] = data_o[37];
  assign data_o[22437] = data_o[37];
  assign data_o[22501] = data_o[37];
  assign data_o[22565] = data_o[37];
  assign data_o[22629] = data_o[37];
  assign data_o[22693] = data_o[37];
  assign data_o[22757] = data_o[37];
  assign data_o[22821] = data_o[37];
  assign data_o[22885] = data_o[37];
  assign data_o[22949] = data_o[37];
  assign data_o[23013] = data_o[37];
  assign data_o[23077] = data_o[37];
  assign data_o[23141] = data_o[37];
  assign data_o[23205] = data_o[37];
  assign data_o[23269] = data_o[37];
  assign data_o[23333] = data_o[37];
  assign data_o[23397] = data_o[37];
  assign data_o[23461] = data_o[37];
  assign data_o[23525] = data_o[37];
  assign data_o[23589] = data_o[37];
  assign data_o[23653] = data_o[37];
  assign data_o[23717] = data_o[37];
  assign data_o[23781] = data_o[37];
  assign data_o[23845] = data_o[37];
  assign data_o[23909] = data_o[37];
  assign data_o[23973] = data_o[37];
  assign data_o[24037] = data_o[37];
  assign data_o[24101] = data_o[37];
  assign data_o[24165] = data_o[37];
  assign data_o[24229] = data_o[37];
  assign data_o[24293] = data_o[37];
  assign data_o[24357] = data_o[37];
  assign data_o[24421] = data_o[37];
  assign data_o[24485] = data_o[37];
  assign data_o[24549] = data_o[37];
  assign data_o[24613] = data_o[37];
  assign data_o[24677] = data_o[37];
  assign data_o[24741] = data_o[37];
  assign data_o[24805] = data_o[37];
  assign data_o[24869] = data_o[37];
  assign data_o[24933] = data_o[37];
  assign data_o[24997] = data_o[37];
  assign data_o[25061] = data_o[37];
  assign data_o[25125] = data_o[37];
  assign data_o[25189] = data_o[37];
  assign data_o[25253] = data_o[37];
  assign data_o[25317] = data_o[37];
  assign data_o[25381] = data_o[37];
  assign data_o[25445] = data_o[37];
  assign data_o[25509] = data_o[37];
  assign data_o[25573] = data_o[37];
  assign data_o[25637] = data_o[37];
  assign data_o[25701] = data_o[37];
  assign data_o[25765] = data_o[37];
  assign data_o[25829] = data_o[37];
  assign data_o[25893] = data_o[37];
  assign data_o[25957] = data_o[37];
  assign data_o[26021] = data_o[37];
  assign data_o[26085] = data_o[37];
  assign data_o[26149] = data_o[37];
  assign data_o[26213] = data_o[37];
  assign data_o[26277] = data_o[37];
  assign data_o[26341] = data_o[37];
  assign data_o[26405] = data_o[37];
  assign data_o[26469] = data_o[37];
  assign data_o[26533] = data_o[37];
  assign data_o[26597] = data_o[37];
  assign data_o[26661] = data_o[37];
  assign data_o[26725] = data_o[37];
  assign data_o[26789] = data_o[37];
  assign data_o[26853] = data_o[37];
  assign data_o[26917] = data_o[37];
  assign data_o[26981] = data_o[37];
  assign data_o[27045] = data_o[37];
  assign data_o[27109] = data_o[37];
  assign data_o[27173] = data_o[37];
  assign data_o[27237] = data_o[37];
  assign data_o[27301] = data_o[37];
  assign data_o[27365] = data_o[37];
  assign data_o[27429] = data_o[37];
  assign data_o[27493] = data_o[37];
  assign data_o[27557] = data_o[37];
  assign data_o[27621] = data_o[37];
  assign data_o[27685] = data_o[37];
  assign data_o[27749] = data_o[37];
  assign data_o[27813] = data_o[37];
  assign data_o[27877] = data_o[37];
  assign data_o[27941] = data_o[37];
  assign data_o[28005] = data_o[37];
  assign data_o[28069] = data_o[37];
  assign data_o[28133] = data_o[37];
  assign data_o[28197] = data_o[37];
  assign data_o[28261] = data_o[37];
  assign data_o[28325] = data_o[37];
  assign data_o[28389] = data_o[37];
  assign data_o[28453] = data_o[37];
  assign data_o[28517] = data_o[37];
  assign data_o[28581] = data_o[37];
  assign data_o[28645] = data_o[37];
  assign data_o[28709] = data_o[37];
  assign data_o[28773] = data_o[37];
  assign data_o[28837] = data_o[37];
  assign data_o[28901] = data_o[37];
  assign data_o[28965] = data_o[37];
  assign data_o[29029] = data_o[37];
  assign data_o[29093] = data_o[37];
  assign data_o[29157] = data_o[37];
  assign data_o[29221] = data_o[37];
  assign data_o[29285] = data_o[37];
  assign data_o[29349] = data_o[37];
  assign data_o[29413] = data_o[37];
  assign data_o[29477] = data_o[37];
  assign data_o[29541] = data_o[37];
  assign data_o[29605] = data_o[37];
  assign data_o[29669] = data_o[37];
  assign data_o[29733] = data_o[37];
  assign data_o[29797] = data_o[37];
  assign data_o[29861] = data_o[37];
  assign data_o[29925] = data_o[37];
  assign data_o[29989] = data_o[37];
  assign data_o[30053] = data_o[37];
  assign data_o[30117] = data_o[37];
  assign data_o[30181] = data_o[37];
  assign data_o[30245] = data_o[37];
  assign data_o[30309] = data_o[37];
  assign data_o[30373] = data_o[37];
  assign data_o[30437] = data_o[37];
  assign data_o[30501] = data_o[37];
  assign data_o[30565] = data_o[37];
  assign data_o[30629] = data_o[37];
  assign data_o[30693] = data_o[37];
  assign data_o[30757] = data_o[37];
  assign data_o[30821] = data_o[37];
  assign data_o[30885] = data_o[37];
  assign data_o[30949] = data_o[37];
  assign data_o[31013] = data_o[37];
  assign data_o[31077] = data_o[37];
  assign data_o[31141] = data_o[37];
  assign data_o[31205] = data_o[37];
  assign data_o[31269] = data_o[37];
  assign data_o[31333] = data_o[37];
  assign data_o[31397] = data_o[37];
  assign data_o[31461] = data_o[37];
  assign data_o[31525] = data_o[37];
  assign data_o[31589] = data_o[37];
  assign data_o[31653] = data_o[37];
  assign data_o[31717] = data_o[37];
  assign data_o[31781] = data_o[37];
  assign data_o[31845] = data_o[37];
  assign data_o[31909] = data_o[37];
  assign data_o[31973] = data_o[37];
  assign data_o[100] = data_o[36];
  assign data_o[164] = data_o[36];
  assign data_o[228] = data_o[36];
  assign data_o[292] = data_o[36];
  assign data_o[356] = data_o[36];
  assign data_o[420] = data_o[36];
  assign data_o[484] = data_o[36];
  assign data_o[548] = data_o[36];
  assign data_o[612] = data_o[36];
  assign data_o[676] = data_o[36];
  assign data_o[740] = data_o[36];
  assign data_o[804] = data_o[36];
  assign data_o[868] = data_o[36];
  assign data_o[932] = data_o[36];
  assign data_o[996] = data_o[36];
  assign data_o[1060] = data_o[36];
  assign data_o[1124] = data_o[36];
  assign data_o[1188] = data_o[36];
  assign data_o[1252] = data_o[36];
  assign data_o[1316] = data_o[36];
  assign data_o[1380] = data_o[36];
  assign data_o[1444] = data_o[36];
  assign data_o[1508] = data_o[36];
  assign data_o[1572] = data_o[36];
  assign data_o[1636] = data_o[36];
  assign data_o[1700] = data_o[36];
  assign data_o[1764] = data_o[36];
  assign data_o[1828] = data_o[36];
  assign data_o[1892] = data_o[36];
  assign data_o[1956] = data_o[36];
  assign data_o[2020] = data_o[36];
  assign data_o[2084] = data_o[36];
  assign data_o[2148] = data_o[36];
  assign data_o[2212] = data_o[36];
  assign data_o[2276] = data_o[36];
  assign data_o[2340] = data_o[36];
  assign data_o[2404] = data_o[36];
  assign data_o[2468] = data_o[36];
  assign data_o[2532] = data_o[36];
  assign data_o[2596] = data_o[36];
  assign data_o[2660] = data_o[36];
  assign data_o[2724] = data_o[36];
  assign data_o[2788] = data_o[36];
  assign data_o[2852] = data_o[36];
  assign data_o[2916] = data_o[36];
  assign data_o[2980] = data_o[36];
  assign data_o[3044] = data_o[36];
  assign data_o[3108] = data_o[36];
  assign data_o[3172] = data_o[36];
  assign data_o[3236] = data_o[36];
  assign data_o[3300] = data_o[36];
  assign data_o[3364] = data_o[36];
  assign data_o[3428] = data_o[36];
  assign data_o[3492] = data_o[36];
  assign data_o[3556] = data_o[36];
  assign data_o[3620] = data_o[36];
  assign data_o[3684] = data_o[36];
  assign data_o[3748] = data_o[36];
  assign data_o[3812] = data_o[36];
  assign data_o[3876] = data_o[36];
  assign data_o[3940] = data_o[36];
  assign data_o[4004] = data_o[36];
  assign data_o[4068] = data_o[36];
  assign data_o[4132] = data_o[36];
  assign data_o[4196] = data_o[36];
  assign data_o[4260] = data_o[36];
  assign data_o[4324] = data_o[36];
  assign data_o[4388] = data_o[36];
  assign data_o[4452] = data_o[36];
  assign data_o[4516] = data_o[36];
  assign data_o[4580] = data_o[36];
  assign data_o[4644] = data_o[36];
  assign data_o[4708] = data_o[36];
  assign data_o[4772] = data_o[36];
  assign data_o[4836] = data_o[36];
  assign data_o[4900] = data_o[36];
  assign data_o[4964] = data_o[36];
  assign data_o[5028] = data_o[36];
  assign data_o[5092] = data_o[36];
  assign data_o[5156] = data_o[36];
  assign data_o[5220] = data_o[36];
  assign data_o[5284] = data_o[36];
  assign data_o[5348] = data_o[36];
  assign data_o[5412] = data_o[36];
  assign data_o[5476] = data_o[36];
  assign data_o[5540] = data_o[36];
  assign data_o[5604] = data_o[36];
  assign data_o[5668] = data_o[36];
  assign data_o[5732] = data_o[36];
  assign data_o[5796] = data_o[36];
  assign data_o[5860] = data_o[36];
  assign data_o[5924] = data_o[36];
  assign data_o[5988] = data_o[36];
  assign data_o[6052] = data_o[36];
  assign data_o[6116] = data_o[36];
  assign data_o[6180] = data_o[36];
  assign data_o[6244] = data_o[36];
  assign data_o[6308] = data_o[36];
  assign data_o[6372] = data_o[36];
  assign data_o[6436] = data_o[36];
  assign data_o[6500] = data_o[36];
  assign data_o[6564] = data_o[36];
  assign data_o[6628] = data_o[36];
  assign data_o[6692] = data_o[36];
  assign data_o[6756] = data_o[36];
  assign data_o[6820] = data_o[36];
  assign data_o[6884] = data_o[36];
  assign data_o[6948] = data_o[36];
  assign data_o[7012] = data_o[36];
  assign data_o[7076] = data_o[36];
  assign data_o[7140] = data_o[36];
  assign data_o[7204] = data_o[36];
  assign data_o[7268] = data_o[36];
  assign data_o[7332] = data_o[36];
  assign data_o[7396] = data_o[36];
  assign data_o[7460] = data_o[36];
  assign data_o[7524] = data_o[36];
  assign data_o[7588] = data_o[36];
  assign data_o[7652] = data_o[36];
  assign data_o[7716] = data_o[36];
  assign data_o[7780] = data_o[36];
  assign data_o[7844] = data_o[36];
  assign data_o[7908] = data_o[36];
  assign data_o[7972] = data_o[36];
  assign data_o[8036] = data_o[36];
  assign data_o[8100] = data_o[36];
  assign data_o[8164] = data_o[36];
  assign data_o[8228] = data_o[36];
  assign data_o[8292] = data_o[36];
  assign data_o[8356] = data_o[36];
  assign data_o[8420] = data_o[36];
  assign data_o[8484] = data_o[36];
  assign data_o[8548] = data_o[36];
  assign data_o[8612] = data_o[36];
  assign data_o[8676] = data_o[36];
  assign data_o[8740] = data_o[36];
  assign data_o[8804] = data_o[36];
  assign data_o[8868] = data_o[36];
  assign data_o[8932] = data_o[36];
  assign data_o[8996] = data_o[36];
  assign data_o[9060] = data_o[36];
  assign data_o[9124] = data_o[36];
  assign data_o[9188] = data_o[36];
  assign data_o[9252] = data_o[36];
  assign data_o[9316] = data_o[36];
  assign data_o[9380] = data_o[36];
  assign data_o[9444] = data_o[36];
  assign data_o[9508] = data_o[36];
  assign data_o[9572] = data_o[36];
  assign data_o[9636] = data_o[36];
  assign data_o[9700] = data_o[36];
  assign data_o[9764] = data_o[36];
  assign data_o[9828] = data_o[36];
  assign data_o[9892] = data_o[36];
  assign data_o[9956] = data_o[36];
  assign data_o[10020] = data_o[36];
  assign data_o[10084] = data_o[36];
  assign data_o[10148] = data_o[36];
  assign data_o[10212] = data_o[36];
  assign data_o[10276] = data_o[36];
  assign data_o[10340] = data_o[36];
  assign data_o[10404] = data_o[36];
  assign data_o[10468] = data_o[36];
  assign data_o[10532] = data_o[36];
  assign data_o[10596] = data_o[36];
  assign data_o[10660] = data_o[36];
  assign data_o[10724] = data_o[36];
  assign data_o[10788] = data_o[36];
  assign data_o[10852] = data_o[36];
  assign data_o[10916] = data_o[36];
  assign data_o[10980] = data_o[36];
  assign data_o[11044] = data_o[36];
  assign data_o[11108] = data_o[36];
  assign data_o[11172] = data_o[36];
  assign data_o[11236] = data_o[36];
  assign data_o[11300] = data_o[36];
  assign data_o[11364] = data_o[36];
  assign data_o[11428] = data_o[36];
  assign data_o[11492] = data_o[36];
  assign data_o[11556] = data_o[36];
  assign data_o[11620] = data_o[36];
  assign data_o[11684] = data_o[36];
  assign data_o[11748] = data_o[36];
  assign data_o[11812] = data_o[36];
  assign data_o[11876] = data_o[36];
  assign data_o[11940] = data_o[36];
  assign data_o[12004] = data_o[36];
  assign data_o[12068] = data_o[36];
  assign data_o[12132] = data_o[36];
  assign data_o[12196] = data_o[36];
  assign data_o[12260] = data_o[36];
  assign data_o[12324] = data_o[36];
  assign data_o[12388] = data_o[36];
  assign data_o[12452] = data_o[36];
  assign data_o[12516] = data_o[36];
  assign data_o[12580] = data_o[36];
  assign data_o[12644] = data_o[36];
  assign data_o[12708] = data_o[36];
  assign data_o[12772] = data_o[36];
  assign data_o[12836] = data_o[36];
  assign data_o[12900] = data_o[36];
  assign data_o[12964] = data_o[36];
  assign data_o[13028] = data_o[36];
  assign data_o[13092] = data_o[36];
  assign data_o[13156] = data_o[36];
  assign data_o[13220] = data_o[36];
  assign data_o[13284] = data_o[36];
  assign data_o[13348] = data_o[36];
  assign data_o[13412] = data_o[36];
  assign data_o[13476] = data_o[36];
  assign data_o[13540] = data_o[36];
  assign data_o[13604] = data_o[36];
  assign data_o[13668] = data_o[36];
  assign data_o[13732] = data_o[36];
  assign data_o[13796] = data_o[36];
  assign data_o[13860] = data_o[36];
  assign data_o[13924] = data_o[36];
  assign data_o[13988] = data_o[36];
  assign data_o[14052] = data_o[36];
  assign data_o[14116] = data_o[36];
  assign data_o[14180] = data_o[36];
  assign data_o[14244] = data_o[36];
  assign data_o[14308] = data_o[36];
  assign data_o[14372] = data_o[36];
  assign data_o[14436] = data_o[36];
  assign data_o[14500] = data_o[36];
  assign data_o[14564] = data_o[36];
  assign data_o[14628] = data_o[36];
  assign data_o[14692] = data_o[36];
  assign data_o[14756] = data_o[36];
  assign data_o[14820] = data_o[36];
  assign data_o[14884] = data_o[36];
  assign data_o[14948] = data_o[36];
  assign data_o[15012] = data_o[36];
  assign data_o[15076] = data_o[36];
  assign data_o[15140] = data_o[36];
  assign data_o[15204] = data_o[36];
  assign data_o[15268] = data_o[36];
  assign data_o[15332] = data_o[36];
  assign data_o[15396] = data_o[36];
  assign data_o[15460] = data_o[36];
  assign data_o[15524] = data_o[36];
  assign data_o[15588] = data_o[36];
  assign data_o[15652] = data_o[36];
  assign data_o[15716] = data_o[36];
  assign data_o[15780] = data_o[36];
  assign data_o[15844] = data_o[36];
  assign data_o[15908] = data_o[36];
  assign data_o[15972] = data_o[36];
  assign data_o[16036] = data_o[36];
  assign data_o[16100] = data_o[36];
  assign data_o[16164] = data_o[36];
  assign data_o[16228] = data_o[36];
  assign data_o[16292] = data_o[36];
  assign data_o[16356] = data_o[36];
  assign data_o[16420] = data_o[36];
  assign data_o[16484] = data_o[36];
  assign data_o[16548] = data_o[36];
  assign data_o[16612] = data_o[36];
  assign data_o[16676] = data_o[36];
  assign data_o[16740] = data_o[36];
  assign data_o[16804] = data_o[36];
  assign data_o[16868] = data_o[36];
  assign data_o[16932] = data_o[36];
  assign data_o[16996] = data_o[36];
  assign data_o[17060] = data_o[36];
  assign data_o[17124] = data_o[36];
  assign data_o[17188] = data_o[36];
  assign data_o[17252] = data_o[36];
  assign data_o[17316] = data_o[36];
  assign data_o[17380] = data_o[36];
  assign data_o[17444] = data_o[36];
  assign data_o[17508] = data_o[36];
  assign data_o[17572] = data_o[36];
  assign data_o[17636] = data_o[36];
  assign data_o[17700] = data_o[36];
  assign data_o[17764] = data_o[36];
  assign data_o[17828] = data_o[36];
  assign data_o[17892] = data_o[36];
  assign data_o[17956] = data_o[36];
  assign data_o[18020] = data_o[36];
  assign data_o[18084] = data_o[36];
  assign data_o[18148] = data_o[36];
  assign data_o[18212] = data_o[36];
  assign data_o[18276] = data_o[36];
  assign data_o[18340] = data_o[36];
  assign data_o[18404] = data_o[36];
  assign data_o[18468] = data_o[36];
  assign data_o[18532] = data_o[36];
  assign data_o[18596] = data_o[36];
  assign data_o[18660] = data_o[36];
  assign data_o[18724] = data_o[36];
  assign data_o[18788] = data_o[36];
  assign data_o[18852] = data_o[36];
  assign data_o[18916] = data_o[36];
  assign data_o[18980] = data_o[36];
  assign data_o[19044] = data_o[36];
  assign data_o[19108] = data_o[36];
  assign data_o[19172] = data_o[36];
  assign data_o[19236] = data_o[36];
  assign data_o[19300] = data_o[36];
  assign data_o[19364] = data_o[36];
  assign data_o[19428] = data_o[36];
  assign data_o[19492] = data_o[36];
  assign data_o[19556] = data_o[36];
  assign data_o[19620] = data_o[36];
  assign data_o[19684] = data_o[36];
  assign data_o[19748] = data_o[36];
  assign data_o[19812] = data_o[36];
  assign data_o[19876] = data_o[36];
  assign data_o[19940] = data_o[36];
  assign data_o[20004] = data_o[36];
  assign data_o[20068] = data_o[36];
  assign data_o[20132] = data_o[36];
  assign data_o[20196] = data_o[36];
  assign data_o[20260] = data_o[36];
  assign data_o[20324] = data_o[36];
  assign data_o[20388] = data_o[36];
  assign data_o[20452] = data_o[36];
  assign data_o[20516] = data_o[36];
  assign data_o[20580] = data_o[36];
  assign data_o[20644] = data_o[36];
  assign data_o[20708] = data_o[36];
  assign data_o[20772] = data_o[36];
  assign data_o[20836] = data_o[36];
  assign data_o[20900] = data_o[36];
  assign data_o[20964] = data_o[36];
  assign data_o[21028] = data_o[36];
  assign data_o[21092] = data_o[36];
  assign data_o[21156] = data_o[36];
  assign data_o[21220] = data_o[36];
  assign data_o[21284] = data_o[36];
  assign data_o[21348] = data_o[36];
  assign data_o[21412] = data_o[36];
  assign data_o[21476] = data_o[36];
  assign data_o[21540] = data_o[36];
  assign data_o[21604] = data_o[36];
  assign data_o[21668] = data_o[36];
  assign data_o[21732] = data_o[36];
  assign data_o[21796] = data_o[36];
  assign data_o[21860] = data_o[36];
  assign data_o[21924] = data_o[36];
  assign data_o[21988] = data_o[36];
  assign data_o[22052] = data_o[36];
  assign data_o[22116] = data_o[36];
  assign data_o[22180] = data_o[36];
  assign data_o[22244] = data_o[36];
  assign data_o[22308] = data_o[36];
  assign data_o[22372] = data_o[36];
  assign data_o[22436] = data_o[36];
  assign data_o[22500] = data_o[36];
  assign data_o[22564] = data_o[36];
  assign data_o[22628] = data_o[36];
  assign data_o[22692] = data_o[36];
  assign data_o[22756] = data_o[36];
  assign data_o[22820] = data_o[36];
  assign data_o[22884] = data_o[36];
  assign data_o[22948] = data_o[36];
  assign data_o[23012] = data_o[36];
  assign data_o[23076] = data_o[36];
  assign data_o[23140] = data_o[36];
  assign data_o[23204] = data_o[36];
  assign data_o[23268] = data_o[36];
  assign data_o[23332] = data_o[36];
  assign data_o[23396] = data_o[36];
  assign data_o[23460] = data_o[36];
  assign data_o[23524] = data_o[36];
  assign data_o[23588] = data_o[36];
  assign data_o[23652] = data_o[36];
  assign data_o[23716] = data_o[36];
  assign data_o[23780] = data_o[36];
  assign data_o[23844] = data_o[36];
  assign data_o[23908] = data_o[36];
  assign data_o[23972] = data_o[36];
  assign data_o[24036] = data_o[36];
  assign data_o[24100] = data_o[36];
  assign data_o[24164] = data_o[36];
  assign data_o[24228] = data_o[36];
  assign data_o[24292] = data_o[36];
  assign data_o[24356] = data_o[36];
  assign data_o[24420] = data_o[36];
  assign data_o[24484] = data_o[36];
  assign data_o[24548] = data_o[36];
  assign data_o[24612] = data_o[36];
  assign data_o[24676] = data_o[36];
  assign data_o[24740] = data_o[36];
  assign data_o[24804] = data_o[36];
  assign data_o[24868] = data_o[36];
  assign data_o[24932] = data_o[36];
  assign data_o[24996] = data_o[36];
  assign data_o[25060] = data_o[36];
  assign data_o[25124] = data_o[36];
  assign data_o[25188] = data_o[36];
  assign data_o[25252] = data_o[36];
  assign data_o[25316] = data_o[36];
  assign data_o[25380] = data_o[36];
  assign data_o[25444] = data_o[36];
  assign data_o[25508] = data_o[36];
  assign data_o[25572] = data_o[36];
  assign data_o[25636] = data_o[36];
  assign data_o[25700] = data_o[36];
  assign data_o[25764] = data_o[36];
  assign data_o[25828] = data_o[36];
  assign data_o[25892] = data_o[36];
  assign data_o[25956] = data_o[36];
  assign data_o[26020] = data_o[36];
  assign data_o[26084] = data_o[36];
  assign data_o[26148] = data_o[36];
  assign data_o[26212] = data_o[36];
  assign data_o[26276] = data_o[36];
  assign data_o[26340] = data_o[36];
  assign data_o[26404] = data_o[36];
  assign data_o[26468] = data_o[36];
  assign data_o[26532] = data_o[36];
  assign data_o[26596] = data_o[36];
  assign data_o[26660] = data_o[36];
  assign data_o[26724] = data_o[36];
  assign data_o[26788] = data_o[36];
  assign data_o[26852] = data_o[36];
  assign data_o[26916] = data_o[36];
  assign data_o[26980] = data_o[36];
  assign data_o[27044] = data_o[36];
  assign data_o[27108] = data_o[36];
  assign data_o[27172] = data_o[36];
  assign data_o[27236] = data_o[36];
  assign data_o[27300] = data_o[36];
  assign data_o[27364] = data_o[36];
  assign data_o[27428] = data_o[36];
  assign data_o[27492] = data_o[36];
  assign data_o[27556] = data_o[36];
  assign data_o[27620] = data_o[36];
  assign data_o[27684] = data_o[36];
  assign data_o[27748] = data_o[36];
  assign data_o[27812] = data_o[36];
  assign data_o[27876] = data_o[36];
  assign data_o[27940] = data_o[36];
  assign data_o[28004] = data_o[36];
  assign data_o[28068] = data_o[36];
  assign data_o[28132] = data_o[36];
  assign data_o[28196] = data_o[36];
  assign data_o[28260] = data_o[36];
  assign data_o[28324] = data_o[36];
  assign data_o[28388] = data_o[36];
  assign data_o[28452] = data_o[36];
  assign data_o[28516] = data_o[36];
  assign data_o[28580] = data_o[36];
  assign data_o[28644] = data_o[36];
  assign data_o[28708] = data_o[36];
  assign data_o[28772] = data_o[36];
  assign data_o[28836] = data_o[36];
  assign data_o[28900] = data_o[36];
  assign data_o[28964] = data_o[36];
  assign data_o[29028] = data_o[36];
  assign data_o[29092] = data_o[36];
  assign data_o[29156] = data_o[36];
  assign data_o[29220] = data_o[36];
  assign data_o[29284] = data_o[36];
  assign data_o[29348] = data_o[36];
  assign data_o[29412] = data_o[36];
  assign data_o[29476] = data_o[36];
  assign data_o[29540] = data_o[36];
  assign data_o[29604] = data_o[36];
  assign data_o[29668] = data_o[36];
  assign data_o[29732] = data_o[36];
  assign data_o[29796] = data_o[36];
  assign data_o[29860] = data_o[36];
  assign data_o[29924] = data_o[36];
  assign data_o[29988] = data_o[36];
  assign data_o[30052] = data_o[36];
  assign data_o[30116] = data_o[36];
  assign data_o[30180] = data_o[36];
  assign data_o[30244] = data_o[36];
  assign data_o[30308] = data_o[36];
  assign data_o[30372] = data_o[36];
  assign data_o[30436] = data_o[36];
  assign data_o[30500] = data_o[36];
  assign data_o[30564] = data_o[36];
  assign data_o[30628] = data_o[36];
  assign data_o[30692] = data_o[36];
  assign data_o[30756] = data_o[36];
  assign data_o[30820] = data_o[36];
  assign data_o[30884] = data_o[36];
  assign data_o[30948] = data_o[36];
  assign data_o[31012] = data_o[36];
  assign data_o[31076] = data_o[36];
  assign data_o[31140] = data_o[36];
  assign data_o[31204] = data_o[36];
  assign data_o[31268] = data_o[36];
  assign data_o[31332] = data_o[36];
  assign data_o[31396] = data_o[36];
  assign data_o[31460] = data_o[36];
  assign data_o[31524] = data_o[36];
  assign data_o[31588] = data_o[36];
  assign data_o[31652] = data_o[36];
  assign data_o[31716] = data_o[36];
  assign data_o[31780] = data_o[36];
  assign data_o[31844] = data_o[36];
  assign data_o[31908] = data_o[36];
  assign data_o[31972] = data_o[36];
  assign data_o[99] = data_o[35];
  assign data_o[163] = data_o[35];
  assign data_o[227] = data_o[35];
  assign data_o[291] = data_o[35];
  assign data_o[355] = data_o[35];
  assign data_o[419] = data_o[35];
  assign data_o[483] = data_o[35];
  assign data_o[547] = data_o[35];
  assign data_o[611] = data_o[35];
  assign data_o[675] = data_o[35];
  assign data_o[739] = data_o[35];
  assign data_o[803] = data_o[35];
  assign data_o[867] = data_o[35];
  assign data_o[931] = data_o[35];
  assign data_o[995] = data_o[35];
  assign data_o[1059] = data_o[35];
  assign data_o[1123] = data_o[35];
  assign data_o[1187] = data_o[35];
  assign data_o[1251] = data_o[35];
  assign data_o[1315] = data_o[35];
  assign data_o[1379] = data_o[35];
  assign data_o[1443] = data_o[35];
  assign data_o[1507] = data_o[35];
  assign data_o[1571] = data_o[35];
  assign data_o[1635] = data_o[35];
  assign data_o[1699] = data_o[35];
  assign data_o[1763] = data_o[35];
  assign data_o[1827] = data_o[35];
  assign data_o[1891] = data_o[35];
  assign data_o[1955] = data_o[35];
  assign data_o[2019] = data_o[35];
  assign data_o[2083] = data_o[35];
  assign data_o[2147] = data_o[35];
  assign data_o[2211] = data_o[35];
  assign data_o[2275] = data_o[35];
  assign data_o[2339] = data_o[35];
  assign data_o[2403] = data_o[35];
  assign data_o[2467] = data_o[35];
  assign data_o[2531] = data_o[35];
  assign data_o[2595] = data_o[35];
  assign data_o[2659] = data_o[35];
  assign data_o[2723] = data_o[35];
  assign data_o[2787] = data_o[35];
  assign data_o[2851] = data_o[35];
  assign data_o[2915] = data_o[35];
  assign data_o[2979] = data_o[35];
  assign data_o[3043] = data_o[35];
  assign data_o[3107] = data_o[35];
  assign data_o[3171] = data_o[35];
  assign data_o[3235] = data_o[35];
  assign data_o[3299] = data_o[35];
  assign data_o[3363] = data_o[35];
  assign data_o[3427] = data_o[35];
  assign data_o[3491] = data_o[35];
  assign data_o[3555] = data_o[35];
  assign data_o[3619] = data_o[35];
  assign data_o[3683] = data_o[35];
  assign data_o[3747] = data_o[35];
  assign data_o[3811] = data_o[35];
  assign data_o[3875] = data_o[35];
  assign data_o[3939] = data_o[35];
  assign data_o[4003] = data_o[35];
  assign data_o[4067] = data_o[35];
  assign data_o[4131] = data_o[35];
  assign data_o[4195] = data_o[35];
  assign data_o[4259] = data_o[35];
  assign data_o[4323] = data_o[35];
  assign data_o[4387] = data_o[35];
  assign data_o[4451] = data_o[35];
  assign data_o[4515] = data_o[35];
  assign data_o[4579] = data_o[35];
  assign data_o[4643] = data_o[35];
  assign data_o[4707] = data_o[35];
  assign data_o[4771] = data_o[35];
  assign data_o[4835] = data_o[35];
  assign data_o[4899] = data_o[35];
  assign data_o[4963] = data_o[35];
  assign data_o[5027] = data_o[35];
  assign data_o[5091] = data_o[35];
  assign data_o[5155] = data_o[35];
  assign data_o[5219] = data_o[35];
  assign data_o[5283] = data_o[35];
  assign data_o[5347] = data_o[35];
  assign data_o[5411] = data_o[35];
  assign data_o[5475] = data_o[35];
  assign data_o[5539] = data_o[35];
  assign data_o[5603] = data_o[35];
  assign data_o[5667] = data_o[35];
  assign data_o[5731] = data_o[35];
  assign data_o[5795] = data_o[35];
  assign data_o[5859] = data_o[35];
  assign data_o[5923] = data_o[35];
  assign data_o[5987] = data_o[35];
  assign data_o[6051] = data_o[35];
  assign data_o[6115] = data_o[35];
  assign data_o[6179] = data_o[35];
  assign data_o[6243] = data_o[35];
  assign data_o[6307] = data_o[35];
  assign data_o[6371] = data_o[35];
  assign data_o[6435] = data_o[35];
  assign data_o[6499] = data_o[35];
  assign data_o[6563] = data_o[35];
  assign data_o[6627] = data_o[35];
  assign data_o[6691] = data_o[35];
  assign data_o[6755] = data_o[35];
  assign data_o[6819] = data_o[35];
  assign data_o[6883] = data_o[35];
  assign data_o[6947] = data_o[35];
  assign data_o[7011] = data_o[35];
  assign data_o[7075] = data_o[35];
  assign data_o[7139] = data_o[35];
  assign data_o[7203] = data_o[35];
  assign data_o[7267] = data_o[35];
  assign data_o[7331] = data_o[35];
  assign data_o[7395] = data_o[35];
  assign data_o[7459] = data_o[35];
  assign data_o[7523] = data_o[35];
  assign data_o[7587] = data_o[35];
  assign data_o[7651] = data_o[35];
  assign data_o[7715] = data_o[35];
  assign data_o[7779] = data_o[35];
  assign data_o[7843] = data_o[35];
  assign data_o[7907] = data_o[35];
  assign data_o[7971] = data_o[35];
  assign data_o[8035] = data_o[35];
  assign data_o[8099] = data_o[35];
  assign data_o[8163] = data_o[35];
  assign data_o[8227] = data_o[35];
  assign data_o[8291] = data_o[35];
  assign data_o[8355] = data_o[35];
  assign data_o[8419] = data_o[35];
  assign data_o[8483] = data_o[35];
  assign data_o[8547] = data_o[35];
  assign data_o[8611] = data_o[35];
  assign data_o[8675] = data_o[35];
  assign data_o[8739] = data_o[35];
  assign data_o[8803] = data_o[35];
  assign data_o[8867] = data_o[35];
  assign data_o[8931] = data_o[35];
  assign data_o[8995] = data_o[35];
  assign data_o[9059] = data_o[35];
  assign data_o[9123] = data_o[35];
  assign data_o[9187] = data_o[35];
  assign data_o[9251] = data_o[35];
  assign data_o[9315] = data_o[35];
  assign data_o[9379] = data_o[35];
  assign data_o[9443] = data_o[35];
  assign data_o[9507] = data_o[35];
  assign data_o[9571] = data_o[35];
  assign data_o[9635] = data_o[35];
  assign data_o[9699] = data_o[35];
  assign data_o[9763] = data_o[35];
  assign data_o[9827] = data_o[35];
  assign data_o[9891] = data_o[35];
  assign data_o[9955] = data_o[35];
  assign data_o[10019] = data_o[35];
  assign data_o[10083] = data_o[35];
  assign data_o[10147] = data_o[35];
  assign data_o[10211] = data_o[35];
  assign data_o[10275] = data_o[35];
  assign data_o[10339] = data_o[35];
  assign data_o[10403] = data_o[35];
  assign data_o[10467] = data_o[35];
  assign data_o[10531] = data_o[35];
  assign data_o[10595] = data_o[35];
  assign data_o[10659] = data_o[35];
  assign data_o[10723] = data_o[35];
  assign data_o[10787] = data_o[35];
  assign data_o[10851] = data_o[35];
  assign data_o[10915] = data_o[35];
  assign data_o[10979] = data_o[35];
  assign data_o[11043] = data_o[35];
  assign data_o[11107] = data_o[35];
  assign data_o[11171] = data_o[35];
  assign data_o[11235] = data_o[35];
  assign data_o[11299] = data_o[35];
  assign data_o[11363] = data_o[35];
  assign data_o[11427] = data_o[35];
  assign data_o[11491] = data_o[35];
  assign data_o[11555] = data_o[35];
  assign data_o[11619] = data_o[35];
  assign data_o[11683] = data_o[35];
  assign data_o[11747] = data_o[35];
  assign data_o[11811] = data_o[35];
  assign data_o[11875] = data_o[35];
  assign data_o[11939] = data_o[35];
  assign data_o[12003] = data_o[35];
  assign data_o[12067] = data_o[35];
  assign data_o[12131] = data_o[35];
  assign data_o[12195] = data_o[35];
  assign data_o[12259] = data_o[35];
  assign data_o[12323] = data_o[35];
  assign data_o[12387] = data_o[35];
  assign data_o[12451] = data_o[35];
  assign data_o[12515] = data_o[35];
  assign data_o[12579] = data_o[35];
  assign data_o[12643] = data_o[35];
  assign data_o[12707] = data_o[35];
  assign data_o[12771] = data_o[35];
  assign data_o[12835] = data_o[35];
  assign data_o[12899] = data_o[35];
  assign data_o[12963] = data_o[35];
  assign data_o[13027] = data_o[35];
  assign data_o[13091] = data_o[35];
  assign data_o[13155] = data_o[35];
  assign data_o[13219] = data_o[35];
  assign data_o[13283] = data_o[35];
  assign data_o[13347] = data_o[35];
  assign data_o[13411] = data_o[35];
  assign data_o[13475] = data_o[35];
  assign data_o[13539] = data_o[35];
  assign data_o[13603] = data_o[35];
  assign data_o[13667] = data_o[35];
  assign data_o[13731] = data_o[35];
  assign data_o[13795] = data_o[35];
  assign data_o[13859] = data_o[35];
  assign data_o[13923] = data_o[35];
  assign data_o[13987] = data_o[35];
  assign data_o[14051] = data_o[35];
  assign data_o[14115] = data_o[35];
  assign data_o[14179] = data_o[35];
  assign data_o[14243] = data_o[35];
  assign data_o[14307] = data_o[35];
  assign data_o[14371] = data_o[35];
  assign data_o[14435] = data_o[35];
  assign data_o[14499] = data_o[35];
  assign data_o[14563] = data_o[35];
  assign data_o[14627] = data_o[35];
  assign data_o[14691] = data_o[35];
  assign data_o[14755] = data_o[35];
  assign data_o[14819] = data_o[35];
  assign data_o[14883] = data_o[35];
  assign data_o[14947] = data_o[35];
  assign data_o[15011] = data_o[35];
  assign data_o[15075] = data_o[35];
  assign data_o[15139] = data_o[35];
  assign data_o[15203] = data_o[35];
  assign data_o[15267] = data_o[35];
  assign data_o[15331] = data_o[35];
  assign data_o[15395] = data_o[35];
  assign data_o[15459] = data_o[35];
  assign data_o[15523] = data_o[35];
  assign data_o[15587] = data_o[35];
  assign data_o[15651] = data_o[35];
  assign data_o[15715] = data_o[35];
  assign data_o[15779] = data_o[35];
  assign data_o[15843] = data_o[35];
  assign data_o[15907] = data_o[35];
  assign data_o[15971] = data_o[35];
  assign data_o[16035] = data_o[35];
  assign data_o[16099] = data_o[35];
  assign data_o[16163] = data_o[35];
  assign data_o[16227] = data_o[35];
  assign data_o[16291] = data_o[35];
  assign data_o[16355] = data_o[35];
  assign data_o[16419] = data_o[35];
  assign data_o[16483] = data_o[35];
  assign data_o[16547] = data_o[35];
  assign data_o[16611] = data_o[35];
  assign data_o[16675] = data_o[35];
  assign data_o[16739] = data_o[35];
  assign data_o[16803] = data_o[35];
  assign data_o[16867] = data_o[35];
  assign data_o[16931] = data_o[35];
  assign data_o[16995] = data_o[35];
  assign data_o[17059] = data_o[35];
  assign data_o[17123] = data_o[35];
  assign data_o[17187] = data_o[35];
  assign data_o[17251] = data_o[35];
  assign data_o[17315] = data_o[35];
  assign data_o[17379] = data_o[35];
  assign data_o[17443] = data_o[35];
  assign data_o[17507] = data_o[35];
  assign data_o[17571] = data_o[35];
  assign data_o[17635] = data_o[35];
  assign data_o[17699] = data_o[35];
  assign data_o[17763] = data_o[35];
  assign data_o[17827] = data_o[35];
  assign data_o[17891] = data_o[35];
  assign data_o[17955] = data_o[35];
  assign data_o[18019] = data_o[35];
  assign data_o[18083] = data_o[35];
  assign data_o[18147] = data_o[35];
  assign data_o[18211] = data_o[35];
  assign data_o[18275] = data_o[35];
  assign data_o[18339] = data_o[35];
  assign data_o[18403] = data_o[35];
  assign data_o[18467] = data_o[35];
  assign data_o[18531] = data_o[35];
  assign data_o[18595] = data_o[35];
  assign data_o[18659] = data_o[35];
  assign data_o[18723] = data_o[35];
  assign data_o[18787] = data_o[35];
  assign data_o[18851] = data_o[35];
  assign data_o[18915] = data_o[35];
  assign data_o[18979] = data_o[35];
  assign data_o[19043] = data_o[35];
  assign data_o[19107] = data_o[35];
  assign data_o[19171] = data_o[35];
  assign data_o[19235] = data_o[35];
  assign data_o[19299] = data_o[35];
  assign data_o[19363] = data_o[35];
  assign data_o[19427] = data_o[35];
  assign data_o[19491] = data_o[35];
  assign data_o[19555] = data_o[35];
  assign data_o[19619] = data_o[35];
  assign data_o[19683] = data_o[35];
  assign data_o[19747] = data_o[35];
  assign data_o[19811] = data_o[35];
  assign data_o[19875] = data_o[35];
  assign data_o[19939] = data_o[35];
  assign data_o[20003] = data_o[35];
  assign data_o[20067] = data_o[35];
  assign data_o[20131] = data_o[35];
  assign data_o[20195] = data_o[35];
  assign data_o[20259] = data_o[35];
  assign data_o[20323] = data_o[35];
  assign data_o[20387] = data_o[35];
  assign data_o[20451] = data_o[35];
  assign data_o[20515] = data_o[35];
  assign data_o[20579] = data_o[35];
  assign data_o[20643] = data_o[35];
  assign data_o[20707] = data_o[35];
  assign data_o[20771] = data_o[35];
  assign data_o[20835] = data_o[35];
  assign data_o[20899] = data_o[35];
  assign data_o[20963] = data_o[35];
  assign data_o[21027] = data_o[35];
  assign data_o[21091] = data_o[35];
  assign data_o[21155] = data_o[35];
  assign data_o[21219] = data_o[35];
  assign data_o[21283] = data_o[35];
  assign data_o[21347] = data_o[35];
  assign data_o[21411] = data_o[35];
  assign data_o[21475] = data_o[35];
  assign data_o[21539] = data_o[35];
  assign data_o[21603] = data_o[35];
  assign data_o[21667] = data_o[35];
  assign data_o[21731] = data_o[35];
  assign data_o[21795] = data_o[35];
  assign data_o[21859] = data_o[35];
  assign data_o[21923] = data_o[35];
  assign data_o[21987] = data_o[35];
  assign data_o[22051] = data_o[35];
  assign data_o[22115] = data_o[35];
  assign data_o[22179] = data_o[35];
  assign data_o[22243] = data_o[35];
  assign data_o[22307] = data_o[35];
  assign data_o[22371] = data_o[35];
  assign data_o[22435] = data_o[35];
  assign data_o[22499] = data_o[35];
  assign data_o[22563] = data_o[35];
  assign data_o[22627] = data_o[35];
  assign data_o[22691] = data_o[35];
  assign data_o[22755] = data_o[35];
  assign data_o[22819] = data_o[35];
  assign data_o[22883] = data_o[35];
  assign data_o[22947] = data_o[35];
  assign data_o[23011] = data_o[35];
  assign data_o[23075] = data_o[35];
  assign data_o[23139] = data_o[35];
  assign data_o[23203] = data_o[35];
  assign data_o[23267] = data_o[35];
  assign data_o[23331] = data_o[35];
  assign data_o[23395] = data_o[35];
  assign data_o[23459] = data_o[35];
  assign data_o[23523] = data_o[35];
  assign data_o[23587] = data_o[35];
  assign data_o[23651] = data_o[35];
  assign data_o[23715] = data_o[35];
  assign data_o[23779] = data_o[35];
  assign data_o[23843] = data_o[35];
  assign data_o[23907] = data_o[35];
  assign data_o[23971] = data_o[35];
  assign data_o[24035] = data_o[35];
  assign data_o[24099] = data_o[35];
  assign data_o[24163] = data_o[35];
  assign data_o[24227] = data_o[35];
  assign data_o[24291] = data_o[35];
  assign data_o[24355] = data_o[35];
  assign data_o[24419] = data_o[35];
  assign data_o[24483] = data_o[35];
  assign data_o[24547] = data_o[35];
  assign data_o[24611] = data_o[35];
  assign data_o[24675] = data_o[35];
  assign data_o[24739] = data_o[35];
  assign data_o[24803] = data_o[35];
  assign data_o[24867] = data_o[35];
  assign data_o[24931] = data_o[35];
  assign data_o[24995] = data_o[35];
  assign data_o[25059] = data_o[35];
  assign data_o[25123] = data_o[35];
  assign data_o[25187] = data_o[35];
  assign data_o[25251] = data_o[35];
  assign data_o[25315] = data_o[35];
  assign data_o[25379] = data_o[35];
  assign data_o[25443] = data_o[35];
  assign data_o[25507] = data_o[35];
  assign data_o[25571] = data_o[35];
  assign data_o[25635] = data_o[35];
  assign data_o[25699] = data_o[35];
  assign data_o[25763] = data_o[35];
  assign data_o[25827] = data_o[35];
  assign data_o[25891] = data_o[35];
  assign data_o[25955] = data_o[35];
  assign data_o[26019] = data_o[35];
  assign data_o[26083] = data_o[35];
  assign data_o[26147] = data_o[35];
  assign data_o[26211] = data_o[35];
  assign data_o[26275] = data_o[35];
  assign data_o[26339] = data_o[35];
  assign data_o[26403] = data_o[35];
  assign data_o[26467] = data_o[35];
  assign data_o[26531] = data_o[35];
  assign data_o[26595] = data_o[35];
  assign data_o[26659] = data_o[35];
  assign data_o[26723] = data_o[35];
  assign data_o[26787] = data_o[35];
  assign data_o[26851] = data_o[35];
  assign data_o[26915] = data_o[35];
  assign data_o[26979] = data_o[35];
  assign data_o[27043] = data_o[35];
  assign data_o[27107] = data_o[35];
  assign data_o[27171] = data_o[35];
  assign data_o[27235] = data_o[35];
  assign data_o[27299] = data_o[35];
  assign data_o[27363] = data_o[35];
  assign data_o[27427] = data_o[35];
  assign data_o[27491] = data_o[35];
  assign data_o[27555] = data_o[35];
  assign data_o[27619] = data_o[35];
  assign data_o[27683] = data_o[35];
  assign data_o[27747] = data_o[35];
  assign data_o[27811] = data_o[35];
  assign data_o[27875] = data_o[35];
  assign data_o[27939] = data_o[35];
  assign data_o[28003] = data_o[35];
  assign data_o[28067] = data_o[35];
  assign data_o[28131] = data_o[35];
  assign data_o[28195] = data_o[35];
  assign data_o[28259] = data_o[35];
  assign data_o[28323] = data_o[35];
  assign data_o[28387] = data_o[35];
  assign data_o[28451] = data_o[35];
  assign data_o[28515] = data_o[35];
  assign data_o[28579] = data_o[35];
  assign data_o[28643] = data_o[35];
  assign data_o[28707] = data_o[35];
  assign data_o[28771] = data_o[35];
  assign data_o[28835] = data_o[35];
  assign data_o[28899] = data_o[35];
  assign data_o[28963] = data_o[35];
  assign data_o[29027] = data_o[35];
  assign data_o[29091] = data_o[35];
  assign data_o[29155] = data_o[35];
  assign data_o[29219] = data_o[35];
  assign data_o[29283] = data_o[35];
  assign data_o[29347] = data_o[35];
  assign data_o[29411] = data_o[35];
  assign data_o[29475] = data_o[35];
  assign data_o[29539] = data_o[35];
  assign data_o[29603] = data_o[35];
  assign data_o[29667] = data_o[35];
  assign data_o[29731] = data_o[35];
  assign data_o[29795] = data_o[35];
  assign data_o[29859] = data_o[35];
  assign data_o[29923] = data_o[35];
  assign data_o[29987] = data_o[35];
  assign data_o[30051] = data_o[35];
  assign data_o[30115] = data_o[35];
  assign data_o[30179] = data_o[35];
  assign data_o[30243] = data_o[35];
  assign data_o[30307] = data_o[35];
  assign data_o[30371] = data_o[35];
  assign data_o[30435] = data_o[35];
  assign data_o[30499] = data_o[35];
  assign data_o[30563] = data_o[35];
  assign data_o[30627] = data_o[35];
  assign data_o[30691] = data_o[35];
  assign data_o[30755] = data_o[35];
  assign data_o[30819] = data_o[35];
  assign data_o[30883] = data_o[35];
  assign data_o[30947] = data_o[35];
  assign data_o[31011] = data_o[35];
  assign data_o[31075] = data_o[35];
  assign data_o[31139] = data_o[35];
  assign data_o[31203] = data_o[35];
  assign data_o[31267] = data_o[35];
  assign data_o[31331] = data_o[35];
  assign data_o[31395] = data_o[35];
  assign data_o[31459] = data_o[35];
  assign data_o[31523] = data_o[35];
  assign data_o[31587] = data_o[35];
  assign data_o[31651] = data_o[35];
  assign data_o[31715] = data_o[35];
  assign data_o[31779] = data_o[35];
  assign data_o[31843] = data_o[35];
  assign data_o[31907] = data_o[35];
  assign data_o[31971] = data_o[35];
  assign data_o[98] = data_o[34];
  assign data_o[162] = data_o[34];
  assign data_o[226] = data_o[34];
  assign data_o[290] = data_o[34];
  assign data_o[354] = data_o[34];
  assign data_o[418] = data_o[34];
  assign data_o[482] = data_o[34];
  assign data_o[546] = data_o[34];
  assign data_o[610] = data_o[34];
  assign data_o[674] = data_o[34];
  assign data_o[738] = data_o[34];
  assign data_o[802] = data_o[34];
  assign data_o[866] = data_o[34];
  assign data_o[930] = data_o[34];
  assign data_o[994] = data_o[34];
  assign data_o[1058] = data_o[34];
  assign data_o[1122] = data_o[34];
  assign data_o[1186] = data_o[34];
  assign data_o[1250] = data_o[34];
  assign data_o[1314] = data_o[34];
  assign data_o[1378] = data_o[34];
  assign data_o[1442] = data_o[34];
  assign data_o[1506] = data_o[34];
  assign data_o[1570] = data_o[34];
  assign data_o[1634] = data_o[34];
  assign data_o[1698] = data_o[34];
  assign data_o[1762] = data_o[34];
  assign data_o[1826] = data_o[34];
  assign data_o[1890] = data_o[34];
  assign data_o[1954] = data_o[34];
  assign data_o[2018] = data_o[34];
  assign data_o[2082] = data_o[34];
  assign data_o[2146] = data_o[34];
  assign data_o[2210] = data_o[34];
  assign data_o[2274] = data_o[34];
  assign data_o[2338] = data_o[34];
  assign data_o[2402] = data_o[34];
  assign data_o[2466] = data_o[34];
  assign data_o[2530] = data_o[34];
  assign data_o[2594] = data_o[34];
  assign data_o[2658] = data_o[34];
  assign data_o[2722] = data_o[34];
  assign data_o[2786] = data_o[34];
  assign data_o[2850] = data_o[34];
  assign data_o[2914] = data_o[34];
  assign data_o[2978] = data_o[34];
  assign data_o[3042] = data_o[34];
  assign data_o[3106] = data_o[34];
  assign data_o[3170] = data_o[34];
  assign data_o[3234] = data_o[34];
  assign data_o[3298] = data_o[34];
  assign data_o[3362] = data_o[34];
  assign data_o[3426] = data_o[34];
  assign data_o[3490] = data_o[34];
  assign data_o[3554] = data_o[34];
  assign data_o[3618] = data_o[34];
  assign data_o[3682] = data_o[34];
  assign data_o[3746] = data_o[34];
  assign data_o[3810] = data_o[34];
  assign data_o[3874] = data_o[34];
  assign data_o[3938] = data_o[34];
  assign data_o[4002] = data_o[34];
  assign data_o[4066] = data_o[34];
  assign data_o[4130] = data_o[34];
  assign data_o[4194] = data_o[34];
  assign data_o[4258] = data_o[34];
  assign data_o[4322] = data_o[34];
  assign data_o[4386] = data_o[34];
  assign data_o[4450] = data_o[34];
  assign data_o[4514] = data_o[34];
  assign data_o[4578] = data_o[34];
  assign data_o[4642] = data_o[34];
  assign data_o[4706] = data_o[34];
  assign data_o[4770] = data_o[34];
  assign data_o[4834] = data_o[34];
  assign data_o[4898] = data_o[34];
  assign data_o[4962] = data_o[34];
  assign data_o[5026] = data_o[34];
  assign data_o[5090] = data_o[34];
  assign data_o[5154] = data_o[34];
  assign data_o[5218] = data_o[34];
  assign data_o[5282] = data_o[34];
  assign data_o[5346] = data_o[34];
  assign data_o[5410] = data_o[34];
  assign data_o[5474] = data_o[34];
  assign data_o[5538] = data_o[34];
  assign data_o[5602] = data_o[34];
  assign data_o[5666] = data_o[34];
  assign data_o[5730] = data_o[34];
  assign data_o[5794] = data_o[34];
  assign data_o[5858] = data_o[34];
  assign data_o[5922] = data_o[34];
  assign data_o[5986] = data_o[34];
  assign data_o[6050] = data_o[34];
  assign data_o[6114] = data_o[34];
  assign data_o[6178] = data_o[34];
  assign data_o[6242] = data_o[34];
  assign data_o[6306] = data_o[34];
  assign data_o[6370] = data_o[34];
  assign data_o[6434] = data_o[34];
  assign data_o[6498] = data_o[34];
  assign data_o[6562] = data_o[34];
  assign data_o[6626] = data_o[34];
  assign data_o[6690] = data_o[34];
  assign data_o[6754] = data_o[34];
  assign data_o[6818] = data_o[34];
  assign data_o[6882] = data_o[34];
  assign data_o[6946] = data_o[34];
  assign data_o[7010] = data_o[34];
  assign data_o[7074] = data_o[34];
  assign data_o[7138] = data_o[34];
  assign data_o[7202] = data_o[34];
  assign data_o[7266] = data_o[34];
  assign data_o[7330] = data_o[34];
  assign data_o[7394] = data_o[34];
  assign data_o[7458] = data_o[34];
  assign data_o[7522] = data_o[34];
  assign data_o[7586] = data_o[34];
  assign data_o[7650] = data_o[34];
  assign data_o[7714] = data_o[34];
  assign data_o[7778] = data_o[34];
  assign data_o[7842] = data_o[34];
  assign data_o[7906] = data_o[34];
  assign data_o[7970] = data_o[34];
  assign data_o[8034] = data_o[34];
  assign data_o[8098] = data_o[34];
  assign data_o[8162] = data_o[34];
  assign data_o[8226] = data_o[34];
  assign data_o[8290] = data_o[34];
  assign data_o[8354] = data_o[34];
  assign data_o[8418] = data_o[34];
  assign data_o[8482] = data_o[34];
  assign data_o[8546] = data_o[34];
  assign data_o[8610] = data_o[34];
  assign data_o[8674] = data_o[34];
  assign data_o[8738] = data_o[34];
  assign data_o[8802] = data_o[34];
  assign data_o[8866] = data_o[34];
  assign data_o[8930] = data_o[34];
  assign data_o[8994] = data_o[34];
  assign data_o[9058] = data_o[34];
  assign data_o[9122] = data_o[34];
  assign data_o[9186] = data_o[34];
  assign data_o[9250] = data_o[34];
  assign data_o[9314] = data_o[34];
  assign data_o[9378] = data_o[34];
  assign data_o[9442] = data_o[34];
  assign data_o[9506] = data_o[34];
  assign data_o[9570] = data_o[34];
  assign data_o[9634] = data_o[34];
  assign data_o[9698] = data_o[34];
  assign data_o[9762] = data_o[34];
  assign data_o[9826] = data_o[34];
  assign data_o[9890] = data_o[34];
  assign data_o[9954] = data_o[34];
  assign data_o[10018] = data_o[34];
  assign data_o[10082] = data_o[34];
  assign data_o[10146] = data_o[34];
  assign data_o[10210] = data_o[34];
  assign data_o[10274] = data_o[34];
  assign data_o[10338] = data_o[34];
  assign data_o[10402] = data_o[34];
  assign data_o[10466] = data_o[34];
  assign data_o[10530] = data_o[34];
  assign data_o[10594] = data_o[34];
  assign data_o[10658] = data_o[34];
  assign data_o[10722] = data_o[34];
  assign data_o[10786] = data_o[34];
  assign data_o[10850] = data_o[34];
  assign data_o[10914] = data_o[34];
  assign data_o[10978] = data_o[34];
  assign data_o[11042] = data_o[34];
  assign data_o[11106] = data_o[34];
  assign data_o[11170] = data_o[34];
  assign data_o[11234] = data_o[34];
  assign data_o[11298] = data_o[34];
  assign data_o[11362] = data_o[34];
  assign data_o[11426] = data_o[34];
  assign data_o[11490] = data_o[34];
  assign data_o[11554] = data_o[34];
  assign data_o[11618] = data_o[34];
  assign data_o[11682] = data_o[34];
  assign data_o[11746] = data_o[34];
  assign data_o[11810] = data_o[34];
  assign data_o[11874] = data_o[34];
  assign data_o[11938] = data_o[34];
  assign data_o[12002] = data_o[34];
  assign data_o[12066] = data_o[34];
  assign data_o[12130] = data_o[34];
  assign data_o[12194] = data_o[34];
  assign data_o[12258] = data_o[34];
  assign data_o[12322] = data_o[34];
  assign data_o[12386] = data_o[34];
  assign data_o[12450] = data_o[34];
  assign data_o[12514] = data_o[34];
  assign data_o[12578] = data_o[34];
  assign data_o[12642] = data_o[34];
  assign data_o[12706] = data_o[34];
  assign data_o[12770] = data_o[34];
  assign data_o[12834] = data_o[34];
  assign data_o[12898] = data_o[34];
  assign data_o[12962] = data_o[34];
  assign data_o[13026] = data_o[34];
  assign data_o[13090] = data_o[34];
  assign data_o[13154] = data_o[34];
  assign data_o[13218] = data_o[34];
  assign data_o[13282] = data_o[34];
  assign data_o[13346] = data_o[34];
  assign data_o[13410] = data_o[34];
  assign data_o[13474] = data_o[34];
  assign data_o[13538] = data_o[34];
  assign data_o[13602] = data_o[34];
  assign data_o[13666] = data_o[34];
  assign data_o[13730] = data_o[34];
  assign data_o[13794] = data_o[34];
  assign data_o[13858] = data_o[34];
  assign data_o[13922] = data_o[34];
  assign data_o[13986] = data_o[34];
  assign data_o[14050] = data_o[34];
  assign data_o[14114] = data_o[34];
  assign data_o[14178] = data_o[34];
  assign data_o[14242] = data_o[34];
  assign data_o[14306] = data_o[34];
  assign data_o[14370] = data_o[34];
  assign data_o[14434] = data_o[34];
  assign data_o[14498] = data_o[34];
  assign data_o[14562] = data_o[34];
  assign data_o[14626] = data_o[34];
  assign data_o[14690] = data_o[34];
  assign data_o[14754] = data_o[34];
  assign data_o[14818] = data_o[34];
  assign data_o[14882] = data_o[34];
  assign data_o[14946] = data_o[34];
  assign data_o[15010] = data_o[34];
  assign data_o[15074] = data_o[34];
  assign data_o[15138] = data_o[34];
  assign data_o[15202] = data_o[34];
  assign data_o[15266] = data_o[34];
  assign data_o[15330] = data_o[34];
  assign data_o[15394] = data_o[34];
  assign data_o[15458] = data_o[34];
  assign data_o[15522] = data_o[34];
  assign data_o[15586] = data_o[34];
  assign data_o[15650] = data_o[34];
  assign data_o[15714] = data_o[34];
  assign data_o[15778] = data_o[34];
  assign data_o[15842] = data_o[34];
  assign data_o[15906] = data_o[34];
  assign data_o[15970] = data_o[34];
  assign data_o[16034] = data_o[34];
  assign data_o[16098] = data_o[34];
  assign data_o[16162] = data_o[34];
  assign data_o[16226] = data_o[34];
  assign data_o[16290] = data_o[34];
  assign data_o[16354] = data_o[34];
  assign data_o[16418] = data_o[34];
  assign data_o[16482] = data_o[34];
  assign data_o[16546] = data_o[34];
  assign data_o[16610] = data_o[34];
  assign data_o[16674] = data_o[34];
  assign data_o[16738] = data_o[34];
  assign data_o[16802] = data_o[34];
  assign data_o[16866] = data_o[34];
  assign data_o[16930] = data_o[34];
  assign data_o[16994] = data_o[34];
  assign data_o[17058] = data_o[34];
  assign data_o[17122] = data_o[34];
  assign data_o[17186] = data_o[34];
  assign data_o[17250] = data_o[34];
  assign data_o[17314] = data_o[34];
  assign data_o[17378] = data_o[34];
  assign data_o[17442] = data_o[34];
  assign data_o[17506] = data_o[34];
  assign data_o[17570] = data_o[34];
  assign data_o[17634] = data_o[34];
  assign data_o[17698] = data_o[34];
  assign data_o[17762] = data_o[34];
  assign data_o[17826] = data_o[34];
  assign data_o[17890] = data_o[34];
  assign data_o[17954] = data_o[34];
  assign data_o[18018] = data_o[34];
  assign data_o[18082] = data_o[34];
  assign data_o[18146] = data_o[34];
  assign data_o[18210] = data_o[34];
  assign data_o[18274] = data_o[34];
  assign data_o[18338] = data_o[34];
  assign data_o[18402] = data_o[34];
  assign data_o[18466] = data_o[34];
  assign data_o[18530] = data_o[34];
  assign data_o[18594] = data_o[34];
  assign data_o[18658] = data_o[34];
  assign data_o[18722] = data_o[34];
  assign data_o[18786] = data_o[34];
  assign data_o[18850] = data_o[34];
  assign data_o[18914] = data_o[34];
  assign data_o[18978] = data_o[34];
  assign data_o[19042] = data_o[34];
  assign data_o[19106] = data_o[34];
  assign data_o[19170] = data_o[34];
  assign data_o[19234] = data_o[34];
  assign data_o[19298] = data_o[34];
  assign data_o[19362] = data_o[34];
  assign data_o[19426] = data_o[34];
  assign data_o[19490] = data_o[34];
  assign data_o[19554] = data_o[34];
  assign data_o[19618] = data_o[34];
  assign data_o[19682] = data_o[34];
  assign data_o[19746] = data_o[34];
  assign data_o[19810] = data_o[34];
  assign data_o[19874] = data_o[34];
  assign data_o[19938] = data_o[34];
  assign data_o[20002] = data_o[34];
  assign data_o[20066] = data_o[34];
  assign data_o[20130] = data_o[34];
  assign data_o[20194] = data_o[34];
  assign data_o[20258] = data_o[34];
  assign data_o[20322] = data_o[34];
  assign data_o[20386] = data_o[34];
  assign data_o[20450] = data_o[34];
  assign data_o[20514] = data_o[34];
  assign data_o[20578] = data_o[34];
  assign data_o[20642] = data_o[34];
  assign data_o[20706] = data_o[34];
  assign data_o[20770] = data_o[34];
  assign data_o[20834] = data_o[34];
  assign data_o[20898] = data_o[34];
  assign data_o[20962] = data_o[34];
  assign data_o[21026] = data_o[34];
  assign data_o[21090] = data_o[34];
  assign data_o[21154] = data_o[34];
  assign data_o[21218] = data_o[34];
  assign data_o[21282] = data_o[34];
  assign data_o[21346] = data_o[34];
  assign data_o[21410] = data_o[34];
  assign data_o[21474] = data_o[34];
  assign data_o[21538] = data_o[34];
  assign data_o[21602] = data_o[34];
  assign data_o[21666] = data_o[34];
  assign data_o[21730] = data_o[34];
  assign data_o[21794] = data_o[34];
  assign data_o[21858] = data_o[34];
  assign data_o[21922] = data_o[34];
  assign data_o[21986] = data_o[34];
  assign data_o[22050] = data_o[34];
  assign data_o[22114] = data_o[34];
  assign data_o[22178] = data_o[34];
  assign data_o[22242] = data_o[34];
  assign data_o[22306] = data_o[34];
  assign data_o[22370] = data_o[34];
  assign data_o[22434] = data_o[34];
  assign data_o[22498] = data_o[34];
  assign data_o[22562] = data_o[34];
  assign data_o[22626] = data_o[34];
  assign data_o[22690] = data_o[34];
  assign data_o[22754] = data_o[34];
  assign data_o[22818] = data_o[34];
  assign data_o[22882] = data_o[34];
  assign data_o[22946] = data_o[34];
  assign data_o[23010] = data_o[34];
  assign data_o[23074] = data_o[34];
  assign data_o[23138] = data_o[34];
  assign data_o[23202] = data_o[34];
  assign data_o[23266] = data_o[34];
  assign data_o[23330] = data_o[34];
  assign data_o[23394] = data_o[34];
  assign data_o[23458] = data_o[34];
  assign data_o[23522] = data_o[34];
  assign data_o[23586] = data_o[34];
  assign data_o[23650] = data_o[34];
  assign data_o[23714] = data_o[34];
  assign data_o[23778] = data_o[34];
  assign data_o[23842] = data_o[34];
  assign data_o[23906] = data_o[34];
  assign data_o[23970] = data_o[34];
  assign data_o[24034] = data_o[34];
  assign data_o[24098] = data_o[34];
  assign data_o[24162] = data_o[34];
  assign data_o[24226] = data_o[34];
  assign data_o[24290] = data_o[34];
  assign data_o[24354] = data_o[34];
  assign data_o[24418] = data_o[34];
  assign data_o[24482] = data_o[34];
  assign data_o[24546] = data_o[34];
  assign data_o[24610] = data_o[34];
  assign data_o[24674] = data_o[34];
  assign data_o[24738] = data_o[34];
  assign data_o[24802] = data_o[34];
  assign data_o[24866] = data_o[34];
  assign data_o[24930] = data_o[34];
  assign data_o[24994] = data_o[34];
  assign data_o[25058] = data_o[34];
  assign data_o[25122] = data_o[34];
  assign data_o[25186] = data_o[34];
  assign data_o[25250] = data_o[34];
  assign data_o[25314] = data_o[34];
  assign data_o[25378] = data_o[34];
  assign data_o[25442] = data_o[34];
  assign data_o[25506] = data_o[34];
  assign data_o[25570] = data_o[34];
  assign data_o[25634] = data_o[34];
  assign data_o[25698] = data_o[34];
  assign data_o[25762] = data_o[34];
  assign data_o[25826] = data_o[34];
  assign data_o[25890] = data_o[34];
  assign data_o[25954] = data_o[34];
  assign data_o[26018] = data_o[34];
  assign data_o[26082] = data_o[34];
  assign data_o[26146] = data_o[34];
  assign data_o[26210] = data_o[34];
  assign data_o[26274] = data_o[34];
  assign data_o[26338] = data_o[34];
  assign data_o[26402] = data_o[34];
  assign data_o[26466] = data_o[34];
  assign data_o[26530] = data_o[34];
  assign data_o[26594] = data_o[34];
  assign data_o[26658] = data_o[34];
  assign data_o[26722] = data_o[34];
  assign data_o[26786] = data_o[34];
  assign data_o[26850] = data_o[34];
  assign data_o[26914] = data_o[34];
  assign data_o[26978] = data_o[34];
  assign data_o[27042] = data_o[34];
  assign data_o[27106] = data_o[34];
  assign data_o[27170] = data_o[34];
  assign data_o[27234] = data_o[34];
  assign data_o[27298] = data_o[34];
  assign data_o[27362] = data_o[34];
  assign data_o[27426] = data_o[34];
  assign data_o[27490] = data_o[34];
  assign data_o[27554] = data_o[34];
  assign data_o[27618] = data_o[34];
  assign data_o[27682] = data_o[34];
  assign data_o[27746] = data_o[34];
  assign data_o[27810] = data_o[34];
  assign data_o[27874] = data_o[34];
  assign data_o[27938] = data_o[34];
  assign data_o[28002] = data_o[34];
  assign data_o[28066] = data_o[34];
  assign data_o[28130] = data_o[34];
  assign data_o[28194] = data_o[34];
  assign data_o[28258] = data_o[34];
  assign data_o[28322] = data_o[34];
  assign data_o[28386] = data_o[34];
  assign data_o[28450] = data_o[34];
  assign data_o[28514] = data_o[34];
  assign data_o[28578] = data_o[34];
  assign data_o[28642] = data_o[34];
  assign data_o[28706] = data_o[34];
  assign data_o[28770] = data_o[34];
  assign data_o[28834] = data_o[34];
  assign data_o[28898] = data_o[34];
  assign data_o[28962] = data_o[34];
  assign data_o[29026] = data_o[34];
  assign data_o[29090] = data_o[34];
  assign data_o[29154] = data_o[34];
  assign data_o[29218] = data_o[34];
  assign data_o[29282] = data_o[34];
  assign data_o[29346] = data_o[34];
  assign data_o[29410] = data_o[34];
  assign data_o[29474] = data_o[34];
  assign data_o[29538] = data_o[34];
  assign data_o[29602] = data_o[34];
  assign data_o[29666] = data_o[34];
  assign data_o[29730] = data_o[34];
  assign data_o[29794] = data_o[34];
  assign data_o[29858] = data_o[34];
  assign data_o[29922] = data_o[34];
  assign data_o[29986] = data_o[34];
  assign data_o[30050] = data_o[34];
  assign data_o[30114] = data_o[34];
  assign data_o[30178] = data_o[34];
  assign data_o[30242] = data_o[34];
  assign data_o[30306] = data_o[34];
  assign data_o[30370] = data_o[34];
  assign data_o[30434] = data_o[34];
  assign data_o[30498] = data_o[34];
  assign data_o[30562] = data_o[34];
  assign data_o[30626] = data_o[34];
  assign data_o[30690] = data_o[34];
  assign data_o[30754] = data_o[34];
  assign data_o[30818] = data_o[34];
  assign data_o[30882] = data_o[34];
  assign data_o[30946] = data_o[34];
  assign data_o[31010] = data_o[34];
  assign data_o[31074] = data_o[34];
  assign data_o[31138] = data_o[34];
  assign data_o[31202] = data_o[34];
  assign data_o[31266] = data_o[34];
  assign data_o[31330] = data_o[34];
  assign data_o[31394] = data_o[34];
  assign data_o[31458] = data_o[34];
  assign data_o[31522] = data_o[34];
  assign data_o[31586] = data_o[34];
  assign data_o[31650] = data_o[34];
  assign data_o[31714] = data_o[34];
  assign data_o[31778] = data_o[34];
  assign data_o[31842] = data_o[34];
  assign data_o[31906] = data_o[34];
  assign data_o[31970] = data_o[34];
  assign data_o[97] = data_o[33];
  assign data_o[161] = data_o[33];
  assign data_o[225] = data_o[33];
  assign data_o[289] = data_o[33];
  assign data_o[353] = data_o[33];
  assign data_o[417] = data_o[33];
  assign data_o[481] = data_o[33];
  assign data_o[545] = data_o[33];
  assign data_o[609] = data_o[33];
  assign data_o[673] = data_o[33];
  assign data_o[737] = data_o[33];
  assign data_o[801] = data_o[33];
  assign data_o[865] = data_o[33];
  assign data_o[929] = data_o[33];
  assign data_o[993] = data_o[33];
  assign data_o[1057] = data_o[33];
  assign data_o[1121] = data_o[33];
  assign data_o[1185] = data_o[33];
  assign data_o[1249] = data_o[33];
  assign data_o[1313] = data_o[33];
  assign data_o[1377] = data_o[33];
  assign data_o[1441] = data_o[33];
  assign data_o[1505] = data_o[33];
  assign data_o[1569] = data_o[33];
  assign data_o[1633] = data_o[33];
  assign data_o[1697] = data_o[33];
  assign data_o[1761] = data_o[33];
  assign data_o[1825] = data_o[33];
  assign data_o[1889] = data_o[33];
  assign data_o[1953] = data_o[33];
  assign data_o[2017] = data_o[33];
  assign data_o[2081] = data_o[33];
  assign data_o[2145] = data_o[33];
  assign data_o[2209] = data_o[33];
  assign data_o[2273] = data_o[33];
  assign data_o[2337] = data_o[33];
  assign data_o[2401] = data_o[33];
  assign data_o[2465] = data_o[33];
  assign data_o[2529] = data_o[33];
  assign data_o[2593] = data_o[33];
  assign data_o[2657] = data_o[33];
  assign data_o[2721] = data_o[33];
  assign data_o[2785] = data_o[33];
  assign data_o[2849] = data_o[33];
  assign data_o[2913] = data_o[33];
  assign data_o[2977] = data_o[33];
  assign data_o[3041] = data_o[33];
  assign data_o[3105] = data_o[33];
  assign data_o[3169] = data_o[33];
  assign data_o[3233] = data_o[33];
  assign data_o[3297] = data_o[33];
  assign data_o[3361] = data_o[33];
  assign data_o[3425] = data_o[33];
  assign data_o[3489] = data_o[33];
  assign data_o[3553] = data_o[33];
  assign data_o[3617] = data_o[33];
  assign data_o[3681] = data_o[33];
  assign data_o[3745] = data_o[33];
  assign data_o[3809] = data_o[33];
  assign data_o[3873] = data_o[33];
  assign data_o[3937] = data_o[33];
  assign data_o[4001] = data_o[33];
  assign data_o[4065] = data_o[33];
  assign data_o[4129] = data_o[33];
  assign data_o[4193] = data_o[33];
  assign data_o[4257] = data_o[33];
  assign data_o[4321] = data_o[33];
  assign data_o[4385] = data_o[33];
  assign data_o[4449] = data_o[33];
  assign data_o[4513] = data_o[33];
  assign data_o[4577] = data_o[33];
  assign data_o[4641] = data_o[33];
  assign data_o[4705] = data_o[33];
  assign data_o[4769] = data_o[33];
  assign data_o[4833] = data_o[33];
  assign data_o[4897] = data_o[33];
  assign data_o[4961] = data_o[33];
  assign data_o[5025] = data_o[33];
  assign data_o[5089] = data_o[33];
  assign data_o[5153] = data_o[33];
  assign data_o[5217] = data_o[33];
  assign data_o[5281] = data_o[33];
  assign data_o[5345] = data_o[33];
  assign data_o[5409] = data_o[33];
  assign data_o[5473] = data_o[33];
  assign data_o[5537] = data_o[33];
  assign data_o[5601] = data_o[33];
  assign data_o[5665] = data_o[33];
  assign data_o[5729] = data_o[33];
  assign data_o[5793] = data_o[33];
  assign data_o[5857] = data_o[33];
  assign data_o[5921] = data_o[33];
  assign data_o[5985] = data_o[33];
  assign data_o[6049] = data_o[33];
  assign data_o[6113] = data_o[33];
  assign data_o[6177] = data_o[33];
  assign data_o[6241] = data_o[33];
  assign data_o[6305] = data_o[33];
  assign data_o[6369] = data_o[33];
  assign data_o[6433] = data_o[33];
  assign data_o[6497] = data_o[33];
  assign data_o[6561] = data_o[33];
  assign data_o[6625] = data_o[33];
  assign data_o[6689] = data_o[33];
  assign data_o[6753] = data_o[33];
  assign data_o[6817] = data_o[33];
  assign data_o[6881] = data_o[33];
  assign data_o[6945] = data_o[33];
  assign data_o[7009] = data_o[33];
  assign data_o[7073] = data_o[33];
  assign data_o[7137] = data_o[33];
  assign data_o[7201] = data_o[33];
  assign data_o[7265] = data_o[33];
  assign data_o[7329] = data_o[33];
  assign data_o[7393] = data_o[33];
  assign data_o[7457] = data_o[33];
  assign data_o[7521] = data_o[33];
  assign data_o[7585] = data_o[33];
  assign data_o[7649] = data_o[33];
  assign data_o[7713] = data_o[33];
  assign data_o[7777] = data_o[33];
  assign data_o[7841] = data_o[33];
  assign data_o[7905] = data_o[33];
  assign data_o[7969] = data_o[33];
  assign data_o[8033] = data_o[33];
  assign data_o[8097] = data_o[33];
  assign data_o[8161] = data_o[33];
  assign data_o[8225] = data_o[33];
  assign data_o[8289] = data_o[33];
  assign data_o[8353] = data_o[33];
  assign data_o[8417] = data_o[33];
  assign data_o[8481] = data_o[33];
  assign data_o[8545] = data_o[33];
  assign data_o[8609] = data_o[33];
  assign data_o[8673] = data_o[33];
  assign data_o[8737] = data_o[33];
  assign data_o[8801] = data_o[33];
  assign data_o[8865] = data_o[33];
  assign data_o[8929] = data_o[33];
  assign data_o[8993] = data_o[33];
  assign data_o[9057] = data_o[33];
  assign data_o[9121] = data_o[33];
  assign data_o[9185] = data_o[33];
  assign data_o[9249] = data_o[33];
  assign data_o[9313] = data_o[33];
  assign data_o[9377] = data_o[33];
  assign data_o[9441] = data_o[33];
  assign data_o[9505] = data_o[33];
  assign data_o[9569] = data_o[33];
  assign data_o[9633] = data_o[33];
  assign data_o[9697] = data_o[33];
  assign data_o[9761] = data_o[33];
  assign data_o[9825] = data_o[33];
  assign data_o[9889] = data_o[33];
  assign data_o[9953] = data_o[33];
  assign data_o[10017] = data_o[33];
  assign data_o[10081] = data_o[33];
  assign data_o[10145] = data_o[33];
  assign data_o[10209] = data_o[33];
  assign data_o[10273] = data_o[33];
  assign data_o[10337] = data_o[33];
  assign data_o[10401] = data_o[33];
  assign data_o[10465] = data_o[33];
  assign data_o[10529] = data_o[33];
  assign data_o[10593] = data_o[33];
  assign data_o[10657] = data_o[33];
  assign data_o[10721] = data_o[33];
  assign data_o[10785] = data_o[33];
  assign data_o[10849] = data_o[33];
  assign data_o[10913] = data_o[33];
  assign data_o[10977] = data_o[33];
  assign data_o[11041] = data_o[33];
  assign data_o[11105] = data_o[33];
  assign data_o[11169] = data_o[33];
  assign data_o[11233] = data_o[33];
  assign data_o[11297] = data_o[33];
  assign data_o[11361] = data_o[33];
  assign data_o[11425] = data_o[33];
  assign data_o[11489] = data_o[33];
  assign data_o[11553] = data_o[33];
  assign data_o[11617] = data_o[33];
  assign data_o[11681] = data_o[33];
  assign data_o[11745] = data_o[33];
  assign data_o[11809] = data_o[33];
  assign data_o[11873] = data_o[33];
  assign data_o[11937] = data_o[33];
  assign data_o[12001] = data_o[33];
  assign data_o[12065] = data_o[33];
  assign data_o[12129] = data_o[33];
  assign data_o[12193] = data_o[33];
  assign data_o[12257] = data_o[33];
  assign data_o[12321] = data_o[33];
  assign data_o[12385] = data_o[33];
  assign data_o[12449] = data_o[33];
  assign data_o[12513] = data_o[33];
  assign data_o[12577] = data_o[33];
  assign data_o[12641] = data_o[33];
  assign data_o[12705] = data_o[33];
  assign data_o[12769] = data_o[33];
  assign data_o[12833] = data_o[33];
  assign data_o[12897] = data_o[33];
  assign data_o[12961] = data_o[33];
  assign data_o[13025] = data_o[33];
  assign data_o[13089] = data_o[33];
  assign data_o[13153] = data_o[33];
  assign data_o[13217] = data_o[33];
  assign data_o[13281] = data_o[33];
  assign data_o[13345] = data_o[33];
  assign data_o[13409] = data_o[33];
  assign data_o[13473] = data_o[33];
  assign data_o[13537] = data_o[33];
  assign data_o[13601] = data_o[33];
  assign data_o[13665] = data_o[33];
  assign data_o[13729] = data_o[33];
  assign data_o[13793] = data_o[33];
  assign data_o[13857] = data_o[33];
  assign data_o[13921] = data_o[33];
  assign data_o[13985] = data_o[33];
  assign data_o[14049] = data_o[33];
  assign data_o[14113] = data_o[33];
  assign data_o[14177] = data_o[33];
  assign data_o[14241] = data_o[33];
  assign data_o[14305] = data_o[33];
  assign data_o[14369] = data_o[33];
  assign data_o[14433] = data_o[33];
  assign data_o[14497] = data_o[33];
  assign data_o[14561] = data_o[33];
  assign data_o[14625] = data_o[33];
  assign data_o[14689] = data_o[33];
  assign data_o[14753] = data_o[33];
  assign data_o[14817] = data_o[33];
  assign data_o[14881] = data_o[33];
  assign data_o[14945] = data_o[33];
  assign data_o[15009] = data_o[33];
  assign data_o[15073] = data_o[33];
  assign data_o[15137] = data_o[33];
  assign data_o[15201] = data_o[33];
  assign data_o[15265] = data_o[33];
  assign data_o[15329] = data_o[33];
  assign data_o[15393] = data_o[33];
  assign data_o[15457] = data_o[33];
  assign data_o[15521] = data_o[33];
  assign data_o[15585] = data_o[33];
  assign data_o[15649] = data_o[33];
  assign data_o[15713] = data_o[33];
  assign data_o[15777] = data_o[33];
  assign data_o[15841] = data_o[33];
  assign data_o[15905] = data_o[33];
  assign data_o[15969] = data_o[33];
  assign data_o[16033] = data_o[33];
  assign data_o[16097] = data_o[33];
  assign data_o[16161] = data_o[33];
  assign data_o[16225] = data_o[33];
  assign data_o[16289] = data_o[33];
  assign data_o[16353] = data_o[33];
  assign data_o[16417] = data_o[33];
  assign data_o[16481] = data_o[33];
  assign data_o[16545] = data_o[33];
  assign data_o[16609] = data_o[33];
  assign data_o[16673] = data_o[33];
  assign data_o[16737] = data_o[33];
  assign data_o[16801] = data_o[33];
  assign data_o[16865] = data_o[33];
  assign data_o[16929] = data_o[33];
  assign data_o[16993] = data_o[33];
  assign data_o[17057] = data_o[33];
  assign data_o[17121] = data_o[33];
  assign data_o[17185] = data_o[33];
  assign data_o[17249] = data_o[33];
  assign data_o[17313] = data_o[33];
  assign data_o[17377] = data_o[33];
  assign data_o[17441] = data_o[33];
  assign data_o[17505] = data_o[33];
  assign data_o[17569] = data_o[33];
  assign data_o[17633] = data_o[33];
  assign data_o[17697] = data_o[33];
  assign data_o[17761] = data_o[33];
  assign data_o[17825] = data_o[33];
  assign data_o[17889] = data_o[33];
  assign data_o[17953] = data_o[33];
  assign data_o[18017] = data_o[33];
  assign data_o[18081] = data_o[33];
  assign data_o[18145] = data_o[33];
  assign data_o[18209] = data_o[33];
  assign data_o[18273] = data_o[33];
  assign data_o[18337] = data_o[33];
  assign data_o[18401] = data_o[33];
  assign data_o[18465] = data_o[33];
  assign data_o[18529] = data_o[33];
  assign data_o[18593] = data_o[33];
  assign data_o[18657] = data_o[33];
  assign data_o[18721] = data_o[33];
  assign data_o[18785] = data_o[33];
  assign data_o[18849] = data_o[33];
  assign data_o[18913] = data_o[33];
  assign data_o[18977] = data_o[33];
  assign data_o[19041] = data_o[33];
  assign data_o[19105] = data_o[33];
  assign data_o[19169] = data_o[33];
  assign data_o[19233] = data_o[33];
  assign data_o[19297] = data_o[33];
  assign data_o[19361] = data_o[33];
  assign data_o[19425] = data_o[33];
  assign data_o[19489] = data_o[33];
  assign data_o[19553] = data_o[33];
  assign data_o[19617] = data_o[33];
  assign data_o[19681] = data_o[33];
  assign data_o[19745] = data_o[33];
  assign data_o[19809] = data_o[33];
  assign data_o[19873] = data_o[33];
  assign data_o[19937] = data_o[33];
  assign data_o[20001] = data_o[33];
  assign data_o[20065] = data_o[33];
  assign data_o[20129] = data_o[33];
  assign data_o[20193] = data_o[33];
  assign data_o[20257] = data_o[33];
  assign data_o[20321] = data_o[33];
  assign data_o[20385] = data_o[33];
  assign data_o[20449] = data_o[33];
  assign data_o[20513] = data_o[33];
  assign data_o[20577] = data_o[33];
  assign data_o[20641] = data_o[33];
  assign data_o[20705] = data_o[33];
  assign data_o[20769] = data_o[33];
  assign data_o[20833] = data_o[33];
  assign data_o[20897] = data_o[33];
  assign data_o[20961] = data_o[33];
  assign data_o[21025] = data_o[33];
  assign data_o[21089] = data_o[33];
  assign data_o[21153] = data_o[33];
  assign data_o[21217] = data_o[33];
  assign data_o[21281] = data_o[33];
  assign data_o[21345] = data_o[33];
  assign data_o[21409] = data_o[33];
  assign data_o[21473] = data_o[33];
  assign data_o[21537] = data_o[33];
  assign data_o[21601] = data_o[33];
  assign data_o[21665] = data_o[33];
  assign data_o[21729] = data_o[33];
  assign data_o[21793] = data_o[33];
  assign data_o[21857] = data_o[33];
  assign data_o[21921] = data_o[33];
  assign data_o[21985] = data_o[33];
  assign data_o[22049] = data_o[33];
  assign data_o[22113] = data_o[33];
  assign data_o[22177] = data_o[33];
  assign data_o[22241] = data_o[33];
  assign data_o[22305] = data_o[33];
  assign data_o[22369] = data_o[33];
  assign data_o[22433] = data_o[33];
  assign data_o[22497] = data_o[33];
  assign data_o[22561] = data_o[33];
  assign data_o[22625] = data_o[33];
  assign data_o[22689] = data_o[33];
  assign data_o[22753] = data_o[33];
  assign data_o[22817] = data_o[33];
  assign data_o[22881] = data_o[33];
  assign data_o[22945] = data_o[33];
  assign data_o[23009] = data_o[33];
  assign data_o[23073] = data_o[33];
  assign data_o[23137] = data_o[33];
  assign data_o[23201] = data_o[33];
  assign data_o[23265] = data_o[33];
  assign data_o[23329] = data_o[33];
  assign data_o[23393] = data_o[33];
  assign data_o[23457] = data_o[33];
  assign data_o[23521] = data_o[33];
  assign data_o[23585] = data_o[33];
  assign data_o[23649] = data_o[33];
  assign data_o[23713] = data_o[33];
  assign data_o[23777] = data_o[33];
  assign data_o[23841] = data_o[33];
  assign data_o[23905] = data_o[33];
  assign data_o[23969] = data_o[33];
  assign data_o[24033] = data_o[33];
  assign data_o[24097] = data_o[33];
  assign data_o[24161] = data_o[33];
  assign data_o[24225] = data_o[33];
  assign data_o[24289] = data_o[33];
  assign data_o[24353] = data_o[33];
  assign data_o[24417] = data_o[33];
  assign data_o[24481] = data_o[33];
  assign data_o[24545] = data_o[33];
  assign data_o[24609] = data_o[33];
  assign data_o[24673] = data_o[33];
  assign data_o[24737] = data_o[33];
  assign data_o[24801] = data_o[33];
  assign data_o[24865] = data_o[33];
  assign data_o[24929] = data_o[33];
  assign data_o[24993] = data_o[33];
  assign data_o[25057] = data_o[33];
  assign data_o[25121] = data_o[33];
  assign data_o[25185] = data_o[33];
  assign data_o[25249] = data_o[33];
  assign data_o[25313] = data_o[33];
  assign data_o[25377] = data_o[33];
  assign data_o[25441] = data_o[33];
  assign data_o[25505] = data_o[33];
  assign data_o[25569] = data_o[33];
  assign data_o[25633] = data_o[33];
  assign data_o[25697] = data_o[33];
  assign data_o[25761] = data_o[33];
  assign data_o[25825] = data_o[33];
  assign data_o[25889] = data_o[33];
  assign data_o[25953] = data_o[33];
  assign data_o[26017] = data_o[33];
  assign data_o[26081] = data_o[33];
  assign data_o[26145] = data_o[33];
  assign data_o[26209] = data_o[33];
  assign data_o[26273] = data_o[33];
  assign data_o[26337] = data_o[33];
  assign data_o[26401] = data_o[33];
  assign data_o[26465] = data_o[33];
  assign data_o[26529] = data_o[33];
  assign data_o[26593] = data_o[33];
  assign data_o[26657] = data_o[33];
  assign data_o[26721] = data_o[33];
  assign data_o[26785] = data_o[33];
  assign data_o[26849] = data_o[33];
  assign data_o[26913] = data_o[33];
  assign data_o[26977] = data_o[33];
  assign data_o[27041] = data_o[33];
  assign data_o[27105] = data_o[33];
  assign data_o[27169] = data_o[33];
  assign data_o[27233] = data_o[33];
  assign data_o[27297] = data_o[33];
  assign data_o[27361] = data_o[33];
  assign data_o[27425] = data_o[33];
  assign data_o[27489] = data_o[33];
  assign data_o[27553] = data_o[33];
  assign data_o[27617] = data_o[33];
  assign data_o[27681] = data_o[33];
  assign data_o[27745] = data_o[33];
  assign data_o[27809] = data_o[33];
  assign data_o[27873] = data_o[33];
  assign data_o[27937] = data_o[33];
  assign data_o[28001] = data_o[33];
  assign data_o[28065] = data_o[33];
  assign data_o[28129] = data_o[33];
  assign data_o[28193] = data_o[33];
  assign data_o[28257] = data_o[33];
  assign data_o[28321] = data_o[33];
  assign data_o[28385] = data_o[33];
  assign data_o[28449] = data_o[33];
  assign data_o[28513] = data_o[33];
  assign data_o[28577] = data_o[33];
  assign data_o[28641] = data_o[33];
  assign data_o[28705] = data_o[33];
  assign data_o[28769] = data_o[33];
  assign data_o[28833] = data_o[33];
  assign data_o[28897] = data_o[33];
  assign data_o[28961] = data_o[33];
  assign data_o[29025] = data_o[33];
  assign data_o[29089] = data_o[33];
  assign data_o[29153] = data_o[33];
  assign data_o[29217] = data_o[33];
  assign data_o[29281] = data_o[33];
  assign data_o[29345] = data_o[33];
  assign data_o[29409] = data_o[33];
  assign data_o[29473] = data_o[33];
  assign data_o[29537] = data_o[33];
  assign data_o[29601] = data_o[33];
  assign data_o[29665] = data_o[33];
  assign data_o[29729] = data_o[33];
  assign data_o[29793] = data_o[33];
  assign data_o[29857] = data_o[33];
  assign data_o[29921] = data_o[33];
  assign data_o[29985] = data_o[33];
  assign data_o[30049] = data_o[33];
  assign data_o[30113] = data_o[33];
  assign data_o[30177] = data_o[33];
  assign data_o[30241] = data_o[33];
  assign data_o[30305] = data_o[33];
  assign data_o[30369] = data_o[33];
  assign data_o[30433] = data_o[33];
  assign data_o[30497] = data_o[33];
  assign data_o[30561] = data_o[33];
  assign data_o[30625] = data_o[33];
  assign data_o[30689] = data_o[33];
  assign data_o[30753] = data_o[33];
  assign data_o[30817] = data_o[33];
  assign data_o[30881] = data_o[33];
  assign data_o[30945] = data_o[33];
  assign data_o[31009] = data_o[33];
  assign data_o[31073] = data_o[33];
  assign data_o[31137] = data_o[33];
  assign data_o[31201] = data_o[33];
  assign data_o[31265] = data_o[33];
  assign data_o[31329] = data_o[33];
  assign data_o[31393] = data_o[33];
  assign data_o[31457] = data_o[33];
  assign data_o[31521] = data_o[33];
  assign data_o[31585] = data_o[33];
  assign data_o[31649] = data_o[33];
  assign data_o[31713] = data_o[33];
  assign data_o[31777] = data_o[33];
  assign data_o[31841] = data_o[33];
  assign data_o[31905] = data_o[33];
  assign data_o[31969] = data_o[33];
  assign data_o[96] = data_o[32];
  assign data_o[160] = data_o[32];
  assign data_o[224] = data_o[32];
  assign data_o[288] = data_o[32];
  assign data_o[352] = data_o[32];
  assign data_o[416] = data_o[32];
  assign data_o[480] = data_o[32];
  assign data_o[544] = data_o[32];
  assign data_o[608] = data_o[32];
  assign data_o[672] = data_o[32];
  assign data_o[736] = data_o[32];
  assign data_o[800] = data_o[32];
  assign data_o[864] = data_o[32];
  assign data_o[928] = data_o[32];
  assign data_o[992] = data_o[32];
  assign data_o[1056] = data_o[32];
  assign data_o[1120] = data_o[32];
  assign data_o[1184] = data_o[32];
  assign data_o[1248] = data_o[32];
  assign data_o[1312] = data_o[32];
  assign data_o[1376] = data_o[32];
  assign data_o[1440] = data_o[32];
  assign data_o[1504] = data_o[32];
  assign data_o[1568] = data_o[32];
  assign data_o[1632] = data_o[32];
  assign data_o[1696] = data_o[32];
  assign data_o[1760] = data_o[32];
  assign data_o[1824] = data_o[32];
  assign data_o[1888] = data_o[32];
  assign data_o[1952] = data_o[32];
  assign data_o[2016] = data_o[32];
  assign data_o[2080] = data_o[32];
  assign data_o[2144] = data_o[32];
  assign data_o[2208] = data_o[32];
  assign data_o[2272] = data_o[32];
  assign data_o[2336] = data_o[32];
  assign data_o[2400] = data_o[32];
  assign data_o[2464] = data_o[32];
  assign data_o[2528] = data_o[32];
  assign data_o[2592] = data_o[32];
  assign data_o[2656] = data_o[32];
  assign data_o[2720] = data_o[32];
  assign data_o[2784] = data_o[32];
  assign data_o[2848] = data_o[32];
  assign data_o[2912] = data_o[32];
  assign data_o[2976] = data_o[32];
  assign data_o[3040] = data_o[32];
  assign data_o[3104] = data_o[32];
  assign data_o[3168] = data_o[32];
  assign data_o[3232] = data_o[32];
  assign data_o[3296] = data_o[32];
  assign data_o[3360] = data_o[32];
  assign data_o[3424] = data_o[32];
  assign data_o[3488] = data_o[32];
  assign data_o[3552] = data_o[32];
  assign data_o[3616] = data_o[32];
  assign data_o[3680] = data_o[32];
  assign data_o[3744] = data_o[32];
  assign data_o[3808] = data_o[32];
  assign data_o[3872] = data_o[32];
  assign data_o[3936] = data_o[32];
  assign data_o[4000] = data_o[32];
  assign data_o[4064] = data_o[32];
  assign data_o[4128] = data_o[32];
  assign data_o[4192] = data_o[32];
  assign data_o[4256] = data_o[32];
  assign data_o[4320] = data_o[32];
  assign data_o[4384] = data_o[32];
  assign data_o[4448] = data_o[32];
  assign data_o[4512] = data_o[32];
  assign data_o[4576] = data_o[32];
  assign data_o[4640] = data_o[32];
  assign data_o[4704] = data_o[32];
  assign data_o[4768] = data_o[32];
  assign data_o[4832] = data_o[32];
  assign data_o[4896] = data_o[32];
  assign data_o[4960] = data_o[32];
  assign data_o[5024] = data_o[32];
  assign data_o[5088] = data_o[32];
  assign data_o[5152] = data_o[32];
  assign data_o[5216] = data_o[32];
  assign data_o[5280] = data_o[32];
  assign data_o[5344] = data_o[32];
  assign data_o[5408] = data_o[32];
  assign data_o[5472] = data_o[32];
  assign data_o[5536] = data_o[32];
  assign data_o[5600] = data_o[32];
  assign data_o[5664] = data_o[32];
  assign data_o[5728] = data_o[32];
  assign data_o[5792] = data_o[32];
  assign data_o[5856] = data_o[32];
  assign data_o[5920] = data_o[32];
  assign data_o[5984] = data_o[32];
  assign data_o[6048] = data_o[32];
  assign data_o[6112] = data_o[32];
  assign data_o[6176] = data_o[32];
  assign data_o[6240] = data_o[32];
  assign data_o[6304] = data_o[32];
  assign data_o[6368] = data_o[32];
  assign data_o[6432] = data_o[32];
  assign data_o[6496] = data_o[32];
  assign data_o[6560] = data_o[32];
  assign data_o[6624] = data_o[32];
  assign data_o[6688] = data_o[32];
  assign data_o[6752] = data_o[32];
  assign data_o[6816] = data_o[32];
  assign data_o[6880] = data_o[32];
  assign data_o[6944] = data_o[32];
  assign data_o[7008] = data_o[32];
  assign data_o[7072] = data_o[32];
  assign data_o[7136] = data_o[32];
  assign data_o[7200] = data_o[32];
  assign data_o[7264] = data_o[32];
  assign data_o[7328] = data_o[32];
  assign data_o[7392] = data_o[32];
  assign data_o[7456] = data_o[32];
  assign data_o[7520] = data_o[32];
  assign data_o[7584] = data_o[32];
  assign data_o[7648] = data_o[32];
  assign data_o[7712] = data_o[32];
  assign data_o[7776] = data_o[32];
  assign data_o[7840] = data_o[32];
  assign data_o[7904] = data_o[32];
  assign data_o[7968] = data_o[32];
  assign data_o[8032] = data_o[32];
  assign data_o[8096] = data_o[32];
  assign data_o[8160] = data_o[32];
  assign data_o[8224] = data_o[32];
  assign data_o[8288] = data_o[32];
  assign data_o[8352] = data_o[32];
  assign data_o[8416] = data_o[32];
  assign data_o[8480] = data_o[32];
  assign data_o[8544] = data_o[32];
  assign data_o[8608] = data_o[32];
  assign data_o[8672] = data_o[32];
  assign data_o[8736] = data_o[32];
  assign data_o[8800] = data_o[32];
  assign data_o[8864] = data_o[32];
  assign data_o[8928] = data_o[32];
  assign data_o[8992] = data_o[32];
  assign data_o[9056] = data_o[32];
  assign data_o[9120] = data_o[32];
  assign data_o[9184] = data_o[32];
  assign data_o[9248] = data_o[32];
  assign data_o[9312] = data_o[32];
  assign data_o[9376] = data_o[32];
  assign data_o[9440] = data_o[32];
  assign data_o[9504] = data_o[32];
  assign data_o[9568] = data_o[32];
  assign data_o[9632] = data_o[32];
  assign data_o[9696] = data_o[32];
  assign data_o[9760] = data_o[32];
  assign data_o[9824] = data_o[32];
  assign data_o[9888] = data_o[32];
  assign data_o[9952] = data_o[32];
  assign data_o[10016] = data_o[32];
  assign data_o[10080] = data_o[32];
  assign data_o[10144] = data_o[32];
  assign data_o[10208] = data_o[32];
  assign data_o[10272] = data_o[32];
  assign data_o[10336] = data_o[32];
  assign data_o[10400] = data_o[32];
  assign data_o[10464] = data_o[32];
  assign data_o[10528] = data_o[32];
  assign data_o[10592] = data_o[32];
  assign data_o[10656] = data_o[32];
  assign data_o[10720] = data_o[32];
  assign data_o[10784] = data_o[32];
  assign data_o[10848] = data_o[32];
  assign data_o[10912] = data_o[32];
  assign data_o[10976] = data_o[32];
  assign data_o[11040] = data_o[32];
  assign data_o[11104] = data_o[32];
  assign data_o[11168] = data_o[32];
  assign data_o[11232] = data_o[32];
  assign data_o[11296] = data_o[32];
  assign data_o[11360] = data_o[32];
  assign data_o[11424] = data_o[32];
  assign data_o[11488] = data_o[32];
  assign data_o[11552] = data_o[32];
  assign data_o[11616] = data_o[32];
  assign data_o[11680] = data_o[32];
  assign data_o[11744] = data_o[32];
  assign data_o[11808] = data_o[32];
  assign data_o[11872] = data_o[32];
  assign data_o[11936] = data_o[32];
  assign data_o[12000] = data_o[32];
  assign data_o[12064] = data_o[32];
  assign data_o[12128] = data_o[32];
  assign data_o[12192] = data_o[32];
  assign data_o[12256] = data_o[32];
  assign data_o[12320] = data_o[32];
  assign data_o[12384] = data_o[32];
  assign data_o[12448] = data_o[32];
  assign data_o[12512] = data_o[32];
  assign data_o[12576] = data_o[32];
  assign data_o[12640] = data_o[32];
  assign data_o[12704] = data_o[32];
  assign data_o[12768] = data_o[32];
  assign data_o[12832] = data_o[32];
  assign data_o[12896] = data_o[32];
  assign data_o[12960] = data_o[32];
  assign data_o[13024] = data_o[32];
  assign data_o[13088] = data_o[32];
  assign data_o[13152] = data_o[32];
  assign data_o[13216] = data_o[32];
  assign data_o[13280] = data_o[32];
  assign data_o[13344] = data_o[32];
  assign data_o[13408] = data_o[32];
  assign data_o[13472] = data_o[32];
  assign data_o[13536] = data_o[32];
  assign data_o[13600] = data_o[32];
  assign data_o[13664] = data_o[32];
  assign data_o[13728] = data_o[32];
  assign data_o[13792] = data_o[32];
  assign data_o[13856] = data_o[32];
  assign data_o[13920] = data_o[32];
  assign data_o[13984] = data_o[32];
  assign data_o[14048] = data_o[32];
  assign data_o[14112] = data_o[32];
  assign data_o[14176] = data_o[32];
  assign data_o[14240] = data_o[32];
  assign data_o[14304] = data_o[32];
  assign data_o[14368] = data_o[32];
  assign data_o[14432] = data_o[32];
  assign data_o[14496] = data_o[32];
  assign data_o[14560] = data_o[32];
  assign data_o[14624] = data_o[32];
  assign data_o[14688] = data_o[32];
  assign data_o[14752] = data_o[32];
  assign data_o[14816] = data_o[32];
  assign data_o[14880] = data_o[32];
  assign data_o[14944] = data_o[32];
  assign data_o[15008] = data_o[32];
  assign data_o[15072] = data_o[32];
  assign data_o[15136] = data_o[32];
  assign data_o[15200] = data_o[32];
  assign data_o[15264] = data_o[32];
  assign data_o[15328] = data_o[32];
  assign data_o[15392] = data_o[32];
  assign data_o[15456] = data_o[32];
  assign data_o[15520] = data_o[32];
  assign data_o[15584] = data_o[32];
  assign data_o[15648] = data_o[32];
  assign data_o[15712] = data_o[32];
  assign data_o[15776] = data_o[32];
  assign data_o[15840] = data_o[32];
  assign data_o[15904] = data_o[32];
  assign data_o[15968] = data_o[32];
  assign data_o[16032] = data_o[32];
  assign data_o[16096] = data_o[32];
  assign data_o[16160] = data_o[32];
  assign data_o[16224] = data_o[32];
  assign data_o[16288] = data_o[32];
  assign data_o[16352] = data_o[32];
  assign data_o[16416] = data_o[32];
  assign data_o[16480] = data_o[32];
  assign data_o[16544] = data_o[32];
  assign data_o[16608] = data_o[32];
  assign data_o[16672] = data_o[32];
  assign data_o[16736] = data_o[32];
  assign data_o[16800] = data_o[32];
  assign data_o[16864] = data_o[32];
  assign data_o[16928] = data_o[32];
  assign data_o[16992] = data_o[32];
  assign data_o[17056] = data_o[32];
  assign data_o[17120] = data_o[32];
  assign data_o[17184] = data_o[32];
  assign data_o[17248] = data_o[32];
  assign data_o[17312] = data_o[32];
  assign data_o[17376] = data_o[32];
  assign data_o[17440] = data_o[32];
  assign data_o[17504] = data_o[32];
  assign data_o[17568] = data_o[32];
  assign data_o[17632] = data_o[32];
  assign data_o[17696] = data_o[32];
  assign data_o[17760] = data_o[32];
  assign data_o[17824] = data_o[32];
  assign data_o[17888] = data_o[32];
  assign data_o[17952] = data_o[32];
  assign data_o[18016] = data_o[32];
  assign data_o[18080] = data_o[32];
  assign data_o[18144] = data_o[32];
  assign data_o[18208] = data_o[32];
  assign data_o[18272] = data_o[32];
  assign data_o[18336] = data_o[32];
  assign data_o[18400] = data_o[32];
  assign data_o[18464] = data_o[32];
  assign data_o[18528] = data_o[32];
  assign data_o[18592] = data_o[32];
  assign data_o[18656] = data_o[32];
  assign data_o[18720] = data_o[32];
  assign data_o[18784] = data_o[32];
  assign data_o[18848] = data_o[32];
  assign data_o[18912] = data_o[32];
  assign data_o[18976] = data_o[32];
  assign data_o[19040] = data_o[32];
  assign data_o[19104] = data_o[32];
  assign data_o[19168] = data_o[32];
  assign data_o[19232] = data_o[32];
  assign data_o[19296] = data_o[32];
  assign data_o[19360] = data_o[32];
  assign data_o[19424] = data_o[32];
  assign data_o[19488] = data_o[32];
  assign data_o[19552] = data_o[32];
  assign data_o[19616] = data_o[32];
  assign data_o[19680] = data_o[32];
  assign data_o[19744] = data_o[32];
  assign data_o[19808] = data_o[32];
  assign data_o[19872] = data_o[32];
  assign data_o[19936] = data_o[32];
  assign data_o[20000] = data_o[32];
  assign data_o[20064] = data_o[32];
  assign data_o[20128] = data_o[32];
  assign data_o[20192] = data_o[32];
  assign data_o[20256] = data_o[32];
  assign data_o[20320] = data_o[32];
  assign data_o[20384] = data_o[32];
  assign data_o[20448] = data_o[32];
  assign data_o[20512] = data_o[32];
  assign data_o[20576] = data_o[32];
  assign data_o[20640] = data_o[32];
  assign data_o[20704] = data_o[32];
  assign data_o[20768] = data_o[32];
  assign data_o[20832] = data_o[32];
  assign data_o[20896] = data_o[32];
  assign data_o[20960] = data_o[32];
  assign data_o[21024] = data_o[32];
  assign data_o[21088] = data_o[32];
  assign data_o[21152] = data_o[32];
  assign data_o[21216] = data_o[32];
  assign data_o[21280] = data_o[32];
  assign data_o[21344] = data_o[32];
  assign data_o[21408] = data_o[32];
  assign data_o[21472] = data_o[32];
  assign data_o[21536] = data_o[32];
  assign data_o[21600] = data_o[32];
  assign data_o[21664] = data_o[32];
  assign data_o[21728] = data_o[32];
  assign data_o[21792] = data_o[32];
  assign data_o[21856] = data_o[32];
  assign data_o[21920] = data_o[32];
  assign data_o[21984] = data_o[32];
  assign data_o[22048] = data_o[32];
  assign data_o[22112] = data_o[32];
  assign data_o[22176] = data_o[32];
  assign data_o[22240] = data_o[32];
  assign data_o[22304] = data_o[32];
  assign data_o[22368] = data_o[32];
  assign data_o[22432] = data_o[32];
  assign data_o[22496] = data_o[32];
  assign data_o[22560] = data_o[32];
  assign data_o[22624] = data_o[32];
  assign data_o[22688] = data_o[32];
  assign data_o[22752] = data_o[32];
  assign data_o[22816] = data_o[32];
  assign data_o[22880] = data_o[32];
  assign data_o[22944] = data_o[32];
  assign data_o[23008] = data_o[32];
  assign data_o[23072] = data_o[32];
  assign data_o[23136] = data_o[32];
  assign data_o[23200] = data_o[32];
  assign data_o[23264] = data_o[32];
  assign data_o[23328] = data_o[32];
  assign data_o[23392] = data_o[32];
  assign data_o[23456] = data_o[32];
  assign data_o[23520] = data_o[32];
  assign data_o[23584] = data_o[32];
  assign data_o[23648] = data_o[32];
  assign data_o[23712] = data_o[32];
  assign data_o[23776] = data_o[32];
  assign data_o[23840] = data_o[32];
  assign data_o[23904] = data_o[32];
  assign data_o[23968] = data_o[32];
  assign data_o[24032] = data_o[32];
  assign data_o[24096] = data_o[32];
  assign data_o[24160] = data_o[32];
  assign data_o[24224] = data_o[32];
  assign data_o[24288] = data_o[32];
  assign data_o[24352] = data_o[32];
  assign data_o[24416] = data_o[32];
  assign data_o[24480] = data_o[32];
  assign data_o[24544] = data_o[32];
  assign data_o[24608] = data_o[32];
  assign data_o[24672] = data_o[32];
  assign data_o[24736] = data_o[32];
  assign data_o[24800] = data_o[32];
  assign data_o[24864] = data_o[32];
  assign data_o[24928] = data_o[32];
  assign data_o[24992] = data_o[32];
  assign data_o[25056] = data_o[32];
  assign data_o[25120] = data_o[32];
  assign data_o[25184] = data_o[32];
  assign data_o[25248] = data_o[32];
  assign data_o[25312] = data_o[32];
  assign data_o[25376] = data_o[32];
  assign data_o[25440] = data_o[32];
  assign data_o[25504] = data_o[32];
  assign data_o[25568] = data_o[32];
  assign data_o[25632] = data_o[32];
  assign data_o[25696] = data_o[32];
  assign data_o[25760] = data_o[32];
  assign data_o[25824] = data_o[32];
  assign data_o[25888] = data_o[32];
  assign data_o[25952] = data_o[32];
  assign data_o[26016] = data_o[32];
  assign data_o[26080] = data_o[32];
  assign data_o[26144] = data_o[32];
  assign data_o[26208] = data_o[32];
  assign data_o[26272] = data_o[32];
  assign data_o[26336] = data_o[32];
  assign data_o[26400] = data_o[32];
  assign data_o[26464] = data_o[32];
  assign data_o[26528] = data_o[32];
  assign data_o[26592] = data_o[32];
  assign data_o[26656] = data_o[32];
  assign data_o[26720] = data_o[32];
  assign data_o[26784] = data_o[32];
  assign data_o[26848] = data_o[32];
  assign data_o[26912] = data_o[32];
  assign data_o[26976] = data_o[32];
  assign data_o[27040] = data_o[32];
  assign data_o[27104] = data_o[32];
  assign data_o[27168] = data_o[32];
  assign data_o[27232] = data_o[32];
  assign data_o[27296] = data_o[32];
  assign data_o[27360] = data_o[32];
  assign data_o[27424] = data_o[32];
  assign data_o[27488] = data_o[32];
  assign data_o[27552] = data_o[32];
  assign data_o[27616] = data_o[32];
  assign data_o[27680] = data_o[32];
  assign data_o[27744] = data_o[32];
  assign data_o[27808] = data_o[32];
  assign data_o[27872] = data_o[32];
  assign data_o[27936] = data_o[32];
  assign data_o[28000] = data_o[32];
  assign data_o[28064] = data_o[32];
  assign data_o[28128] = data_o[32];
  assign data_o[28192] = data_o[32];
  assign data_o[28256] = data_o[32];
  assign data_o[28320] = data_o[32];
  assign data_o[28384] = data_o[32];
  assign data_o[28448] = data_o[32];
  assign data_o[28512] = data_o[32];
  assign data_o[28576] = data_o[32];
  assign data_o[28640] = data_o[32];
  assign data_o[28704] = data_o[32];
  assign data_o[28768] = data_o[32];
  assign data_o[28832] = data_o[32];
  assign data_o[28896] = data_o[32];
  assign data_o[28960] = data_o[32];
  assign data_o[29024] = data_o[32];
  assign data_o[29088] = data_o[32];
  assign data_o[29152] = data_o[32];
  assign data_o[29216] = data_o[32];
  assign data_o[29280] = data_o[32];
  assign data_o[29344] = data_o[32];
  assign data_o[29408] = data_o[32];
  assign data_o[29472] = data_o[32];
  assign data_o[29536] = data_o[32];
  assign data_o[29600] = data_o[32];
  assign data_o[29664] = data_o[32];
  assign data_o[29728] = data_o[32];
  assign data_o[29792] = data_o[32];
  assign data_o[29856] = data_o[32];
  assign data_o[29920] = data_o[32];
  assign data_o[29984] = data_o[32];
  assign data_o[30048] = data_o[32];
  assign data_o[30112] = data_o[32];
  assign data_o[30176] = data_o[32];
  assign data_o[30240] = data_o[32];
  assign data_o[30304] = data_o[32];
  assign data_o[30368] = data_o[32];
  assign data_o[30432] = data_o[32];
  assign data_o[30496] = data_o[32];
  assign data_o[30560] = data_o[32];
  assign data_o[30624] = data_o[32];
  assign data_o[30688] = data_o[32];
  assign data_o[30752] = data_o[32];
  assign data_o[30816] = data_o[32];
  assign data_o[30880] = data_o[32];
  assign data_o[30944] = data_o[32];
  assign data_o[31008] = data_o[32];
  assign data_o[31072] = data_o[32];
  assign data_o[31136] = data_o[32];
  assign data_o[31200] = data_o[32];
  assign data_o[31264] = data_o[32];
  assign data_o[31328] = data_o[32];
  assign data_o[31392] = data_o[32];
  assign data_o[31456] = data_o[32];
  assign data_o[31520] = data_o[32];
  assign data_o[31584] = data_o[32];
  assign data_o[31648] = data_o[32];
  assign data_o[31712] = data_o[32];
  assign data_o[31776] = data_o[32];
  assign data_o[31840] = data_o[32];
  assign data_o[31904] = data_o[32];
  assign data_o[31968] = data_o[32];
  assign data_o[95] = data_o[31];
  assign data_o[159] = data_o[31];
  assign data_o[223] = data_o[31];
  assign data_o[287] = data_o[31];
  assign data_o[351] = data_o[31];
  assign data_o[415] = data_o[31];
  assign data_o[479] = data_o[31];
  assign data_o[543] = data_o[31];
  assign data_o[607] = data_o[31];
  assign data_o[671] = data_o[31];
  assign data_o[735] = data_o[31];
  assign data_o[799] = data_o[31];
  assign data_o[863] = data_o[31];
  assign data_o[927] = data_o[31];
  assign data_o[991] = data_o[31];
  assign data_o[1055] = data_o[31];
  assign data_o[1119] = data_o[31];
  assign data_o[1183] = data_o[31];
  assign data_o[1247] = data_o[31];
  assign data_o[1311] = data_o[31];
  assign data_o[1375] = data_o[31];
  assign data_o[1439] = data_o[31];
  assign data_o[1503] = data_o[31];
  assign data_o[1567] = data_o[31];
  assign data_o[1631] = data_o[31];
  assign data_o[1695] = data_o[31];
  assign data_o[1759] = data_o[31];
  assign data_o[1823] = data_o[31];
  assign data_o[1887] = data_o[31];
  assign data_o[1951] = data_o[31];
  assign data_o[2015] = data_o[31];
  assign data_o[2079] = data_o[31];
  assign data_o[2143] = data_o[31];
  assign data_o[2207] = data_o[31];
  assign data_o[2271] = data_o[31];
  assign data_o[2335] = data_o[31];
  assign data_o[2399] = data_o[31];
  assign data_o[2463] = data_o[31];
  assign data_o[2527] = data_o[31];
  assign data_o[2591] = data_o[31];
  assign data_o[2655] = data_o[31];
  assign data_o[2719] = data_o[31];
  assign data_o[2783] = data_o[31];
  assign data_o[2847] = data_o[31];
  assign data_o[2911] = data_o[31];
  assign data_o[2975] = data_o[31];
  assign data_o[3039] = data_o[31];
  assign data_o[3103] = data_o[31];
  assign data_o[3167] = data_o[31];
  assign data_o[3231] = data_o[31];
  assign data_o[3295] = data_o[31];
  assign data_o[3359] = data_o[31];
  assign data_o[3423] = data_o[31];
  assign data_o[3487] = data_o[31];
  assign data_o[3551] = data_o[31];
  assign data_o[3615] = data_o[31];
  assign data_o[3679] = data_o[31];
  assign data_o[3743] = data_o[31];
  assign data_o[3807] = data_o[31];
  assign data_o[3871] = data_o[31];
  assign data_o[3935] = data_o[31];
  assign data_o[3999] = data_o[31];
  assign data_o[4063] = data_o[31];
  assign data_o[4127] = data_o[31];
  assign data_o[4191] = data_o[31];
  assign data_o[4255] = data_o[31];
  assign data_o[4319] = data_o[31];
  assign data_o[4383] = data_o[31];
  assign data_o[4447] = data_o[31];
  assign data_o[4511] = data_o[31];
  assign data_o[4575] = data_o[31];
  assign data_o[4639] = data_o[31];
  assign data_o[4703] = data_o[31];
  assign data_o[4767] = data_o[31];
  assign data_o[4831] = data_o[31];
  assign data_o[4895] = data_o[31];
  assign data_o[4959] = data_o[31];
  assign data_o[5023] = data_o[31];
  assign data_o[5087] = data_o[31];
  assign data_o[5151] = data_o[31];
  assign data_o[5215] = data_o[31];
  assign data_o[5279] = data_o[31];
  assign data_o[5343] = data_o[31];
  assign data_o[5407] = data_o[31];
  assign data_o[5471] = data_o[31];
  assign data_o[5535] = data_o[31];
  assign data_o[5599] = data_o[31];
  assign data_o[5663] = data_o[31];
  assign data_o[5727] = data_o[31];
  assign data_o[5791] = data_o[31];
  assign data_o[5855] = data_o[31];
  assign data_o[5919] = data_o[31];
  assign data_o[5983] = data_o[31];
  assign data_o[6047] = data_o[31];
  assign data_o[6111] = data_o[31];
  assign data_o[6175] = data_o[31];
  assign data_o[6239] = data_o[31];
  assign data_o[6303] = data_o[31];
  assign data_o[6367] = data_o[31];
  assign data_o[6431] = data_o[31];
  assign data_o[6495] = data_o[31];
  assign data_o[6559] = data_o[31];
  assign data_o[6623] = data_o[31];
  assign data_o[6687] = data_o[31];
  assign data_o[6751] = data_o[31];
  assign data_o[6815] = data_o[31];
  assign data_o[6879] = data_o[31];
  assign data_o[6943] = data_o[31];
  assign data_o[7007] = data_o[31];
  assign data_o[7071] = data_o[31];
  assign data_o[7135] = data_o[31];
  assign data_o[7199] = data_o[31];
  assign data_o[7263] = data_o[31];
  assign data_o[7327] = data_o[31];
  assign data_o[7391] = data_o[31];
  assign data_o[7455] = data_o[31];
  assign data_o[7519] = data_o[31];
  assign data_o[7583] = data_o[31];
  assign data_o[7647] = data_o[31];
  assign data_o[7711] = data_o[31];
  assign data_o[7775] = data_o[31];
  assign data_o[7839] = data_o[31];
  assign data_o[7903] = data_o[31];
  assign data_o[7967] = data_o[31];
  assign data_o[8031] = data_o[31];
  assign data_o[8095] = data_o[31];
  assign data_o[8159] = data_o[31];
  assign data_o[8223] = data_o[31];
  assign data_o[8287] = data_o[31];
  assign data_o[8351] = data_o[31];
  assign data_o[8415] = data_o[31];
  assign data_o[8479] = data_o[31];
  assign data_o[8543] = data_o[31];
  assign data_o[8607] = data_o[31];
  assign data_o[8671] = data_o[31];
  assign data_o[8735] = data_o[31];
  assign data_o[8799] = data_o[31];
  assign data_o[8863] = data_o[31];
  assign data_o[8927] = data_o[31];
  assign data_o[8991] = data_o[31];
  assign data_o[9055] = data_o[31];
  assign data_o[9119] = data_o[31];
  assign data_o[9183] = data_o[31];
  assign data_o[9247] = data_o[31];
  assign data_o[9311] = data_o[31];
  assign data_o[9375] = data_o[31];
  assign data_o[9439] = data_o[31];
  assign data_o[9503] = data_o[31];
  assign data_o[9567] = data_o[31];
  assign data_o[9631] = data_o[31];
  assign data_o[9695] = data_o[31];
  assign data_o[9759] = data_o[31];
  assign data_o[9823] = data_o[31];
  assign data_o[9887] = data_o[31];
  assign data_o[9951] = data_o[31];
  assign data_o[10015] = data_o[31];
  assign data_o[10079] = data_o[31];
  assign data_o[10143] = data_o[31];
  assign data_o[10207] = data_o[31];
  assign data_o[10271] = data_o[31];
  assign data_o[10335] = data_o[31];
  assign data_o[10399] = data_o[31];
  assign data_o[10463] = data_o[31];
  assign data_o[10527] = data_o[31];
  assign data_o[10591] = data_o[31];
  assign data_o[10655] = data_o[31];
  assign data_o[10719] = data_o[31];
  assign data_o[10783] = data_o[31];
  assign data_o[10847] = data_o[31];
  assign data_o[10911] = data_o[31];
  assign data_o[10975] = data_o[31];
  assign data_o[11039] = data_o[31];
  assign data_o[11103] = data_o[31];
  assign data_o[11167] = data_o[31];
  assign data_o[11231] = data_o[31];
  assign data_o[11295] = data_o[31];
  assign data_o[11359] = data_o[31];
  assign data_o[11423] = data_o[31];
  assign data_o[11487] = data_o[31];
  assign data_o[11551] = data_o[31];
  assign data_o[11615] = data_o[31];
  assign data_o[11679] = data_o[31];
  assign data_o[11743] = data_o[31];
  assign data_o[11807] = data_o[31];
  assign data_o[11871] = data_o[31];
  assign data_o[11935] = data_o[31];
  assign data_o[11999] = data_o[31];
  assign data_o[12063] = data_o[31];
  assign data_o[12127] = data_o[31];
  assign data_o[12191] = data_o[31];
  assign data_o[12255] = data_o[31];
  assign data_o[12319] = data_o[31];
  assign data_o[12383] = data_o[31];
  assign data_o[12447] = data_o[31];
  assign data_o[12511] = data_o[31];
  assign data_o[12575] = data_o[31];
  assign data_o[12639] = data_o[31];
  assign data_o[12703] = data_o[31];
  assign data_o[12767] = data_o[31];
  assign data_o[12831] = data_o[31];
  assign data_o[12895] = data_o[31];
  assign data_o[12959] = data_o[31];
  assign data_o[13023] = data_o[31];
  assign data_o[13087] = data_o[31];
  assign data_o[13151] = data_o[31];
  assign data_o[13215] = data_o[31];
  assign data_o[13279] = data_o[31];
  assign data_o[13343] = data_o[31];
  assign data_o[13407] = data_o[31];
  assign data_o[13471] = data_o[31];
  assign data_o[13535] = data_o[31];
  assign data_o[13599] = data_o[31];
  assign data_o[13663] = data_o[31];
  assign data_o[13727] = data_o[31];
  assign data_o[13791] = data_o[31];
  assign data_o[13855] = data_o[31];
  assign data_o[13919] = data_o[31];
  assign data_o[13983] = data_o[31];
  assign data_o[14047] = data_o[31];
  assign data_o[14111] = data_o[31];
  assign data_o[14175] = data_o[31];
  assign data_o[14239] = data_o[31];
  assign data_o[14303] = data_o[31];
  assign data_o[14367] = data_o[31];
  assign data_o[14431] = data_o[31];
  assign data_o[14495] = data_o[31];
  assign data_o[14559] = data_o[31];
  assign data_o[14623] = data_o[31];
  assign data_o[14687] = data_o[31];
  assign data_o[14751] = data_o[31];
  assign data_o[14815] = data_o[31];
  assign data_o[14879] = data_o[31];
  assign data_o[14943] = data_o[31];
  assign data_o[15007] = data_o[31];
  assign data_o[15071] = data_o[31];
  assign data_o[15135] = data_o[31];
  assign data_o[15199] = data_o[31];
  assign data_o[15263] = data_o[31];
  assign data_o[15327] = data_o[31];
  assign data_o[15391] = data_o[31];
  assign data_o[15455] = data_o[31];
  assign data_o[15519] = data_o[31];
  assign data_o[15583] = data_o[31];
  assign data_o[15647] = data_o[31];
  assign data_o[15711] = data_o[31];
  assign data_o[15775] = data_o[31];
  assign data_o[15839] = data_o[31];
  assign data_o[15903] = data_o[31];
  assign data_o[15967] = data_o[31];
  assign data_o[16031] = data_o[31];
  assign data_o[16095] = data_o[31];
  assign data_o[16159] = data_o[31];
  assign data_o[16223] = data_o[31];
  assign data_o[16287] = data_o[31];
  assign data_o[16351] = data_o[31];
  assign data_o[16415] = data_o[31];
  assign data_o[16479] = data_o[31];
  assign data_o[16543] = data_o[31];
  assign data_o[16607] = data_o[31];
  assign data_o[16671] = data_o[31];
  assign data_o[16735] = data_o[31];
  assign data_o[16799] = data_o[31];
  assign data_o[16863] = data_o[31];
  assign data_o[16927] = data_o[31];
  assign data_o[16991] = data_o[31];
  assign data_o[17055] = data_o[31];
  assign data_o[17119] = data_o[31];
  assign data_o[17183] = data_o[31];
  assign data_o[17247] = data_o[31];
  assign data_o[17311] = data_o[31];
  assign data_o[17375] = data_o[31];
  assign data_o[17439] = data_o[31];
  assign data_o[17503] = data_o[31];
  assign data_o[17567] = data_o[31];
  assign data_o[17631] = data_o[31];
  assign data_o[17695] = data_o[31];
  assign data_o[17759] = data_o[31];
  assign data_o[17823] = data_o[31];
  assign data_o[17887] = data_o[31];
  assign data_o[17951] = data_o[31];
  assign data_o[18015] = data_o[31];
  assign data_o[18079] = data_o[31];
  assign data_o[18143] = data_o[31];
  assign data_o[18207] = data_o[31];
  assign data_o[18271] = data_o[31];
  assign data_o[18335] = data_o[31];
  assign data_o[18399] = data_o[31];
  assign data_o[18463] = data_o[31];
  assign data_o[18527] = data_o[31];
  assign data_o[18591] = data_o[31];
  assign data_o[18655] = data_o[31];
  assign data_o[18719] = data_o[31];
  assign data_o[18783] = data_o[31];
  assign data_o[18847] = data_o[31];
  assign data_o[18911] = data_o[31];
  assign data_o[18975] = data_o[31];
  assign data_o[19039] = data_o[31];
  assign data_o[19103] = data_o[31];
  assign data_o[19167] = data_o[31];
  assign data_o[19231] = data_o[31];
  assign data_o[19295] = data_o[31];
  assign data_o[19359] = data_o[31];
  assign data_o[19423] = data_o[31];
  assign data_o[19487] = data_o[31];
  assign data_o[19551] = data_o[31];
  assign data_o[19615] = data_o[31];
  assign data_o[19679] = data_o[31];
  assign data_o[19743] = data_o[31];
  assign data_o[19807] = data_o[31];
  assign data_o[19871] = data_o[31];
  assign data_o[19935] = data_o[31];
  assign data_o[19999] = data_o[31];
  assign data_o[20063] = data_o[31];
  assign data_o[20127] = data_o[31];
  assign data_o[20191] = data_o[31];
  assign data_o[20255] = data_o[31];
  assign data_o[20319] = data_o[31];
  assign data_o[20383] = data_o[31];
  assign data_o[20447] = data_o[31];
  assign data_o[20511] = data_o[31];
  assign data_o[20575] = data_o[31];
  assign data_o[20639] = data_o[31];
  assign data_o[20703] = data_o[31];
  assign data_o[20767] = data_o[31];
  assign data_o[20831] = data_o[31];
  assign data_o[20895] = data_o[31];
  assign data_o[20959] = data_o[31];
  assign data_o[21023] = data_o[31];
  assign data_o[21087] = data_o[31];
  assign data_o[21151] = data_o[31];
  assign data_o[21215] = data_o[31];
  assign data_o[21279] = data_o[31];
  assign data_o[21343] = data_o[31];
  assign data_o[21407] = data_o[31];
  assign data_o[21471] = data_o[31];
  assign data_o[21535] = data_o[31];
  assign data_o[21599] = data_o[31];
  assign data_o[21663] = data_o[31];
  assign data_o[21727] = data_o[31];
  assign data_o[21791] = data_o[31];
  assign data_o[21855] = data_o[31];
  assign data_o[21919] = data_o[31];
  assign data_o[21983] = data_o[31];
  assign data_o[22047] = data_o[31];
  assign data_o[22111] = data_o[31];
  assign data_o[22175] = data_o[31];
  assign data_o[22239] = data_o[31];
  assign data_o[22303] = data_o[31];
  assign data_o[22367] = data_o[31];
  assign data_o[22431] = data_o[31];
  assign data_o[22495] = data_o[31];
  assign data_o[22559] = data_o[31];
  assign data_o[22623] = data_o[31];
  assign data_o[22687] = data_o[31];
  assign data_o[22751] = data_o[31];
  assign data_o[22815] = data_o[31];
  assign data_o[22879] = data_o[31];
  assign data_o[22943] = data_o[31];
  assign data_o[23007] = data_o[31];
  assign data_o[23071] = data_o[31];
  assign data_o[23135] = data_o[31];
  assign data_o[23199] = data_o[31];
  assign data_o[23263] = data_o[31];
  assign data_o[23327] = data_o[31];
  assign data_o[23391] = data_o[31];
  assign data_o[23455] = data_o[31];
  assign data_o[23519] = data_o[31];
  assign data_o[23583] = data_o[31];
  assign data_o[23647] = data_o[31];
  assign data_o[23711] = data_o[31];
  assign data_o[23775] = data_o[31];
  assign data_o[23839] = data_o[31];
  assign data_o[23903] = data_o[31];
  assign data_o[23967] = data_o[31];
  assign data_o[24031] = data_o[31];
  assign data_o[24095] = data_o[31];
  assign data_o[24159] = data_o[31];
  assign data_o[24223] = data_o[31];
  assign data_o[24287] = data_o[31];
  assign data_o[24351] = data_o[31];
  assign data_o[24415] = data_o[31];
  assign data_o[24479] = data_o[31];
  assign data_o[24543] = data_o[31];
  assign data_o[24607] = data_o[31];
  assign data_o[24671] = data_o[31];
  assign data_o[24735] = data_o[31];
  assign data_o[24799] = data_o[31];
  assign data_o[24863] = data_o[31];
  assign data_o[24927] = data_o[31];
  assign data_o[24991] = data_o[31];
  assign data_o[25055] = data_o[31];
  assign data_o[25119] = data_o[31];
  assign data_o[25183] = data_o[31];
  assign data_o[25247] = data_o[31];
  assign data_o[25311] = data_o[31];
  assign data_o[25375] = data_o[31];
  assign data_o[25439] = data_o[31];
  assign data_o[25503] = data_o[31];
  assign data_o[25567] = data_o[31];
  assign data_o[25631] = data_o[31];
  assign data_o[25695] = data_o[31];
  assign data_o[25759] = data_o[31];
  assign data_o[25823] = data_o[31];
  assign data_o[25887] = data_o[31];
  assign data_o[25951] = data_o[31];
  assign data_o[26015] = data_o[31];
  assign data_o[26079] = data_o[31];
  assign data_o[26143] = data_o[31];
  assign data_o[26207] = data_o[31];
  assign data_o[26271] = data_o[31];
  assign data_o[26335] = data_o[31];
  assign data_o[26399] = data_o[31];
  assign data_o[26463] = data_o[31];
  assign data_o[26527] = data_o[31];
  assign data_o[26591] = data_o[31];
  assign data_o[26655] = data_o[31];
  assign data_o[26719] = data_o[31];
  assign data_o[26783] = data_o[31];
  assign data_o[26847] = data_o[31];
  assign data_o[26911] = data_o[31];
  assign data_o[26975] = data_o[31];
  assign data_o[27039] = data_o[31];
  assign data_o[27103] = data_o[31];
  assign data_o[27167] = data_o[31];
  assign data_o[27231] = data_o[31];
  assign data_o[27295] = data_o[31];
  assign data_o[27359] = data_o[31];
  assign data_o[27423] = data_o[31];
  assign data_o[27487] = data_o[31];
  assign data_o[27551] = data_o[31];
  assign data_o[27615] = data_o[31];
  assign data_o[27679] = data_o[31];
  assign data_o[27743] = data_o[31];
  assign data_o[27807] = data_o[31];
  assign data_o[27871] = data_o[31];
  assign data_o[27935] = data_o[31];
  assign data_o[27999] = data_o[31];
  assign data_o[28063] = data_o[31];
  assign data_o[28127] = data_o[31];
  assign data_o[28191] = data_o[31];
  assign data_o[28255] = data_o[31];
  assign data_o[28319] = data_o[31];
  assign data_o[28383] = data_o[31];
  assign data_o[28447] = data_o[31];
  assign data_o[28511] = data_o[31];
  assign data_o[28575] = data_o[31];
  assign data_o[28639] = data_o[31];
  assign data_o[28703] = data_o[31];
  assign data_o[28767] = data_o[31];
  assign data_o[28831] = data_o[31];
  assign data_o[28895] = data_o[31];
  assign data_o[28959] = data_o[31];
  assign data_o[29023] = data_o[31];
  assign data_o[29087] = data_o[31];
  assign data_o[29151] = data_o[31];
  assign data_o[29215] = data_o[31];
  assign data_o[29279] = data_o[31];
  assign data_o[29343] = data_o[31];
  assign data_o[29407] = data_o[31];
  assign data_o[29471] = data_o[31];
  assign data_o[29535] = data_o[31];
  assign data_o[29599] = data_o[31];
  assign data_o[29663] = data_o[31];
  assign data_o[29727] = data_o[31];
  assign data_o[29791] = data_o[31];
  assign data_o[29855] = data_o[31];
  assign data_o[29919] = data_o[31];
  assign data_o[29983] = data_o[31];
  assign data_o[30047] = data_o[31];
  assign data_o[30111] = data_o[31];
  assign data_o[30175] = data_o[31];
  assign data_o[30239] = data_o[31];
  assign data_o[30303] = data_o[31];
  assign data_o[30367] = data_o[31];
  assign data_o[30431] = data_o[31];
  assign data_o[30495] = data_o[31];
  assign data_o[30559] = data_o[31];
  assign data_o[30623] = data_o[31];
  assign data_o[30687] = data_o[31];
  assign data_o[30751] = data_o[31];
  assign data_o[30815] = data_o[31];
  assign data_o[30879] = data_o[31];
  assign data_o[30943] = data_o[31];
  assign data_o[31007] = data_o[31];
  assign data_o[31071] = data_o[31];
  assign data_o[31135] = data_o[31];
  assign data_o[31199] = data_o[31];
  assign data_o[31263] = data_o[31];
  assign data_o[31327] = data_o[31];
  assign data_o[31391] = data_o[31];
  assign data_o[31455] = data_o[31];
  assign data_o[31519] = data_o[31];
  assign data_o[31583] = data_o[31];
  assign data_o[31647] = data_o[31];
  assign data_o[31711] = data_o[31];
  assign data_o[31775] = data_o[31];
  assign data_o[31839] = data_o[31];
  assign data_o[31903] = data_o[31];
  assign data_o[31967] = data_o[31];
  assign data_o[94] = data_o[30];
  assign data_o[158] = data_o[30];
  assign data_o[222] = data_o[30];
  assign data_o[286] = data_o[30];
  assign data_o[350] = data_o[30];
  assign data_o[414] = data_o[30];
  assign data_o[478] = data_o[30];
  assign data_o[542] = data_o[30];
  assign data_o[606] = data_o[30];
  assign data_o[670] = data_o[30];
  assign data_o[734] = data_o[30];
  assign data_o[798] = data_o[30];
  assign data_o[862] = data_o[30];
  assign data_o[926] = data_o[30];
  assign data_o[990] = data_o[30];
  assign data_o[1054] = data_o[30];
  assign data_o[1118] = data_o[30];
  assign data_o[1182] = data_o[30];
  assign data_o[1246] = data_o[30];
  assign data_o[1310] = data_o[30];
  assign data_o[1374] = data_o[30];
  assign data_o[1438] = data_o[30];
  assign data_o[1502] = data_o[30];
  assign data_o[1566] = data_o[30];
  assign data_o[1630] = data_o[30];
  assign data_o[1694] = data_o[30];
  assign data_o[1758] = data_o[30];
  assign data_o[1822] = data_o[30];
  assign data_o[1886] = data_o[30];
  assign data_o[1950] = data_o[30];
  assign data_o[2014] = data_o[30];
  assign data_o[2078] = data_o[30];
  assign data_o[2142] = data_o[30];
  assign data_o[2206] = data_o[30];
  assign data_o[2270] = data_o[30];
  assign data_o[2334] = data_o[30];
  assign data_o[2398] = data_o[30];
  assign data_o[2462] = data_o[30];
  assign data_o[2526] = data_o[30];
  assign data_o[2590] = data_o[30];
  assign data_o[2654] = data_o[30];
  assign data_o[2718] = data_o[30];
  assign data_o[2782] = data_o[30];
  assign data_o[2846] = data_o[30];
  assign data_o[2910] = data_o[30];
  assign data_o[2974] = data_o[30];
  assign data_o[3038] = data_o[30];
  assign data_o[3102] = data_o[30];
  assign data_o[3166] = data_o[30];
  assign data_o[3230] = data_o[30];
  assign data_o[3294] = data_o[30];
  assign data_o[3358] = data_o[30];
  assign data_o[3422] = data_o[30];
  assign data_o[3486] = data_o[30];
  assign data_o[3550] = data_o[30];
  assign data_o[3614] = data_o[30];
  assign data_o[3678] = data_o[30];
  assign data_o[3742] = data_o[30];
  assign data_o[3806] = data_o[30];
  assign data_o[3870] = data_o[30];
  assign data_o[3934] = data_o[30];
  assign data_o[3998] = data_o[30];
  assign data_o[4062] = data_o[30];
  assign data_o[4126] = data_o[30];
  assign data_o[4190] = data_o[30];
  assign data_o[4254] = data_o[30];
  assign data_o[4318] = data_o[30];
  assign data_o[4382] = data_o[30];
  assign data_o[4446] = data_o[30];
  assign data_o[4510] = data_o[30];
  assign data_o[4574] = data_o[30];
  assign data_o[4638] = data_o[30];
  assign data_o[4702] = data_o[30];
  assign data_o[4766] = data_o[30];
  assign data_o[4830] = data_o[30];
  assign data_o[4894] = data_o[30];
  assign data_o[4958] = data_o[30];
  assign data_o[5022] = data_o[30];
  assign data_o[5086] = data_o[30];
  assign data_o[5150] = data_o[30];
  assign data_o[5214] = data_o[30];
  assign data_o[5278] = data_o[30];
  assign data_o[5342] = data_o[30];
  assign data_o[5406] = data_o[30];
  assign data_o[5470] = data_o[30];
  assign data_o[5534] = data_o[30];
  assign data_o[5598] = data_o[30];
  assign data_o[5662] = data_o[30];
  assign data_o[5726] = data_o[30];
  assign data_o[5790] = data_o[30];
  assign data_o[5854] = data_o[30];
  assign data_o[5918] = data_o[30];
  assign data_o[5982] = data_o[30];
  assign data_o[6046] = data_o[30];
  assign data_o[6110] = data_o[30];
  assign data_o[6174] = data_o[30];
  assign data_o[6238] = data_o[30];
  assign data_o[6302] = data_o[30];
  assign data_o[6366] = data_o[30];
  assign data_o[6430] = data_o[30];
  assign data_o[6494] = data_o[30];
  assign data_o[6558] = data_o[30];
  assign data_o[6622] = data_o[30];
  assign data_o[6686] = data_o[30];
  assign data_o[6750] = data_o[30];
  assign data_o[6814] = data_o[30];
  assign data_o[6878] = data_o[30];
  assign data_o[6942] = data_o[30];
  assign data_o[7006] = data_o[30];
  assign data_o[7070] = data_o[30];
  assign data_o[7134] = data_o[30];
  assign data_o[7198] = data_o[30];
  assign data_o[7262] = data_o[30];
  assign data_o[7326] = data_o[30];
  assign data_o[7390] = data_o[30];
  assign data_o[7454] = data_o[30];
  assign data_o[7518] = data_o[30];
  assign data_o[7582] = data_o[30];
  assign data_o[7646] = data_o[30];
  assign data_o[7710] = data_o[30];
  assign data_o[7774] = data_o[30];
  assign data_o[7838] = data_o[30];
  assign data_o[7902] = data_o[30];
  assign data_o[7966] = data_o[30];
  assign data_o[8030] = data_o[30];
  assign data_o[8094] = data_o[30];
  assign data_o[8158] = data_o[30];
  assign data_o[8222] = data_o[30];
  assign data_o[8286] = data_o[30];
  assign data_o[8350] = data_o[30];
  assign data_o[8414] = data_o[30];
  assign data_o[8478] = data_o[30];
  assign data_o[8542] = data_o[30];
  assign data_o[8606] = data_o[30];
  assign data_o[8670] = data_o[30];
  assign data_o[8734] = data_o[30];
  assign data_o[8798] = data_o[30];
  assign data_o[8862] = data_o[30];
  assign data_o[8926] = data_o[30];
  assign data_o[8990] = data_o[30];
  assign data_o[9054] = data_o[30];
  assign data_o[9118] = data_o[30];
  assign data_o[9182] = data_o[30];
  assign data_o[9246] = data_o[30];
  assign data_o[9310] = data_o[30];
  assign data_o[9374] = data_o[30];
  assign data_o[9438] = data_o[30];
  assign data_o[9502] = data_o[30];
  assign data_o[9566] = data_o[30];
  assign data_o[9630] = data_o[30];
  assign data_o[9694] = data_o[30];
  assign data_o[9758] = data_o[30];
  assign data_o[9822] = data_o[30];
  assign data_o[9886] = data_o[30];
  assign data_o[9950] = data_o[30];
  assign data_o[10014] = data_o[30];
  assign data_o[10078] = data_o[30];
  assign data_o[10142] = data_o[30];
  assign data_o[10206] = data_o[30];
  assign data_o[10270] = data_o[30];
  assign data_o[10334] = data_o[30];
  assign data_o[10398] = data_o[30];
  assign data_o[10462] = data_o[30];
  assign data_o[10526] = data_o[30];
  assign data_o[10590] = data_o[30];
  assign data_o[10654] = data_o[30];
  assign data_o[10718] = data_o[30];
  assign data_o[10782] = data_o[30];
  assign data_o[10846] = data_o[30];
  assign data_o[10910] = data_o[30];
  assign data_o[10974] = data_o[30];
  assign data_o[11038] = data_o[30];
  assign data_o[11102] = data_o[30];
  assign data_o[11166] = data_o[30];
  assign data_o[11230] = data_o[30];
  assign data_o[11294] = data_o[30];
  assign data_o[11358] = data_o[30];
  assign data_o[11422] = data_o[30];
  assign data_o[11486] = data_o[30];
  assign data_o[11550] = data_o[30];
  assign data_o[11614] = data_o[30];
  assign data_o[11678] = data_o[30];
  assign data_o[11742] = data_o[30];
  assign data_o[11806] = data_o[30];
  assign data_o[11870] = data_o[30];
  assign data_o[11934] = data_o[30];
  assign data_o[11998] = data_o[30];
  assign data_o[12062] = data_o[30];
  assign data_o[12126] = data_o[30];
  assign data_o[12190] = data_o[30];
  assign data_o[12254] = data_o[30];
  assign data_o[12318] = data_o[30];
  assign data_o[12382] = data_o[30];
  assign data_o[12446] = data_o[30];
  assign data_o[12510] = data_o[30];
  assign data_o[12574] = data_o[30];
  assign data_o[12638] = data_o[30];
  assign data_o[12702] = data_o[30];
  assign data_o[12766] = data_o[30];
  assign data_o[12830] = data_o[30];
  assign data_o[12894] = data_o[30];
  assign data_o[12958] = data_o[30];
  assign data_o[13022] = data_o[30];
  assign data_o[13086] = data_o[30];
  assign data_o[13150] = data_o[30];
  assign data_o[13214] = data_o[30];
  assign data_o[13278] = data_o[30];
  assign data_o[13342] = data_o[30];
  assign data_o[13406] = data_o[30];
  assign data_o[13470] = data_o[30];
  assign data_o[13534] = data_o[30];
  assign data_o[13598] = data_o[30];
  assign data_o[13662] = data_o[30];
  assign data_o[13726] = data_o[30];
  assign data_o[13790] = data_o[30];
  assign data_o[13854] = data_o[30];
  assign data_o[13918] = data_o[30];
  assign data_o[13982] = data_o[30];
  assign data_o[14046] = data_o[30];
  assign data_o[14110] = data_o[30];
  assign data_o[14174] = data_o[30];
  assign data_o[14238] = data_o[30];
  assign data_o[14302] = data_o[30];
  assign data_o[14366] = data_o[30];
  assign data_o[14430] = data_o[30];
  assign data_o[14494] = data_o[30];
  assign data_o[14558] = data_o[30];
  assign data_o[14622] = data_o[30];
  assign data_o[14686] = data_o[30];
  assign data_o[14750] = data_o[30];
  assign data_o[14814] = data_o[30];
  assign data_o[14878] = data_o[30];
  assign data_o[14942] = data_o[30];
  assign data_o[15006] = data_o[30];
  assign data_o[15070] = data_o[30];
  assign data_o[15134] = data_o[30];
  assign data_o[15198] = data_o[30];
  assign data_o[15262] = data_o[30];
  assign data_o[15326] = data_o[30];
  assign data_o[15390] = data_o[30];
  assign data_o[15454] = data_o[30];
  assign data_o[15518] = data_o[30];
  assign data_o[15582] = data_o[30];
  assign data_o[15646] = data_o[30];
  assign data_o[15710] = data_o[30];
  assign data_o[15774] = data_o[30];
  assign data_o[15838] = data_o[30];
  assign data_o[15902] = data_o[30];
  assign data_o[15966] = data_o[30];
  assign data_o[16030] = data_o[30];
  assign data_o[16094] = data_o[30];
  assign data_o[16158] = data_o[30];
  assign data_o[16222] = data_o[30];
  assign data_o[16286] = data_o[30];
  assign data_o[16350] = data_o[30];
  assign data_o[16414] = data_o[30];
  assign data_o[16478] = data_o[30];
  assign data_o[16542] = data_o[30];
  assign data_o[16606] = data_o[30];
  assign data_o[16670] = data_o[30];
  assign data_o[16734] = data_o[30];
  assign data_o[16798] = data_o[30];
  assign data_o[16862] = data_o[30];
  assign data_o[16926] = data_o[30];
  assign data_o[16990] = data_o[30];
  assign data_o[17054] = data_o[30];
  assign data_o[17118] = data_o[30];
  assign data_o[17182] = data_o[30];
  assign data_o[17246] = data_o[30];
  assign data_o[17310] = data_o[30];
  assign data_o[17374] = data_o[30];
  assign data_o[17438] = data_o[30];
  assign data_o[17502] = data_o[30];
  assign data_o[17566] = data_o[30];
  assign data_o[17630] = data_o[30];
  assign data_o[17694] = data_o[30];
  assign data_o[17758] = data_o[30];
  assign data_o[17822] = data_o[30];
  assign data_o[17886] = data_o[30];
  assign data_o[17950] = data_o[30];
  assign data_o[18014] = data_o[30];
  assign data_o[18078] = data_o[30];
  assign data_o[18142] = data_o[30];
  assign data_o[18206] = data_o[30];
  assign data_o[18270] = data_o[30];
  assign data_o[18334] = data_o[30];
  assign data_o[18398] = data_o[30];
  assign data_o[18462] = data_o[30];
  assign data_o[18526] = data_o[30];
  assign data_o[18590] = data_o[30];
  assign data_o[18654] = data_o[30];
  assign data_o[18718] = data_o[30];
  assign data_o[18782] = data_o[30];
  assign data_o[18846] = data_o[30];
  assign data_o[18910] = data_o[30];
  assign data_o[18974] = data_o[30];
  assign data_o[19038] = data_o[30];
  assign data_o[19102] = data_o[30];
  assign data_o[19166] = data_o[30];
  assign data_o[19230] = data_o[30];
  assign data_o[19294] = data_o[30];
  assign data_o[19358] = data_o[30];
  assign data_o[19422] = data_o[30];
  assign data_o[19486] = data_o[30];
  assign data_o[19550] = data_o[30];
  assign data_o[19614] = data_o[30];
  assign data_o[19678] = data_o[30];
  assign data_o[19742] = data_o[30];
  assign data_o[19806] = data_o[30];
  assign data_o[19870] = data_o[30];
  assign data_o[19934] = data_o[30];
  assign data_o[19998] = data_o[30];
  assign data_o[20062] = data_o[30];
  assign data_o[20126] = data_o[30];
  assign data_o[20190] = data_o[30];
  assign data_o[20254] = data_o[30];
  assign data_o[20318] = data_o[30];
  assign data_o[20382] = data_o[30];
  assign data_o[20446] = data_o[30];
  assign data_o[20510] = data_o[30];
  assign data_o[20574] = data_o[30];
  assign data_o[20638] = data_o[30];
  assign data_o[20702] = data_o[30];
  assign data_o[20766] = data_o[30];
  assign data_o[20830] = data_o[30];
  assign data_o[20894] = data_o[30];
  assign data_o[20958] = data_o[30];
  assign data_o[21022] = data_o[30];
  assign data_o[21086] = data_o[30];
  assign data_o[21150] = data_o[30];
  assign data_o[21214] = data_o[30];
  assign data_o[21278] = data_o[30];
  assign data_o[21342] = data_o[30];
  assign data_o[21406] = data_o[30];
  assign data_o[21470] = data_o[30];
  assign data_o[21534] = data_o[30];
  assign data_o[21598] = data_o[30];
  assign data_o[21662] = data_o[30];
  assign data_o[21726] = data_o[30];
  assign data_o[21790] = data_o[30];
  assign data_o[21854] = data_o[30];
  assign data_o[21918] = data_o[30];
  assign data_o[21982] = data_o[30];
  assign data_o[22046] = data_o[30];
  assign data_o[22110] = data_o[30];
  assign data_o[22174] = data_o[30];
  assign data_o[22238] = data_o[30];
  assign data_o[22302] = data_o[30];
  assign data_o[22366] = data_o[30];
  assign data_o[22430] = data_o[30];
  assign data_o[22494] = data_o[30];
  assign data_o[22558] = data_o[30];
  assign data_o[22622] = data_o[30];
  assign data_o[22686] = data_o[30];
  assign data_o[22750] = data_o[30];
  assign data_o[22814] = data_o[30];
  assign data_o[22878] = data_o[30];
  assign data_o[22942] = data_o[30];
  assign data_o[23006] = data_o[30];
  assign data_o[23070] = data_o[30];
  assign data_o[23134] = data_o[30];
  assign data_o[23198] = data_o[30];
  assign data_o[23262] = data_o[30];
  assign data_o[23326] = data_o[30];
  assign data_o[23390] = data_o[30];
  assign data_o[23454] = data_o[30];
  assign data_o[23518] = data_o[30];
  assign data_o[23582] = data_o[30];
  assign data_o[23646] = data_o[30];
  assign data_o[23710] = data_o[30];
  assign data_o[23774] = data_o[30];
  assign data_o[23838] = data_o[30];
  assign data_o[23902] = data_o[30];
  assign data_o[23966] = data_o[30];
  assign data_o[24030] = data_o[30];
  assign data_o[24094] = data_o[30];
  assign data_o[24158] = data_o[30];
  assign data_o[24222] = data_o[30];
  assign data_o[24286] = data_o[30];
  assign data_o[24350] = data_o[30];
  assign data_o[24414] = data_o[30];
  assign data_o[24478] = data_o[30];
  assign data_o[24542] = data_o[30];
  assign data_o[24606] = data_o[30];
  assign data_o[24670] = data_o[30];
  assign data_o[24734] = data_o[30];
  assign data_o[24798] = data_o[30];
  assign data_o[24862] = data_o[30];
  assign data_o[24926] = data_o[30];
  assign data_o[24990] = data_o[30];
  assign data_o[25054] = data_o[30];
  assign data_o[25118] = data_o[30];
  assign data_o[25182] = data_o[30];
  assign data_o[25246] = data_o[30];
  assign data_o[25310] = data_o[30];
  assign data_o[25374] = data_o[30];
  assign data_o[25438] = data_o[30];
  assign data_o[25502] = data_o[30];
  assign data_o[25566] = data_o[30];
  assign data_o[25630] = data_o[30];
  assign data_o[25694] = data_o[30];
  assign data_o[25758] = data_o[30];
  assign data_o[25822] = data_o[30];
  assign data_o[25886] = data_o[30];
  assign data_o[25950] = data_o[30];
  assign data_o[26014] = data_o[30];
  assign data_o[26078] = data_o[30];
  assign data_o[26142] = data_o[30];
  assign data_o[26206] = data_o[30];
  assign data_o[26270] = data_o[30];
  assign data_o[26334] = data_o[30];
  assign data_o[26398] = data_o[30];
  assign data_o[26462] = data_o[30];
  assign data_o[26526] = data_o[30];
  assign data_o[26590] = data_o[30];
  assign data_o[26654] = data_o[30];
  assign data_o[26718] = data_o[30];
  assign data_o[26782] = data_o[30];
  assign data_o[26846] = data_o[30];
  assign data_o[26910] = data_o[30];
  assign data_o[26974] = data_o[30];
  assign data_o[27038] = data_o[30];
  assign data_o[27102] = data_o[30];
  assign data_o[27166] = data_o[30];
  assign data_o[27230] = data_o[30];
  assign data_o[27294] = data_o[30];
  assign data_o[27358] = data_o[30];
  assign data_o[27422] = data_o[30];
  assign data_o[27486] = data_o[30];
  assign data_o[27550] = data_o[30];
  assign data_o[27614] = data_o[30];
  assign data_o[27678] = data_o[30];
  assign data_o[27742] = data_o[30];
  assign data_o[27806] = data_o[30];
  assign data_o[27870] = data_o[30];
  assign data_o[27934] = data_o[30];
  assign data_o[27998] = data_o[30];
  assign data_o[28062] = data_o[30];
  assign data_o[28126] = data_o[30];
  assign data_o[28190] = data_o[30];
  assign data_o[28254] = data_o[30];
  assign data_o[28318] = data_o[30];
  assign data_o[28382] = data_o[30];
  assign data_o[28446] = data_o[30];
  assign data_o[28510] = data_o[30];
  assign data_o[28574] = data_o[30];
  assign data_o[28638] = data_o[30];
  assign data_o[28702] = data_o[30];
  assign data_o[28766] = data_o[30];
  assign data_o[28830] = data_o[30];
  assign data_o[28894] = data_o[30];
  assign data_o[28958] = data_o[30];
  assign data_o[29022] = data_o[30];
  assign data_o[29086] = data_o[30];
  assign data_o[29150] = data_o[30];
  assign data_o[29214] = data_o[30];
  assign data_o[29278] = data_o[30];
  assign data_o[29342] = data_o[30];
  assign data_o[29406] = data_o[30];
  assign data_o[29470] = data_o[30];
  assign data_o[29534] = data_o[30];
  assign data_o[29598] = data_o[30];
  assign data_o[29662] = data_o[30];
  assign data_o[29726] = data_o[30];
  assign data_o[29790] = data_o[30];
  assign data_o[29854] = data_o[30];
  assign data_o[29918] = data_o[30];
  assign data_o[29982] = data_o[30];
  assign data_o[30046] = data_o[30];
  assign data_o[30110] = data_o[30];
  assign data_o[30174] = data_o[30];
  assign data_o[30238] = data_o[30];
  assign data_o[30302] = data_o[30];
  assign data_o[30366] = data_o[30];
  assign data_o[30430] = data_o[30];
  assign data_o[30494] = data_o[30];
  assign data_o[30558] = data_o[30];
  assign data_o[30622] = data_o[30];
  assign data_o[30686] = data_o[30];
  assign data_o[30750] = data_o[30];
  assign data_o[30814] = data_o[30];
  assign data_o[30878] = data_o[30];
  assign data_o[30942] = data_o[30];
  assign data_o[31006] = data_o[30];
  assign data_o[31070] = data_o[30];
  assign data_o[31134] = data_o[30];
  assign data_o[31198] = data_o[30];
  assign data_o[31262] = data_o[30];
  assign data_o[31326] = data_o[30];
  assign data_o[31390] = data_o[30];
  assign data_o[31454] = data_o[30];
  assign data_o[31518] = data_o[30];
  assign data_o[31582] = data_o[30];
  assign data_o[31646] = data_o[30];
  assign data_o[31710] = data_o[30];
  assign data_o[31774] = data_o[30];
  assign data_o[31838] = data_o[30];
  assign data_o[31902] = data_o[30];
  assign data_o[31966] = data_o[30];
  assign data_o[93] = data_o[29];
  assign data_o[157] = data_o[29];
  assign data_o[221] = data_o[29];
  assign data_o[285] = data_o[29];
  assign data_o[349] = data_o[29];
  assign data_o[413] = data_o[29];
  assign data_o[477] = data_o[29];
  assign data_o[541] = data_o[29];
  assign data_o[605] = data_o[29];
  assign data_o[669] = data_o[29];
  assign data_o[733] = data_o[29];
  assign data_o[797] = data_o[29];
  assign data_o[861] = data_o[29];
  assign data_o[925] = data_o[29];
  assign data_o[989] = data_o[29];
  assign data_o[1053] = data_o[29];
  assign data_o[1117] = data_o[29];
  assign data_o[1181] = data_o[29];
  assign data_o[1245] = data_o[29];
  assign data_o[1309] = data_o[29];
  assign data_o[1373] = data_o[29];
  assign data_o[1437] = data_o[29];
  assign data_o[1501] = data_o[29];
  assign data_o[1565] = data_o[29];
  assign data_o[1629] = data_o[29];
  assign data_o[1693] = data_o[29];
  assign data_o[1757] = data_o[29];
  assign data_o[1821] = data_o[29];
  assign data_o[1885] = data_o[29];
  assign data_o[1949] = data_o[29];
  assign data_o[2013] = data_o[29];
  assign data_o[2077] = data_o[29];
  assign data_o[2141] = data_o[29];
  assign data_o[2205] = data_o[29];
  assign data_o[2269] = data_o[29];
  assign data_o[2333] = data_o[29];
  assign data_o[2397] = data_o[29];
  assign data_o[2461] = data_o[29];
  assign data_o[2525] = data_o[29];
  assign data_o[2589] = data_o[29];
  assign data_o[2653] = data_o[29];
  assign data_o[2717] = data_o[29];
  assign data_o[2781] = data_o[29];
  assign data_o[2845] = data_o[29];
  assign data_o[2909] = data_o[29];
  assign data_o[2973] = data_o[29];
  assign data_o[3037] = data_o[29];
  assign data_o[3101] = data_o[29];
  assign data_o[3165] = data_o[29];
  assign data_o[3229] = data_o[29];
  assign data_o[3293] = data_o[29];
  assign data_o[3357] = data_o[29];
  assign data_o[3421] = data_o[29];
  assign data_o[3485] = data_o[29];
  assign data_o[3549] = data_o[29];
  assign data_o[3613] = data_o[29];
  assign data_o[3677] = data_o[29];
  assign data_o[3741] = data_o[29];
  assign data_o[3805] = data_o[29];
  assign data_o[3869] = data_o[29];
  assign data_o[3933] = data_o[29];
  assign data_o[3997] = data_o[29];
  assign data_o[4061] = data_o[29];
  assign data_o[4125] = data_o[29];
  assign data_o[4189] = data_o[29];
  assign data_o[4253] = data_o[29];
  assign data_o[4317] = data_o[29];
  assign data_o[4381] = data_o[29];
  assign data_o[4445] = data_o[29];
  assign data_o[4509] = data_o[29];
  assign data_o[4573] = data_o[29];
  assign data_o[4637] = data_o[29];
  assign data_o[4701] = data_o[29];
  assign data_o[4765] = data_o[29];
  assign data_o[4829] = data_o[29];
  assign data_o[4893] = data_o[29];
  assign data_o[4957] = data_o[29];
  assign data_o[5021] = data_o[29];
  assign data_o[5085] = data_o[29];
  assign data_o[5149] = data_o[29];
  assign data_o[5213] = data_o[29];
  assign data_o[5277] = data_o[29];
  assign data_o[5341] = data_o[29];
  assign data_o[5405] = data_o[29];
  assign data_o[5469] = data_o[29];
  assign data_o[5533] = data_o[29];
  assign data_o[5597] = data_o[29];
  assign data_o[5661] = data_o[29];
  assign data_o[5725] = data_o[29];
  assign data_o[5789] = data_o[29];
  assign data_o[5853] = data_o[29];
  assign data_o[5917] = data_o[29];
  assign data_o[5981] = data_o[29];
  assign data_o[6045] = data_o[29];
  assign data_o[6109] = data_o[29];
  assign data_o[6173] = data_o[29];
  assign data_o[6237] = data_o[29];
  assign data_o[6301] = data_o[29];
  assign data_o[6365] = data_o[29];
  assign data_o[6429] = data_o[29];
  assign data_o[6493] = data_o[29];
  assign data_o[6557] = data_o[29];
  assign data_o[6621] = data_o[29];
  assign data_o[6685] = data_o[29];
  assign data_o[6749] = data_o[29];
  assign data_o[6813] = data_o[29];
  assign data_o[6877] = data_o[29];
  assign data_o[6941] = data_o[29];
  assign data_o[7005] = data_o[29];
  assign data_o[7069] = data_o[29];
  assign data_o[7133] = data_o[29];
  assign data_o[7197] = data_o[29];
  assign data_o[7261] = data_o[29];
  assign data_o[7325] = data_o[29];
  assign data_o[7389] = data_o[29];
  assign data_o[7453] = data_o[29];
  assign data_o[7517] = data_o[29];
  assign data_o[7581] = data_o[29];
  assign data_o[7645] = data_o[29];
  assign data_o[7709] = data_o[29];
  assign data_o[7773] = data_o[29];
  assign data_o[7837] = data_o[29];
  assign data_o[7901] = data_o[29];
  assign data_o[7965] = data_o[29];
  assign data_o[8029] = data_o[29];
  assign data_o[8093] = data_o[29];
  assign data_o[8157] = data_o[29];
  assign data_o[8221] = data_o[29];
  assign data_o[8285] = data_o[29];
  assign data_o[8349] = data_o[29];
  assign data_o[8413] = data_o[29];
  assign data_o[8477] = data_o[29];
  assign data_o[8541] = data_o[29];
  assign data_o[8605] = data_o[29];
  assign data_o[8669] = data_o[29];
  assign data_o[8733] = data_o[29];
  assign data_o[8797] = data_o[29];
  assign data_o[8861] = data_o[29];
  assign data_o[8925] = data_o[29];
  assign data_o[8989] = data_o[29];
  assign data_o[9053] = data_o[29];
  assign data_o[9117] = data_o[29];
  assign data_o[9181] = data_o[29];
  assign data_o[9245] = data_o[29];
  assign data_o[9309] = data_o[29];
  assign data_o[9373] = data_o[29];
  assign data_o[9437] = data_o[29];
  assign data_o[9501] = data_o[29];
  assign data_o[9565] = data_o[29];
  assign data_o[9629] = data_o[29];
  assign data_o[9693] = data_o[29];
  assign data_o[9757] = data_o[29];
  assign data_o[9821] = data_o[29];
  assign data_o[9885] = data_o[29];
  assign data_o[9949] = data_o[29];
  assign data_o[10013] = data_o[29];
  assign data_o[10077] = data_o[29];
  assign data_o[10141] = data_o[29];
  assign data_o[10205] = data_o[29];
  assign data_o[10269] = data_o[29];
  assign data_o[10333] = data_o[29];
  assign data_o[10397] = data_o[29];
  assign data_o[10461] = data_o[29];
  assign data_o[10525] = data_o[29];
  assign data_o[10589] = data_o[29];
  assign data_o[10653] = data_o[29];
  assign data_o[10717] = data_o[29];
  assign data_o[10781] = data_o[29];
  assign data_o[10845] = data_o[29];
  assign data_o[10909] = data_o[29];
  assign data_o[10973] = data_o[29];
  assign data_o[11037] = data_o[29];
  assign data_o[11101] = data_o[29];
  assign data_o[11165] = data_o[29];
  assign data_o[11229] = data_o[29];
  assign data_o[11293] = data_o[29];
  assign data_o[11357] = data_o[29];
  assign data_o[11421] = data_o[29];
  assign data_o[11485] = data_o[29];
  assign data_o[11549] = data_o[29];
  assign data_o[11613] = data_o[29];
  assign data_o[11677] = data_o[29];
  assign data_o[11741] = data_o[29];
  assign data_o[11805] = data_o[29];
  assign data_o[11869] = data_o[29];
  assign data_o[11933] = data_o[29];
  assign data_o[11997] = data_o[29];
  assign data_o[12061] = data_o[29];
  assign data_o[12125] = data_o[29];
  assign data_o[12189] = data_o[29];
  assign data_o[12253] = data_o[29];
  assign data_o[12317] = data_o[29];
  assign data_o[12381] = data_o[29];
  assign data_o[12445] = data_o[29];
  assign data_o[12509] = data_o[29];
  assign data_o[12573] = data_o[29];
  assign data_o[12637] = data_o[29];
  assign data_o[12701] = data_o[29];
  assign data_o[12765] = data_o[29];
  assign data_o[12829] = data_o[29];
  assign data_o[12893] = data_o[29];
  assign data_o[12957] = data_o[29];
  assign data_o[13021] = data_o[29];
  assign data_o[13085] = data_o[29];
  assign data_o[13149] = data_o[29];
  assign data_o[13213] = data_o[29];
  assign data_o[13277] = data_o[29];
  assign data_o[13341] = data_o[29];
  assign data_o[13405] = data_o[29];
  assign data_o[13469] = data_o[29];
  assign data_o[13533] = data_o[29];
  assign data_o[13597] = data_o[29];
  assign data_o[13661] = data_o[29];
  assign data_o[13725] = data_o[29];
  assign data_o[13789] = data_o[29];
  assign data_o[13853] = data_o[29];
  assign data_o[13917] = data_o[29];
  assign data_o[13981] = data_o[29];
  assign data_o[14045] = data_o[29];
  assign data_o[14109] = data_o[29];
  assign data_o[14173] = data_o[29];
  assign data_o[14237] = data_o[29];
  assign data_o[14301] = data_o[29];
  assign data_o[14365] = data_o[29];
  assign data_o[14429] = data_o[29];
  assign data_o[14493] = data_o[29];
  assign data_o[14557] = data_o[29];
  assign data_o[14621] = data_o[29];
  assign data_o[14685] = data_o[29];
  assign data_o[14749] = data_o[29];
  assign data_o[14813] = data_o[29];
  assign data_o[14877] = data_o[29];
  assign data_o[14941] = data_o[29];
  assign data_o[15005] = data_o[29];
  assign data_o[15069] = data_o[29];
  assign data_o[15133] = data_o[29];
  assign data_o[15197] = data_o[29];
  assign data_o[15261] = data_o[29];
  assign data_o[15325] = data_o[29];
  assign data_o[15389] = data_o[29];
  assign data_o[15453] = data_o[29];
  assign data_o[15517] = data_o[29];
  assign data_o[15581] = data_o[29];
  assign data_o[15645] = data_o[29];
  assign data_o[15709] = data_o[29];
  assign data_o[15773] = data_o[29];
  assign data_o[15837] = data_o[29];
  assign data_o[15901] = data_o[29];
  assign data_o[15965] = data_o[29];
  assign data_o[16029] = data_o[29];
  assign data_o[16093] = data_o[29];
  assign data_o[16157] = data_o[29];
  assign data_o[16221] = data_o[29];
  assign data_o[16285] = data_o[29];
  assign data_o[16349] = data_o[29];
  assign data_o[16413] = data_o[29];
  assign data_o[16477] = data_o[29];
  assign data_o[16541] = data_o[29];
  assign data_o[16605] = data_o[29];
  assign data_o[16669] = data_o[29];
  assign data_o[16733] = data_o[29];
  assign data_o[16797] = data_o[29];
  assign data_o[16861] = data_o[29];
  assign data_o[16925] = data_o[29];
  assign data_o[16989] = data_o[29];
  assign data_o[17053] = data_o[29];
  assign data_o[17117] = data_o[29];
  assign data_o[17181] = data_o[29];
  assign data_o[17245] = data_o[29];
  assign data_o[17309] = data_o[29];
  assign data_o[17373] = data_o[29];
  assign data_o[17437] = data_o[29];
  assign data_o[17501] = data_o[29];
  assign data_o[17565] = data_o[29];
  assign data_o[17629] = data_o[29];
  assign data_o[17693] = data_o[29];
  assign data_o[17757] = data_o[29];
  assign data_o[17821] = data_o[29];
  assign data_o[17885] = data_o[29];
  assign data_o[17949] = data_o[29];
  assign data_o[18013] = data_o[29];
  assign data_o[18077] = data_o[29];
  assign data_o[18141] = data_o[29];
  assign data_o[18205] = data_o[29];
  assign data_o[18269] = data_o[29];
  assign data_o[18333] = data_o[29];
  assign data_o[18397] = data_o[29];
  assign data_o[18461] = data_o[29];
  assign data_o[18525] = data_o[29];
  assign data_o[18589] = data_o[29];
  assign data_o[18653] = data_o[29];
  assign data_o[18717] = data_o[29];
  assign data_o[18781] = data_o[29];
  assign data_o[18845] = data_o[29];
  assign data_o[18909] = data_o[29];
  assign data_o[18973] = data_o[29];
  assign data_o[19037] = data_o[29];
  assign data_o[19101] = data_o[29];
  assign data_o[19165] = data_o[29];
  assign data_o[19229] = data_o[29];
  assign data_o[19293] = data_o[29];
  assign data_o[19357] = data_o[29];
  assign data_o[19421] = data_o[29];
  assign data_o[19485] = data_o[29];
  assign data_o[19549] = data_o[29];
  assign data_o[19613] = data_o[29];
  assign data_o[19677] = data_o[29];
  assign data_o[19741] = data_o[29];
  assign data_o[19805] = data_o[29];
  assign data_o[19869] = data_o[29];
  assign data_o[19933] = data_o[29];
  assign data_o[19997] = data_o[29];
  assign data_o[20061] = data_o[29];
  assign data_o[20125] = data_o[29];
  assign data_o[20189] = data_o[29];
  assign data_o[20253] = data_o[29];
  assign data_o[20317] = data_o[29];
  assign data_o[20381] = data_o[29];
  assign data_o[20445] = data_o[29];
  assign data_o[20509] = data_o[29];
  assign data_o[20573] = data_o[29];
  assign data_o[20637] = data_o[29];
  assign data_o[20701] = data_o[29];
  assign data_o[20765] = data_o[29];
  assign data_o[20829] = data_o[29];
  assign data_o[20893] = data_o[29];
  assign data_o[20957] = data_o[29];
  assign data_o[21021] = data_o[29];
  assign data_o[21085] = data_o[29];
  assign data_o[21149] = data_o[29];
  assign data_o[21213] = data_o[29];
  assign data_o[21277] = data_o[29];
  assign data_o[21341] = data_o[29];
  assign data_o[21405] = data_o[29];
  assign data_o[21469] = data_o[29];
  assign data_o[21533] = data_o[29];
  assign data_o[21597] = data_o[29];
  assign data_o[21661] = data_o[29];
  assign data_o[21725] = data_o[29];
  assign data_o[21789] = data_o[29];
  assign data_o[21853] = data_o[29];
  assign data_o[21917] = data_o[29];
  assign data_o[21981] = data_o[29];
  assign data_o[22045] = data_o[29];
  assign data_o[22109] = data_o[29];
  assign data_o[22173] = data_o[29];
  assign data_o[22237] = data_o[29];
  assign data_o[22301] = data_o[29];
  assign data_o[22365] = data_o[29];
  assign data_o[22429] = data_o[29];
  assign data_o[22493] = data_o[29];
  assign data_o[22557] = data_o[29];
  assign data_o[22621] = data_o[29];
  assign data_o[22685] = data_o[29];
  assign data_o[22749] = data_o[29];
  assign data_o[22813] = data_o[29];
  assign data_o[22877] = data_o[29];
  assign data_o[22941] = data_o[29];
  assign data_o[23005] = data_o[29];
  assign data_o[23069] = data_o[29];
  assign data_o[23133] = data_o[29];
  assign data_o[23197] = data_o[29];
  assign data_o[23261] = data_o[29];
  assign data_o[23325] = data_o[29];
  assign data_o[23389] = data_o[29];
  assign data_o[23453] = data_o[29];
  assign data_o[23517] = data_o[29];
  assign data_o[23581] = data_o[29];
  assign data_o[23645] = data_o[29];
  assign data_o[23709] = data_o[29];
  assign data_o[23773] = data_o[29];
  assign data_o[23837] = data_o[29];
  assign data_o[23901] = data_o[29];
  assign data_o[23965] = data_o[29];
  assign data_o[24029] = data_o[29];
  assign data_o[24093] = data_o[29];
  assign data_o[24157] = data_o[29];
  assign data_o[24221] = data_o[29];
  assign data_o[24285] = data_o[29];
  assign data_o[24349] = data_o[29];
  assign data_o[24413] = data_o[29];
  assign data_o[24477] = data_o[29];
  assign data_o[24541] = data_o[29];
  assign data_o[24605] = data_o[29];
  assign data_o[24669] = data_o[29];
  assign data_o[24733] = data_o[29];
  assign data_o[24797] = data_o[29];
  assign data_o[24861] = data_o[29];
  assign data_o[24925] = data_o[29];
  assign data_o[24989] = data_o[29];
  assign data_o[25053] = data_o[29];
  assign data_o[25117] = data_o[29];
  assign data_o[25181] = data_o[29];
  assign data_o[25245] = data_o[29];
  assign data_o[25309] = data_o[29];
  assign data_o[25373] = data_o[29];
  assign data_o[25437] = data_o[29];
  assign data_o[25501] = data_o[29];
  assign data_o[25565] = data_o[29];
  assign data_o[25629] = data_o[29];
  assign data_o[25693] = data_o[29];
  assign data_o[25757] = data_o[29];
  assign data_o[25821] = data_o[29];
  assign data_o[25885] = data_o[29];
  assign data_o[25949] = data_o[29];
  assign data_o[26013] = data_o[29];
  assign data_o[26077] = data_o[29];
  assign data_o[26141] = data_o[29];
  assign data_o[26205] = data_o[29];
  assign data_o[26269] = data_o[29];
  assign data_o[26333] = data_o[29];
  assign data_o[26397] = data_o[29];
  assign data_o[26461] = data_o[29];
  assign data_o[26525] = data_o[29];
  assign data_o[26589] = data_o[29];
  assign data_o[26653] = data_o[29];
  assign data_o[26717] = data_o[29];
  assign data_o[26781] = data_o[29];
  assign data_o[26845] = data_o[29];
  assign data_o[26909] = data_o[29];
  assign data_o[26973] = data_o[29];
  assign data_o[27037] = data_o[29];
  assign data_o[27101] = data_o[29];
  assign data_o[27165] = data_o[29];
  assign data_o[27229] = data_o[29];
  assign data_o[27293] = data_o[29];
  assign data_o[27357] = data_o[29];
  assign data_o[27421] = data_o[29];
  assign data_o[27485] = data_o[29];
  assign data_o[27549] = data_o[29];
  assign data_o[27613] = data_o[29];
  assign data_o[27677] = data_o[29];
  assign data_o[27741] = data_o[29];
  assign data_o[27805] = data_o[29];
  assign data_o[27869] = data_o[29];
  assign data_o[27933] = data_o[29];
  assign data_o[27997] = data_o[29];
  assign data_o[28061] = data_o[29];
  assign data_o[28125] = data_o[29];
  assign data_o[28189] = data_o[29];
  assign data_o[28253] = data_o[29];
  assign data_o[28317] = data_o[29];
  assign data_o[28381] = data_o[29];
  assign data_o[28445] = data_o[29];
  assign data_o[28509] = data_o[29];
  assign data_o[28573] = data_o[29];
  assign data_o[28637] = data_o[29];
  assign data_o[28701] = data_o[29];
  assign data_o[28765] = data_o[29];
  assign data_o[28829] = data_o[29];
  assign data_o[28893] = data_o[29];
  assign data_o[28957] = data_o[29];
  assign data_o[29021] = data_o[29];
  assign data_o[29085] = data_o[29];
  assign data_o[29149] = data_o[29];
  assign data_o[29213] = data_o[29];
  assign data_o[29277] = data_o[29];
  assign data_o[29341] = data_o[29];
  assign data_o[29405] = data_o[29];
  assign data_o[29469] = data_o[29];
  assign data_o[29533] = data_o[29];
  assign data_o[29597] = data_o[29];
  assign data_o[29661] = data_o[29];
  assign data_o[29725] = data_o[29];
  assign data_o[29789] = data_o[29];
  assign data_o[29853] = data_o[29];
  assign data_o[29917] = data_o[29];
  assign data_o[29981] = data_o[29];
  assign data_o[30045] = data_o[29];
  assign data_o[30109] = data_o[29];
  assign data_o[30173] = data_o[29];
  assign data_o[30237] = data_o[29];
  assign data_o[30301] = data_o[29];
  assign data_o[30365] = data_o[29];
  assign data_o[30429] = data_o[29];
  assign data_o[30493] = data_o[29];
  assign data_o[30557] = data_o[29];
  assign data_o[30621] = data_o[29];
  assign data_o[30685] = data_o[29];
  assign data_o[30749] = data_o[29];
  assign data_o[30813] = data_o[29];
  assign data_o[30877] = data_o[29];
  assign data_o[30941] = data_o[29];
  assign data_o[31005] = data_o[29];
  assign data_o[31069] = data_o[29];
  assign data_o[31133] = data_o[29];
  assign data_o[31197] = data_o[29];
  assign data_o[31261] = data_o[29];
  assign data_o[31325] = data_o[29];
  assign data_o[31389] = data_o[29];
  assign data_o[31453] = data_o[29];
  assign data_o[31517] = data_o[29];
  assign data_o[31581] = data_o[29];
  assign data_o[31645] = data_o[29];
  assign data_o[31709] = data_o[29];
  assign data_o[31773] = data_o[29];
  assign data_o[31837] = data_o[29];
  assign data_o[31901] = data_o[29];
  assign data_o[31965] = data_o[29];
  assign data_o[92] = data_o[28];
  assign data_o[156] = data_o[28];
  assign data_o[220] = data_o[28];
  assign data_o[284] = data_o[28];
  assign data_o[348] = data_o[28];
  assign data_o[412] = data_o[28];
  assign data_o[476] = data_o[28];
  assign data_o[540] = data_o[28];
  assign data_o[604] = data_o[28];
  assign data_o[668] = data_o[28];
  assign data_o[732] = data_o[28];
  assign data_o[796] = data_o[28];
  assign data_o[860] = data_o[28];
  assign data_o[924] = data_o[28];
  assign data_o[988] = data_o[28];
  assign data_o[1052] = data_o[28];
  assign data_o[1116] = data_o[28];
  assign data_o[1180] = data_o[28];
  assign data_o[1244] = data_o[28];
  assign data_o[1308] = data_o[28];
  assign data_o[1372] = data_o[28];
  assign data_o[1436] = data_o[28];
  assign data_o[1500] = data_o[28];
  assign data_o[1564] = data_o[28];
  assign data_o[1628] = data_o[28];
  assign data_o[1692] = data_o[28];
  assign data_o[1756] = data_o[28];
  assign data_o[1820] = data_o[28];
  assign data_o[1884] = data_o[28];
  assign data_o[1948] = data_o[28];
  assign data_o[2012] = data_o[28];
  assign data_o[2076] = data_o[28];
  assign data_o[2140] = data_o[28];
  assign data_o[2204] = data_o[28];
  assign data_o[2268] = data_o[28];
  assign data_o[2332] = data_o[28];
  assign data_o[2396] = data_o[28];
  assign data_o[2460] = data_o[28];
  assign data_o[2524] = data_o[28];
  assign data_o[2588] = data_o[28];
  assign data_o[2652] = data_o[28];
  assign data_o[2716] = data_o[28];
  assign data_o[2780] = data_o[28];
  assign data_o[2844] = data_o[28];
  assign data_o[2908] = data_o[28];
  assign data_o[2972] = data_o[28];
  assign data_o[3036] = data_o[28];
  assign data_o[3100] = data_o[28];
  assign data_o[3164] = data_o[28];
  assign data_o[3228] = data_o[28];
  assign data_o[3292] = data_o[28];
  assign data_o[3356] = data_o[28];
  assign data_o[3420] = data_o[28];
  assign data_o[3484] = data_o[28];
  assign data_o[3548] = data_o[28];
  assign data_o[3612] = data_o[28];
  assign data_o[3676] = data_o[28];
  assign data_o[3740] = data_o[28];
  assign data_o[3804] = data_o[28];
  assign data_o[3868] = data_o[28];
  assign data_o[3932] = data_o[28];
  assign data_o[3996] = data_o[28];
  assign data_o[4060] = data_o[28];
  assign data_o[4124] = data_o[28];
  assign data_o[4188] = data_o[28];
  assign data_o[4252] = data_o[28];
  assign data_o[4316] = data_o[28];
  assign data_o[4380] = data_o[28];
  assign data_o[4444] = data_o[28];
  assign data_o[4508] = data_o[28];
  assign data_o[4572] = data_o[28];
  assign data_o[4636] = data_o[28];
  assign data_o[4700] = data_o[28];
  assign data_o[4764] = data_o[28];
  assign data_o[4828] = data_o[28];
  assign data_o[4892] = data_o[28];
  assign data_o[4956] = data_o[28];
  assign data_o[5020] = data_o[28];
  assign data_o[5084] = data_o[28];
  assign data_o[5148] = data_o[28];
  assign data_o[5212] = data_o[28];
  assign data_o[5276] = data_o[28];
  assign data_o[5340] = data_o[28];
  assign data_o[5404] = data_o[28];
  assign data_o[5468] = data_o[28];
  assign data_o[5532] = data_o[28];
  assign data_o[5596] = data_o[28];
  assign data_o[5660] = data_o[28];
  assign data_o[5724] = data_o[28];
  assign data_o[5788] = data_o[28];
  assign data_o[5852] = data_o[28];
  assign data_o[5916] = data_o[28];
  assign data_o[5980] = data_o[28];
  assign data_o[6044] = data_o[28];
  assign data_o[6108] = data_o[28];
  assign data_o[6172] = data_o[28];
  assign data_o[6236] = data_o[28];
  assign data_o[6300] = data_o[28];
  assign data_o[6364] = data_o[28];
  assign data_o[6428] = data_o[28];
  assign data_o[6492] = data_o[28];
  assign data_o[6556] = data_o[28];
  assign data_o[6620] = data_o[28];
  assign data_o[6684] = data_o[28];
  assign data_o[6748] = data_o[28];
  assign data_o[6812] = data_o[28];
  assign data_o[6876] = data_o[28];
  assign data_o[6940] = data_o[28];
  assign data_o[7004] = data_o[28];
  assign data_o[7068] = data_o[28];
  assign data_o[7132] = data_o[28];
  assign data_o[7196] = data_o[28];
  assign data_o[7260] = data_o[28];
  assign data_o[7324] = data_o[28];
  assign data_o[7388] = data_o[28];
  assign data_o[7452] = data_o[28];
  assign data_o[7516] = data_o[28];
  assign data_o[7580] = data_o[28];
  assign data_o[7644] = data_o[28];
  assign data_o[7708] = data_o[28];
  assign data_o[7772] = data_o[28];
  assign data_o[7836] = data_o[28];
  assign data_o[7900] = data_o[28];
  assign data_o[7964] = data_o[28];
  assign data_o[8028] = data_o[28];
  assign data_o[8092] = data_o[28];
  assign data_o[8156] = data_o[28];
  assign data_o[8220] = data_o[28];
  assign data_o[8284] = data_o[28];
  assign data_o[8348] = data_o[28];
  assign data_o[8412] = data_o[28];
  assign data_o[8476] = data_o[28];
  assign data_o[8540] = data_o[28];
  assign data_o[8604] = data_o[28];
  assign data_o[8668] = data_o[28];
  assign data_o[8732] = data_o[28];
  assign data_o[8796] = data_o[28];
  assign data_o[8860] = data_o[28];
  assign data_o[8924] = data_o[28];
  assign data_o[8988] = data_o[28];
  assign data_o[9052] = data_o[28];
  assign data_o[9116] = data_o[28];
  assign data_o[9180] = data_o[28];
  assign data_o[9244] = data_o[28];
  assign data_o[9308] = data_o[28];
  assign data_o[9372] = data_o[28];
  assign data_o[9436] = data_o[28];
  assign data_o[9500] = data_o[28];
  assign data_o[9564] = data_o[28];
  assign data_o[9628] = data_o[28];
  assign data_o[9692] = data_o[28];
  assign data_o[9756] = data_o[28];
  assign data_o[9820] = data_o[28];
  assign data_o[9884] = data_o[28];
  assign data_o[9948] = data_o[28];
  assign data_o[10012] = data_o[28];
  assign data_o[10076] = data_o[28];
  assign data_o[10140] = data_o[28];
  assign data_o[10204] = data_o[28];
  assign data_o[10268] = data_o[28];
  assign data_o[10332] = data_o[28];
  assign data_o[10396] = data_o[28];
  assign data_o[10460] = data_o[28];
  assign data_o[10524] = data_o[28];
  assign data_o[10588] = data_o[28];
  assign data_o[10652] = data_o[28];
  assign data_o[10716] = data_o[28];
  assign data_o[10780] = data_o[28];
  assign data_o[10844] = data_o[28];
  assign data_o[10908] = data_o[28];
  assign data_o[10972] = data_o[28];
  assign data_o[11036] = data_o[28];
  assign data_o[11100] = data_o[28];
  assign data_o[11164] = data_o[28];
  assign data_o[11228] = data_o[28];
  assign data_o[11292] = data_o[28];
  assign data_o[11356] = data_o[28];
  assign data_o[11420] = data_o[28];
  assign data_o[11484] = data_o[28];
  assign data_o[11548] = data_o[28];
  assign data_o[11612] = data_o[28];
  assign data_o[11676] = data_o[28];
  assign data_o[11740] = data_o[28];
  assign data_o[11804] = data_o[28];
  assign data_o[11868] = data_o[28];
  assign data_o[11932] = data_o[28];
  assign data_o[11996] = data_o[28];
  assign data_o[12060] = data_o[28];
  assign data_o[12124] = data_o[28];
  assign data_o[12188] = data_o[28];
  assign data_o[12252] = data_o[28];
  assign data_o[12316] = data_o[28];
  assign data_o[12380] = data_o[28];
  assign data_o[12444] = data_o[28];
  assign data_o[12508] = data_o[28];
  assign data_o[12572] = data_o[28];
  assign data_o[12636] = data_o[28];
  assign data_o[12700] = data_o[28];
  assign data_o[12764] = data_o[28];
  assign data_o[12828] = data_o[28];
  assign data_o[12892] = data_o[28];
  assign data_o[12956] = data_o[28];
  assign data_o[13020] = data_o[28];
  assign data_o[13084] = data_o[28];
  assign data_o[13148] = data_o[28];
  assign data_o[13212] = data_o[28];
  assign data_o[13276] = data_o[28];
  assign data_o[13340] = data_o[28];
  assign data_o[13404] = data_o[28];
  assign data_o[13468] = data_o[28];
  assign data_o[13532] = data_o[28];
  assign data_o[13596] = data_o[28];
  assign data_o[13660] = data_o[28];
  assign data_o[13724] = data_o[28];
  assign data_o[13788] = data_o[28];
  assign data_o[13852] = data_o[28];
  assign data_o[13916] = data_o[28];
  assign data_o[13980] = data_o[28];
  assign data_o[14044] = data_o[28];
  assign data_o[14108] = data_o[28];
  assign data_o[14172] = data_o[28];
  assign data_o[14236] = data_o[28];
  assign data_o[14300] = data_o[28];
  assign data_o[14364] = data_o[28];
  assign data_o[14428] = data_o[28];
  assign data_o[14492] = data_o[28];
  assign data_o[14556] = data_o[28];
  assign data_o[14620] = data_o[28];
  assign data_o[14684] = data_o[28];
  assign data_o[14748] = data_o[28];
  assign data_o[14812] = data_o[28];
  assign data_o[14876] = data_o[28];
  assign data_o[14940] = data_o[28];
  assign data_o[15004] = data_o[28];
  assign data_o[15068] = data_o[28];
  assign data_o[15132] = data_o[28];
  assign data_o[15196] = data_o[28];
  assign data_o[15260] = data_o[28];
  assign data_o[15324] = data_o[28];
  assign data_o[15388] = data_o[28];
  assign data_o[15452] = data_o[28];
  assign data_o[15516] = data_o[28];
  assign data_o[15580] = data_o[28];
  assign data_o[15644] = data_o[28];
  assign data_o[15708] = data_o[28];
  assign data_o[15772] = data_o[28];
  assign data_o[15836] = data_o[28];
  assign data_o[15900] = data_o[28];
  assign data_o[15964] = data_o[28];
  assign data_o[16028] = data_o[28];
  assign data_o[16092] = data_o[28];
  assign data_o[16156] = data_o[28];
  assign data_o[16220] = data_o[28];
  assign data_o[16284] = data_o[28];
  assign data_o[16348] = data_o[28];
  assign data_o[16412] = data_o[28];
  assign data_o[16476] = data_o[28];
  assign data_o[16540] = data_o[28];
  assign data_o[16604] = data_o[28];
  assign data_o[16668] = data_o[28];
  assign data_o[16732] = data_o[28];
  assign data_o[16796] = data_o[28];
  assign data_o[16860] = data_o[28];
  assign data_o[16924] = data_o[28];
  assign data_o[16988] = data_o[28];
  assign data_o[17052] = data_o[28];
  assign data_o[17116] = data_o[28];
  assign data_o[17180] = data_o[28];
  assign data_o[17244] = data_o[28];
  assign data_o[17308] = data_o[28];
  assign data_o[17372] = data_o[28];
  assign data_o[17436] = data_o[28];
  assign data_o[17500] = data_o[28];
  assign data_o[17564] = data_o[28];
  assign data_o[17628] = data_o[28];
  assign data_o[17692] = data_o[28];
  assign data_o[17756] = data_o[28];
  assign data_o[17820] = data_o[28];
  assign data_o[17884] = data_o[28];
  assign data_o[17948] = data_o[28];
  assign data_o[18012] = data_o[28];
  assign data_o[18076] = data_o[28];
  assign data_o[18140] = data_o[28];
  assign data_o[18204] = data_o[28];
  assign data_o[18268] = data_o[28];
  assign data_o[18332] = data_o[28];
  assign data_o[18396] = data_o[28];
  assign data_o[18460] = data_o[28];
  assign data_o[18524] = data_o[28];
  assign data_o[18588] = data_o[28];
  assign data_o[18652] = data_o[28];
  assign data_o[18716] = data_o[28];
  assign data_o[18780] = data_o[28];
  assign data_o[18844] = data_o[28];
  assign data_o[18908] = data_o[28];
  assign data_o[18972] = data_o[28];
  assign data_o[19036] = data_o[28];
  assign data_o[19100] = data_o[28];
  assign data_o[19164] = data_o[28];
  assign data_o[19228] = data_o[28];
  assign data_o[19292] = data_o[28];
  assign data_o[19356] = data_o[28];
  assign data_o[19420] = data_o[28];
  assign data_o[19484] = data_o[28];
  assign data_o[19548] = data_o[28];
  assign data_o[19612] = data_o[28];
  assign data_o[19676] = data_o[28];
  assign data_o[19740] = data_o[28];
  assign data_o[19804] = data_o[28];
  assign data_o[19868] = data_o[28];
  assign data_o[19932] = data_o[28];
  assign data_o[19996] = data_o[28];
  assign data_o[20060] = data_o[28];
  assign data_o[20124] = data_o[28];
  assign data_o[20188] = data_o[28];
  assign data_o[20252] = data_o[28];
  assign data_o[20316] = data_o[28];
  assign data_o[20380] = data_o[28];
  assign data_o[20444] = data_o[28];
  assign data_o[20508] = data_o[28];
  assign data_o[20572] = data_o[28];
  assign data_o[20636] = data_o[28];
  assign data_o[20700] = data_o[28];
  assign data_o[20764] = data_o[28];
  assign data_o[20828] = data_o[28];
  assign data_o[20892] = data_o[28];
  assign data_o[20956] = data_o[28];
  assign data_o[21020] = data_o[28];
  assign data_o[21084] = data_o[28];
  assign data_o[21148] = data_o[28];
  assign data_o[21212] = data_o[28];
  assign data_o[21276] = data_o[28];
  assign data_o[21340] = data_o[28];
  assign data_o[21404] = data_o[28];
  assign data_o[21468] = data_o[28];
  assign data_o[21532] = data_o[28];
  assign data_o[21596] = data_o[28];
  assign data_o[21660] = data_o[28];
  assign data_o[21724] = data_o[28];
  assign data_o[21788] = data_o[28];
  assign data_o[21852] = data_o[28];
  assign data_o[21916] = data_o[28];
  assign data_o[21980] = data_o[28];
  assign data_o[22044] = data_o[28];
  assign data_o[22108] = data_o[28];
  assign data_o[22172] = data_o[28];
  assign data_o[22236] = data_o[28];
  assign data_o[22300] = data_o[28];
  assign data_o[22364] = data_o[28];
  assign data_o[22428] = data_o[28];
  assign data_o[22492] = data_o[28];
  assign data_o[22556] = data_o[28];
  assign data_o[22620] = data_o[28];
  assign data_o[22684] = data_o[28];
  assign data_o[22748] = data_o[28];
  assign data_o[22812] = data_o[28];
  assign data_o[22876] = data_o[28];
  assign data_o[22940] = data_o[28];
  assign data_o[23004] = data_o[28];
  assign data_o[23068] = data_o[28];
  assign data_o[23132] = data_o[28];
  assign data_o[23196] = data_o[28];
  assign data_o[23260] = data_o[28];
  assign data_o[23324] = data_o[28];
  assign data_o[23388] = data_o[28];
  assign data_o[23452] = data_o[28];
  assign data_o[23516] = data_o[28];
  assign data_o[23580] = data_o[28];
  assign data_o[23644] = data_o[28];
  assign data_o[23708] = data_o[28];
  assign data_o[23772] = data_o[28];
  assign data_o[23836] = data_o[28];
  assign data_o[23900] = data_o[28];
  assign data_o[23964] = data_o[28];
  assign data_o[24028] = data_o[28];
  assign data_o[24092] = data_o[28];
  assign data_o[24156] = data_o[28];
  assign data_o[24220] = data_o[28];
  assign data_o[24284] = data_o[28];
  assign data_o[24348] = data_o[28];
  assign data_o[24412] = data_o[28];
  assign data_o[24476] = data_o[28];
  assign data_o[24540] = data_o[28];
  assign data_o[24604] = data_o[28];
  assign data_o[24668] = data_o[28];
  assign data_o[24732] = data_o[28];
  assign data_o[24796] = data_o[28];
  assign data_o[24860] = data_o[28];
  assign data_o[24924] = data_o[28];
  assign data_o[24988] = data_o[28];
  assign data_o[25052] = data_o[28];
  assign data_o[25116] = data_o[28];
  assign data_o[25180] = data_o[28];
  assign data_o[25244] = data_o[28];
  assign data_o[25308] = data_o[28];
  assign data_o[25372] = data_o[28];
  assign data_o[25436] = data_o[28];
  assign data_o[25500] = data_o[28];
  assign data_o[25564] = data_o[28];
  assign data_o[25628] = data_o[28];
  assign data_o[25692] = data_o[28];
  assign data_o[25756] = data_o[28];
  assign data_o[25820] = data_o[28];
  assign data_o[25884] = data_o[28];
  assign data_o[25948] = data_o[28];
  assign data_o[26012] = data_o[28];
  assign data_o[26076] = data_o[28];
  assign data_o[26140] = data_o[28];
  assign data_o[26204] = data_o[28];
  assign data_o[26268] = data_o[28];
  assign data_o[26332] = data_o[28];
  assign data_o[26396] = data_o[28];
  assign data_o[26460] = data_o[28];
  assign data_o[26524] = data_o[28];
  assign data_o[26588] = data_o[28];
  assign data_o[26652] = data_o[28];
  assign data_o[26716] = data_o[28];
  assign data_o[26780] = data_o[28];
  assign data_o[26844] = data_o[28];
  assign data_o[26908] = data_o[28];
  assign data_o[26972] = data_o[28];
  assign data_o[27036] = data_o[28];
  assign data_o[27100] = data_o[28];
  assign data_o[27164] = data_o[28];
  assign data_o[27228] = data_o[28];
  assign data_o[27292] = data_o[28];
  assign data_o[27356] = data_o[28];
  assign data_o[27420] = data_o[28];
  assign data_o[27484] = data_o[28];
  assign data_o[27548] = data_o[28];
  assign data_o[27612] = data_o[28];
  assign data_o[27676] = data_o[28];
  assign data_o[27740] = data_o[28];
  assign data_o[27804] = data_o[28];
  assign data_o[27868] = data_o[28];
  assign data_o[27932] = data_o[28];
  assign data_o[27996] = data_o[28];
  assign data_o[28060] = data_o[28];
  assign data_o[28124] = data_o[28];
  assign data_o[28188] = data_o[28];
  assign data_o[28252] = data_o[28];
  assign data_o[28316] = data_o[28];
  assign data_o[28380] = data_o[28];
  assign data_o[28444] = data_o[28];
  assign data_o[28508] = data_o[28];
  assign data_o[28572] = data_o[28];
  assign data_o[28636] = data_o[28];
  assign data_o[28700] = data_o[28];
  assign data_o[28764] = data_o[28];
  assign data_o[28828] = data_o[28];
  assign data_o[28892] = data_o[28];
  assign data_o[28956] = data_o[28];
  assign data_o[29020] = data_o[28];
  assign data_o[29084] = data_o[28];
  assign data_o[29148] = data_o[28];
  assign data_o[29212] = data_o[28];
  assign data_o[29276] = data_o[28];
  assign data_o[29340] = data_o[28];
  assign data_o[29404] = data_o[28];
  assign data_o[29468] = data_o[28];
  assign data_o[29532] = data_o[28];
  assign data_o[29596] = data_o[28];
  assign data_o[29660] = data_o[28];
  assign data_o[29724] = data_o[28];
  assign data_o[29788] = data_o[28];
  assign data_o[29852] = data_o[28];
  assign data_o[29916] = data_o[28];
  assign data_o[29980] = data_o[28];
  assign data_o[30044] = data_o[28];
  assign data_o[30108] = data_o[28];
  assign data_o[30172] = data_o[28];
  assign data_o[30236] = data_o[28];
  assign data_o[30300] = data_o[28];
  assign data_o[30364] = data_o[28];
  assign data_o[30428] = data_o[28];
  assign data_o[30492] = data_o[28];
  assign data_o[30556] = data_o[28];
  assign data_o[30620] = data_o[28];
  assign data_o[30684] = data_o[28];
  assign data_o[30748] = data_o[28];
  assign data_o[30812] = data_o[28];
  assign data_o[30876] = data_o[28];
  assign data_o[30940] = data_o[28];
  assign data_o[31004] = data_o[28];
  assign data_o[31068] = data_o[28];
  assign data_o[31132] = data_o[28];
  assign data_o[31196] = data_o[28];
  assign data_o[31260] = data_o[28];
  assign data_o[31324] = data_o[28];
  assign data_o[31388] = data_o[28];
  assign data_o[31452] = data_o[28];
  assign data_o[31516] = data_o[28];
  assign data_o[31580] = data_o[28];
  assign data_o[31644] = data_o[28];
  assign data_o[31708] = data_o[28];
  assign data_o[31772] = data_o[28];
  assign data_o[31836] = data_o[28];
  assign data_o[31900] = data_o[28];
  assign data_o[31964] = data_o[28];
  assign data_o[91] = data_o[27];
  assign data_o[155] = data_o[27];
  assign data_o[219] = data_o[27];
  assign data_o[283] = data_o[27];
  assign data_o[347] = data_o[27];
  assign data_o[411] = data_o[27];
  assign data_o[475] = data_o[27];
  assign data_o[539] = data_o[27];
  assign data_o[603] = data_o[27];
  assign data_o[667] = data_o[27];
  assign data_o[731] = data_o[27];
  assign data_o[795] = data_o[27];
  assign data_o[859] = data_o[27];
  assign data_o[923] = data_o[27];
  assign data_o[987] = data_o[27];
  assign data_o[1051] = data_o[27];
  assign data_o[1115] = data_o[27];
  assign data_o[1179] = data_o[27];
  assign data_o[1243] = data_o[27];
  assign data_o[1307] = data_o[27];
  assign data_o[1371] = data_o[27];
  assign data_o[1435] = data_o[27];
  assign data_o[1499] = data_o[27];
  assign data_o[1563] = data_o[27];
  assign data_o[1627] = data_o[27];
  assign data_o[1691] = data_o[27];
  assign data_o[1755] = data_o[27];
  assign data_o[1819] = data_o[27];
  assign data_o[1883] = data_o[27];
  assign data_o[1947] = data_o[27];
  assign data_o[2011] = data_o[27];
  assign data_o[2075] = data_o[27];
  assign data_o[2139] = data_o[27];
  assign data_o[2203] = data_o[27];
  assign data_o[2267] = data_o[27];
  assign data_o[2331] = data_o[27];
  assign data_o[2395] = data_o[27];
  assign data_o[2459] = data_o[27];
  assign data_o[2523] = data_o[27];
  assign data_o[2587] = data_o[27];
  assign data_o[2651] = data_o[27];
  assign data_o[2715] = data_o[27];
  assign data_o[2779] = data_o[27];
  assign data_o[2843] = data_o[27];
  assign data_o[2907] = data_o[27];
  assign data_o[2971] = data_o[27];
  assign data_o[3035] = data_o[27];
  assign data_o[3099] = data_o[27];
  assign data_o[3163] = data_o[27];
  assign data_o[3227] = data_o[27];
  assign data_o[3291] = data_o[27];
  assign data_o[3355] = data_o[27];
  assign data_o[3419] = data_o[27];
  assign data_o[3483] = data_o[27];
  assign data_o[3547] = data_o[27];
  assign data_o[3611] = data_o[27];
  assign data_o[3675] = data_o[27];
  assign data_o[3739] = data_o[27];
  assign data_o[3803] = data_o[27];
  assign data_o[3867] = data_o[27];
  assign data_o[3931] = data_o[27];
  assign data_o[3995] = data_o[27];
  assign data_o[4059] = data_o[27];
  assign data_o[4123] = data_o[27];
  assign data_o[4187] = data_o[27];
  assign data_o[4251] = data_o[27];
  assign data_o[4315] = data_o[27];
  assign data_o[4379] = data_o[27];
  assign data_o[4443] = data_o[27];
  assign data_o[4507] = data_o[27];
  assign data_o[4571] = data_o[27];
  assign data_o[4635] = data_o[27];
  assign data_o[4699] = data_o[27];
  assign data_o[4763] = data_o[27];
  assign data_o[4827] = data_o[27];
  assign data_o[4891] = data_o[27];
  assign data_o[4955] = data_o[27];
  assign data_o[5019] = data_o[27];
  assign data_o[5083] = data_o[27];
  assign data_o[5147] = data_o[27];
  assign data_o[5211] = data_o[27];
  assign data_o[5275] = data_o[27];
  assign data_o[5339] = data_o[27];
  assign data_o[5403] = data_o[27];
  assign data_o[5467] = data_o[27];
  assign data_o[5531] = data_o[27];
  assign data_o[5595] = data_o[27];
  assign data_o[5659] = data_o[27];
  assign data_o[5723] = data_o[27];
  assign data_o[5787] = data_o[27];
  assign data_o[5851] = data_o[27];
  assign data_o[5915] = data_o[27];
  assign data_o[5979] = data_o[27];
  assign data_o[6043] = data_o[27];
  assign data_o[6107] = data_o[27];
  assign data_o[6171] = data_o[27];
  assign data_o[6235] = data_o[27];
  assign data_o[6299] = data_o[27];
  assign data_o[6363] = data_o[27];
  assign data_o[6427] = data_o[27];
  assign data_o[6491] = data_o[27];
  assign data_o[6555] = data_o[27];
  assign data_o[6619] = data_o[27];
  assign data_o[6683] = data_o[27];
  assign data_o[6747] = data_o[27];
  assign data_o[6811] = data_o[27];
  assign data_o[6875] = data_o[27];
  assign data_o[6939] = data_o[27];
  assign data_o[7003] = data_o[27];
  assign data_o[7067] = data_o[27];
  assign data_o[7131] = data_o[27];
  assign data_o[7195] = data_o[27];
  assign data_o[7259] = data_o[27];
  assign data_o[7323] = data_o[27];
  assign data_o[7387] = data_o[27];
  assign data_o[7451] = data_o[27];
  assign data_o[7515] = data_o[27];
  assign data_o[7579] = data_o[27];
  assign data_o[7643] = data_o[27];
  assign data_o[7707] = data_o[27];
  assign data_o[7771] = data_o[27];
  assign data_o[7835] = data_o[27];
  assign data_o[7899] = data_o[27];
  assign data_o[7963] = data_o[27];
  assign data_o[8027] = data_o[27];
  assign data_o[8091] = data_o[27];
  assign data_o[8155] = data_o[27];
  assign data_o[8219] = data_o[27];
  assign data_o[8283] = data_o[27];
  assign data_o[8347] = data_o[27];
  assign data_o[8411] = data_o[27];
  assign data_o[8475] = data_o[27];
  assign data_o[8539] = data_o[27];
  assign data_o[8603] = data_o[27];
  assign data_o[8667] = data_o[27];
  assign data_o[8731] = data_o[27];
  assign data_o[8795] = data_o[27];
  assign data_o[8859] = data_o[27];
  assign data_o[8923] = data_o[27];
  assign data_o[8987] = data_o[27];
  assign data_o[9051] = data_o[27];
  assign data_o[9115] = data_o[27];
  assign data_o[9179] = data_o[27];
  assign data_o[9243] = data_o[27];
  assign data_o[9307] = data_o[27];
  assign data_o[9371] = data_o[27];
  assign data_o[9435] = data_o[27];
  assign data_o[9499] = data_o[27];
  assign data_o[9563] = data_o[27];
  assign data_o[9627] = data_o[27];
  assign data_o[9691] = data_o[27];
  assign data_o[9755] = data_o[27];
  assign data_o[9819] = data_o[27];
  assign data_o[9883] = data_o[27];
  assign data_o[9947] = data_o[27];
  assign data_o[10011] = data_o[27];
  assign data_o[10075] = data_o[27];
  assign data_o[10139] = data_o[27];
  assign data_o[10203] = data_o[27];
  assign data_o[10267] = data_o[27];
  assign data_o[10331] = data_o[27];
  assign data_o[10395] = data_o[27];
  assign data_o[10459] = data_o[27];
  assign data_o[10523] = data_o[27];
  assign data_o[10587] = data_o[27];
  assign data_o[10651] = data_o[27];
  assign data_o[10715] = data_o[27];
  assign data_o[10779] = data_o[27];
  assign data_o[10843] = data_o[27];
  assign data_o[10907] = data_o[27];
  assign data_o[10971] = data_o[27];
  assign data_o[11035] = data_o[27];
  assign data_o[11099] = data_o[27];
  assign data_o[11163] = data_o[27];
  assign data_o[11227] = data_o[27];
  assign data_o[11291] = data_o[27];
  assign data_o[11355] = data_o[27];
  assign data_o[11419] = data_o[27];
  assign data_o[11483] = data_o[27];
  assign data_o[11547] = data_o[27];
  assign data_o[11611] = data_o[27];
  assign data_o[11675] = data_o[27];
  assign data_o[11739] = data_o[27];
  assign data_o[11803] = data_o[27];
  assign data_o[11867] = data_o[27];
  assign data_o[11931] = data_o[27];
  assign data_o[11995] = data_o[27];
  assign data_o[12059] = data_o[27];
  assign data_o[12123] = data_o[27];
  assign data_o[12187] = data_o[27];
  assign data_o[12251] = data_o[27];
  assign data_o[12315] = data_o[27];
  assign data_o[12379] = data_o[27];
  assign data_o[12443] = data_o[27];
  assign data_o[12507] = data_o[27];
  assign data_o[12571] = data_o[27];
  assign data_o[12635] = data_o[27];
  assign data_o[12699] = data_o[27];
  assign data_o[12763] = data_o[27];
  assign data_o[12827] = data_o[27];
  assign data_o[12891] = data_o[27];
  assign data_o[12955] = data_o[27];
  assign data_o[13019] = data_o[27];
  assign data_o[13083] = data_o[27];
  assign data_o[13147] = data_o[27];
  assign data_o[13211] = data_o[27];
  assign data_o[13275] = data_o[27];
  assign data_o[13339] = data_o[27];
  assign data_o[13403] = data_o[27];
  assign data_o[13467] = data_o[27];
  assign data_o[13531] = data_o[27];
  assign data_o[13595] = data_o[27];
  assign data_o[13659] = data_o[27];
  assign data_o[13723] = data_o[27];
  assign data_o[13787] = data_o[27];
  assign data_o[13851] = data_o[27];
  assign data_o[13915] = data_o[27];
  assign data_o[13979] = data_o[27];
  assign data_o[14043] = data_o[27];
  assign data_o[14107] = data_o[27];
  assign data_o[14171] = data_o[27];
  assign data_o[14235] = data_o[27];
  assign data_o[14299] = data_o[27];
  assign data_o[14363] = data_o[27];
  assign data_o[14427] = data_o[27];
  assign data_o[14491] = data_o[27];
  assign data_o[14555] = data_o[27];
  assign data_o[14619] = data_o[27];
  assign data_o[14683] = data_o[27];
  assign data_o[14747] = data_o[27];
  assign data_o[14811] = data_o[27];
  assign data_o[14875] = data_o[27];
  assign data_o[14939] = data_o[27];
  assign data_o[15003] = data_o[27];
  assign data_o[15067] = data_o[27];
  assign data_o[15131] = data_o[27];
  assign data_o[15195] = data_o[27];
  assign data_o[15259] = data_o[27];
  assign data_o[15323] = data_o[27];
  assign data_o[15387] = data_o[27];
  assign data_o[15451] = data_o[27];
  assign data_o[15515] = data_o[27];
  assign data_o[15579] = data_o[27];
  assign data_o[15643] = data_o[27];
  assign data_o[15707] = data_o[27];
  assign data_o[15771] = data_o[27];
  assign data_o[15835] = data_o[27];
  assign data_o[15899] = data_o[27];
  assign data_o[15963] = data_o[27];
  assign data_o[16027] = data_o[27];
  assign data_o[16091] = data_o[27];
  assign data_o[16155] = data_o[27];
  assign data_o[16219] = data_o[27];
  assign data_o[16283] = data_o[27];
  assign data_o[16347] = data_o[27];
  assign data_o[16411] = data_o[27];
  assign data_o[16475] = data_o[27];
  assign data_o[16539] = data_o[27];
  assign data_o[16603] = data_o[27];
  assign data_o[16667] = data_o[27];
  assign data_o[16731] = data_o[27];
  assign data_o[16795] = data_o[27];
  assign data_o[16859] = data_o[27];
  assign data_o[16923] = data_o[27];
  assign data_o[16987] = data_o[27];
  assign data_o[17051] = data_o[27];
  assign data_o[17115] = data_o[27];
  assign data_o[17179] = data_o[27];
  assign data_o[17243] = data_o[27];
  assign data_o[17307] = data_o[27];
  assign data_o[17371] = data_o[27];
  assign data_o[17435] = data_o[27];
  assign data_o[17499] = data_o[27];
  assign data_o[17563] = data_o[27];
  assign data_o[17627] = data_o[27];
  assign data_o[17691] = data_o[27];
  assign data_o[17755] = data_o[27];
  assign data_o[17819] = data_o[27];
  assign data_o[17883] = data_o[27];
  assign data_o[17947] = data_o[27];
  assign data_o[18011] = data_o[27];
  assign data_o[18075] = data_o[27];
  assign data_o[18139] = data_o[27];
  assign data_o[18203] = data_o[27];
  assign data_o[18267] = data_o[27];
  assign data_o[18331] = data_o[27];
  assign data_o[18395] = data_o[27];
  assign data_o[18459] = data_o[27];
  assign data_o[18523] = data_o[27];
  assign data_o[18587] = data_o[27];
  assign data_o[18651] = data_o[27];
  assign data_o[18715] = data_o[27];
  assign data_o[18779] = data_o[27];
  assign data_o[18843] = data_o[27];
  assign data_o[18907] = data_o[27];
  assign data_o[18971] = data_o[27];
  assign data_o[19035] = data_o[27];
  assign data_o[19099] = data_o[27];
  assign data_o[19163] = data_o[27];
  assign data_o[19227] = data_o[27];
  assign data_o[19291] = data_o[27];
  assign data_o[19355] = data_o[27];
  assign data_o[19419] = data_o[27];
  assign data_o[19483] = data_o[27];
  assign data_o[19547] = data_o[27];
  assign data_o[19611] = data_o[27];
  assign data_o[19675] = data_o[27];
  assign data_o[19739] = data_o[27];
  assign data_o[19803] = data_o[27];
  assign data_o[19867] = data_o[27];
  assign data_o[19931] = data_o[27];
  assign data_o[19995] = data_o[27];
  assign data_o[20059] = data_o[27];
  assign data_o[20123] = data_o[27];
  assign data_o[20187] = data_o[27];
  assign data_o[20251] = data_o[27];
  assign data_o[20315] = data_o[27];
  assign data_o[20379] = data_o[27];
  assign data_o[20443] = data_o[27];
  assign data_o[20507] = data_o[27];
  assign data_o[20571] = data_o[27];
  assign data_o[20635] = data_o[27];
  assign data_o[20699] = data_o[27];
  assign data_o[20763] = data_o[27];
  assign data_o[20827] = data_o[27];
  assign data_o[20891] = data_o[27];
  assign data_o[20955] = data_o[27];
  assign data_o[21019] = data_o[27];
  assign data_o[21083] = data_o[27];
  assign data_o[21147] = data_o[27];
  assign data_o[21211] = data_o[27];
  assign data_o[21275] = data_o[27];
  assign data_o[21339] = data_o[27];
  assign data_o[21403] = data_o[27];
  assign data_o[21467] = data_o[27];
  assign data_o[21531] = data_o[27];
  assign data_o[21595] = data_o[27];
  assign data_o[21659] = data_o[27];
  assign data_o[21723] = data_o[27];
  assign data_o[21787] = data_o[27];
  assign data_o[21851] = data_o[27];
  assign data_o[21915] = data_o[27];
  assign data_o[21979] = data_o[27];
  assign data_o[22043] = data_o[27];
  assign data_o[22107] = data_o[27];
  assign data_o[22171] = data_o[27];
  assign data_o[22235] = data_o[27];
  assign data_o[22299] = data_o[27];
  assign data_o[22363] = data_o[27];
  assign data_o[22427] = data_o[27];
  assign data_o[22491] = data_o[27];
  assign data_o[22555] = data_o[27];
  assign data_o[22619] = data_o[27];
  assign data_o[22683] = data_o[27];
  assign data_o[22747] = data_o[27];
  assign data_o[22811] = data_o[27];
  assign data_o[22875] = data_o[27];
  assign data_o[22939] = data_o[27];
  assign data_o[23003] = data_o[27];
  assign data_o[23067] = data_o[27];
  assign data_o[23131] = data_o[27];
  assign data_o[23195] = data_o[27];
  assign data_o[23259] = data_o[27];
  assign data_o[23323] = data_o[27];
  assign data_o[23387] = data_o[27];
  assign data_o[23451] = data_o[27];
  assign data_o[23515] = data_o[27];
  assign data_o[23579] = data_o[27];
  assign data_o[23643] = data_o[27];
  assign data_o[23707] = data_o[27];
  assign data_o[23771] = data_o[27];
  assign data_o[23835] = data_o[27];
  assign data_o[23899] = data_o[27];
  assign data_o[23963] = data_o[27];
  assign data_o[24027] = data_o[27];
  assign data_o[24091] = data_o[27];
  assign data_o[24155] = data_o[27];
  assign data_o[24219] = data_o[27];
  assign data_o[24283] = data_o[27];
  assign data_o[24347] = data_o[27];
  assign data_o[24411] = data_o[27];
  assign data_o[24475] = data_o[27];
  assign data_o[24539] = data_o[27];
  assign data_o[24603] = data_o[27];
  assign data_o[24667] = data_o[27];
  assign data_o[24731] = data_o[27];
  assign data_o[24795] = data_o[27];
  assign data_o[24859] = data_o[27];
  assign data_o[24923] = data_o[27];
  assign data_o[24987] = data_o[27];
  assign data_o[25051] = data_o[27];
  assign data_o[25115] = data_o[27];
  assign data_o[25179] = data_o[27];
  assign data_o[25243] = data_o[27];
  assign data_o[25307] = data_o[27];
  assign data_o[25371] = data_o[27];
  assign data_o[25435] = data_o[27];
  assign data_o[25499] = data_o[27];
  assign data_o[25563] = data_o[27];
  assign data_o[25627] = data_o[27];
  assign data_o[25691] = data_o[27];
  assign data_o[25755] = data_o[27];
  assign data_o[25819] = data_o[27];
  assign data_o[25883] = data_o[27];
  assign data_o[25947] = data_o[27];
  assign data_o[26011] = data_o[27];
  assign data_o[26075] = data_o[27];
  assign data_o[26139] = data_o[27];
  assign data_o[26203] = data_o[27];
  assign data_o[26267] = data_o[27];
  assign data_o[26331] = data_o[27];
  assign data_o[26395] = data_o[27];
  assign data_o[26459] = data_o[27];
  assign data_o[26523] = data_o[27];
  assign data_o[26587] = data_o[27];
  assign data_o[26651] = data_o[27];
  assign data_o[26715] = data_o[27];
  assign data_o[26779] = data_o[27];
  assign data_o[26843] = data_o[27];
  assign data_o[26907] = data_o[27];
  assign data_o[26971] = data_o[27];
  assign data_o[27035] = data_o[27];
  assign data_o[27099] = data_o[27];
  assign data_o[27163] = data_o[27];
  assign data_o[27227] = data_o[27];
  assign data_o[27291] = data_o[27];
  assign data_o[27355] = data_o[27];
  assign data_o[27419] = data_o[27];
  assign data_o[27483] = data_o[27];
  assign data_o[27547] = data_o[27];
  assign data_o[27611] = data_o[27];
  assign data_o[27675] = data_o[27];
  assign data_o[27739] = data_o[27];
  assign data_o[27803] = data_o[27];
  assign data_o[27867] = data_o[27];
  assign data_o[27931] = data_o[27];
  assign data_o[27995] = data_o[27];
  assign data_o[28059] = data_o[27];
  assign data_o[28123] = data_o[27];
  assign data_o[28187] = data_o[27];
  assign data_o[28251] = data_o[27];
  assign data_o[28315] = data_o[27];
  assign data_o[28379] = data_o[27];
  assign data_o[28443] = data_o[27];
  assign data_o[28507] = data_o[27];
  assign data_o[28571] = data_o[27];
  assign data_o[28635] = data_o[27];
  assign data_o[28699] = data_o[27];
  assign data_o[28763] = data_o[27];
  assign data_o[28827] = data_o[27];
  assign data_o[28891] = data_o[27];
  assign data_o[28955] = data_o[27];
  assign data_o[29019] = data_o[27];
  assign data_o[29083] = data_o[27];
  assign data_o[29147] = data_o[27];
  assign data_o[29211] = data_o[27];
  assign data_o[29275] = data_o[27];
  assign data_o[29339] = data_o[27];
  assign data_o[29403] = data_o[27];
  assign data_o[29467] = data_o[27];
  assign data_o[29531] = data_o[27];
  assign data_o[29595] = data_o[27];
  assign data_o[29659] = data_o[27];
  assign data_o[29723] = data_o[27];
  assign data_o[29787] = data_o[27];
  assign data_o[29851] = data_o[27];
  assign data_o[29915] = data_o[27];
  assign data_o[29979] = data_o[27];
  assign data_o[30043] = data_o[27];
  assign data_o[30107] = data_o[27];
  assign data_o[30171] = data_o[27];
  assign data_o[30235] = data_o[27];
  assign data_o[30299] = data_o[27];
  assign data_o[30363] = data_o[27];
  assign data_o[30427] = data_o[27];
  assign data_o[30491] = data_o[27];
  assign data_o[30555] = data_o[27];
  assign data_o[30619] = data_o[27];
  assign data_o[30683] = data_o[27];
  assign data_o[30747] = data_o[27];
  assign data_o[30811] = data_o[27];
  assign data_o[30875] = data_o[27];
  assign data_o[30939] = data_o[27];
  assign data_o[31003] = data_o[27];
  assign data_o[31067] = data_o[27];
  assign data_o[31131] = data_o[27];
  assign data_o[31195] = data_o[27];
  assign data_o[31259] = data_o[27];
  assign data_o[31323] = data_o[27];
  assign data_o[31387] = data_o[27];
  assign data_o[31451] = data_o[27];
  assign data_o[31515] = data_o[27];
  assign data_o[31579] = data_o[27];
  assign data_o[31643] = data_o[27];
  assign data_o[31707] = data_o[27];
  assign data_o[31771] = data_o[27];
  assign data_o[31835] = data_o[27];
  assign data_o[31899] = data_o[27];
  assign data_o[31963] = data_o[27];
  assign data_o[90] = data_o[26];
  assign data_o[154] = data_o[26];
  assign data_o[218] = data_o[26];
  assign data_o[282] = data_o[26];
  assign data_o[346] = data_o[26];
  assign data_o[410] = data_o[26];
  assign data_o[474] = data_o[26];
  assign data_o[538] = data_o[26];
  assign data_o[602] = data_o[26];
  assign data_o[666] = data_o[26];
  assign data_o[730] = data_o[26];
  assign data_o[794] = data_o[26];
  assign data_o[858] = data_o[26];
  assign data_o[922] = data_o[26];
  assign data_o[986] = data_o[26];
  assign data_o[1050] = data_o[26];
  assign data_o[1114] = data_o[26];
  assign data_o[1178] = data_o[26];
  assign data_o[1242] = data_o[26];
  assign data_o[1306] = data_o[26];
  assign data_o[1370] = data_o[26];
  assign data_o[1434] = data_o[26];
  assign data_o[1498] = data_o[26];
  assign data_o[1562] = data_o[26];
  assign data_o[1626] = data_o[26];
  assign data_o[1690] = data_o[26];
  assign data_o[1754] = data_o[26];
  assign data_o[1818] = data_o[26];
  assign data_o[1882] = data_o[26];
  assign data_o[1946] = data_o[26];
  assign data_o[2010] = data_o[26];
  assign data_o[2074] = data_o[26];
  assign data_o[2138] = data_o[26];
  assign data_o[2202] = data_o[26];
  assign data_o[2266] = data_o[26];
  assign data_o[2330] = data_o[26];
  assign data_o[2394] = data_o[26];
  assign data_o[2458] = data_o[26];
  assign data_o[2522] = data_o[26];
  assign data_o[2586] = data_o[26];
  assign data_o[2650] = data_o[26];
  assign data_o[2714] = data_o[26];
  assign data_o[2778] = data_o[26];
  assign data_o[2842] = data_o[26];
  assign data_o[2906] = data_o[26];
  assign data_o[2970] = data_o[26];
  assign data_o[3034] = data_o[26];
  assign data_o[3098] = data_o[26];
  assign data_o[3162] = data_o[26];
  assign data_o[3226] = data_o[26];
  assign data_o[3290] = data_o[26];
  assign data_o[3354] = data_o[26];
  assign data_o[3418] = data_o[26];
  assign data_o[3482] = data_o[26];
  assign data_o[3546] = data_o[26];
  assign data_o[3610] = data_o[26];
  assign data_o[3674] = data_o[26];
  assign data_o[3738] = data_o[26];
  assign data_o[3802] = data_o[26];
  assign data_o[3866] = data_o[26];
  assign data_o[3930] = data_o[26];
  assign data_o[3994] = data_o[26];
  assign data_o[4058] = data_o[26];
  assign data_o[4122] = data_o[26];
  assign data_o[4186] = data_o[26];
  assign data_o[4250] = data_o[26];
  assign data_o[4314] = data_o[26];
  assign data_o[4378] = data_o[26];
  assign data_o[4442] = data_o[26];
  assign data_o[4506] = data_o[26];
  assign data_o[4570] = data_o[26];
  assign data_o[4634] = data_o[26];
  assign data_o[4698] = data_o[26];
  assign data_o[4762] = data_o[26];
  assign data_o[4826] = data_o[26];
  assign data_o[4890] = data_o[26];
  assign data_o[4954] = data_o[26];
  assign data_o[5018] = data_o[26];
  assign data_o[5082] = data_o[26];
  assign data_o[5146] = data_o[26];
  assign data_o[5210] = data_o[26];
  assign data_o[5274] = data_o[26];
  assign data_o[5338] = data_o[26];
  assign data_o[5402] = data_o[26];
  assign data_o[5466] = data_o[26];
  assign data_o[5530] = data_o[26];
  assign data_o[5594] = data_o[26];
  assign data_o[5658] = data_o[26];
  assign data_o[5722] = data_o[26];
  assign data_o[5786] = data_o[26];
  assign data_o[5850] = data_o[26];
  assign data_o[5914] = data_o[26];
  assign data_o[5978] = data_o[26];
  assign data_o[6042] = data_o[26];
  assign data_o[6106] = data_o[26];
  assign data_o[6170] = data_o[26];
  assign data_o[6234] = data_o[26];
  assign data_o[6298] = data_o[26];
  assign data_o[6362] = data_o[26];
  assign data_o[6426] = data_o[26];
  assign data_o[6490] = data_o[26];
  assign data_o[6554] = data_o[26];
  assign data_o[6618] = data_o[26];
  assign data_o[6682] = data_o[26];
  assign data_o[6746] = data_o[26];
  assign data_o[6810] = data_o[26];
  assign data_o[6874] = data_o[26];
  assign data_o[6938] = data_o[26];
  assign data_o[7002] = data_o[26];
  assign data_o[7066] = data_o[26];
  assign data_o[7130] = data_o[26];
  assign data_o[7194] = data_o[26];
  assign data_o[7258] = data_o[26];
  assign data_o[7322] = data_o[26];
  assign data_o[7386] = data_o[26];
  assign data_o[7450] = data_o[26];
  assign data_o[7514] = data_o[26];
  assign data_o[7578] = data_o[26];
  assign data_o[7642] = data_o[26];
  assign data_o[7706] = data_o[26];
  assign data_o[7770] = data_o[26];
  assign data_o[7834] = data_o[26];
  assign data_o[7898] = data_o[26];
  assign data_o[7962] = data_o[26];
  assign data_o[8026] = data_o[26];
  assign data_o[8090] = data_o[26];
  assign data_o[8154] = data_o[26];
  assign data_o[8218] = data_o[26];
  assign data_o[8282] = data_o[26];
  assign data_o[8346] = data_o[26];
  assign data_o[8410] = data_o[26];
  assign data_o[8474] = data_o[26];
  assign data_o[8538] = data_o[26];
  assign data_o[8602] = data_o[26];
  assign data_o[8666] = data_o[26];
  assign data_o[8730] = data_o[26];
  assign data_o[8794] = data_o[26];
  assign data_o[8858] = data_o[26];
  assign data_o[8922] = data_o[26];
  assign data_o[8986] = data_o[26];
  assign data_o[9050] = data_o[26];
  assign data_o[9114] = data_o[26];
  assign data_o[9178] = data_o[26];
  assign data_o[9242] = data_o[26];
  assign data_o[9306] = data_o[26];
  assign data_o[9370] = data_o[26];
  assign data_o[9434] = data_o[26];
  assign data_o[9498] = data_o[26];
  assign data_o[9562] = data_o[26];
  assign data_o[9626] = data_o[26];
  assign data_o[9690] = data_o[26];
  assign data_o[9754] = data_o[26];
  assign data_o[9818] = data_o[26];
  assign data_o[9882] = data_o[26];
  assign data_o[9946] = data_o[26];
  assign data_o[10010] = data_o[26];
  assign data_o[10074] = data_o[26];
  assign data_o[10138] = data_o[26];
  assign data_o[10202] = data_o[26];
  assign data_o[10266] = data_o[26];
  assign data_o[10330] = data_o[26];
  assign data_o[10394] = data_o[26];
  assign data_o[10458] = data_o[26];
  assign data_o[10522] = data_o[26];
  assign data_o[10586] = data_o[26];
  assign data_o[10650] = data_o[26];
  assign data_o[10714] = data_o[26];
  assign data_o[10778] = data_o[26];
  assign data_o[10842] = data_o[26];
  assign data_o[10906] = data_o[26];
  assign data_o[10970] = data_o[26];
  assign data_o[11034] = data_o[26];
  assign data_o[11098] = data_o[26];
  assign data_o[11162] = data_o[26];
  assign data_o[11226] = data_o[26];
  assign data_o[11290] = data_o[26];
  assign data_o[11354] = data_o[26];
  assign data_o[11418] = data_o[26];
  assign data_o[11482] = data_o[26];
  assign data_o[11546] = data_o[26];
  assign data_o[11610] = data_o[26];
  assign data_o[11674] = data_o[26];
  assign data_o[11738] = data_o[26];
  assign data_o[11802] = data_o[26];
  assign data_o[11866] = data_o[26];
  assign data_o[11930] = data_o[26];
  assign data_o[11994] = data_o[26];
  assign data_o[12058] = data_o[26];
  assign data_o[12122] = data_o[26];
  assign data_o[12186] = data_o[26];
  assign data_o[12250] = data_o[26];
  assign data_o[12314] = data_o[26];
  assign data_o[12378] = data_o[26];
  assign data_o[12442] = data_o[26];
  assign data_o[12506] = data_o[26];
  assign data_o[12570] = data_o[26];
  assign data_o[12634] = data_o[26];
  assign data_o[12698] = data_o[26];
  assign data_o[12762] = data_o[26];
  assign data_o[12826] = data_o[26];
  assign data_o[12890] = data_o[26];
  assign data_o[12954] = data_o[26];
  assign data_o[13018] = data_o[26];
  assign data_o[13082] = data_o[26];
  assign data_o[13146] = data_o[26];
  assign data_o[13210] = data_o[26];
  assign data_o[13274] = data_o[26];
  assign data_o[13338] = data_o[26];
  assign data_o[13402] = data_o[26];
  assign data_o[13466] = data_o[26];
  assign data_o[13530] = data_o[26];
  assign data_o[13594] = data_o[26];
  assign data_o[13658] = data_o[26];
  assign data_o[13722] = data_o[26];
  assign data_o[13786] = data_o[26];
  assign data_o[13850] = data_o[26];
  assign data_o[13914] = data_o[26];
  assign data_o[13978] = data_o[26];
  assign data_o[14042] = data_o[26];
  assign data_o[14106] = data_o[26];
  assign data_o[14170] = data_o[26];
  assign data_o[14234] = data_o[26];
  assign data_o[14298] = data_o[26];
  assign data_o[14362] = data_o[26];
  assign data_o[14426] = data_o[26];
  assign data_o[14490] = data_o[26];
  assign data_o[14554] = data_o[26];
  assign data_o[14618] = data_o[26];
  assign data_o[14682] = data_o[26];
  assign data_o[14746] = data_o[26];
  assign data_o[14810] = data_o[26];
  assign data_o[14874] = data_o[26];
  assign data_o[14938] = data_o[26];
  assign data_o[15002] = data_o[26];
  assign data_o[15066] = data_o[26];
  assign data_o[15130] = data_o[26];
  assign data_o[15194] = data_o[26];
  assign data_o[15258] = data_o[26];
  assign data_o[15322] = data_o[26];
  assign data_o[15386] = data_o[26];
  assign data_o[15450] = data_o[26];
  assign data_o[15514] = data_o[26];
  assign data_o[15578] = data_o[26];
  assign data_o[15642] = data_o[26];
  assign data_o[15706] = data_o[26];
  assign data_o[15770] = data_o[26];
  assign data_o[15834] = data_o[26];
  assign data_o[15898] = data_o[26];
  assign data_o[15962] = data_o[26];
  assign data_o[16026] = data_o[26];
  assign data_o[16090] = data_o[26];
  assign data_o[16154] = data_o[26];
  assign data_o[16218] = data_o[26];
  assign data_o[16282] = data_o[26];
  assign data_o[16346] = data_o[26];
  assign data_o[16410] = data_o[26];
  assign data_o[16474] = data_o[26];
  assign data_o[16538] = data_o[26];
  assign data_o[16602] = data_o[26];
  assign data_o[16666] = data_o[26];
  assign data_o[16730] = data_o[26];
  assign data_o[16794] = data_o[26];
  assign data_o[16858] = data_o[26];
  assign data_o[16922] = data_o[26];
  assign data_o[16986] = data_o[26];
  assign data_o[17050] = data_o[26];
  assign data_o[17114] = data_o[26];
  assign data_o[17178] = data_o[26];
  assign data_o[17242] = data_o[26];
  assign data_o[17306] = data_o[26];
  assign data_o[17370] = data_o[26];
  assign data_o[17434] = data_o[26];
  assign data_o[17498] = data_o[26];
  assign data_o[17562] = data_o[26];
  assign data_o[17626] = data_o[26];
  assign data_o[17690] = data_o[26];
  assign data_o[17754] = data_o[26];
  assign data_o[17818] = data_o[26];
  assign data_o[17882] = data_o[26];
  assign data_o[17946] = data_o[26];
  assign data_o[18010] = data_o[26];
  assign data_o[18074] = data_o[26];
  assign data_o[18138] = data_o[26];
  assign data_o[18202] = data_o[26];
  assign data_o[18266] = data_o[26];
  assign data_o[18330] = data_o[26];
  assign data_o[18394] = data_o[26];
  assign data_o[18458] = data_o[26];
  assign data_o[18522] = data_o[26];
  assign data_o[18586] = data_o[26];
  assign data_o[18650] = data_o[26];
  assign data_o[18714] = data_o[26];
  assign data_o[18778] = data_o[26];
  assign data_o[18842] = data_o[26];
  assign data_o[18906] = data_o[26];
  assign data_o[18970] = data_o[26];
  assign data_o[19034] = data_o[26];
  assign data_o[19098] = data_o[26];
  assign data_o[19162] = data_o[26];
  assign data_o[19226] = data_o[26];
  assign data_o[19290] = data_o[26];
  assign data_o[19354] = data_o[26];
  assign data_o[19418] = data_o[26];
  assign data_o[19482] = data_o[26];
  assign data_o[19546] = data_o[26];
  assign data_o[19610] = data_o[26];
  assign data_o[19674] = data_o[26];
  assign data_o[19738] = data_o[26];
  assign data_o[19802] = data_o[26];
  assign data_o[19866] = data_o[26];
  assign data_o[19930] = data_o[26];
  assign data_o[19994] = data_o[26];
  assign data_o[20058] = data_o[26];
  assign data_o[20122] = data_o[26];
  assign data_o[20186] = data_o[26];
  assign data_o[20250] = data_o[26];
  assign data_o[20314] = data_o[26];
  assign data_o[20378] = data_o[26];
  assign data_o[20442] = data_o[26];
  assign data_o[20506] = data_o[26];
  assign data_o[20570] = data_o[26];
  assign data_o[20634] = data_o[26];
  assign data_o[20698] = data_o[26];
  assign data_o[20762] = data_o[26];
  assign data_o[20826] = data_o[26];
  assign data_o[20890] = data_o[26];
  assign data_o[20954] = data_o[26];
  assign data_o[21018] = data_o[26];
  assign data_o[21082] = data_o[26];
  assign data_o[21146] = data_o[26];
  assign data_o[21210] = data_o[26];
  assign data_o[21274] = data_o[26];
  assign data_o[21338] = data_o[26];
  assign data_o[21402] = data_o[26];
  assign data_o[21466] = data_o[26];
  assign data_o[21530] = data_o[26];
  assign data_o[21594] = data_o[26];
  assign data_o[21658] = data_o[26];
  assign data_o[21722] = data_o[26];
  assign data_o[21786] = data_o[26];
  assign data_o[21850] = data_o[26];
  assign data_o[21914] = data_o[26];
  assign data_o[21978] = data_o[26];
  assign data_o[22042] = data_o[26];
  assign data_o[22106] = data_o[26];
  assign data_o[22170] = data_o[26];
  assign data_o[22234] = data_o[26];
  assign data_o[22298] = data_o[26];
  assign data_o[22362] = data_o[26];
  assign data_o[22426] = data_o[26];
  assign data_o[22490] = data_o[26];
  assign data_o[22554] = data_o[26];
  assign data_o[22618] = data_o[26];
  assign data_o[22682] = data_o[26];
  assign data_o[22746] = data_o[26];
  assign data_o[22810] = data_o[26];
  assign data_o[22874] = data_o[26];
  assign data_o[22938] = data_o[26];
  assign data_o[23002] = data_o[26];
  assign data_o[23066] = data_o[26];
  assign data_o[23130] = data_o[26];
  assign data_o[23194] = data_o[26];
  assign data_o[23258] = data_o[26];
  assign data_o[23322] = data_o[26];
  assign data_o[23386] = data_o[26];
  assign data_o[23450] = data_o[26];
  assign data_o[23514] = data_o[26];
  assign data_o[23578] = data_o[26];
  assign data_o[23642] = data_o[26];
  assign data_o[23706] = data_o[26];
  assign data_o[23770] = data_o[26];
  assign data_o[23834] = data_o[26];
  assign data_o[23898] = data_o[26];
  assign data_o[23962] = data_o[26];
  assign data_o[24026] = data_o[26];
  assign data_o[24090] = data_o[26];
  assign data_o[24154] = data_o[26];
  assign data_o[24218] = data_o[26];
  assign data_o[24282] = data_o[26];
  assign data_o[24346] = data_o[26];
  assign data_o[24410] = data_o[26];
  assign data_o[24474] = data_o[26];
  assign data_o[24538] = data_o[26];
  assign data_o[24602] = data_o[26];
  assign data_o[24666] = data_o[26];
  assign data_o[24730] = data_o[26];
  assign data_o[24794] = data_o[26];
  assign data_o[24858] = data_o[26];
  assign data_o[24922] = data_o[26];
  assign data_o[24986] = data_o[26];
  assign data_o[25050] = data_o[26];
  assign data_o[25114] = data_o[26];
  assign data_o[25178] = data_o[26];
  assign data_o[25242] = data_o[26];
  assign data_o[25306] = data_o[26];
  assign data_o[25370] = data_o[26];
  assign data_o[25434] = data_o[26];
  assign data_o[25498] = data_o[26];
  assign data_o[25562] = data_o[26];
  assign data_o[25626] = data_o[26];
  assign data_o[25690] = data_o[26];
  assign data_o[25754] = data_o[26];
  assign data_o[25818] = data_o[26];
  assign data_o[25882] = data_o[26];
  assign data_o[25946] = data_o[26];
  assign data_o[26010] = data_o[26];
  assign data_o[26074] = data_o[26];
  assign data_o[26138] = data_o[26];
  assign data_o[26202] = data_o[26];
  assign data_o[26266] = data_o[26];
  assign data_o[26330] = data_o[26];
  assign data_o[26394] = data_o[26];
  assign data_o[26458] = data_o[26];
  assign data_o[26522] = data_o[26];
  assign data_o[26586] = data_o[26];
  assign data_o[26650] = data_o[26];
  assign data_o[26714] = data_o[26];
  assign data_o[26778] = data_o[26];
  assign data_o[26842] = data_o[26];
  assign data_o[26906] = data_o[26];
  assign data_o[26970] = data_o[26];
  assign data_o[27034] = data_o[26];
  assign data_o[27098] = data_o[26];
  assign data_o[27162] = data_o[26];
  assign data_o[27226] = data_o[26];
  assign data_o[27290] = data_o[26];
  assign data_o[27354] = data_o[26];
  assign data_o[27418] = data_o[26];
  assign data_o[27482] = data_o[26];
  assign data_o[27546] = data_o[26];
  assign data_o[27610] = data_o[26];
  assign data_o[27674] = data_o[26];
  assign data_o[27738] = data_o[26];
  assign data_o[27802] = data_o[26];
  assign data_o[27866] = data_o[26];
  assign data_o[27930] = data_o[26];
  assign data_o[27994] = data_o[26];
  assign data_o[28058] = data_o[26];
  assign data_o[28122] = data_o[26];
  assign data_o[28186] = data_o[26];
  assign data_o[28250] = data_o[26];
  assign data_o[28314] = data_o[26];
  assign data_o[28378] = data_o[26];
  assign data_o[28442] = data_o[26];
  assign data_o[28506] = data_o[26];
  assign data_o[28570] = data_o[26];
  assign data_o[28634] = data_o[26];
  assign data_o[28698] = data_o[26];
  assign data_o[28762] = data_o[26];
  assign data_o[28826] = data_o[26];
  assign data_o[28890] = data_o[26];
  assign data_o[28954] = data_o[26];
  assign data_o[29018] = data_o[26];
  assign data_o[29082] = data_o[26];
  assign data_o[29146] = data_o[26];
  assign data_o[29210] = data_o[26];
  assign data_o[29274] = data_o[26];
  assign data_o[29338] = data_o[26];
  assign data_o[29402] = data_o[26];
  assign data_o[29466] = data_o[26];
  assign data_o[29530] = data_o[26];
  assign data_o[29594] = data_o[26];
  assign data_o[29658] = data_o[26];
  assign data_o[29722] = data_o[26];
  assign data_o[29786] = data_o[26];
  assign data_o[29850] = data_o[26];
  assign data_o[29914] = data_o[26];
  assign data_o[29978] = data_o[26];
  assign data_o[30042] = data_o[26];
  assign data_o[30106] = data_o[26];
  assign data_o[30170] = data_o[26];
  assign data_o[30234] = data_o[26];
  assign data_o[30298] = data_o[26];
  assign data_o[30362] = data_o[26];
  assign data_o[30426] = data_o[26];
  assign data_o[30490] = data_o[26];
  assign data_o[30554] = data_o[26];
  assign data_o[30618] = data_o[26];
  assign data_o[30682] = data_o[26];
  assign data_o[30746] = data_o[26];
  assign data_o[30810] = data_o[26];
  assign data_o[30874] = data_o[26];
  assign data_o[30938] = data_o[26];
  assign data_o[31002] = data_o[26];
  assign data_o[31066] = data_o[26];
  assign data_o[31130] = data_o[26];
  assign data_o[31194] = data_o[26];
  assign data_o[31258] = data_o[26];
  assign data_o[31322] = data_o[26];
  assign data_o[31386] = data_o[26];
  assign data_o[31450] = data_o[26];
  assign data_o[31514] = data_o[26];
  assign data_o[31578] = data_o[26];
  assign data_o[31642] = data_o[26];
  assign data_o[31706] = data_o[26];
  assign data_o[31770] = data_o[26];
  assign data_o[31834] = data_o[26];
  assign data_o[31898] = data_o[26];
  assign data_o[31962] = data_o[26];
  assign data_o[89] = data_o[25];
  assign data_o[153] = data_o[25];
  assign data_o[217] = data_o[25];
  assign data_o[281] = data_o[25];
  assign data_o[345] = data_o[25];
  assign data_o[409] = data_o[25];
  assign data_o[473] = data_o[25];
  assign data_o[537] = data_o[25];
  assign data_o[601] = data_o[25];
  assign data_o[665] = data_o[25];
  assign data_o[729] = data_o[25];
  assign data_o[793] = data_o[25];
  assign data_o[857] = data_o[25];
  assign data_o[921] = data_o[25];
  assign data_o[985] = data_o[25];
  assign data_o[1049] = data_o[25];
  assign data_o[1113] = data_o[25];
  assign data_o[1177] = data_o[25];
  assign data_o[1241] = data_o[25];
  assign data_o[1305] = data_o[25];
  assign data_o[1369] = data_o[25];
  assign data_o[1433] = data_o[25];
  assign data_o[1497] = data_o[25];
  assign data_o[1561] = data_o[25];
  assign data_o[1625] = data_o[25];
  assign data_o[1689] = data_o[25];
  assign data_o[1753] = data_o[25];
  assign data_o[1817] = data_o[25];
  assign data_o[1881] = data_o[25];
  assign data_o[1945] = data_o[25];
  assign data_o[2009] = data_o[25];
  assign data_o[2073] = data_o[25];
  assign data_o[2137] = data_o[25];
  assign data_o[2201] = data_o[25];
  assign data_o[2265] = data_o[25];
  assign data_o[2329] = data_o[25];
  assign data_o[2393] = data_o[25];
  assign data_o[2457] = data_o[25];
  assign data_o[2521] = data_o[25];
  assign data_o[2585] = data_o[25];
  assign data_o[2649] = data_o[25];
  assign data_o[2713] = data_o[25];
  assign data_o[2777] = data_o[25];
  assign data_o[2841] = data_o[25];
  assign data_o[2905] = data_o[25];
  assign data_o[2969] = data_o[25];
  assign data_o[3033] = data_o[25];
  assign data_o[3097] = data_o[25];
  assign data_o[3161] = data_o[25];
  assign data_o[3225] = data_o[25];
  assign data_o[3289] = data_o[25];
  assign data_o[3353] = data_o[25];
  assign data_o[3417] = data_o[25];
  assign data_o[3481] = data_o[25];
  assign data_o[3545] = data_o[25];
  assign data_o[3609] = data_o[25];
  assign data_o[3673] = data_o[25];
  assign data_o[3737] = data_o[25];
  assign data_o[3801] = data_o[25];
  assign data_o[3865] = data_o[25];
  assign data_o[3929] = data_o[25];
  assign data_o[3993] = data_o[25];
  assign data_o[4057] = data_o[25];
  assign data_o[4121] = data_o[25];
  assign data_o[4185] = data_o[25];
  assign data_o[4249] = data_o[25];
  assign data_o[4313] = data_o[25];
  assign data_o[4377] = data_o[25];
  assign data_o[4441] = data_o[25];
  assign data_o[4505] = data_o[25];
  assign data_o[4569] = data_o[25];
  assign data_o[4633] = data_o[25];
  assign data_o[4697] = data_o[25];
  assign data_o[4761] = data_o[25];
  assign data_o[4825] = data_o[25];
  assign data_o[4889] = data_o[25];
  assign data_o[4953] = data_o[25];
  assign data_o[5017] = data_o[25];
  assign data_o[5081] = data_o[25];
  assign data_o[5145] = data_o[25];
  assign data_o[5209] = data_o[25];
  assign data_o[5273] = data_o[25];
  assign data_o[5337] = data_o[25];
  assign data_o[5401] = data_o[25];
  assign data_o[5465] = data_o[25];
  assign data_o[5529] = data_o[25];
  assign data_o[5593] = data_o[25];
  assign data_o[5657] = data_o[25];
  assign data_o[5721] = data_o[25];
  assign data_o[5785] = data_o[25];
  assign data_o[5849] = data_o[25];
  assign data_o[5913] = data_o[25];
  assign data_o[5977] = data_o[25];
  assign data_o[6041] = data_o[25];
  assign data_o[6105] = data_o[25];
  assign data_o[6169] = data_o[25];
  assign data_o[6233] = data_o[25];
  assign data_o[6297] = data_o[25];
  assign data_o[6361] = data_o[25];
  assign data_o[6425] = data_o[25];
  assign data_o[6489] = data_o[25];
  assign data_o[6553] = data_o[25];
  assign data_o[6617] = data_o[25];
  assign data_o[6681] = data_o[25];
  assign data_o[6745] = data_o[25];
  assign data_o[6809] = data_o[25];
  assign data_o[6873] = data_o[25];
  assign data_o[6937] = data_o[25];
  assign data_o[7001] = data_o[25];
  assign data_o[7065] = data_o[25];
  assign data_o[7129] = data_o[25];
  assign data_o[7193] = data_o[25];
  assign data_o[7257] = data_o[25];
  assign data_o[7321] = data_o[25];
  assign data_o[7385] = data_o[25];
  assign data_o[7449] = data_o[25];
  assign data_o[7513] = data_o[25];
  assign data_o[7577] = data_o[25];
  assign data_o[7641] = data_o[25];
  assign data_o[7705] = data_o[25];
  assign data_o[7769] = data_o[25];
  assign data_o[7833] = data_o[25];
  assign data_o[7897] = data_o[25];
  assign data_o[7961] = data_o[25];
  assign data_o[8025] = data_o[25];
  assign data_o[8089] = data_o[25];
  assign data_o[8153] = data_o[25];
  assign data_o[8217] = data_o[25];
  assign data_o[8281] = data_o[25];
  assign data_o[8345] = data_o[25];
  assign data_o[8409] = data_o[25];
  assign data_o[8473] = data_o[25];
  assign data_o[8537] = data_o[25];
  assign data_o[8601] = data_o[25];
  assign data_o[8665] = data_o[25];
  assign data_o[8729] = data_o[25];
  assign data_o[8793] = data_o[25];
  assign data_o[8857] = data_o[25];
  assign data_o[8921] = data_o[25];
  assign data_o[8985] = data_o[25];
  assign data_o[9049] = data_o[25];
  assign data_o[9113] = data_o[25];
  assign data_o[9177] = data_o[25];
  assign data_o[9241] = data_o[25];
  assign data_o[9305] = data_o[25];
  assign data_o[9369] = data_o[25];
  assign data_o[9433] = data_o[25];
  assign data_o[9497] = data_o[25];
  assign data_o[9561] = data_o[25];
  assign data_o[9625] = data_o[25];
  assign data_o[9689] = data_o[25];
  assign data_o[9753] = data_o[25];
  assign data_o[9817] = data_o[25];
  assign data_o[9881] = data_o[25];
  assign data_o[9945] = data_o[25];
  assign data_o[10009] = data_o[25];
  assign data_o[10073] = data_o[25];
  assign data_o[10137] = data_o[25];
  assign data_o[10201] = data_o[25];
  assign data_o[10265] = data_o[25];
  assign data_o[10329] = data_o[25];
  assign data_o[10393] = data_o[25];
  assign data_o[10457] = data_o[25];
  assign data_o[10521] = data_o[25];
  assign data_o[10585] = data_o[25];
  assign data_o[10649] = data_o[25];
  assign data_o[10713] = data_o[25];
  assign data_o[10777] = data_o[25];
  assign data_o[10841] = data_o[25];
  assign data_o[10905] = data_o[25];
  assign data_o[10969] = data_o[25];
  assign data_o[11033] = data_o[25];
  assign data_o[11097] = data_o[25];
  assign data_o[11161] = data_o[25];
  assign data_o[11225] = data_o[25];
  assign data_o[11289] = data_o[25];
  assign data_o[11353] = data_o[25];
  assign data_o[11417] = data_o[25];
  assign data_o[11481] = data_o[25];
  assign data_o[11545] = data_o[25];
  assign data_o[11609] = data_o[25];
  assign data_o[11673] = data_o[25];
  assign data_o[11737] = data_o[25];
  assign data_o[11801] = data_o[25];
  assign data_o[11865] = data_o[25];
  assign data_o[11929] = data_o[25];
  assign data_o[11993] = data_o[25];
  assign data_o[12057] = data_o[25];
  assign data_o[12121] = data_o[25];
  assign data_o[12185] = data_o[25];
  assign data_o[12249] = data_o[25];
  assign data_o[12313] = data_o[25];
  assign data_o[12377] = data_o[25];
  assign data_o[12441] = data_o[25];
  assign data_o[12505] = data_o[25];
  assign data_o[12569] = data_o[25];
  assign data_o[12633] = data_o[25];
  assign data_o[12697] = data_o[25];
  assign data_o[12761] = data_o[25];
  assign data_o[12825] = data_o[25];
  assign data_o[12889] = data_o[25];
  assign data_o[12953] = data_o[25];
  assign data_o[13017] = data_o[25];
  assign data_o[13081] = data_o[25];
  assign data_o[13145] = data_o[25];
  assign data_o[13209] = data_o[25];
  assign data_o[13273] = data_o[25];
  assign data_o[13337] = data_o[25];
  assign data_o[13401] = data_o[25];
  assign data_o[13465] = data_o[25];
  assign data_o[13529] = data_o[25];
  assign data_o[13593] = data_o[25];
  assign data_o[13657] = data_o[25];
  assign data_o[13721] = data_o[25];
  assign data_o[13785] = data_o[25];
  assign data_o[13849] = data_o[25];
  assign data_o[13913] = data_o[25];
  assign data_o[13977] = data_o[25];
  assign data_o[14041] = data_o[25];
  assign data_o[14105] = data_o[25];
  assign data_o[14169] = data_o[25];
  assign data_o[14233] = data_o[25];
  assign data_o[14297] = data_o[25];
  assign data_o[14361] = data_o[25];
  assign data_o[14425] = data_o[25];
  assign data_o[14489] = data_o[25];
  assign data_o[14553] = data_o[25];
  assign data_o[14617] = data_o[25];
  assign data_o[14681] = data_o[25];
  assign data_o[14745] = data_o[25];
  assign data_o[14809] = data_o[25];
  assign data_o[14873] = data_o[25];
  assign data_o[14937] = data_o[25];
  assign data_o[15001] = data_o[25];
  assign data_o[15065] = data_o[25];
  assign data_o[15129] = data_o[25];
  assign data_o[15193] = data_o[25];
  assign data_o[15257] = data_o[25];
  assign data_o[15321] = data_o[25];
  assign data_o[15385] = data_o[25];
  assign data_o[15449] = data_o[25];
  assign data_o[15513] = data_o[25];
  assign data_o[15577] = data_o[25];
  assign data_o[15641] = data_o[25];
  assign data_o[15705] = data_o[25];
  assign data_o[15769] = data_o[25];
  assign data_o[15833] = data_o[25];
  assign data_o[15897] = data_o[25];
  assign data_o[15961] = data_o[25];
  assign data_o[16025] = data_o[25];
  assign data_o[16089] = data_o[25];
  assign data_o[16153] = data_o[25];
  assign data_o[16217] = data_o[25];
  assign data_o[16281] = data_o[25];
  assign data_o[16345] = data_o[25];
  assign data_o[16409] = data_o[25];
  assign data_o[16473] = data_o[25];
  assign data_o[16537] = data_o[25];
  assign data_o[16601] = data_o[25];
  assign data_o[16665] = data_o[25];
  assign data_o[16729] = data_o[25];
  assign data_o[16793] = data_o[25];
  assign data_o[16857] = data_o[25];
  assign data_o[16921] = data_o[25];
  assign data_o[16985] = data_o[25];
  assign data_o[17049] = data_o[25];
  assign data_o[17113] = data_o[25];
  assign data_o[17177] = data_o[25];
  assign data_o[17241] = data_o[25];
  assign data_o[17305] = data_o[25];
  assign data_o[17369] = data_o[25];
  assign data_o[17433] = data_o[25];
  assign data_o[17497] = data_o[25];
  assign data_o[17561] = data_o[25];
  assign data_o[17625] = data_o[25];
  assign data_o[17689] = data_o[25];
  assign data_o[17753] = data_o[25];
  assign data_o[17817] = data_o[25];
  assign data_o[17881] = data_o[25];
  assign data_o[17945] = data_o[25];
  assign data_o[18009] = data_o[25];
  assign data_o[18073] = data_o[25];
  assign data_o[18137] = data_o[25];
  assign data_o[18201] = data_o[25];
  assign data_o[18265] = data_o[25];
  assign data_o[18329] = data_o[25];
  assign data_o[18393] = data_o[25];
  assign data_o[18457] = data_o[25];
  assign data_o[18521] = data_o[25];
  assign data_o[18585] = data_o[25];
  assign data_o[18649] = data_o[25];
  assign data_o[18713] = data_o[25];
  assign data_o[18777] = data_o[25];
  assign data_o[18841] = data_o[25];
  assign data_o[18905] = data_o[25];
  assign data_o[18969] = data_o[25];
  assign data_o[19033] = data_o[25];
  assign data_o[19097] = data_o[25];
  assign data_o[19161] = data_o[25];
  assign data_o[19225] = data_o[25];
  assign data_o[19289] = data_o[25];
  assign data_o[19353] = data_o[25];
  assign data_o[19417] = data_o[25];
  assign data_o[19481] = data_o[25];
  assign data_o[19545] = data_o[25];
  assign data_o[19609] = data_o[25];
  assign data_o[19673] = data_o[25];
  assign data_o[19737] = data_o[25];
  assign data_o[19801] = data_o[25];
  assign data_o[19865] = data_o[25];
  assign data_o[19929] = data_o[25];
  assign data_o[19993] = data_o[25];
  assign data_o[20057] = data_o[25];
  assign data_o[20121] = data_o[25];
  assign data_o[20185] = data_o[25];
  assign data_o[20249] = data_o[25];
  assign data_o[20313] = data_o[25];
  assign data_o[20377] = data_o[25];
  assign data_o[20441] = data_o[25];
  assign data_o[20505] = data_o[25];
  assign data_o[20569] = data_o[25];
  assign data_o[20633] = data_o[25];
  assign data_o[20697] = data_o[25];
  assign data_o[20761] = data_o[25];
  assign data_o[20825] = data_o[25];
  assign data_o[20889] = data_o[25];
  assign data_o[20953] = data_o[25];
  assign data_o[21017] = data_o[25];
  assign data_o[21081] = data_o[25];
  assign data_o[21145] = data_o[25];
  assign data_o[21209] = data_o[25];
  assign data_o[21273] = data_o[25];
  assign data_o[21337] = data_o[25];
  assign data_o[21401] = data_o[25];
  assign data_o[21465] = data_o[25];
  assign data_o[21529] = data_o[25];
  assign data_o[21593] = data_o[25];
  assign data_o[21657] = data_o[25];
  assign data_o[21721] = data_o[25];
  assign data_o[21785] = data_o[25];
  assign data_o[21849] = data_o[25];
  assign data_o[21913] = data_o[25];
  assign data_o[21977] = data_o[25];
  assign data_o[22041] = data_o[25];
  assign data_o[22105] = data_o[25];
  assign data_o[22169] = data_o[25];
  assign data_o[22233] = data_o[25];
  assign data_o[22297] = data_o[25];
  assign data_o[22361] = data_o[25];
  assign data_o[22425] = data_o[25];
  assign data_o[22489] = data_o[25];
  assign data_o[22553] = data_o[25];
  assign data_o[22617] = data_o[25];
  assign data_o[22681] = data_o[25];
  assign data_o[22745] = data_o[25];
  assign data_o[22809] = data_o[25];
  assign data_o[22873] = data_o[25];
  assign data_o[22937] = data_o[25];
  assign data_o[23001] = data_o[25];
  assign data_o[23065] = data_o[25];
  assign data_o[23129] = data_o[25];
  assign data_o[23193] = data_o[25];
  assign data_o[23257] = data_o[25];
  assign data_o[23321] = data_o[25];
  assign data_o[23385] = data_o[25];
  assign data_o[23449] = data_o[25];
  assign data_o[23513] = data_o[25];
  assign data_o[23577] = data_o[25];
  assign data_o[23641] = data_o[25];
  assign data_o[23705] = data_o[25];
  assign data_o[23769] = data_o[25];
  assign data_o[23833] = data_o[25];
  assign data_o[23897] = data_o[25];
  assign data_o[23961] = data_o[25];
  assign data_o[24025] = data_o[25];
  assign data_o[24089] = data_o[25];
  assign data_o[24153] = data_o[25];
  assign data_o[24217] = data_o[25];
  assign data_o[24281] = data_o[25];
  assign data_o[24345] = data_o[25];
  assign data_o[24409] = data_o[25];
  assign data_o[24473] = data_o[25];
  assign data_o[24537] = data_o[25];
  assign data_o[24601] = data_o[25];
  assign data_o[24665] = data_o[25];
  assign data_o[24729] = data_o[25];
  assign data_o[24793] = data_o[25];
  assign data_o[24857] = data_o[25];
  assign data_o[24921] = data_o[25];
  assign data_o[24985] = data_o[25];
  assign data_o[25049] = data_o[25];
  assign data_o[25113] = data_o[25];
  assign data_o[25177] = data_o[25];
  assign data_o[25241] = data_o[25];
  assign data_o[25305] = data_o[25];
  assign data_o[25369] = data_o[25];
  assign data_o[25433] = data_o[25];
  assign data_o[25497] = data_o[25];
  assign data_o[25561] = data_o[25];
  assign data_o[25625] = data_o[25];
  assign data_o[25689] = data_o[25];
  assign data_o[25753] = data_o[25];
  assign data_o[25817] = data_o[25];
  assign data_o[25881] = data_o[25];
  assign data_o[25945] = data_o[25];
  assign data_o[26009] = data_o[25];
  assign data_o[26073] = data_o[25];
  assign data_o[26137] = data_o[25];
  assign data_o[26201] = data_o[25];
  assign data_o[26265] = data_o[25];
  assign data_o[26329] = data_o[25];
  assign data_o[26393] = data_o[25];
  assign data_o[26457] = data_o[25];
  assign data_o[26521] = data_o[25];
  assign data_o[26585] = data_o[25];
  assign data_o[26649] = data_o[25];
  assign data_o[26713] = data_o[25];
  assign data_o[26777] = data_o[25];
  assign data_o[26841] = data_o[25];
  assign data_o[26905] = data_o[25];
  assign data_o[26969] = data_o[25];
  assign data_o[27033] = data_o[25];
  assign data_o[27097] = data_o[25];
  assign data_o[27161] = data_o[25];
  assign data_o[27225] = data_o[25];
  assign data_o[27289] = data_o[25];
  assign data_o[27353] = data_o[25];
  assign data_o[27417] = data_o[25];
  assign data_o[27481] = data_o[25];
  assign data_o[27545] = data_o[25];
  assign data_o[27609] = data_o[25];
  assign data_o[27673] = data_o[25];
  assign data_o[27737] = data_o[25];
  assign data_o[27801] = data_o[25];
  assign data_o[27865] = data_o[25];
  assign data_o[27929] = data_o[25];
  assign data_o[27993] = data_o[25];
  assign data_o[28057] = data_o[25];
  assign data_o[28121] = data_o[25];
  assign data_o[28185] = data_o[25];
  assign data_o[28249] = data_o[25];
  assign data_o[28313] = data_o[25];
  assign data_o[28377] = data_o[25];
  assign data_o[28441] = data_o[25];
  assign data_o[28505] = data_o[25];
  assign data_o[28569] = data_o[25];
  assign data_o[28633] = data_o[25];
  assign data_o[28697] = data_o[25];
  assign data_o[28761] = data_o[25];
  assign data_o[28825] = data_o[25];
  assign data_o[28889] = data_o[25];
  assign data_o[28953] = data_o[25];
  assign data_o[29017] = data_o[25];
  assign data_o[29081] = data_o[25];
  assign data_o[29145] = data_o[25];
  assign data_o[29209] = data_o[25];
  assign data_o[29273] = data_o[25];
  assign data_o[29337] = data_o[25];
  assign data_o[29401] = data_o[25];
  assign data_o[29465] = data_o[25];
  assign data_o[29529] = data_o[25];
  assign data_o[29593] = data_o[25];
  assign data_o[29657] = data_o[25];
  assign data_o[29721] = data_o[25];
  assign data_o[29785] = data_o[25];
  assign data_o[29849] = data_o[25];
  assign data_o[29913] = data_o[25];
  assign data_o[29977] = data_o[25];
  assign data_o[30041] = data_o[25];
  assign data_o[30105] = data_o[25];
  assign data_o[30169] = data_o[25];
  assign data_o[30233] = data_o[25];
  assign data_o[30297] = data_o[25];
  assign data_o[30361] = data_o[25];
  assign data_o[30425] = data_o[25];
  assign data_o[30489] = data_o[25];
  assign data_o[30553] = data_o[25];
  assign data_o[30617] = data_o[25];
  assign data_o[30681] = data_o[25];
  assign data_o[30745] = data_o[25];
  assign data_o[30809] = data_o[25];
  assign data_o[30873] = data_o[25];
  assign data_o[30937] = data_o[25];
  assign data_o[31001] = data_o[25];
  assign data_o[31065] = data_o[25];
  assign data_o[31129] = data_o[25];
  assign data_o[31193] = data_o[25];
  assign data_o[31257] = data_o[25];
  assign data_o[31321] = data_o[25];
  assign data_o[31385] = data_o[25];
  assign data_o[31449] = data_o[25];
  assign data_o[31513] = data_o[25];
  assign data_o[31577] = data_o[25];
  assign data_o[31641] = data_o[25];
  assign data_o[31705] = data_o[25];
  assign data_o[31769] = data_o[25];
  assign data_o[31833] = data_o[25];
  assign data_o[31897] = data_o[25];
  assign data_o[31961] = data_o[25];
  assign data_o[88] = data_o[24];
  assign data_o[152] = data_o[24];
  assign data_o[216] = data_o[24];
  assign data_o[280] = data_o[24];
  assign data_o[344] = data_o[24];
  assign data_o[408] = data_o[24];
  assign data_o[472] = data_o[24];
  assign data_o[536] = data_o[24];
  assign data_o[600] = data_o[24];
  assign data_o[664] = data_o[24];
  assign data_o[728] = data_o[24];
  assign data_o[792] = data_o[24];
  assign data_o[856] = data_o[24];
  assign data_o[920] = data_o[24];
  assign data_o[984] = data_o[24];
  assign data_o[1048] = data_o[24];
  assign data_o[1112] = data_o[24];
  assign data_o[1176] = data_o[24];
  assign data_o[1240] = data_o[24];
  assign data_o[1304] = data_o[24];
  assign data_o[1368] = data_o[24];
  assign data_o[1432] = data_o[24];
  assign data_o[1496] = data_o[24];
  assign data_o[1560] = data_o[24];
  assign data_o[1624] = data_o[24];
  assign data_o[1688] = data_o[24];
  assign data_o[1752] = data_o[24];
  assign data_o[1816] = data_o[24];
  assign data_o[1880] = data_o[24];
  assign data_o[1944] = data_o[24];
  assign data_o[2008] = data_o[24];
  assign data_o[2072] = data_o[24];
  assign data_o[2136] = data_o[24];
  assign data_o[2200] = data_o[24];
  assign data_o[2264] = data_o[24];
  assign data_o[2328] = data_o[24];
  assign data_o[2392] = data_o[24];
  assign data_o[2456] = data_o[24];
  assign data_o[2520] = data_o[24];
  assign data_o[2584] = data_o[24];
  assign data_o[2648] = data_o[24];
  assign data_o[2712] = data_o[24];
  assign data_o[2776] = data_o[24];
  assign data_o[2840] = data_o[24];
  assign data_o[2904] = data_o[24];
  assign data_o[2968] = data_o[24];
  assign data_o[3032] = data_o[24];
  assign data_o[3096] = data_o[24];
  assign data_o[3160] = data_o[24];
  assign data_o[3224] = data_o[24];
  assign data_o[3288] = data_o[24];
  assign data_o[3352] = data_o[24];
  assign data_o[3416] = data_o[24];
  assign data_o[3480] = data_o[24];
  assign data_o[3544] = data_o[24];
  assign data_o[3608] = data_o[24];
  assign data_o[3672] = data_o[24];
  assign data_o[3736] = data_o[24];
  assign data_o[3800] = data_o[24];
  assign data_o[3864] = data_o[24];
  assign data_o[3928] = data_o[24];
  assign data_o[3992] = data_o[24];
  assign data_o[4056] = data_o[24];
  assign data_o[4120] = data_o[24];
  assign data_o[4184] = data_o[24];
  assign data_o[4248] = data_o[24];
  assign data_o[4312] = data_o[24];
  assign data_o[4376] = data_o[24];
  assign data_o[4440] = data_o[24];
  assign data_o[4504] = data_o[24];
  assign data_o[4568] = data_o[24];
  assign data_o[4632] = data_o[24];
  assign data_o[4696] = data_o[24];
  assign data_o[4760] = data_o[24];
  assign data_o[4824] = data_o[24];
  assign data_o[4888] = data_o[24];
  assign data_o[4952] = data_o[24];
  assign data_o[5016] = data_o[24];
  assign data_o[5080] = data_o[24];
  assign data_o[5144] = data_o[24];
  assign data_o[5208] = data_o[24];
  assign data_o[5272] = data_o[24];
  assign data_o[5336] = data_o[24];
  assign data_o[5400] = data_o[24];
  assign data_o[5464] = data_o[24];
  assign data_o[5528] = data_o[24];
  assign data_o[5592] = data_o[24];
  assign data_o[5656] = data_o[24];
  assign data_o[5720] = data_o[24];
  assign data_o[5784] = data_o[24];
  assign data_o[5848] = data_o[24];
  assign data_o[5912] = data_o[24];
  assign data_o[5976] = data_o[24];
  assign data_o[6040] = data_o[24];
  assign data_o[6104] = data_o[24];
  assign data_o[6168] = data_o[24];
  assign data_o[6232] = data_o[24];
  assign data_o[6296] = data_o[24];
  assign data_o[6360] = data_o[24];
  assign data_o[6424] = data_o[24];
  assign data_o[6488] = data_o[24];
  assign data_o[6552] = data_o[24];
  assign data_o[6616] = data_o[24];
  assign data_o[6680] = data_o[24];
  assign data_o[6744] = data_o[24];
  assign data_o[6808] = data_o[24];
  assign data_o[6872] = data_o[24];
  assign data_o[6936] = data_o[24];
  assign data_o[7000] = data_o[24];
  assign data_o[7064] = data_o[24];
  assign data_o[7128] = data_o[24];
  assign data_o[7192] = data_o[24];
  assign data_o[7256] = data_o[24];
  assign data_o[7320] = data_o[24];
  assign data_o[7384] = data_o[24];
  assign data_o[7448] = data_o[24];
  assign data_o[7512] = data_o[24];
  assign data_o[7576] = data_o[24];
  assign data_o[7640] = data_o[24];
  assign data_o[7704] = data_o[24];
  assign data_o[7768] = data_o[24];
  assign data_o[7832] = data_o[24];
  assign data_o[7896] = data_o[24];
  assign data_o[7960] = data_o[24];
  assign data_o[8024] = data_o[24];
  assign data_o[8088] = data_o[24];
  assign data_o[8152] = data_o[24];
  assign data_o[8216] = data_o[24];
  assign data_o[8280] = data_o[24];
  assign data_o[8344] = data_o[24];
  assign data_o[8408] = data_o[24];
  assign data_o[8472] = data_o[24];
  assign data_o[8536] = data_o[24];
  assign data_o[8600] = data_o[24];
  assign data_o[8664] = data_o[24];
  assign data_o[8728] = data_o[24];
  assign data_o[8792] = data_o[24];
  assign data_o[8856] = data_o[24];
  assign data_o[8920] = data_o[24];
  assign data_o[8984] = data_o[24];
  assign data_o[9048] = data_o[24];
  assign data_o[9112] = data_o[24];
  assign data_o[9176] = data_o[24];
  assign data_o[9240] = data_o[24];
  assign data_o[9304] = data_o[24];
  assign data_o[9368] = data_o[24];
  assign data_o[9432] = data_o[24];
  assign data_o[9496] = data_o[24];
  assign data_o[9560] = data_o[24];
  assign data_o[9624] = data_o[24];
  assign data_o[9688] = data_o[24];
  assign data_o[9752] = data_o[24];
  assign data_o[9816] = data_o[24];
  assign data_o[9880] = data_o[24];
  assign data_o[9944] = data_o[24];
  assign data_o[10008] = data_o[24];
  assign data_o[10072] = data_o[24];
  assign data_o[10136] = data_o[24];
  assign data_o[10200] = data_o[24];
  assign data_o[10264] = data_o[24];
  assign data_o[10328] = data_o[24];
  assign data_o[10392] = data_o[24];
  assign data_o[10456] = data_o[24];
  assign data_o[10520] = data_o[24];
  assign data_o[10584] = data_o[24];
  assign data_o[10648] = data_o[24];
  assign data_o[10712] = data_o[24];
  assign data_o[10776] = data_o[24];
  assign data_o[10840] = data_o[24];
  assign data_o[10904] = data_o[24];
  assign data_o[10968] = data_o[24];
  assign data_o[11032] = data_o[24];
  assign data_o[11096] = data_o[24];
  assign data_o[11160] = data_o[24];
  assign data_o[11224] = data_o[24];
  assign data_o[11288] = data_o[24];
  assign data_o[11352] = data_o[24];
  assign data_o[11416] = data_o[24];
  assign data_o[11480] = data_o[24];
  assign data_o[11544] = data_o[24];
  assign data_o[11608] = data_o[24];
  assign data_o[11672] = data_o[24];
  assign data_o[11736] = data_o[24];
  assign data_o[11800] = data_o[24];
  assign data_o[11864] = data_o[24];
  assign data_o[11928] = data_o[24];
  assign data_o[11992] = data_o[24];
  assign data_o[12056] = data_o[24];
  assign data_o[12120] = data_o[24];
  assign data_o[12184] = data_o[24];
  assign data_o[12248] = data_o[24];
  assign data_o[12312] = data_o[24];
  assign data_o[12376] = data_o[24];
  assign data_o[12440] = data_o[24];
  assign data_o[12504] = data_o[24];
  assign data_o[12568] = data_o[24];
  assign data_o[12632] = data_o[24];
  assign data_o[12696] = data_o[24];
  assign data_o[12760] = data_o[24];
  assign data_o[12824] = data_o[24];
  assign data_o[12888] = data_o[24];
  assign data_o[12952] = data_o[24];
  assign data_o[13016] = data_o[24];
  assign data_o[13080] = data_o[24];
  assign data_o[13144] = data_o[24];
  assign data_o[13208] = data_o[24];
  assign data_o[13272] = data_o[24];
  assign data_o[13336] = data_o[24];
  assign data_o[13400] = data_o[24];
  assign data_o[13464] = data_o[24];
  assign data_o[13528] = data_o[24];
  assign data_o[13592] = data_o[24];
  assign data_o[13656] = data_o[24];
  assign data_o[13720] = data_o[24];
  assign data_o[13784] = data_o[24];
  assign data_o[13848] = data_o[24];
  assign data_o[13912] = data_o[24];
  assign data_o[13976] = data_o[24];
  assign data_o[14040] = data_o[24];
  assign data_o[14104] = data_o[24];
  assign data_o[14168] = data_o[24];
  assign data_o[14232] = data_o[24];
  assign data_o[14296] = data_o[24];
  assign data_o[14360] = data_o[24];
  assign data_o[14424] = data_o[24];
  assign data_o[14488] = data_o[24];
  assign data_o[14552] = data_o[24];
  assign data_o[14616] = data_o[24];
  assign data_o[14680] = data_o[24];
  assign data_o[14744] = data_o[24];
  assign data_o[14808] = data_o[24];
  assign data_o[14872] = data_o[24];
  assign data_o[14936] = data_o[24];
  assign data_o[15000] = data_o[24];
  assign data_o[15064] = data_o[24];
  assign data_o[15128] = data_o[24];
  assign data_o[15192] = data_o[24];
  assign data_o[15256] = data_o[24];
  assign data_o[15320] = data_o[24];
  assign data_o[15384] = data_o[24];
  assign data_o[15448] = data_o[24];
  assign data_o[15512] = data_o[24];
  assign data_o[15576] = data_o[24];
  assign data_o[15640] = data_o[24];
  assign data_o[15704] = data_o[24];
  assign data_o[15768] = data_o[24];
  assign data_o[15832] = data_o[24];
  assign data_o[15896] = data_o[24];
  assign data_o[15960] = data_o[24];
  assign data_o[16024] = data_o[24];
  assign data_o[16088] = data_o[24];
  assign data_o[16152] = data_o[24];
  assign data_o[16216] = data_o[24];
  assign data_o[16280] = data_o[24];
  assign data_o[16344] = data_o[24];
  assign data_o[16408] = data_o[24];
  assign data_o[16472] = data_o[24];
  assign data_o[16536] = data_o[24];
  assign data_o[16600] = data_o[24];
  assign data_o[16664] = data_o[24];
  assign data_o[16728] = data_o[24];
  assign data_o[16792] = data_o[24];
  assign data_o[16856] = data_o[24];
  assign data_o[16920] = data_o[24];
  assign data_o[16984] = data_o[24];
  assign data_o[17048] = data_o[24];
  assign data_o[17112] = data_o[24];
  assign data_o[17176] = data_o[24];
  assign data_o[17240] = data_o[24];
  assign data_o[17304] = data_o[24];
  assign data_o[17368] = data_o[24];
  assign data_o[17432] = data_o[24];
  assign data_o[17496] = data_o[24];
  assign data_o[17560] = data_o[24];
  assign data_o[17624] = data_o[24];
  assign data_o[17688] = data_o[24];
  assign data_o[17752] = data_o[24];
  assign data_o[17816] = data_o[24];
  assign data_o[17880] = data_o[24];
  assign data_o[17944] = data_o[24];
  assign data_o[18008] = data_o[24];
  assign data_o[18072] = data_o[24];
  assign data_o[18136] = data_o[24];
  assign data_o[18200] = data_o[24];
  assign data_o[18264] = data_o[24];
  assign data_o[18328] = data_o[24];
  assign data_o[18392] = data_o[24];
  assign data_o[18456] = data_o[24];
  assign data_o[18520] = data_o[24];
  assign data_o[18584] = data_o[24];
  assign data_o[18648] = data_o[24];
  assign data_o[18712] = data_o[24];
  assign data_o[18776] = data_o[24];
  assign data_o[18840] = data_o[24];
  assign data_o[18904] = data_o[24];
  assign data_o[18968] = data_o[24];
  assign data_o[19032] = data_o[24];
  assign data_o[19096] = data_o[24];
  assign data_o[19160] = data_o[24];
  assign data_o[19224] = data_o[24];
  assign data_o[19288] = data_o[24];
  assign data_o[19352] = data_o[24];
  assign data_o[19416] = data_o[24];
  assign data_o[19480] = data_o[24];
  assign data_o[19544] = data_o[24];
  assign data_o[19608] = data_o[24];
  assign data_o[19672] = data_o[24];
  assign data_o[19736] = data_o[24];
  assign data_o[19800] = data_o[24];
  assign data_o[19864] = data_o[24];
  assign data_o[19928] = data_o[24];
  assign data_o[19992] = data_o[24];
  assign data_o[20056] = data_o[24];
  assign data_o[20120] = data_o[24];
  assign data_o[20184] = data_o[24];
  assign data_o[20248] = data_o[24];
  assign data_o[20312] = data_o[24];
  assign data_o[20376] = data_o[24];
  assign data_o[20440] = data_o[24];
  assign data_o[20504] = data_o[24];
  assign data_o[20568] = data_o[24];
  assign data_o[20632] = data_o[24];
  assign data_o[20696] = data_o[24];
  assign data_o[20760] = data_o[24];
  assign data_o[20824] = data_o[24];
  assign data_o[20888] = data_o[24];
  assign data_o[20952] = data_o[24];
  assign data_o[21016] = data_o[24];
  assign data_o[21080] = data_o[24];
  assign data_o[21144] = data_o[24];
  assign data_o[21208] = data_o[24];
  assign data_o[21272] = data_o[24];
  assign data_o[21336] = data_o[24];
  assign data_o[21400] = data_o[24];
  assign data_o[21464] = data_o[24];
  assign data_o[21528] = data_o[24];
  assign data_o[21592] = data_o[24];
  assign data_o[21656] = data_o[24];
  assign data_o[21720] = data_o[24];
  assign data_o[21784] = data_o[24];
  assign data_o[21848] = data_o[24];
  assign data_o[21912] = data_o[24];
  assign data_o[21976] = data_o[24];
  assign data_o[22040] = data_o[24];
  assign data_o[22104] = data_o[24];
  assign data_o[22168] = data_o[24];
  assign data_o[22232] = data_o[24];
  assign data_o[22296] = data_o[24];
  assign data_o[22360] = data_o[24];
  assign data_o[22424] = data_o[24];
  assign data_o[22488] = data_o[24];
  assign data_o[22552] = data_o[24];
  assign data_o[22616] = data_o[24];
  assign data_o[22680] = data_o[24];
  assign data_o[22744] = data_o[24];
  assign data_o[22808] = data_o[24];
  assign data_o[22872] = data_o[24];
  assign data_o[22936] = data_o[24];
  assign data_o[23000] = data_o[24];
  assign data_o[23064] = data_o[24];
  assign data_o[23128] = data_o[24];
  assign data_o[23192] = data_o[24];
  assign data_o[23256] = data_o[24];
  assign data_o[23320] = data_o[24];
  assign data_o[23384] = data_o[24];
  assign data_o[23448] = data_o[24];
  assign data_o[23512] = data_o[24];
  assign data_o[23576] = data_o[24];
  assign data_o[23640] = data_o[24];
  assign data_o[23704] = data_o[24];
  assign data_o[23768] = data_o[24];
  assign data_o[23832] = data_o[24];
  assign data_o[23896] = data_o[24];
  assign data_o[23960] = data_o[24];
  assign data_o[24024] = data_o[24];
  assign data_o[24088] = data_o[24];
  assign data_o[24152] = data_o[24];
  assign data_o[24216] = data_o[24];
  assign data_o[24280] = data_o[24];
  assign data_o[24344] = data_o[24];
  assign data_o[24408] = data_o[24];
  assign data_o[24472] = data_o[24];
  assign data_o[24536] = data_o[24];
  assign data_o[24600] = data_o[24];
  assign data_o[24664] = data_o[24];
  assign data_o[24728] = data_o[24];
  assign data_o[24792] = data_o[24];
  assign data_o[24856] = data_o[24];
  assign data_o[24920] = data_o[24];
  assign data_o[24984] = data_o[24];
  assign data_o[25048] = data_o[24];
  assign data_o[25112] = data_o[24];
  assign data_o[25176] = data_o[24];
  assign data_o[25240] = data_o[24];
  assign data_o[25304] = data_o[24];
  assign data_o[25368] = data_o[24];
  assign data_o[25432] = data_o[24];
  assign data_o[25496] = data_o[24];
  assign data_o[25560] = data_o[24];
  assign data_o[25624] = data_o[24];
  assign data_o[25688] = data_o[24];
  assign data_o[25752] = data_o[24];
  assign data_o[25816] = data_o[24];
  assign data_o[25880] = data_o[24];
  assign data_o[25944] = data_o[24];
  assign data_o[26008] = data_o[24];
  assign data_o[26072] = data_o[24];
  assign data_o[26136] = data_o[24];
  assign data_o[26200] = data_o[24];
  assign data_o[26264] = data_o[24];
  assign data_o[26328] = data_o[24];
  assign data_o[26392] = data_o[24];
  assign data_o[26456] = data_o[24];
  assign data_o[26520] = data_o[24];
  assign data_o[26584] = data_o[24];
  assign data_o[26648] = data_o[24];
  assign data_o[26712] = data_o[24];
  assign data_o[26776] = data_o[24];
  assign data_o[26840] = data_o[24];
  assign data_o[26904] = data_o[24];
  assign data_o[26968] = data_o[24];
  assign data_o[27032] = data_o[24];
  assign data_o[27096] = data_o[24];
  assign data_o[27160] = data_o[24];
  assign data_o[27224] = data_o[24];
  assign data_o[27288] = data_o[24];
  assign data_o[27352] = data_o[24];
  assign data_o[27416] = data_o[24];
  assign data_o[27480] = data_o[24];
  assign data_o[27544] = data_o[24];
  assign data_o[27608] = data_o[24];
  assign data_o[27672] = data_o[24];
  assign data_o[27736] = data_o[24];
  assign data_o[27800] = data_o[24];
  assign data_o[27864] = data_o[24];
  assign data_o[27928] = data_o[24];
  assign data_o[27992] = data_o[24];
  assign data_o[28056] = data_o[24];
  assign data_o[28120] = data_o[24];
  assign data_o[28184] = data_o[24];
  assign data_o[28248] = data_o[24];
  assign data_o[28312] = data_o[24];
  assign data_o[28376] = data_o[24];
  assign data_o[28440] = data_o[24];
  assign data_o[28504] = data_o[24];
  assign data_o[28568] = data_o[24];
  assign data_o[28632] = data_o[24];
  assign data_o[28696] = data_o[24];
  assign data_o[28760] = data_o[24];
  assign data_o[28824] = data_o[24];
  assign data_o[28888] = data_o[24];
  assign data_o[28952] = data_o[24];
  assign data_o[29016] = data_o[24];
  assign data_o[29080] = data_o[24];
  assign data_o[29144] = data_o[24];
  assign data_o[29208] = data_o[24];
  assign data_o[29272] = data_o[24];
  assign data_o[29336] = data_o[24];
  assign data_o[29400] = data_o[24];
  assign data_o[29464] = data_o[24];
  assign data_o[29528] = data_o[24];
  assign data_o[29592] = data_o[24];
  assign data_o[29656] = data_o[24];
  assign data_o[29720] = data_o[24];
  assign data_o[29784] = data_o[24];
  assign data_o[29848] = data_o[24];
  assign data_o[29912] = data_o[24];
  assign data_o[29976] = data_o[24];
  assign data_o[30040] = data_o[24];
  assign data_o[30104] = data_o[24];
  assign data_o[30168] = data_o[24];
  assign data_o[30232] = data_o[24];
  assign data_o[30296] = data_o[24];
  assign data_o[30360] = data_o[24];
  assign data_o[30424] = data_o[24];
  assign data_o[30488] = data_o[24];
  assign data_o[30552] = data_o[24];
  assign data_o[30616] = data_o[24];
  assign data_o[30680] = data_o[24];
  assign data_o[30744] = data_o[24];
  assign data_o[30808] = data_o[24];
  assign data_o[30872] = data_o[24];
  assign data_o[30936] = data_o[24];
  assign data_o[31000] = data_o[24];
  assign data_o[31064] = data_o[24];
  assign data_o[31128] = data_o[24];
  assign data_o[31192] = data_o[24];
  assign data_o[31256] = data_o[24];
  assign data_o[31320] = data_o[24];
  assign data_o[31384] = data_o[24];
  assign data_o[31448] = data_o[24];
  assign data_o[31512] = data_o[24];
  assign data_o[31576] = data_o[24];
  assign data_o[31640] = data_o[24];
  assign data_o[31704] = data_o[24];
  assign data_o[31768] = data_o[24];
  assign data_o[31832] = data_o[24];
  assign data_o[31896] = data_o[24];
  assign data_o[31960] = data_o[24];
  assign data_o[87] = data_o[23];
  assign data_o[151] = data_o[23];
  assign data_o[215] = data_o[23];
  assign data_o[279] = data_o[23];
  assign data_o[343] = data_o[23];
  assign data_o[407] = data_o[23];
  assign data_o[471] = data_o[23];
  assign data_o[535] = data_o[23];
  assign data_o[599] = data_o[23];
  assign data_o[663] = data_o[23];
  assign data_o[727] = data_o[23];
  assign data_o[791] = data_o[23];
  assign data_o[855] = data_o[23];
  assign data_o[919] = data_o[23];
  assign data_o[983] = data_o[23];
  assign data_o[1047] = data_o[23];
  assign data_o[1111] = data_o[23];
  assign data_o[1175] = data_o[23];
  assign data_o[1239] = data_o[23];
  assign data_o[1303] = data_o[23];
  assign data_o[1367] = data_o[23];
  assign data_o[1431] = data_o[23];
  assign data_o[1495] = data_o[23];
  assign data_o[1559] = data_o[23];
  assign data_o[1623] = data_o[23];
  assign data_o[1687] = data_o[23];
  assign data_o[1751] = data_o[23];
  assign data_o[1815] = data_o[23];
  assign data_o[1879] = data_o[23];
  assign data_o[1943] = data_o[23];
  assign data_o[2007] = data_o[23];
  assign data_o[2071] = data_o[23];
  assign data_o[2135] = data_o[23];
  assign data_o[2199] = data_o[23];
  assign data_o[2263] = data_o[23];
  assign data_o[2327] = data_o[23];
  assign data_o[2391] = data_o[23];
  assign data_o[2455] = data_o[23];
  assign data_o[2519] = data_o[23];
  assign data_o[2583] = data_o[23];
  assign data_o[2647] = data_o[23];
  assign data_o[2711] = data_o[23];
  assign data_o[2775] = data_o[23];
  assign data_o[2839] = data_o[23];
  assign data_o[2903] = data_o[23];
  assign data_o[2967] = data_o[23];
  assign data_o[3031] = data_o[23];
  assign data_o[3095] = data_o[23];
  assign data_o[3159] = data_o[23];
  assign data_o[3223] = data_o[23];
  assign data_o[3287] = data_o[23];
  assign data_o[3351] = data_o[23];
  assign data_o[3415] = data_o[23];
  assign data_o[3479] = data_o[23];
  assign data_o[3543] = data_o[23];
  assign data_o[3607] = data_o[23];
  assign data_o[3671] = data_o[23];
  assign data_o[3735] = data_o[23];
  assign data_o[3799] = data_o[23];
  assign data_o[3863] = data_o[23];
  assign data_o[3927] = data_o[23];
  assign data_o[3991] = data_o[23];
  assign data_o[4055] = data_o[23];
  assign data_o[4119] = data_o[23];
  assign data_o[4183] = data_o[23];
  assign data_o[4247] = data_o[23];
  assign data_o[4311] = data_o[23];
  assign data_o[4375] = data_o[23];
  assign data_o[4439] = data_o[23];
  assign data_o[4503] = data_o[23];
  assign data_o[4567] = data_o[23];
  assign data_o[4631] = data_o[23];
  assign data_o[4695] = data_o[23];
  assign data_o[4759] = data_o[23];
  assign data_o[4823] = data_o[23];
  assign data_o[4887] = data_o[23];
  assign data_o[4951] = data_o[23];
  assign data_o[5015] = data_o[23];
  assign data_o[5079] = data_o[23];
  assign data_o[5143] = data_o[23];
  assign data_o[5207] = data_o[23];
  assign data_o[5271] = data_o[23];
  assign data_o[5335] = data_o[23];
  assign data_o[5399] = data_o[23];
  assign data_o[5463] = data_o[23];
  assign data_o[5527] = data_o[23];
  assign data_o[5591] = data_o[23];
  assign data_o[5655] = data_o[23];
  assign data_o[5719] = data_o[23];
  assign data_o[5783] = data_o[23];
  assign data_o[5847] = data_o[23];
  assign data_o[5911] = data_o[23];
  assign data_o[5975] = data_o[23];
  assign data_o[6039] = data_o[23];
  assign data_o[6103] = data_o[23];
  assign data_o[6167] = data_o[23];
  assign data_o[6231] = data_o[23];
  assign data_o[6295] = data_o[23];
  assign data_o[6359] = data_o[23];
  assign data_o[6423] = data_o[23];
  assign data_o[6487] = data_o[23];
  assign data_o[6551] = data_o[23];
  assign data_o[6615] = data_o[23];
  assign data_o[6679] = data_o[23];
  assign data_o[6743] = data_o[23];
  assign data_o[6807] = data_o[23];
  assign data_o[6871] = data_o[23];
  assign data_o[6935] = data_o[23];
  assign data_o[6999] = data_o[23];
  assign data_o[7063] = data_o[23];
  assign data_o[7127] = data_o[23];
  assign data_o[7191] = data_o[23];
  assign data_o[7255] = data_o[23];
  assign data_o[7319] = data_o[23];
  assign data_o[7383] = data_o[23];
  assign data_o[7447] = data_o[23];
  assign data_o[7511] = data_o[23];
  assign data_o[7575] = data_o[23];
  assign data_o[7639] = data_o[23];
  assign data_o[7703] = data_o[23];
  assign data_o[7767] = data_o[23];
  assign data_o[7831] = data_o[23];
  assign data_o[7895] = data_o[23];
  assign data_o[7959] = data_o[23];
  assign data_o[8023] = data_o[23];
  assign data_o[8087] = data_o[23];
  assign data_o[8151] = data_o[23];
  assign data_o[8215] = data_o[23];
  assign data_o[8279] = data_o[23];
  assign data_o[8343] = data_o[23];
  assign data_o[8407] = data_o[23];
  assign data_o[8471] = data_o[23];
  assign data_o[8535] = data_o[23];
  assign data_o[8599] = data_o[23];
  assign data_o[8663] = data_o[23];
  assign data_o[8727] = data_o[23];
  assign data_o[8791] = data_o[23];
  assign data_o[8855] = data_o[23];
  assign data_o[8919] = data_o[23];
  assign data_o[8983] = data_o[23];
  assign data_o[9047] = data_o[23];
  assign data_o[9111] = data_o[23];
  assign data_o[9175] = data_o[23];
  assign data_o[9239] = data_o[23];
  assign data_o[9303] = data_o[23];
  assign data_o[9367] = data_o[23];
  assign data_o[9431] = data_o[23];
  assign data_o[9495] = data_o[23];
  assign data_o[9559] = data_o[23];
  assign data_o[9623] = data_o[23];
  assign data_o[9687] = data_o[23];
  assign data_o[9751] = data_o[23];
  assign data_o[9815] = data_o[23];
  assign data_o[9879] = data_o[23];
  assign data_o[9943] = data_o[23];
  assign data_o[10007] = data_o[23];
  assign data_o[10071] = data_o[23];
  assign data_o[10135] = data_o[23];
  assign data_o[10199] = data_o[23];
  assign data_o[10263] = data_o[23];
  assign data_o[10327] = data_o[23];
  assign data_o[10391] = data_o[23];
  assign data_o[10455] = data_o[23];
  assign data_o[10519] = data_o[23];
  assign data_o[10583] = data_o[23];
  assign data_o[10647] = data_o[23];
  assign data_o[10711] = data_o[23];
  assign data_o[10775] = data_o[23];
  assign data_o[10839] = data_o[23];
  assign data_o[10903] = data_o[23];
  assign data_o[10967] = data_o[23];
  assign data_o[11031] = data_o[23];
  assign data_o[11095] = data_o[23];
  assign data_o[11159] = data_o[23];
  assign data_o[11223] = data_o[23];
  assign data_o[11287] = data_o[23];
  assign data_o[11351] = data_o[23];
  assign data_o[11415] = data_o[23];
  assign data_o[11479] = data_o[23];
  assign data_o[11543] = data_o[23];
  assign data_o[11607] = data_o[23];
  assign data_o[11671] = data_o[23];
  assign data_o[11735] = data_o[23];
  assign data_o[11799] = data_o[23];
  assign data_o[11863] = data_o[23];
  assign data_o[11927] = data_o[23];
  assign data_o[11991] = data_o[23];
  assign data_o[12055] = data_o[23];
  assign data_o[12119] = data_o[23];
  assign data_o[12183] = data_o[23];
  assign data_o[12247] = data_o[23];
  assign data_o[12311] = data_o[23];
  assign data_o[12375] = data_o[23];
  assign data_o[12439] = data_o[23];
  assign data_o[12503] = data_o[23];
  assign data_o[12567] = data_o[23];
  assign data_o[12631] = data_o[23];
  assign data_o[12695] = data_o[23];
  assign data_o[12759] = data_o[23];
  assign data_o[12823] = data_o[23];
  assign data_o[12887] = data_o[23];
  assign data_o[12951] = data_o[23];
  assign data_o[13015] = data_o[23];
  assign data_o[13079] = data_o[23];
  assign data_o[13143] = data_o[23];
  assign data_o[13207] = data_o[23];
  assign data_o[13271] = data_o[23];
  assign data_o[13335] = data_o[23];
  assign data_o[13399] = data_o[23];
  assign data_o[13463] = data_o[23];
  assign data_o[13527] = data_o[23];
  assign data_o[13591] = data_o[23];
  assign data_o[13655] = data_o[23];
  assign data_o[13719] = data_o[23];
  assign data_o[13783] = data_o[23];
  assign data_o[13847] = data_o[23];
  assign data_o[13911] = data_o[23];
  assign data_o[13975] = data_o[23];
  assign data_o[14039] = data_o[23];
  assign data_o[14103] = data_o[23];
  assign data_o[14167] = data_o[23];
  assign data_o[14231] = data_o[23];
  assign data_o[14295] = data_o[23];
  assign data_o[14359] = data_o[23];
  assign data_o[14423] = data_o[23];
  assign data_o[14487] = data_o[23];
  assign data_o[14551] = data_o[23];
  assign data_o[14615] = data_o[23];
  assign data_o[14679] = data_o[23];
  assign data_o[14743] = data_o[23];
  assign data_o[14807] = data_o[23];
  assign data_o[14871] = data_o[23];
  assign data_o[14935] = data_o[23];
  assign data_o[14999] = data_o[23];
  assign data_o[15063] = data_o[23];
  assign data_o[15127] = data_o[23];
  assign data_o[15191] = data_o[23];
  assign data_o[15255] = data_o[23];
  assign data_o[15319] = data_o[23];
  assign data_o[15383] = data_o[23];
  assign data_o[15447] = data_o[23];
  assign data_o[15511] = data_o[23];
  assign data_o[15575] = data_o[23];
  assign data_o[15639] = data_o[23];
  assign data_o[15703] = data_o[23];
  assign data_o[15767] = data_o[23];
  assign data_o[15831] = data_o[23];
  assign data_o[15895] = data_o[23];
  assign data_o[15959] = data_o[23];
  assign data_o[16023] = data_o[23];
  assign data_o[16087] = data_o[23];
  assign data_o[16151] = data_o[23];
  assign data_o[16215] = data_o[23];
  assign data_o[16279] = data_o[23];
  assign data_o[16343] = data_o[23];
  assign data_o[16407] = data_o[23];
  assign data_o[16471] = data_o[23];
  assign data_o[16535] = data_o[23];
  assign data_o[16599] = data_o[23];
  assign data_o[16663] = data_o[23];
  assign data_o[16727] = data_o[23];
  assign data_o[16791] = data_o[23];
  assign data_o[16855] = data_o[23];
  assign data_o[16919] = data_o[23];
  assign data_o[16983] = data_o[23];
  assign data_o[17047] = data_o[23];
  assign data_o[17111] = data_o[23];
  assign data_o[17175] = data_o[23];
  assign data_o[17239] = data_o[23];
  assign data_o[17303] = data_o[23];
  assign data_o[17367] = data_o[23];
  assign data_o[17431] = data_o[23];
  assign data_o[17495] = data_o[23];
  assign data_o[17559] = data_o[23];
  assign data_o[17623] = data_o[23];
  assign data_o[17687] = data_o[23];
  assign data_o[17751] = data_o[23];
  assign data_o[17815] = data_o[23];
  assign data_o[17879] = data_o[23];
  assign data_o[17943] = data_o[23];
  assign data_o[18007] = data_o[23];
  assign data_o[18071] = data_o[23];
  assign data_o[18135] = data_o[23];
  assign data_o[18199] = data_o[23];
  assign data_o[18263] = data_o[23];
  assign data_o[18327] = data_o[23];
  assign data_o[18391] = data_o[23];
  assign data_o[18455] = data_o[23];
  assign data_o[18519] = data_o[23];
  assign data_o[18583] = data_o[23];
  assign data_o[18647] = data_o[23];
  assign data_o[18711] = data_o[23];
  assign data_o[18775] = data_o[23];
  assign data_o[18839] = data_o[23];
  assign data_o[18903] = data_o[23];
  assign data_o[18967] = data_o[23];
  assign data_o[19031] = data_o[23];
  assign data_o[19095] = data_o[23];
  assign data_o[19159] = data_o[23];
  assign data_o[19223] = data_o[23];
  assign data_o[19287] = data_o[23];
  assign data_o[19351] = data_o[23];
  assign data_o[19415] = data_o[23];
  assign data_o[19479] = data_o[23];
  assign data_o[19543] = data_o[23];
  assign data_o[19607] = data_o[23];
  assign data_o[19671] = data_o[23];
  assign data_o[19735] = data_o[23];
  assign data_o[19799] = data_o[23];
  assign data_o[19863] = data_o[23];
  assign data_o[19927] = data_o[23];
  assign data_o[19991] = data_o[23];
  assign data_o[20055] = data_o[23];
  assign data_o[20119] = data_o[23];
  assign data_o[20183] = data_o[23];
  assign data_o[20247] = data_o[23];
  assign data_o[20311] = data_o[23];
  assign data_o[20375] = data_o[23];
  assign data_o[20439] = data_o[23];
  assign data_o[20503] = data_o[23];
  assign data_o[20567] = data_o[23];
  assign data_o[20631] = data_o[23];
  assign data_o[20695] = data_o[23];
  assign data_o[20759] = data_o[23];
  assign data_o[20823] = data_o[23];
  assign data_o[20887] = data_o[23];
  assign data_o[20951] = data_o[23];
  assign data_o[21015] = data_o[23];
  assign data_o[21079] = data_o[23];
  assign data_o[21143] = data_o[23];
  assign data_o[21207] = data_o[23];
  assign data_o[21271] = data_o[23];
  assign data_o[21335] = data_o[23];
  assign data_o[21399] = data_o[23];
  assign data_o[21463] = data_o[23];
  assign data_o[21527] = data_o[23];
  assign data_o[21591] = data_o[23];
  assign data_o[21655] = data_o[23];
  assign data_o[21719] = data_o[23];
  assign data_o[21783] = data_o[23];
  assign data_o[21847] = data_o[23];
  assign data_o[21911] = data_o[23];
  assign data_o[21975] = data_o[23];
  assign data_o[22039] = data_o[23];
  assign data_o[22103] = data_o[23];
  assign data_o[22167] = data_o[23];
  assign data_o[22231] = data_o[23];
  assign data_o[22295] = data_o[23];
  assign data_o[22359] = data_o[23];
  assign data_o[22423] = data_o[23];
  assign data_o[22487] = data_o[23];
  assign data_o[22551] = data_o[23];
  assign data_o[22615] = data_o[23];
  assign data_o[22679] = data_o[23];
  assign data_o[22743] = data_o[23];
  assign data_o[22807] = data_o[23];
  assign data_o[22871] = data_o[23];
  assign data_o[22935] = data_o[23];
  assign data_o[22999] = data_o[23];
  assign data_o[23063] = data_o[23];
  assign data_o[23127] = data_o[23];
  assign data_o[23191] = data_o[23];
  assign data_o[23255] = data_o[23];
  assign data_o[23319] = data_o[23];
  assign data_o[23383] = data_o[23];
  assign data_o[23447] = data_o[23];
  assign data_o[23511] = data_o[23];
  assign data_o[23575] = data_o[23];
  assign data_o[23639] = data_o[23];
  assign data_o[23703] = data_o[23];
  assign data_o[23767] = data_o[23];
  assign data_o[23831] = data_o[23];
  assign data_o[23895] = data_o[23];
  assign data_o[23959] = data_o[23];
  assign data_o[24023] = data_o[23];
  assign data_o[24087] = data_o[23];
  assign data_o[24151] = data_o[23];
  assign data_o[24215] = data_o[23];
  assign data_o[24279] = data_o[23];
  assign data_o[24343] = data_o[23];
  assign data_o[24407] = data_o[23];
  assign data_o[24471] = data_o[23];
  assign data_o[24535] = data_o[23];
  assign data_o[24599] = data_o[23];
  assign data_o[24663] = data_o[23];
  assign data_o[24727] = data_o[23];
  assign data_o[24791] = data_o[23];
  assign data_o[24855] = data_o[23];
  assign data_o[24919] = data_o[23];
  assign data_o[24983] = data_o[23];
  assign data_o[25047] = data_o[23];
  assign data_o[25111] = data_o[23];
  assign data_o[25175] = data_o[23];
  assign data_o[25239] = data_o[23];
  assign data_o[25303] = data_o[23];
  assign data_o[25367] = data_o[23];
  assign data_o[25431] = data_o[23];
  assign data_o[25495] = data_o[23];
  assign data_o[25559] = data_o[23];
  assign data_o[25623] = data_o[23];
  assign data_o[25687] = data_o[23];
  assign data_o[25751] = data_o[23];
  assign data_o[25815] = data_o[23];
  assign data_o[25879] = data_o[23];
  assign data_o[25943] = data_o[23];
  assign data_o[26007] = data_o[23];
  assign data_o[26071] = data_o[23];
  assign data_o[26135] = data_o[23];
  assign data_o[26199] = data_o[23];
  assign data_o[26263] = data_o[23];
  assign data_o[26327] = data_o[23];
  assign data_o[26391] = data_o[23];
  assign data_o[26455] = data_o[23];
  assign data_o[26519] = data_o[23];
  assign data_o[26583] = data_o[23];
  assign data_o[26647] = data_o[23];
  assign data_o[26711] = data_o[23];
  assign data_o[26775] = data_o[23];
  assign data_o[26839] = data_o[23];
  assign data_o[26903] = data_o[23];
  assign data_o[26967] = data_o[23];
  assign data_o[27031] = data_o[23];
  assign data_o[27095] = data_o[23];
  assign data_o[27159] = data_o[23];
  assign data_o[27223] = data_o[23];
  assign data_o[27287] = data_o[23];
  assign data_o[27351] = data_o[23];
  assign data_o[27415] = data_o[23];
  assign data_o[27479] = data_o[23];
  assign data_o[27543] = data_o[23];
  assign data_o[27607] = data_o[23];
  assign data_o[27671] = data_o[23];
  assign data_o[27735] = data_o[23];
  assign data_o[27799] = data_o[23];
  assign data_o[27863] = data_o[23];
  assign data_o[27927] = data_o[23];
  assign data_o[27991] = data_o[23];
  assign data_o[28055] = data_o[23];
  assign data_o[28119] = data_o[23];
  assign data_o[28183] = data_o[23];
  assign data_o[28247] = data_o[23];
  assign data_o[28311] = data_o[23];
  assign data_o[28375] = data_o[23];
  assign data_o[28439] = data_o[23];
  assign data_o[28503] = data_o[23];
  assign data_o[28567] = data_o[23];
  assign data_o[28631] = data_o[23];
  assign data_o[28695] = data_o[23];
  assign data_o[28759] = data_o[23];
  assign data_o[28823] = data_o[23];
  assign data_o[28887] = data_o[23];
  assign data_o[28951] = data_o[23];
  assign data_o[29015] = data_o[23];
  assign data_o[29079] = data_o[23];
  assign data_o[29143] = data_o[23];
  assign data_o[29207] = data_o[23];
  assign data_o[29271] = data_o[23];
  assign data_o[29335] = data_o[23];
  assign data_o[29399] = data_o[23];
  assign data_o[29463] = data_o[23];
  assign data_o[29527] = data_o[23];
  assign data_o[29591] = data_o[23];
  assign data_o[29655] = data_o[23];
  assign data_o[29719] = data_o[23];
  assign data_o[29783] = data_o[23];
  assign data_o[29847] = data_o[23];
  assign data_o[29911] = data_o[23];
  assign data_o[29975] = data_o[23];
  assign data_o[30039] = data_o[23];
  assign data_o[30103] = data_o[23];
  assign data_o[30167] = data_o[23];
  assign data_o[30231] = data_o[23];
  assign data_o[30295] = data_o[23];
  assign data_o[30359] = data_o[23];
  assign data_o[30423] = data_o[23];
  assign data_o[30487] = data_o[23];
  assign data_o[30551] = data_o[23];
  assign data_o[30615] = data_o[23];
  assign data_o[30679] = data_o[23];
  assign data_o[30743] = data_o[23];
  assign data_o[30807] = data_o[23];
  assign data_o[30871] = data_o[23];
  assign data_o[30935] = data_o[23];
  assign data_o[30999] = data_o[23];
  assign data_o[31063] = data_o[23];
  assign data_o[31127] = data_o[23];
  assign data_o[31191] = data_o[23];
  assign data_o[31255] = data_o[23];
  assign data_o[31319] = data_o[23];
  assign data_o[31383] = data_o[23];
  assign data_o[31447] = data_o[23];
  assign data_o[31511] = data_o[23];
  assign data_o[31575] = data_o[23];
  assign data_o[31639] = data_o[23];
  assign data_o[31703] = data_o[23];
  assign data_o[31767] = data_o[23];
  assign data_o[31831] = data_o[23];
  assign data_o[31895] = data_o[23];
  assign data_o[31959] = data_o[23];
  assign data_o[86] = data_o[22];
  assign data_o[150] = data_o[22];
  assign data_o[214] = data_o[22];
  assign data_o[278] = data_o[22];
  assign data_o[342] = data_o[22];
  assign data_o[406] = data_o[22];
  assign data_o[470] = data_o[22];
  assign data_o[534] = data_o[22];
  assign data_o[598] = data_o[22];
  assign data_o[662] = data_o[22];
  assign data_o[726] = data_o[22];
  assign data_o[790] = data_o[22];
  assign data_o[854] = data_o[22];
  assign data_o[918] = data_o[22];
  assign data_o[982] = data_o[22];
  assign data_o[1046] = data_o[22];
  assign data_o[1110] = data_o[22];
  assign data_o[1174] = data_o[22];
  assign data_o[1238] = data_o[22];
  assign data_o[1302] = data_o[22];
  assign data_o[1366] = data_o[22];
  assign data_o[1430] = data_o[22];
  assign data_o[1494] = data_o[22];
  assign data_o[1558] = data_o[22];
  assign data_o[1622] = data_o[22];
  assign data_o[1686] = data_o[22];
  assign data_o[1750] = data_o[22];
  assign data_o[1814] = data_o[22];
  assign data_o[1878] = data_o[22];
  assign data_o[1942] = data_o[22];
  assign data_o[2006] = data_o[22];
  assign data_o[2070] = data_o[22];
  assign data_o[2134] = data_o[22];
  assign data_o[2198] = data_o[22];
  assign data_o[2262] = data_o[22];
  assign data_o[2326] = data_o[22];
  assign data_o[2390] = data_o[22];
  assign data_o[2454] = data_o[22];
  assign data_o[2518] = data_o[22];
  assign data_o[2582] = data_o[22];
  assign data_o[2646] = data_o[22];
  assign data_o[2710] = data_o[22];
  assign data_o[2774] = data_o[22];
  assign data_o[2838] = data_o[22];
  assign data_o[2902] = data_o[22];
  assign data_o[2966] = data_o[22];
  assign data_o[3030] = data_o[22];
  assign data_o[3094] = data_o[22];
  assign data_o[3158] = data_o[22];
  assign data_o[3222] = data_o[22];
  assign data_o[3286] = data_o[22];
  assign data_o[3350] = data_o[22];
  assign data_o[3414] = data_o[22];
  assign data_o[3478] = data_o[22];
  assign data_o[3542] = data_o[22];
  assign data_o[3606] = data_o[22];
  assign data_o[3670] = data_o[22];
  assign data_o[3734] = data_o[22];
  assign data_o[3798] = data_o[22];
  assign data_o[3862] = data_o[22];
  assign data_o[3926] = data_o[22];
  assign data_o[3990] = data_o[22];
  assign data_o[4054] = data_o[22];
  assign data_o[4118] = data_o[22];
  assign data_o[4182] = data_o[22];
  assign data_o[4246] = data_o[22];
  assign data_o[4310] = data_o[22];
  assign data_o[4374] = data_o[22];
  assign data_o[4438] = data_o[22];
  assign data_o[4502] = data_o[22];
  assign data_o[4566] = data_o[22];
  assign data_o[4630] = data_o[22];
  assign data_o[4694] = data_o[22];
  assign data_o[4758] = data_o[22];
  assign data_o[4822] = data_o[22];
  assign data_o[4886] = data_o[22];
  assign data_o[4950] = data_o[22];
  assign data_o[5014] = data_o[22];
  assign data_o[5078] = data_o[22];
  assign data_o[5142] = data_o[22];
  assign data_o[5206] = data_o[22];
  assign data_o[5270] = data_o[22];
  assign data_o[5334] = data_o[22];
  assign data_o[5398] = data_o[22];
  assign data_o[5462] = data_o[22];
  assign data_o[5526] = data_o[22];
  assign data_o[5590] = data_o[22];
  assign data_o[5654] = data_o[22];
  assign data_o[5718] = data_o[22];
  assign data_o[5782] = data_o[22];
  assign data_o[5846] = data_o[22];
  assign data_o[5910] = data_o[22];
  assign data_o[5974] = data_o[22];
  assign data_o[6038] = data_o[22];
  assign data_o[6102] = data_o[22];
  assign data_o[6166] = data_o[22];
  assign data_o[6230] = data_o[22];
  assign data_o[6294] = data_o[22];
  assign data_o[6358] = data_o[22];
  assign data_o[6422] = data_o[22];
  assign data_o[6486] = data_o[22];
  assign data_o[6550] = data_o[22];
  assign data_o[6614] = data_o[22];
  assign data_o[6678] = data_o[22];
  assign data_o[6742] = data_o[22];
  assign data_o[6806] = data_o[22];
  assign data_o[6870] = data_o[22];
  assign data_o[6934] = data_o[22];
  assign data_o[6998] = data_o[22];
  assign data_o[7062] = data_o[22];
  assign data_o[7126] = data_o[22];
  assign data_o[7190] = data_o[22];
  assign data_o[7254] = data_o[22];
  assign data_o[7318] = data_o[22];
  assign data_o[7382] = data_o[22];
  assign data_o[7446] = data_o[22];
  assign data_o[7510] = data_o[22];
  assign data_o[7574] = data_o[22];
  assign data_o[7638] = data_o[22];
  assign data_o[7702] = data_o[22];
  assign data_o[7766] = data_o[22];
  assign data_o[7830] = data_o[22];
  assign data_o[7894] = data_o[22];
  assign data_o[7958] = data_o[22];
  assign data_o[8022] = data_o[22];
  assign data_o[8086] = data_o[22];
  assign data_o[8150] = data_o[22];
  assign data_o[8214] = data_o[22];
  assign data_o[8278] = data_o[22];
  assign data_o[8342] = data_o[22];
  assign data_o[8406] = data_o[22];
  assign data_o[8470] = data_o[22];
  assign data_o[8534] = data_o[22];
  assign data_o[8598] = data_o[22];
  assign data_o[8662] = data_o[22];
  assign data_o[8726] = data_o[22];
  assign data_o[8790] = data_o[22];
  assign data_o[8854] = data_o[22];
  assign data_o[8918] = data_o[22];
  assign data_o[8982] = data_o[22];
  assign data_o[9046] = data_o[22];
  assign data_o[9110] = data_o[22];
  assign data_o[9174] = data_o[22];
  assign data_o[9238] = data_o[22];
  assign data_o[9302] = data_o[22];
  assign data_o[9366] = data_o[22];
  assign data_o[9430] = data_o[22];
  assign data_o[9494] = data_o[22];
  assign data_o[9558] = data_o[22];
  assign data_o[9622] = data_o[22];
  assign data_o[9686] = data_o[22];
  assign data_o[9750] = data_o[22];
  assign data_o[9814] = data_o[22];
  assign data_o[9878] = data_o[22];
  assign data_o[9942] = data_o[22];
  assign data_o[10006] = data_o[22];
  assign data_o[10070] = data_o[22];
  assign data_o[10134] = data_o[22];
  assign data_o[10198] = data_o[22];
  assign data_o[10262] = data_o[22];
  assign data_o[10326] = data_o[22];
  assign data_o[10390] = data_o[22];
  assign data_o[10454] = data_o[22];
  assign data_o[10518] = data_o[22];
  assign data_o[10582] = data_o[22];
  assign data_o[10646] = data_o[22];
  assign data_o[10710] = data_o[22];
  assign data_o[10774] = data_o[22];
  assign data_o[10838] = data_o[22];
  assign data_o[10902] = data_o[22];
  assign data_o[10966] = data_o[22];
  assign data_o[11030] = data_o[22];
  assign data_o[11094] = data_o[22];
  assign data_o[11158] = data_o[22];
  assign data_o[11222] = data_o[22];
  assign data_o[11286] = data_o[22];
  assign data_o[11350] = data_o[22];
  assign data_o[11414] = data_o[22];
  assign data_o[11478] = data_o[22];
  assign data_o[11542] = data_o[22];
  assign data_o[11606] = data_o[22];
  assign data_o[11670] = data_o[22];
  assign data_o[11734] = data_o[22];
  assign data_o[11798] = data_o[22];
  assign data_o[11862] = data_o[22];
  assign data_o[11926] = data_o[22];
  assign data_o[11990] = data_o[22];
  assign data_o[12054] = data_o[22];
  assign data_o[12118] = data_o[22];
  assign data_o[12182] = data_o[22];
  assign data_o[12246] = data_o[22];
  assign data_o[12310] = data_o[22];
  assign data_o[12374] = data_o[22];
  assign data_o[12438] = data_o[22];
  assign data_o[12502] = data_o[22];
  assign data_o[12566] = data_o[22];
  assign data_o[12630] = data_o[22];
  assign data_o[12694] = data_o[22];
  assign data_o[12758] = data_o[22];
  assign data_o[12822] = data_o[22];
  assign data_o[12886] = data_o[22];
  assign data_o[12950] = data_o[22];
  assign data_o[13014] = data_o[22];
  assign data_o[13078] = data_o[22];
  assign data_o[13142] = data_o[22];
  assign data_o[13206] = data_o[22];
  assign data_o[13270] = data_o[22];
  assign data_o[13334] = data_o[22];
  assign data_o[13398] = data_o[22];
  assign data_o[13462] = data_o[22];
  assign data_o[13526] = data_o[22];
  assign data_o[13590] = data_o[22];
  assign data_o[13654] = data_o[22];
  assign data_o[13718] = data_o[22];
  assign data_o[13782] = data_o[22];
  assign data_o[13846] = data_o[22];
  assign data_o[13910] = data_o[22];
  assign data_o[13974] = data_o[22];
  assign data_o[14038] = data_o[22];
  assign data_o[14102] = data_o[22];
  assign data_o[14166] = data_o[22];
  assign data_o[14230] = data_o[22];
  assign data_o[14294] = data_o[22];
  assign data_o[14358] = data_o[22];
  assign data_o[14422] = data_o[22];
  assign data_o[14486] = data_o[22];
  assign data_o[14550] = data_o[22];
  assign data_o[14614] = data_o[22];
  assign data_o[14678] = data_o[22];
  assign data_o[14742] = data_o[22];
  assign data_o[14806] = data_o[22];
  assign data_o[14870] = data_o[22];
  assign data_o[14934] = data_o[22];
  assign data_o[14998] = data_o[22];
  assign data_o[15062] = data_o[22];
  assign data_o[15126] = data_o[22];
  assign data_o[15190] = data_o[22];
  assign data_o[15254] = data_o[22];
  assign data_o[15318] = data_o[22];
  assign data_o[15382] = data_o[22];
  assign data_o[15446] = data_o[22];
  assign data_o[15510] = data_o[22];
  assign data_o[15574] = data_o[22];
  assign data_o[15638] = data_o[22];
  assign data_o[15702] = data_o[22];
  assign data_o[15766] = data_o[22];
  assign data_o[15830] = data_o[22];
  assign data_o[15894] = data_o[22];
  assign data_o[15958] = data_o[22];
  assign data_o[16022] = data_o[22];
  assign data_o[16086] = data_o[22];
  assign data_o[16150] = data_o[22];
  assign data_o[16214] = data_o[22];
  assign data_o[16278] = data_o[22];
  assign data_o[16342] = data_o[22];
  assign data_o[16406] = data_o[22];
  assign data_o[16470] = data_o[22];
  assign data_o[16534] = data_o[22];
  assign data_o[16598] = data_o[22];
  assign data_o[16662] = data_o[22];
  assign data_o[16726] = data_o[22];
  assign data_o[16790] = data_o[22];
  assign data_o[16854] = data_o[22];
  assign data_o[16918] = data_o[22];
  assign data_o[16982] = data_o[22];
  assign data_o[17046] = data_o[22];
  assign data_o[17110] = data_o[22];
  assign data_o[17174] = data_o[22];
  assign data_o[17238] = data_o[22];
  assign data_o[17302] = data_o[22];
  assign data_o[17366] = data_o[22];
  assign data_o[17430] = data_o[22];
  assign data_o[17494] = data_o[22];
  assign data_o[17558] = data_o[22];
  assign data_o[17622] = data_o[22];
  assign data_o[17686] = data_o[22];
  assign data_o[17750] = data_o[22];
  assign data_o[17814] = data_o[22];
  assign data_o[17878] = data_o[22];
  assign data_o[17942] = data_o[22];
  assign data_o[18006] = data_o[22];
  assign data_o[18070] = data_o[22];
  assign data_o[18134] = data_o[22];
  assign data_o[18198] = data_o[22];
  assign data_o[18262] = data_o[22];
  assign data_o[18326] = data_o[22];
  assign data_o[18390] = data_o[22];
  assign data_o[18454] = data_o[22];
  assign data_o[18518] = data_o[22];
  assign data_o[18582] = data_o[22];
  assign data_o[18646] = data_o[22];
  assign data_o[18710] = data_o[22];
  assign data_o[18774] = data_o[22];
  assign data_o[18838] = data_o[22];
  assign data_o[18902] = data_o[22];
  assign data_o[18966] = data_o[22];
  assign data_o[19030] = data_o[22];
  assign data_o[19094] = data_o[22];
  assign data_o[19158] = data_o[22];
  assign data_o[19222] = data_o[22];
  assign data_o[19286] = data_o[22];
  assign data_o[19350] = data_o[22];
  assign data_o[19414] = data_o[22];
  assign data_o[19478] = data_o[22];
  assign data_o[19542] = data_o[22];
  assign data_o[19606] = data_o[22];
  assign data_o[19670] = data_o[22];
  assign data_o[19734] = data_o[22];
  assign data_o[19798] = data_o[22];
  assign data_o[19862] = data_o[22];
  assign data_o[19926] = data_o[22];
  assign data_o[19990] = data_o[22];
  assign data_o[20054] = data_o[22];
  assign data_o[20118] = data_o[22];
  assign data_o[20182] = data_o[22];
  assign data_o[20246] = data_o[22];
  assign data_o[20310] = data_o[22];
  assign data_o[20374] = data_o[22];
  assign data_o[20438] = data_o[22];
  assign data_o[20502] = data_o[22];
  assign data_o[20566] = data_o[22];
  assign data_o[20630] = data_o[22];
  assign data_o[20694] = data_o[22];
  assign data_o[20758] = data_o[22];
  assign data_o[20822] = data_o[22];
  assign data_o[20886] = data_o[22];
  assign data_o[20950] = data_o[22];
  assign data_o[21014] = data_o[22];
  assign data_o[21078] = data_o[22];
  assign data_o[21142] = data_o[22];
  assign data_o[21206] = data_o[22];
  assign data_o[21270] = data_o[22];
  assign data_o[21334] = data_o[22];
  assign data_o[21398] = data_o[22];
  assign data_o[21462] = data_o[22];
  assign data_o[21526] = data_o[22];
  assign data_o[21590] = data_o[22];
  assign data_o[21654] = data_o[22];
  assign data_o[21718] = data_o[22];
  assign data_o[21782] = data_o[22];
  assign data_o[21846] = data_o[22];
  assign data_o[21910] = data_o[22];
  assign data_o[21974] = data_o[22];
  assign data_o[22038] = data_o[22];
  assign data_o[22102] = data_o[22];
  assign data_o[22166] = data_o[22];
  assign data_o[22230] = data_o[22];
  assign data_o[22294] = data_o[22];
  assign data_o[22358] = data_o[22];
  assign data_o[22422] = data_o[22];
  assign data_o[22486] = data_o[22];
  assign data_o[22550] = data_o[22];
  assign data_o[22614] = data_o[22];
  assign data_o[22678] = data_o[22];
  assign data_o[22742] = data_o[22];
  assign data_o[22806] = data_o[22];
  assign data_o[22870] = data_o[22];
  assign data_o[22934] = data_o[22];
  assign data_o[22998] = data_o[22];
  assign data_o[23062] = data_o[22];
  assign data_o[23126] = data_o[22];
  assign data_o[23190] = data_o[22];
  assign data_o[23254] = data_o[22];
  assign data_o[23318] = data_o[22];
  assign data_o[23382] = data_o[22];
  assign data_o[23446] = data_o[22];
  assign data_o[23510] = data_o[22];
  assign data_o[23574] = data_o[22];
  assign data_o[23638] = data_o[22];
  assign data_o[23702] = data_o[22];
  assign data_o[23766] = data_o[22];
  assign data_o[23830] = data_o[22];
  assign data_o[23894] = data_o[22];
  assign data_o[23958] = data_o[22];
  assign data_o[24022] = data_o[22];
  assign data_o[24086] = data_o[22];
  assign data_o[24150] = data_o[22];
  assign data_o[24214] = data_o[22];
  assign data_o[24278] = data_o[22];
  assign data_o[24342] = data_o[22];
  assign data_o[24406] = data_o[22];
  assign data_o[24470] = data_o[22];
  assign data_o[24534] = data_o[22];
  assign data_o[24598] = data_o[22];
  assign data_o[24662] = data_o[22];
  assign data_o[24726] = data_o[22];
  assign data_o[24790] = data_o[22];
  assign data_o[24854] = data_o[22];
  assign data_o[24918] = data_o[22];
  assign data_o[24982] = data_o[22];
  assign data_o[25046] = data_o[22];
  assign data_o[25110] = data_o[22];
  assign data_o[25174] = data_o[22];
  assign data_o[25238] = data_o[22];
  assign data_o[25302] = data_o[22];
  assign data_o[25366] = data_o[22];
  assign data_o[25430] = data_o[22];
  assign data_o[25494] = data_o[22];
  assign data_o[25558] = data_o[22];
  assign data_o[25622] = data_o[22];
  assign data_o[25686] = data_o[22];
  assign data_o[25750] = data_o[22];
  assign data_o[25814] = data_o[22];
  assign data_o[25878] = data_o[22];
  assign data_o[25942] = data_o[22];
  assign data_o[26006] = data_o[22];
  assign data_o[26070] = data_o[22];
  assign data_o[26134] = data_o[22];
  assign data_o[26198] = data_o[22];
  assign data_o[26262] = data_o[22];
  assign data_o[26326] = data_o[22];
  assign data_o[26390] = data_o[22];
  assign data_o[26454] = data_o[22];
  assign data_o[26518] = data_o[22];
  assign data_o[26582] = data_o[22];
  assign data_o[26646] = data_o[22];
  assign data_o[26710] = data_o[22];
  assign data_o[26774] = data_o[22];
  assign data_o[26838] = data_o[22];
  assign data_o[26902] = data_o[22];
  assign data_o[26966] = data_o[22];
  assign data_o[27030] = data_o[22];
  assign data_o[27094] = data_o[22];
  assign data_o[27158] = data_o[22];
  assign data_o[27222] = data_o[22];
  assign data_o[27286] = data_o[22];
  assign data_o[27350] = data_o[22];
  assign data_o[27414] = data_o[22];
  assign data_o[27478] = data_o[22];
  assign data_o[27542] = data_o[22];
  assign data_o[27606] = data_o[22];
  assign data_o[27670] = data_o[22];
  assign data_o[27734] = data_o[22];
  assign data_o[27798] = data_o[22];
  assign data_o[27862] = data_o[22];
  assign data_o[27926] = data_o[22];
  assign data_o[27990] = data_o[22];
  assign data_o[28054] = data_o[22];
  assign data_o[28118] = data_o[22];
  assign data_o[28182] = data_o[22];
  assign data_o[28246] = data_o[22];
  assign data_o[28310] = data_o[22];
  assign data_o[28374] = data_o[22];
  assign data_o[28438] = data_o[22];
  assign data_o[28502] = data_o[22];
  assign data_o[28566] = data_o[22];
  assign data_o[28630] = data_o[22];
  assign data_o[28694] = data_o[22];
  assign data_o[28758] = data_o[22];
  assign data_o[28822] = data_o[22];
  assign data_o[28886] = data_o[22];
  assign data_o[28950] = data_o[22];
  assign data_o[29014] = data_o[22];
  assign data_o[29078] = data_o[22];
  assign data_o[29142] = data_o[22];
  assign data_o[29206] = data_o[22];
  assign data_o[29270] = data_o[22];
  assign data_o[29334] = data_o[22];
  assign data_o[29398] = data_o[22];
  assign data_o[29462] = data_o[22];
  assign data_o[29526] = data_o[22];
  assign data_o[29590] = data_o[22];
  assign data_o[29654] = data_o[22];
  assign data_o[29718] = data_o[22];
  assign data_o[29782] = data_o[22];
  assign data_o[29846] = data_o[22];
  assign data_o[29910] = data_o[22];
  assign data_o[29974] = data_o[22];
  assign data_o[30038] = data_o[22];
  assign data_o[30102] = data_o[22];
  assign data_o[30166] = data_o[22];
  assign data_o[30230] = data_o[22];
  assign data_o[30294] = data_o[22];
  assign data_o[30358] = data_o[22];
  assign data_o[30422] = data_o[22];
  assign data_o[30486] = data_o[22];
  assign data_o[30550] = data_o[22];
  assign data_o[30614] = data_o[22];
  assign data_o[30678] = data_o[22];
  assign data_o[30742] = data_o[22];
  assign data_o[30806] = data_o[22];
  assign data_o[30870] = data_o[22];
  assign data_o[30934] = data_o[22];
  assign data_o[30998] = data_o[22];
  assign data_o[31062] = data_o[22];
  assign data_o[31126] = data_o[22];
  assign data_o[31190] = data_o[22];
  assign data_o[31254] = data_o[22];
  assign data_o[31318] = data_o[22];
  assign data_o[31382] = data_o[22];
  assign data_o[31446] = data_o[22];
  assign data_o[31510] = data_o[22];
  assign data_o[31574] = data_o[22];
  assign data_o[31638] = data_o[22];
  assign data_o[31702] = data_o[22];
  assign data_o[31766] = data_o[22];
  assign data_o[31830] = data_o[22];
  assign data_o[31894] = data_o[22];
  assign data_o[31958] = data_o[22];
  assign data_o[85] = data_o[21];
  assign data_o[149] = data_o[21];
  assign data_o[213] = data_o[21];
  assign data_o[277] = data_o[21];
  assign data_o[341] = data_o[21];
  assign data_o[405] = data_o[21];
  assign data_o[469] = data_o[21];
  assign data_o[533] = data_o[21];
  assign data_o[597] = data_o[21];
  assign data_o[661] = data_o[21];
  assign data_o[725] = data_o[21];
  assign data_o[789] = data_o[21];
  assign data_o[853] = data_o[21];
  assign data_o[917] = data_o[21];
  assign data_o[981] = data_o[21];
  assign data_o[1045] = data_o[21];
  assign data_o[1109] = data_o[21];
  assign data_o[1173] = data_o[21];
  assign data_o[1237] = data_o[21];
  assign data_o[1301] = data_o[21];
  assign data_o[1365] = data_o[21];
  assign data_o[1429] = data_o[21];
  assign data_o[1493] = data_o[21];
  assign data_o[1557] = data_o[21];
  assign data_o[1621] = data_o[21];
  assign data_o[1685] = data_o[21];
  assign data_o[1749] = data_o[21];
  assign data_o[1813] = data_o[21];
  assign data_o[1877] = data_o[21];
  assign data_o[1941] = data_o[21];
  assign data_o[2005] = data_o[21];
  assign data_o[2069] = data_o[21];
  assign data_o[2133] = data_o[21];
  assign data_o[2197] = data_o[21];
  assign data_o[2261] = data_o[21];
  assign data_o[2325] = data_o[21];
  assign data_o[2389] = data_o[21];
  assign data_o[2453] = data_o[21];
  assign data_o[2517] = data_o[21];
  assign data_o[2581] = data_o[21];
  assign data_o[2645] = data_o[21];
  assign data_o[2709] = data_o[21];
  assign data_o[2773] = data_o[21];
  assign data_o[2837] = data_o[21];
  assign data_o[2901] = data_o[21];
  assign data_o[2965] = data_o[21];
  assign data_o[3029] = data_o[21];
  assign data_o[3093] = data_o[21];
  assign data_o[3157] = data_o[21];
  assign data_o[3221] = data_o[21];
  assign data_o[3285] = data_o[21];
  assign data_o[3349] = data_o[21];
  assign data_o[3413] = data_o[21];
  assign data_o[3477] = data_o[21];
  assign data_o[3541] = data_o[21];
  assign data_o[3605] = data_o[21];
  assign data_o[3669] = data_o[21];
  assign data_o[3733] = data_o[21];
  assign data_o[3797] = data_o[21];
  assign data_o[3861] = data_o[21];
  assign data_o[3925] = data_o[21];
  assign data_o[3989] = data_o[21];
  assign data_o[4053] = data_o[21];
  assign data_o[4117] = data_o[21];
  assign data_o[4181] = data_o[21];
  assign data_o[4245] = data_o[21];
  assign data_o[4309] = data_o[21];
  assign data_o[4373] = data_o[21];
  assign data_o[4437] = data_o[21];
  assign data_o[4501] = data_o[21];
  assign data_o[4565] = data_o[21];
  assign data_o[4629] = data_o[21];
  assign data_o[4693] = data_o[21];
  assign data_o[4757] = data_o[21];
  assign data_o[4821] = data_o[21];
  assign data_o[4885] = data_o[21];
  assign data_o[4949] = data_o[21];
  assign data_o[5013] = data_o[21];
  assign data_o[5077] = data_o[21];
  assign data_o[5141] = data_o[21];
  assign data_o[5205] = data_o[21];
  assign data_o[5269] = data_o[21];
  assign data_o[5333] = data_o[21];
  assign data_o[5397] = data_o[21];
  assign data_o[5461] = data_o[21];
  assign data_o[5525] = data_o[21];
  assign data_o[5589] = data_o[21];
  assign data_o[5653] = data_o[21];
  assign data_o[5717] = data_o[21];
  assign data_o[5781] = data_o[21];
  assign data_o[5845] = data_o[21];
  assign data_o[5909] = data_o[21];
  assign data_o[5973] = data_o[21];
  assign data_o[6037] = data_o[21];
  assign data_o[6101] = data_o[21];
  assign data_o[6165] = data_o[21];
  assign data_o[6229] = data_o[21];
  assign data_o[6293] = data_o[21];
  assign data_o[6357] = data_o[21];
  assign data_o[6421] = data_o[21];
  assign data_o[6485] = data_o[21];
  assign data_o[6549] = data_o[21];
  assign data_o[6613] = data_o[21];
  assign data_o[6677] = data_o[21];
  assign data_o[6741] = data_o[21];
  assign data_o[6805] = data_o[21];
  assign data_o[6869] = data_o[21];
  assign data_o[6933] = data_o[21];
  assign data_o[6997] = data_o[21];
  assign data_o[7061] = data_o[21];
  assign data_o[7125] = data_o[21];
  assign data_o[7189] = data_o[21];
  assign data_o[7253] = data_o[21];
  assign data_o[7317] = data_o[21];
  assign data_o[7381] = data_o[21];
  assign data_o[7445] = data_o[21];
  assign data_o[7509] = data_o[21];
  assign data_o[7573] = data_o[21];
  assign data_o[7637] = data_o[21];
  assign data_o[7701] = data_o[21];
  assign data_o[7765] = data_o[21];
  assign data_o[7829] = data_o[21];
  assign data_o[7893] = data_o[21];
  assign data_o[7957] = data_o[21];
  assign data_o[8021] = data_o[21];
  assign data_o[8085] = data_o[21];
  assign data_o[8149] = data_o[21];
  assign data_o[8213] = data_o[21];
  assign data_o[8277] = data_o[21];
  assign data_o[8341] = data_o[21];
  assign data_o[8405] = data_o[21];
  assign data_o[8469] = data_o[21];
  assign data_o[8533] = data_o[21];
  assign data_o[8597] = data_o[21];
  assign data_o[8661] = data_o[21];
  assign data_o[8725] = data_o[21];
  assign data_o[8789] = data_o[21];
  assign data_o[8853] = data_o[21];
  assign data_o[8917] = data_o[21];
  assign data_o[8981] = data_o[21];
  assign data_o[9045] = data_o[21];
  assign data_o[9109] = data_o[21];
  assign data_o[9173] = data_o[21];
  assign data_o[9237] = data_o[21];
  assign data_o[9301] = data_o[21];
  assign data_o[9365] = data_o[21];
  assign data_o[9429] = data_o[21];
  assign data_o[9493] = data_o[21];
  assign data_o[9557] = data_o[21];
  assign data_o[9621] = data_o[21];
  assign data_o[9685] = data_o[21];
  assign data_o[9749] = data_o[21];
  assign data_o[9813] = data_o[21];
  assign data_o[9877] = data_o[21];
  assign data_o[9941] = data_o[21];
  assign data_o[10005] = data_o[21];
  assign data_o[10069] = data_o[21];
  assign data_o[10133] = data_o[21];
  assign data_o[10197] = data_o[21];
  assign data_o[10261] = data_o[21];
  assign data_o[10325] = data_o[21];
  assign data_o[10389] = data_o[21];
  assign data_o[10453] = data_o[21];
  assign data_o[10517] = data_o[21];
  assign data_o[10581] = data_o[21];
  assign data_o[10645] = data_o[21];
  assign data_o[10709] = data_o[21];
  assign data_o[10773] = data_o[21];
  assign data_o[10837] = data_o[21];
  assign data_o[10901] = data_o[21];
  assign data_o[10965] = data_o[21];
  assign data_o[11029] = data_o[21];
  assign data_o[11093] = data_o[21];
  assign data_o[11157] = data_o[21];
  assign data_o[11221] = data_o[21];
  assign data_o[11285] = data_o[21];
  assign data_o[11349] = data_o[21];
  assign data_o[11413] = data_o[21];
  assign data_o[11477] = data_o[21];
  assign data_o[11541] = data_o[21];
  assign data_o[11605] = data_o[21];
  assign data_o[11669] = data_o[21];
  assign data_o[11733] = data_o[21];
  assign data_o[11797] = data_o[21];
  assign data_o[11861] = data_o[21];
  assign data_o[11925] = data_o[21];
  assign data_o[11989] = data_o[21];
  assign data_o[12053] = data_o[21];
  assign data_o[12117] = data_o[21];
  assign data_o[12181] = data_o[21];
  assign data_o[12245] = data_o[21];
  assign data_o[12309] = data_o[21];
  assign data_o[12373] = data_o[21];
  assign data_o[12437] = data_o[21];
  assign data_o[12501] = data_o[21];
  assign data_o[12565] = data_o[21];
  assign data_o[12629] = data_o[21];
  assign data_o[12693] = data_o[21];
  assign data_o[12757] = data_o[21];
  assign data_o[12821] = data_o[21];
  assign data_o[12885] = data_o[21];
  assign data_o[12949] = data_o[21];
  assign data_o[13013] = data_o[21];
  assign data_o[13077] = data_o[21];
  assign data_o[13141] = data_o[21];
  assign data_o[13205] = data_o[21];
  assign data_o[13269] = data_o[21];
  assign data_o[13333] = data_o[21];
  assign data_o[13397] = data_o[21];
  assign data_o[13461] = data_o[21];
  assign data_o[13525] = data_o[21];
  assign data_o[13589] = data_o[21];
  assign data_o[13653] = data_o[21];
  assign data_o[13717] = data_o[21];
  assign data_o[13781] = data_o[21];
  assign data_o[13845] = data_o[21];
  assign data_o[13909] = data_o[21];
  assign data_o[13973] = data_o[21];
  assign data_o[14037] = data_o[21];
  assign data_o[14101] = data_o[21];
  assign data_o[14165] = data_o[21];
  assign data_o[14229] = data_o[21];
  assign data_o[14293] = data_o[21];
  assign data_o[14357] = data_o[21];
  assign data_o[14421] = data_o[21];
  assign data_o[14485] = data_o[21];
  assign data_o[14549] = data_o[21];
  assign data_o[14613] = data_o[21];
  assign data_o[14677] = data_o[21];
  assign data_o[14741] = data_o[21];
  assign data_o[14805] = data_o[21];
  assign data_o[14869] = data_o[21];
  assign data_o[14933] = data_o[21];
  assign data_o[14997] = data_o[21];
  assign data_o[15061] = data_o[21];
  assign data_o[15125] = data_o[21];
  assign data_o[15189] = data_o[21];
  assign data_o[15253] = data_o[21];
  assign data_o[15317] = data_o[21];
  assign data_o[15381] = data_o[21];
  assign data_o[15445] = data_o[21];
  assign data_o[15509] = data_o[21];
  assign data_o[15573] = data_o[21];
  assign data_o[15637] = data_o[21];
  assign data_o[15701] = data_o[21];
  assign data_o[15765] = data_o[21];
  assign data_o[15829] = data_o[21];
  assign data_o[15893] = data_o[21];
  assign data_o[15957] = data_o[21];
  assign data_o[16021] = data_o[21];
  assign data_o[16085] = data_o[21];
  assign data_o[16149] = data_o[21];
  assign data_o[16213] = data_o[21];
  assign data_o[16277] = data_o[21];
  assign data_o[16341] = data_o[21];
  assign data_o[16405] = data_o[21];
  assign data_o[16469] = data_o[21];
  assign data_o[16533] = data_o[21];
  assign data_o[16597] = data_o[21];
  assign data_o[16661] = data_o[21];
  assign data_o[16725] = data_o[21];
  assign data_o[16789] = data_o[21];
  assign data_o[16853] = data_o[21];
  assign data_o[16917] = data_o[21];
  assign data_o[16981] = data_o[21];
  assign data_o[17045] = data_o[21];
  assign data_o[17109] = data_o[21];
  assign data_o[17173] = data_o[21];
  assign data_o[17237] = data_o[21];
  assign data_o[17301] = data_o[21];
  assign data_o[17365] = data_o[21];
  assign data_o[17429] = data_o[21];
  assign data_o[17493] = data_o[21];
  assign data_o[17557] = data_o[21];
  assign data_o[17621] = data_o[21];
  assign data_o[17685] = data_o[21];
  assign data_o[17749] = data_o[21];
  assign data_o[17813] = data_o[21];
  assign data_o[17877] = data_o[21];
  assign data_o[17941] = data_o[21];
  assign data_o[18005] = data_o[21];
  assign data_o[18069] = data_o[21];
  assign data_o[18133] = data_o[21];
  assign data_o[18197] = data_o[21];
  assign data_o[18261] = data_o[21];
  assign data_o[18325] = data_o[21];
  assign data_o[18389] = data_o[21];
  assign data_o[18453] = data_o[21];
  assign data_o[18517] = data_o[21];
  assign data_o[18581] = data_o[21];
  assign data_o[18645] = data_o[21];
  assign data_o[18709] = data_o[21];
  assign data_o[18773] = data_o[21];
  assign data_o[18837] = data_o[21];
  assign data_o[18901] = data_o[21];
  assign data_o[18965] = data_o[21];
  assign data_o[19029] = data_o[21];
  assign data_o[19093] = data_o[21];
  assign data_o[19157] = data_o[21];
  assign data_o[19221] = data_o[21];
  assign data_o[19285] = data_o[21];
  assign data_o[19349] = data_o[21];
  assign data_o[19413] = data_o[21];
  assign data_o[19477] = data_o[21];
  assign data_o[19541] = data_o[21];
  assign data_o[19605] = data_o[21];
  assign data_o[19669] = data_o[21];
  assign data_o[19733] = data_o[21];
  assign data_o[19797] = data_o[21];
  assign data_o[19861] = data_o[21];
  assign data_o[19925] = data_o[21];
  assign data_o[19989] = data_o[21];
  assign data_o[20053] = data_o[21];
  assign data_o[20117] = data_o[21];
  assign data_o[20181] = data_o[21];
  assign data_o[20245] = data_o[21];
  assign data_o[20309] = data_o[21];
  assign data_o[20373] = data_o[21];
  assign data_o[20437] = data_o[21];
  assign data_o[20501] = data_o[21];
  assign data_o[20565] = data_o[21];
  assign data_o[20629] = data_o[21];
  assign data_o[20693] = data_o[21];
  assign data_o[20757] = data_o[21];
  assign data_o[20821] = data_o[21];
  assign data_o[20885] = data_o[21];
  assign data_o[20949] = data_o[21];
  assign data_o[21013] = data_o[21];
  assign data_o[21077] = data_o[21];
  assign data_o[21141] = data_o[21];
  assign data_o[21205] = data_o[21];
  assign data_o[21269] = data_o[21];
  assign data_o[21333] = data_o[21];
  assign data_o[21397] = data_o[21];
  assign data_o[21461] = data_o[21];
  assign data_o[21525] = data_o[21];
  assign data_o[21589] = data_o[21];
  assign data_o[21653] = data_o[21];
  assign data_o[21717] = data_o[21];
  assign data_o[21781] = data_o[21];
  assign data_o[21845] = data_o[21];
  assign data_o[21909] = data_o[21];
  assign data_o[21973] = data_o[21];
  assign data_o[22037] = data_o[21];
  assign data_o[22101] = data_o[21];
  assign data_o[22165] = data_o[21];
  assign data_o[22229] = data_o[21];
  assign data_o[22293] = data_o[21];
  assign data_o[22357] = data_o[21];
  assign data_o[22421] = data_o[21];
  assign data_o[22485] = data_o[21];
  assign data_o[22549] = data_o[21];
  assign data_o[22613] = data_o[21];
  assign data_o[22677] = data_o[21];
  assign data_o[22741] = data_o[21];
  assign data_o[22805] = data_o[21];
  assign data_o[22869] = data_o[21];
  assign data_o[22933] = data_o[21];
  assign data_o[22997] = data_o[21];
  assign data_o[23061] = data_o[21];
  assign data_o[23125] = data_o[21];
  assign data_o[23189] = data_o[21];
  assign data_o[23253] = data_o[21];
  assign data_o[23317] = data_o[21];
  assign data_o[23381] = data_o[21];
  assign data_o[23445] = data_o[21];
  assign data_o[23509] = data_o[21];
  assign data_o[23573] = data_o[21];
  assign data_o[23637] = data_o[21];
  assign data_o[23701] = data_o[21];
  assign data_o[23765] = data_o[21];
  assign data_o[23829] = data_o[21];
  assign data_o[23893] = data_o[21];
  assign data_o[23957] = data_o[21];
  assign data_o[24021] = data_o[21];
  assign data_o[24085] = data_o[21];
  assign data_o[24149] = data_o[21];
  assign data_o[24213] = data_o[21];
  assign data_o[24277] = data_o[21];
  assign data_o[24341] = data_o[21];
  assign data_o[24405] = data_o[21];
  assign data_o[24469] = data_o[21];
  assign data_o[24533] = data_o[21];
  assign data_o[24597] = data_o[21];
  assign data_o[24661] = data_o[21];
  assign data_o[24725] = data_o[21];
  assign data_o[24789] = data_o[21];
  assign data_o[24853] = data_o[21];
  assign data_o[24917] = data_o[21];
  assign data_o[24981] = data_o[21];
  assign data_o[25045] = data_o[21];
  assign data_o[25109] = data_o[21];
  assign data_o[25173] = data_o[21];
  assign data_o[25237] = data_o[21];
  assign data_o[25301] = data_o[21];
  assign data_o[25365] = data_o[21];
  assign data_o[25429] = data_o[21];
  assign data_o[25493] = data_o[21];
  assign data_o[25557] = data_o[21];
  assign data_o[25621] = data_o[21];
  assign data_o[25685] = data_o[21];
  assign data_o[25749] = data_o[21];
  assign data_o[25813] = data_o[21];
  assign data_o[25877] = data_o[21];
  assign data_o[25941] = data_o[21];
  assign data_o[26005] = data_o[21];
  assign data_o[26069] = data_o[21];
  assign data_o[26133] = data_o[21];
  assign data_o[26197] = data_o[21];
  assign data_o[26261] = data_o[21];
  assign data_o[26325] = data_o[21];
  assign data_o[26389] = data_o[21];
  assign data_o[26453] = data_o[21];
  assign data_o[26517] = data_o[21];
  assign data_o[26581] = data_o[21];
  assign data_o[26645] = data_o[21];
  assign data_o[26709] = data_o[21];
  assign data_o[26773] = data_o[21];
  assign data_o[26837] = data_o[21];
  assign data_o[26901] = data_o[21];
  assign data_o[26965] = data_o[21];
  assign data_o[27029] = data_o[21];
  assign data_o[27093] = data_o[21];
  assign data_o[27157] = data_o[21];
  assign data_o[27221] = data_o[21];
  assign data_o[27285] = data_o[21];
  assign data_o[27349] = data_o[21];
  assign data_o[27413] = data_o[21];
  assign data_o[27477] = data_o[21];
  assign data_o[27541] = data_o[21];
  assign data_o[27605] = data_o[21];
  assign data_o[27669] = data_o[21];
  assign data_o[27733] = data_o[21];
  assign data_o[27797] = data_o[21];
  assign data_o[27861] = data_o[21];
  assign data_o[27925] = data_o[21];
  assign data_o[27989] = data_o[21];
  assign data_o[28053] = data_o[21];
  assign data_o[28117] = data_o[21];
  assign data_o[28181] = data_o[21];
  assign data_o[28245] = data_o[21];
  assign data_o[28309] = data_o[21];
  assign data_o[28373] = data_o[21];
  assign data_o[28437] = data_o[21];
  assign data_o[28501] = data_o[21];
  assign data_o[28565] = data_o[21];
  assign data_o[28629] = data_o[21];
  assign data_o[28693] = data_o[21];
  assign data_o[28757] = data_o[21];
  assign data_o[28821] = data_o[21];
  assign data_o[28885] = data_o[21];
  assign data_o[28949] = data_o[21];
  assign data_o[29013] = data_o[21];
  assign data_o[29077] = data_o[21];
  assign data_o[29141] = data_o[21];
  assign data_o[29205] = data_o[21];
  assign data_o[29269] = data_o[21];
  assign data_o[29333] = data_o[21];
  assign data_o[29397] = data_o[21];
  assign data_o[29461] = data_o[21];
  assign data_o[29525] = data_o[21];
  assign data_o[29589] = data_o[21];
  assign data_o[29653] = data_o[21];
  assign data_o[29717] = data_o[21];
  assign data_o[29781] = data_o[21];
  assign data_o[29845] = data_o[21];
  assign data_o[29909] = data_o[21];
  assign data_o[29973] = data_o[21];
  assign data_o[30037] = data_o[21];
  assign data_o[30101] = data_o[21];
  assign data_o[30165] = data_o[21];
  assign data_o[30229] = data_o[21];
  assign data_o[30293] = data_o[21];
  assign data_o[30357] = data_o[21];
  assign data_o[30421] = data_o[21];
  assign data_o[30485] = data_o[21];
  assign data_o[30549] = data_o[21];
  assign data_o[30613] = data_o[21];
  assign data_o[30677] = data_o[21];
  assign data_o[30741] = data_o[21];
  assign data_o[30805] = data_o[21];
  assign data_o[30869] = data_o[21];
  assign data_o[30933] = data_o[21];
  assign data_o[30997] = data_o[21];
  assign data_o[31061] = data_o[21];
  assign data_o[31125] = data_o[21];
  assign data_o[31189] = data_o[21];
  assign data_o[31253] = data_o[21];
  assign data_o[31317] = data_o[21];
  assign data_o[31381] = data_o[21];
  assign data_o[31445] = data_o[21];
  assign data_o[31509] = data_o[21];
  assign data_o[31573] = data_o[21];
  assign data_o[31637] = data_o[21];
  assign data_o[31701] = data_o[21];
  assign data_o[31765] = data_o[21];
  assign data_o[31829] = data_o[21];
  assign data_o[31893] = data_o[21];
  assign data_o[31957] = data_o[21];
  assign data_o[84] = data_o[20];
  assign data_o[148] = data_o[20];
  assign data_o[212] = data_o[20];
  assign data_o[276] = data_o[20];
  assign data_o[340] = data_o[20];
  assign data_o[404] = data_o[20];
  assign data_o[468] = data_o[20];
  assign data_o[532] = data_o[20];
  assign data_o[596] = data_o[20];
  assign data_o[660] = data_o[20];
  assign data_o[724] = data_o[20];
  assign data_o[788] = data_o[20];
  assign data_o[852] = data_o[20];
  assign data_o[916] = data_o[20];
  assign data_o[980] = data_o[20];
  assign data_o[1044] = data_o[20];
  assign data_o[1108] = data_o[20];
  assign data_o[1172] = data_o[20];
  assign data_o[1236] = data_o[20];
  assign data_o[1300] = data_o[20];
  assign data_o[1364] = data_o[20];
  assign data_o[1428] = data_o[20];
  assign data_o[1492] = data_o[20];
  assign data_o[1556] = data_o[20];
  assign data_o[1620] = data_o[20];
  assign data_o[1684] = data_o[20];
  assign data_o[1748] = data_o[20];
  assign data_o[1812] = data_o[20];
  assign data_o[1876] = data_o[20];
  assign data_o[1940] = data_o[20];
  assign data_o[2004] = data_o[20];
  assign data_o[2068] = data_o[20];
  assign data_o[2132] = data_o[20];
  assign data_o[2196] = data_o[20];
  assign data_o[2260] = data_o[20];
  assign data_o[2324] = data_o[20];
  assign data_o[2388] = data_o[20];
  assign data_o[2452] = data_o[20];
  assign data_o[2516] = data_o[20];
  assign data_o[2580] = data_o[20];
  assign data_o[2644] = data_o[20];
  assign data_o[2708] = data_o[20];
  assign data_o[2772] = data_o[20];
  assign data_o[2836] = data_o[20];
  assign data_o[2900] = data_o[20];
  assign data_o[2964] = data_o[20];
  assign data_o[3028] = data_o[20];
  assign data_o[3092] = data_o[20];
  assign data_o[3156] = data_o[20];
  assign data_o[3220] = data_o[20];
  assign data_o[3284] = data_o[20];
  assign data_o[3348] = data_o[20];
  assign data_o[3412] = data_o[20];
  assign data_o[3476] = data_o[20];
  assign data_o[3540] = data_o[20];
  assign data_o[3604] = data_o[20];
  assign data_o[3668] = data_o[20];
  assign data_o[3732] = data_o[20];
  assign data_o[3796] = data_o[20];
  assign data_o[3860] = data_o[20];
  assign data_o[3924] = data_o[20];
  assign data_o[3988] = data_o[20];
  assign data_o[4052] = data_o[20];
  assign data_o[4116] = data_o[20];
  assign data_o[4180] = data_o[20];
  assign data_o[4244] = data_o[20];
  assign data_o[4308] = data_o[20];
  assign data_o[4372] = data_o[20];
  assign data_o[4436] = data_o[20];
  assign data_o[4500] = data_o[20];
  assign data_o[4564] = data_o[20];
  assign data_o[4628] = data_o[20];
  assign data_o[4692] = data_o[20];
  assign data_o[4756] = data_o[20];
  assign data_o[4820] = data_o[20];
  assign data_o[4884] = data_o[20];
  assign data_o[4948] = data_o[20];
  assign data_o[5012] = data_o[20];
  assign data_o[5076] = data_o[20];
  assign data_o[5140] = data_o[20];
  assign data_o[5204] = data_o[20];
  assign data_o[5268] = data_o[20];
  assign data_o[5332] = data_o[20];
  assign data_o[5396] = data_o[20];
  assign data_o[5460] = data_o[20];
  assign data_o[5524] = data_o[20];
  assign data_o[5588] = data_o[20];
  assign data_o[5652] = data_o[20];
  assign data_o[5716] = data_o[20];
  assign data_o[5780] = data_o[20];
  assign data_o[5844] = data_o[20];
  assign data_o[5908] = data_o[20];
  assign data_o[5972] = data_o[20];
  assign data_o[6036] = data_o[20];
  assign data_o[6100] = data_o[20];
  assign data_o[6164] = data_o[20];
  assign data_o[6228] = data_o[20];
  assign data_o[6292] = data_o[20];
  assign data_o[6356] = data_o[20];
  assign data_o[6420] = data_o[20];
  assign data_o[6484] = data_o[20];
  assign data_o[6548] = data_o[20];
  assign data_o[6612] = data_o[20];
  assign data_o[6676] = data_o[20];
  assign data_o[6740] = data_o[20];
  assign data_o[6804] = data_o[20];
  assign data_o[6868] = data_o[20];
  assign data_o[6932] = data_o[20];
  assign data_o[6996] = data_o[20];
  assign data_o[7060] = data_o[20];
  assign data_o[7124] = data_o[20];
  assign data_o[7188] = data_o[20];
  assign data_o[7252] = data_o[20];
  assign data_o[7316] = data_o[20];
  assign data_o[7380] = data_o[20];
  assign data_o[7444] = data_o[20];
  assign data_o[7508] = data_o[20];
  assign data_o[7572] = data_o[20];
  assign data_o[7636] = data_o[20];
  assign data_o[7700] = data_o[20];
  assign data_o[7764] = data_o[20];
  assign data_o[7828] = data_o[20];
  assign data_o[7892] = data_o[20];
  assign data_o[7956] = data_o[20];
  assign data_o[8020] = data_o[20];
  assign data_o[8084] = data_o[20];
  assign data_o[8148] = data_o[20];
  assign data_o[8212] = data_o[20];
  assign data_o[8276] = data_o[20];
  assign data_o[8340] = data_o[20];
  assign data_o[8404] = data_o[20];
  assign data_o[8468] = data_o[20];
  assign data_o[8532] = data_o[20];
  assign data_o[8596] = data_o[20];
  assign data_o[8660] = data_o[20];
  assign data_o[8724] = data_o[20];
  assign data_o[8788] = data_o[20];
  assign data_o[8852] = data_o[20];
  assign data_o[8916] = data_o[20];
  assign data_o[8980] = data_o[20];
  assign data_o[9044] = data_o[20];
  assign data_o[9108] = data_o[20];
  assign data_o[9172] = data_o[20];
  assign data_o[9236] = data_o[20];
  assign data_o[9300] = data_o[20];
  assign data_o[9364] = data_o[20];
  assign data_o[9428] = data_o[20];
  assign data_o[9492] = data_o[20];
  assign data_o[9556] = data_o[20];
  assign data_o[9620] = data_o[20];
  assign data_o[9684] = data_o[20];
  assign data_o[9748] = data_o[20];
  assign data_o[9812] = data_o[20];
  assign data_o[9876] = data_o[20];
  assign data_o[9940] = data_o[20];
  assign data_o[10004] = data_o[20];
  assign data_o[10068] = data_o[20];
  assign data_o[10132] = data_o[20];
  assign data_o[10196] = data_o[20];
  assign data_o[10260] = data_o[20];
  assign data_o[10324] = data_o[20];
  assign data_o[10388] = data_o[20];
  assign data_o[10452] = data_o[20];
  assign data_o[10516] = data_o[20];
  assign data_o[10580] = data_o[20];
  assign data_o[10644] = data_o[20];
  assign data_o[10708] = data_o[20];
  assign data_o[10772] = data_o[20];
  assign data_o[10836] = data_o[20];
  assign data_o[10900] = data_o[20];
  assign data_o[10964] = data_o[20];
  assign data_o[11028] = data_o[20];
  assign data_o[11092] = data_o[20];
  assign data_o[11156] = data_o[20];
  assign data_o[11220] = data_o[20];
  assign data_o[11284] = data_o[20];
  assign data_o[11348] = data_o[20];
  assign data_o[11412] = data_o[20];
  assign data_o[11476] = data_o[20];
  assign data_o[11540] = data_o[20];
  assign data_o[11604] = data_o[20];
  assign data_o[11668] = data_o[20];
  assign data_o[11732] = data_o[20];
  assign data_o[11796] = data_o[20];
  assign data_o[11860] = data_o[20];
  assign data_o[11924] = data_o[20];
  assign data_o[11988] = data_o[20];
  assign data_o[12052] = data_o[20];
  assign data_o[12116] = data_o[20];
  assign data_o[12180] = data_o[20];
  assign data_o[12244] = data_o[20];
  assign data_o[12308] = data_o[20];
  assign data_o[12372] = data_o[20];
  assign data_o[12436] = data_o[20];
  assign data_o[12500] = data_o[20];
  assign data_o[12564] = data_o[20];
  assign data_o[12628] = data_o[20];
  assign data_o[12692] = data_o[20];
  assign data_o[12756] = data_o[20];
  assign data_o[12820] = data_o[20];
  assign data_o[12884] = data_o[20];
  assign data_o[12948] = data_o[20];
  assign data_o[13012] = data_o[20];
  assign data_o[13076] = data_o[20];
  assign data_o[13140] = data_o[20];
  assign data_o[13204] = data_o[20];
  assign data_o[13268] = data_o[20];
  assign data_o[13332] = data_o[20];
  assign data_o[13396] = data_o[20];
  assign data_o[13460] = data_o[20];
  assign data_o[13524] = data_o[20];
  assign data_o[13588] = data_o[20];
  assign data_o[13652] = data_o[20];
  assign data_o[13716] = data_o[20];
  assign data_o[13780] = data_o[20];
  assign data_o[13844] = data_o[20];
  assign data_o[13908] = data_o[20];
  assign data_o[13972] = data_o[20];
  assign data_o[14036] = data_o[20];
  assign data_o[14100] = data_o[20];
  assign data_o[14164] = data_o[20];
  assign data_o[14228] = data_o[20];
  assign data_o[14292] = data_o[20];
  assign data_o[14356] = data_o[20];
  assign data_o[14420] = data_o[20];
  assign data_o[14484] = data_o[20];
  assign data_o[14548] = data_o[20];
  assign data_o[14612] = data_o[20];
  assign data_o[14676] = data_o[20];
  assign data_o[14740] = data_o[20];
  assign data_o[14804] = data_o[20];
  assign data_o[14868] = data_o[20];
  assign data_o[14932] = data_o[20];
  assign data_o[14996] = data_o[20];
  assign data_o[15060] = data_o[20];
  assign data_o[15124] = data_o[20];
  assign data_o[15188] = data_o[20];
  assign data_o[15252] = data_o[20];
  assign data_o[15316] = data_o[20];
  assign data_o[15380] = data_o[20];
  assign data_o[15444] = data_o[20];
  assign data_o[15508] = data_o[20];
  assign data_o[15572] = data_o[20];
  assign data_o[15636] = data_o[20];
  assign data_o[15700] = data_o[20];
  assign data_o[15764] = data_o[20];
  assign data_o[15828] = data_o[20];
  assign data_o[15892] = data_o[20];
  assign data_o[15956] = data_o[20];
  assign data_o[16020] = data_o[20];
  assign data_o[16084] = data_o[20];
  assign data_o[16148] = data_o[20];
  assign data_o[16212] = data_o[20];
  assign data_o[16276] = data_o[20];
  assign data_o[16340] = data_o[20];
  assign data_o[16404] = data_o[20];
  assign data_o[16468] = data_o[20];
  assign data_o[16532] = data_o[20];
  assign data_o[16596] = data_o[20];
  assign data_o[16660] = data_o[20];
  assign data_o[16724] = data_o[20];
  assign data_o[16788] = data_o[20];
  assign data_o[16852] = data_o[20];
  assign data_o[16916] = data_o[20];
  assign data_o[16980] = data_o[20];
  assign data_o[17044] = data_o[20];
  assign data_o[17108] = data_o[20];
  assign data_o[17172] = data_o[20];
  assign data_o[17236] = data_o[20];
  assign data_o[17300] = data_o[20];
  assign data_o[17364] = data_o[20];
  assign data_o[17428] = data_o[20];
  assign data_o[17492] = data_o[20];
  assign data_o[17556] = data_o[20];
  assign data_o[17620] = data_o[20];
  assign data_o[17684] = data_o[20];
  assign data_o[17748] = data_o[20];
  assign data_o[17812] = data_o[20];
  assign data_o[17876] = data_o[20];
  assign data_o[17940] = data_o[20];
  assign data_o[18004] = data_o[20];
  assign data_o[18068] = data_o[20];
  assign data_o[18132] = data_o[20];
  assign data_o[18196] = data_o[20];
  assign data_o[18260] = data_o[20];
  assign data_o[18324] = data_o[20];
  assign data_o[18388] = data_o[20];
  assign data_o[18452] = data_o[20];
  assign data_o[18516] = data_o[20];
  assign data_o[18580] = data_o[20];
  assign data_o[18644] = data_o[20];
  assign data_o[18708] = data_o[20];
  assign data_o[18772] = data_o[20];
  assign data_o[18836] = data_o[20];
  assign data_o[18900] = data_o[20];
  assign data_o[18964] = data_o[20];
  assign data_o[19028] = data_o[20];
  assign data_o[19092] = data_o[20];
  assign data_o[19156] = data_o[20];
  assign data_o[19220] = data_o[20];
  assign data_o[19284] = data_o[20];
  assign data_o[19348] = data_o[20];
  assign data_o[19412] = data_o[20];
  assign data_o[19476] = data_o[20];
  assign data_o[19540] = data_o[20];
  assign data_o[19604] = data_o[20];
  assign data_o[19668] = data_o[20];
  assign data_o[19732] = data_o[20];
  assign data_o[19796] = data_o[20];
  assign data_o[19860] = data_o[20];
  assign data_o[19924] = data_o[20];
  assign data_o[19988] = data_o[20];
  assign data_o[20052] = data_o[20];
  assign data_o[20116] = data_o[20];
  assign data_o[20180] = data_o[20];
  assign data_o[20244] = data_o[20];
  assign data_o[20308] = data_o[20];
  assign data_o[20372] = data_o[20];
  assign data_o[20436] = data_o[20];
  assign data_o[20500] = data_o[20];
  assign data_o[20564] = data_o[20];
  assign data_o[20628] = data_o[20];
  assign data_o[20692] = data_o[20];
  assign data_o[20756] = data_o[20];
  assign data_o[20820] = data_o[20];
  assign data_o[20884] = data_o[20];
  assign data_o[20948] = data_o[20];
  assign data_o[21012] = data_o[20];
  assign data_o[21076] = data_o[20];
  assign data_o[21140] = data_o[20];
  assign data_o[21204] = data_o[20];
  assign data_o[21268] = data_o[20];
  assign data_o[21332] = data_o[20];
  assign data_o[21396] = data_o[20];
  assign data_o[21460] = data_o[20];
  assign data_o[21524] = data_o[20];
  assign data_o[21588] = data_o[20];
  assign data_o[21652] = data_o[20];
  assign data_o[21716] = data_o[20];
  assign data_o[21780] = data_o[20];
  assign data_o[21844] = data_o[20];
  assign data_o[21908] = data_o[20];
  assign data_o[21972] = data_o[20];
  assign data_o[22036] = data_o[20];
  assign data_o[22100] = data_o[20];
  assign data_o[22164] = data_o[20];
  assign data_o[22228] = data_o[20];
  assign data_o[22292] = data_o[20];
  assign data_o[22356] = data_o[20];
  assign data_o[22420] = data_o[20];
  assign data_o[22484] = data_o[20];
  assign data_o[22548] = data_o[20];
  assign data_o[22612] = data_o[20];
  assign data_o[22676] = data_o[20];
  assign data_o[22740] = data_o[20];
  assign data_o[22804] = data_o[20];
  assign data_o[22868] = data_o[20];
  assign data_o[22932] = data_o[20];
  assign data_o[22996] = data_o[20];
  assign data_o[23060] = data_o[20];
  assign data_o[23124] = data_o[20];
  assign data_o[23188] = data_o[20];
  assign data_o[23252] = data_o[20];
  assign data_o[23316] = data_o[20];
  assign data_o[23380] = data_o[20];
  assign data_o[23444] = data_o[20];
  assign data_o[23508] = data_o[20];
  assign data_o[23572] = data_o[20];
  assign data_o[23636] = data_o[20];
  assign data_o[23700] = data_o[20];
  assign data_o[23764] = data_o[20];
  assign data_o[23828] = data_o[20];
  assign data_o[23892] = data_o[20];
  assign data_o[23956] = data_o[20];
  assign data_o[24020] = data_o[20];
  assign data_o[24084] = data_o[20];
  assign data_o[24148] = data_o[20];
  assign data_o[24212] = data_o[20];
  assign data_o[24276] = data_o[20];
  assign data_o[24340] = data_o[20];
  assign data_o[24404] = data_o[20];
  assign data_o[24468] = data_o[20];
  assign data_o[24532] = data_o[20];
  assign data_o[24596] = data_o[20];
  assign data_o[24660] = data_o[20];
  assign data_o[24724] = data_o[20];
  assign data_o[24788] = data_o[20];
  assign data_o[24852] = data_o[20];
  assign data_o[24916] = data_o[20];
  assign data_o[24980] = data_o[20];
  assign data_o[25044] = data_o[20];
  assign data_o[25108] = data_o[20];
  assign data_o[25172] = data_o[20];
  assign data_o[25236] = data_o[20];
  assign data_o[25300] = data_o[20];
  assign data_o[25364] = data_o[20];
  assign data_o[25428] = data_o[20];
  assign data_o[25492] = data_o[20];
  assign data_o[25556] = data_o[20];
  assign data_o[25620] = data_o[20];
  assign data_o[25684] = data_o[20];
  assign data_o[25748] = data_o[20];
  assign data_o[25812] = data_o[20];
  assign data_o[25876] = data_o[20];
  assign data_o[25940] = data_o[20];
  assign data_o[26004] = data_o[20];
  assign data_o[26068] = data_o[20];
  assign data_o[26132] = data_o[20];
  assign data_o[26196] = data_o[20];
  assign data_o[26260] = data_o[20];
  assign data_o[26324] = data_o[20];
  assign data_o[26388] = data_o[20];
  assign data_o[26452] = data_o[20];
  assign data_o[26516] = data_o[20];
  assign data_o[26580] = data_o[20];
  assign data_o[26644] = data_o[20];
  assign data_o[26708] = data_o[20];
  assign data_o[26772] = data_o[20];
  assign data_o[26836] = data_o[20];
  assign data_o[26900] = data_o[20];
  assign data_o[26964] = data_o[20];
  assign data_o[27028] = data_o[20];
  assign data_o[27092] = data_o[20];
  assign data_o[27156] = data_o[20];
  assign data_o[27220] = data_o[20];
  assign data_o[27284] = data_o[20];
  assign data_o[27348] = data_o[20];
  assign data_o[27412] = data_o[20];
  assign data_o[27476] = data_o[20];
  assign data_o[27540] = data_o[20];
  assign data_o[27604] = data_o[20];
  assign data_o[27668] = data_o[20];
  assign data_o[27732] = data_o[20];
  assign data_o[27796] = data_o[20];
  assign data_o[27860] = data_o[20];
  assign data_o[27924] = data_o[20];
  assign data_o[27988] = data_o[20];
  assign data_o[28052] = data_o[20];
  assign data_o[28116] = data_o[20];
  assign data_o[28180] = data_o[20];
  assign data_o[28244] = data_o[20];
  assign data_o[28308] = data_o[20];
  assign data_o[28372] = data_o[20];
  assign data_o[28436] = data_o[20];
  assign data_o[28500] = data_o[20];
  assign data_o[28564] = data_o[20];
  assign data_o[28628] = data_o[20];
  assign data_o[28692] = data_o[20];
  assign data_o[28756] = data_o[20];
  assign data_o[28820] = data_o[20];
  assign data_o[28884] = data_o[20];
  assign data_o[28948] = data_o[20];
  assign data_o[29012] = data_o[20];
  assign data_o[29076] = data_o[20];
  assign data_o[29140] = data_o[20];
  assign data_o[29204] = data_o[20];
  assign data_o[29268] = data_o[20];
  assign data_o[29332] = data_o[20];
  assign data_o[29396] = data_o[20];
  assign data_o[29460] = data_o[20];
  assign data_o[29524] = data_o[20];
  assign data_o[29588] = data_o[20];
  assign data_o[29652] = data_o[20];
  assign data_o[29716] = data_o[20];
  assign data_o[29780] = data_o[20];
  assign data_o[29844] = data_o[20];
  assign data_o[29908] = data_o[20];
  assign data_o[29972] = data_o[20];
  assign data_o[30036] = data_o[20];
  assign data_o[30100] = data_o[20];
  assign data_o[30164] = data_o[20];
  assign data_o[30228] = data_o[20];
  assign data_o[30292] = data_o[20];
  assign data_o[30356] = data_o[20];
  assign data_o[30420] = data_o[20];
  assign data_o[30484] = data_o[20];
  assign data_o[30548] = data_o[20];
  assign data_o[30612] = data_o[20];
  assign data_o[30676] = data_o[20];
  assign data_o[30740] = data_o[20];
  assign data_o[30804] = data_o[20];
  assign data_o[30868] = data_o[20];
  assign data_o[30932] = data_o[20];
  assign data_o[30996] = data_o[20];
  assign data_o[31060] = data_o[20];
  assign data_o[31124] = data_o[20];
  assign data_o[31188] = data_o[20];
  assign data_o[31252] = data_o[20];
  assign data_o[31316] = data_o[20];
  assign data_o[31380] = data_o[20];
  assign data_o[31444] = data_o[20];
  assign data_o[31508] = data_o[20];
  assign data_o[31572] = data_o[20];
  assign data_o[31636] = data_o[20];
  assign data_o[31700] = data_o[20];
  assign data_o[31764] = data_o[20];
  assign data_o[31828] = data_o[20];
  assign data_o[31892] = data_o[20];
  assign data_o[31956] = data_o[20];
  assign data_o[83] = data_o[19];
  assign data_o[147] = data_o[19];
  assign data_o[211] = data_o[19];
  assign data_o[275] = data_o[19];
  assign data_o[339] = data_o[19];
  assign data_o[403] = data_o[19];
  assign data_o[467] = data_o[19];
  assign data_o[531] = data_o[19];
  assign data_o[595] = data_o[19];
  assign data_o[659] = data_o[19];
  assign data_o[723] = data_o[19];
  assign data_o[787] = data_o[19];
  assign data_o[851] = data_o[19];
  assign data_o[915] = data_o[19];
  assign data_o[979] = data_o[19];
  assign data_o[1043] = data_o[19];
  assign data_o[1107] = data_o[19];
  assign data_o[1171] = data_o[19];
  assign data_o[1235] = data_o[19];
  assign data_o[1299] = data_o[19];
  assign data_o[1363] = data_o[19];
  assign data_o[1427] = data_o[19];
  assign data_o[1491] = data_o[19];
  assign data_o[1555] = data_o[19];
  assign data_o[1619] = data_o[19];
  assign data_o[1683] = data_o[19];
  assign data_o[1747] = data_o[19];
  assign data_o[1811] = data_o[19];
  assign data_o[1875] = data_o[19];
  assign data_o[1939] = data_o[19];
  assign data_o[2003] = data_o[19];
  assign data_o[2067] = data_o[19];
  assign data_o[2131] = data_o[19];
  assign data_o[2195] = data_o[19];
  assign data_o[2259] = data_o[19];
  assign data_o[2323] = data_o[19];
  assign data_o[2387] = data_o[19];
  assign data_o[2451] = data_o[19];
  assign data_o[2515] = data_o[19];
  assign data_o[2579] = data_o[19];
  assign data_o[2643] = data_o[19];
  assign data_o[2707] = data_o[19];
  assign data_o[2771] = data_o[19];
  assign data_o[2835] = data_o[19];
  assign data_o[2899] = data_o[19];
  assign data_o[2963] = data_o[19];
  assign data_o[3027] = data_o[19];
  assign data_o[3091] = data_o[19];
  assign data_o[3155] = data_o[19];
  assign data_o[3219] = data_o[19];
  assign data_o[3283] = data_o[19];
  assign data_o[3347] = data_o[19];
  assign data_o[3411] = data_o[19];
  assign data_o[3475] = data_o[19];
  assign data_o[3539] = data_o[19];
  assign data_o[3603] = data_o[19];
  assign data_o[3667] = data_o[19];
  assign data_o[3731] = data_o[19];
  assign data_o[3795] = data_o[19];
  assign data_o[3859] = data_o[19];
  assign data_o[3923] = data_o[19];
  assign data_o[3987] = data_o[19];
  assign data_o[4051] = data_o[19];
  assign data_o[4115] = data_o[19];
  assign data_o[4179] = data_o[19];
  assign data_o[4243] = data_o[19];
  assign data_o[4307] = data_o[19];
  assign data_o[4371] = data_o[19];
  assign data_o[4435] = data_o[19];
  assign data_o[4499] = data_o[19];
  assign data_o[4563] = data_o[19];
  assign data_o[4627] = data_o[19];
  assign data_o[4691] = data_o[19];
  assign data_o[4755] = data_o[19];
  assign data_o[4819] = data_o[19];
  assign data_o[4883] = data_o[19];
  assign data_o[4947] = data_o[19];
  assign data_o[5011] = data_o[19];
  assign data_o[5075] = data_o[19];
  assign data_o[5139] = data_o[19];
  assign data_o[5203] = data_o[19];
  assign data_o[5267] = data_o[19];
  assign data_o[5331] = data_o[19];
  assign data_o[5395] = data_o[19];
  assign data_o[5459] = data_o[19];
  assign data_o[5523] = data_o[19];
  assign data_o[5587] = data_o[19];
  assign data_o[5651] = data_o[19];
  assign data_o[5715] = data_o[19];
  assign data_o[5779] = data_o[19];
  assign data_o[5843] = data_o[19];
  assign data_o[5907] = data_o[19];
  assign data_o[5971] = data_o[19];
  assign data_o[6035] = data_o[19];
  assign data_o[6099] = data_o[19];
  assign data_o[6163] = data_o[19];
  assign data_o[6227] = data_o[19];
  assign data_o[6291] = data_o[19];
  assign data_o[6355] = data_o[19];
  assign data_o[6419] = data_o[19];
  assign data_o[6483] = data_o[19];
  assign data_o[6547] = data_o[19];
  assign data_o[6611] = data_o[19];
  assign data_o[6675] = data_o[19];
  assign data_o[6739] = data_o[19];
  assign data_o[6803] = data_o[19];
  assign data_o[6867] = data_o[19];
  assign data_o[6931] = data_o[19];
  assign data_o[6995] = data_o[19];
  assign data_o[7059] = data_o[19];
  assign data_o[7123] = data_o[19];
  assign data_o[7187] = data_o[19];
  assign data_o[7251] = data_o[19];
  assign data_o[7315] = data_o[19];
  assign data_o[7379] = data_o[19];
  assign data_o[7443] = data_o[19];
  assign data_o[7507] = data_o[19];
  assign data_o[7571] = data_o[19];
  assign data_o[7635] = data_o[19];
  assign data_o[7699] = data_o[19];
  assign data_o[7763] = data_o[19];
  assign data_o[7827] = data_o[19];
  assign data_o[7891] = data_o[19];
  assign data_o[7955] = data_o[19];
  assign data_o[8019] = data_o[19];
  assign data_o[8083] = data_o[19];
  assign data_o[8147] = data_o[19];
  assign data_o[8211] = data_o[19];
  assign data_o[8275] = data_o[19];
  assign data_o[8339] = data_o[19];
  assign data_o[8403] = data_o[19];
  assign data_o[8467] = data_o[19];
  assign data_o[8531] = data_o[19];
  assign data_o[8595] = data_o[19];
  assign data_o[8659] = data_o[19];
  assign data_o[8723] = data_o[19];
  assign data_o[8787] = data_o[19];
  assign data_o[8851] = data_o[19];
  assign data_o[8915] = data_o[19];
  assign data_o[8979] = data_o[19];
  assign data_o[9043] = data_o[19];
  assign data_o[9107] = data_o[19];
  assign data_o[9171] = data_o[19];
  assign data_o[9235] = data_o[19];
  assign data_o[9299] = data_o[19];
  assign data_o[9363] = data_o[19];
  assign data_o[9427] = data_o[19];
  assign data_o[9491] = data_o[19];
  assign data_o[9555] = data_o[19];
  assign data_o[9619] = data_o[19];
  assign data_o[9683] = data_o[19];
  assign data_o[9747] = data_o[19];
  assign data_o[9811] = data_o[19];
  assign data_o[9875] = data_o[19];
  assign data_o[9939] = data_o[19];
  assign data_o[10003] = data_o[19];
  assign data_o[10067] = data_o[19];
  assign data_o[10131] = data_o[19];
  assign data_o[10195] = data_o[19];
  assign data_o[10259] = data_o[19];
  assign data_o[10323] = data_o[19];
  assign data_o[10387] = data_o[19];
  assign data_o[10451] = data_o[19];
  assign data_o[10515] = data_o[19];
  assign data_o[10579] = data_o[19];
  assign data_o[10643] = data_o[19];
  assign data_o[10707] = data_o[19];
  assign data_o[10771] = data_o[19];
  assign data_o[10835] = data_o[19];
  assign data_o[10899] = data_o[19];
  assign data_o[10963] = data_o[19];
  assign data_o[11027] = data_o[19];
  assign data_o[11091] = data_o[19];
  assign data_o[11155] = data_o[19];
  assign data_o[11219] = data_o[19];
  assign data_o[11283] = data_o[19];
  assign data_o[11347] = data_o[19];
  assign data_o[11411] = data_o[19];
  assign data_o[11475] = data_o[19];
  assign data_o[11539] = data_o[19];
  assign data_o[11603] = data_o[19];
  assign data_o[11667] = data_o[19];
  assign data_o[11731] = data_o[19];
  assign data_o[11795] = data_o[19];
  assign data_o[11859] = data_o[19];
  assign data_o[11923] = data_o[19];
  assign data_o[11987] = data_o[19];
  assign data_o[12051] = data_o[19];
  assign data_o[12115] = data_o[19];
  assign data_o[12179] = data_o[19];
  assign data_o[12243] = data_o[19];
  assign data_o[12307] = data_o[19];
  assign data_o[12371] = data_o[19];
  assign data_o[12435] = data_o[19];
  assign data_o[12499] = data_o[19];
  assign data_o[12563] = data_o[19];
  assign data_o[12627] = data_o[19];
  assign data_o[12691] = data_o[19];
  assign data_o[12755] = data_o[19];
  assign data_o[12819] = data_o[19];
  assign data_o[12883] = data_o[19];
  assign data_o[12947] = data_o[19];
  assign data_o[13011] = data_o[19];
  assign data_o[13075] = data_o[19];
  assign data_o[13139] = data_o[19];
  assign data_o[13203] = data_o[19];
  assign data_o[13267] = data_o[19];
  assign data_o[13331] = data_o[19];
  assign data_o[13395] = data_o[19];
  assign data_o[13459] = data_o[19];
  assign data_o[13523] = data_o[19];
  assign data_o[13587] = data_o[19];
  assign data_o[13651] = data_o[19];
  assign data_o[13715] = data_o[19];
  assign data_o[13779] = data_o[19];
  assign data_o[13843] = data_o[19];
  assign data_o[13907] = data_o[19];
  assign data_o[13971] = data_o[19];
  assign data_o[14035] = data_o[19];
  assign data_o[14099] = data_o[19];
  assign data_o[14163] = data_o[19];
  assign data_o[14227] = data_o[19];
  assign data_o[14291] = data_o[19];
  assign data_o[14355] = data_o[19];
  assign data_o[14419] = data_o[19];
  assign data_o[14483] = data_o[19];
  assign data_o[14547] = data_o[19];
  assign data_o[14611] = data_o[19];
  assign data_o[14675] = data_o[19];
  assign data_o[14739] = data_o[19];
  assign data_o[14803] = data_o[19];
  assign data_o[14867] = data_o[19];
  assign data_o[14931] = data_o[19];
  assign data_o[14995] = data_o[19];
  assign data_o[15059] = data_o[19];
  assign data_o[15123] = data_o[19];
  assign data_o[15187] = data_o[19];
  assign data_o[15251] = data_o[19];
  assign data_o[15315] = data_o[19];
  assign data_o[15379] = data_o[19];
  assign data_o[15443] = data_o[19];
  assign data_o[15507] = data_o[19];
  assign data_o[15571] = data_o[19];
  assign data_o[15635] = data_o[19];
  assign data_o[15699] = data_o[19];
  assign data_o[15763] = data_o[19];
  assign data_o[15827] = data_o[19];
  assign data_o[15891] = data_o[19];
  assign data_o[15955] = data_o[19];
  assign data_o[16019] = data_o[19];
  assign data_o[16083] = data_o[19];
  assign data_o[16147] = data_o[19];
  assign data_o[16211] = data_o[19];
  assign data_o[16275] = data_o[19];
  assign data_o[16339] = data_o[19];
  assign data_o[16403] = data_o[19];
  assign data_o[16467] = data_o[19];
  assign data_o[16531] = data_o[19];
  assign data_o[16595] = data_o[19];
  assign data_o[16659] = data_o[19];
  assign data_o[16723] = data_o[19];
  assign data_o[16787] = data_o[19];
  assign data_o[16851] = data_o[19];
  assign data_o[16915] = data_o[19];
  assign data_o[16979] = data_o[19];
  assign data_o[17043] = data_o[19];
  assign data_o[17107] = data_o[19];
  assign data_o[17171] = data_o[19];
  assign data_o[17235] = data_o[19];
  assign data_o[17299] = data_o[19];
  assign data_o[17363] = data_o[19];
  assign data_o[17427] = data_o[19];
  assign data_o[17491] = data_o[19];
  assign data_o[17555] = data_o[19];
  assign data_o[17619] = data_o[19];
  assign data_o[17683] = data_o[19];
  assign data_o[17747] = data_o[19];
  assign data_o[17811] = data_o[19];
  assign data_o[17875] = data_o[19];
  assign data_o[17939] = data_o[19];
  assign data_o[18003] = data_o[19];
  assign data_o[18067] = data_o[19];
  assign data_o[18131] = data_o[19];
  assign data_o[18195] = data_o[19];
  assign data_o[18259] = data_o[19];
  assign data_o[18323] = data_o[19];
  assign data_o[18387] = data_o[19];
  assign data_o[18451] = data_o[19];
  assign data_o[18515] = data_o[19];
  assign data_o[18579] = data_o[19];
  assign data_o[18643] = data_o[19];
  assign data_o[18707] = data_o[19];
  assign data_o[18771] = data_o[19];
  assign data_o[18835] = data_o[19];
  assign data_o[18899] = data_o[19];
  assign data_o[18963] = data_o[19];
  assign data_o[19027] = data_o[19];
  assign data_o[19091] = data_o[19];
  assign data_o[19155] = data_o[19];
  assign data_o[19219] = data_o[19];
  assign data_o[19283] = data_o[19];
  assign data_o[19347] = data_o[19];
  assign data_o[19411] = data_o[19];
  assign data_o[19475] = data_o[19];
  assign data_o[19539] = data_o[19];
  assign data_o[19603] = data_o[19];
  assign data_o[19667] = data_o[19];
  assign data_o[19731] = data_o[19];
  assign data_o[19795] = data_o[19];
  assign data_o[19859] = data_o[19];
  assign data_o[19923] = data_o[19];
  assign data_o[19987] = data_o[19];
  assign data_o[20051] = data_o[19];
  assign data_o[20115] = data_o[19];
  assign data_o[20179] = data_o[19];
  assign data_o[20243] = data_o[19];
  assign data_o[20307] = data_o[19];
  assign data_o[20371] = data_o[19];
  assign data_o[20435] = data_o[19];
  assign data_o[20499] = data_o[19];
  assign data_o[20563] = data_o[19];
  assign data_o[20627] = data_o[19];
  assign data_o[20691] = data_o[19];
  assign data_o[20755] = data_o[19];
  assign data_o[20819] = data_o[19];
  assign data_o[20883] = data_o[19];
  assign data_o[20947] = data_o[19];
  assign data_o[21011] = data_o[19];
  assign data_o[21075] = data_o[19];
  assign data_o[21139] = data_o[19];
  assign data_o[21203] = data_o[19];
  assign data_o[21267] = data_o[19];
  assign data_o[21331] = data_o[19];
  assign data_o[21395] = data_o[19];
  assign data_o[21459] = data_o[19];
  assign data_o[21523] = data_o[19];
  assign data_o[21587] = data_o[19];
  assign data_o[21651] = data_o[19];
  assign data_o[21715] = data_o[19];
  assign data_o[21779] = data_o[19];
  assign data_o[21843] = data_o[19];
  assign data_o[21907] = data_o[19];
  assign data_o[21971] = data_o[19];
  assign data_o[22035] = data_o[19];
  assign data_o[22099] = data_o[19];
  assign data_o[22163] = data_o[19];
  assign data_o[22227] = data_o[19];
  assign data_o[22291] = data_o[19];
  assign data_o[22355] = data_o[19];
  assign data_o[22419] = data_o[19];
  assign data_o[22483] = data_o[19];
  assign data_o[22547] = data_o[19];
  assign data_o[22611] = data_o[19];
  assign data_o[22675] = data_o[19];
  assign data_o[22739] = data_o[19];
  assign data_o[22803] = data_o[19];
  assign data_o[22867] = data_o[19];
  assign data_o[22931] = data_o[19];
  assign data_o[22995] = data_o[19];
  assign data_o[23059] = data_o[19];
  assign data_o[23123] = data_o[19];
  assign data_o[23187] = data_o[19];
  assign data_o[23251] = data_o[19];
  assign data_o[23315] = data_o[19];
  assign data_o[23379] = data_o[19];
  assign data_o[23443] = data_o[19];
  assign data_o[23507] = data_o[19];
  assign data_o[23571] = data_o[19];
  assign data_o[23635] = data_o[19];
  assign data_o[23699] = data_o[19];
  assign data_o[23763] = data_o[19];
  assign data_o[23827] = data_o[19];
  assign data_o[23891] = data_o[19];
  assign data_o[23955] = data_o[19];
  assign data_o[24019] = data_o[19];
  assign data_o[24083] = data_o[19];
  assign data_o[24147] = data_o[19];
  assign data_o[24211] = data_o[19];
  assign data_o[24275] = data_o[19];
  assign data_o[24339] = data_o[19];
  assign data_o[24403] = data_o[19];
  assign data_o[24467] = data_o[19];
  assign data_o[24531] = data_o[19];
  assign data_o[24595] = data_o[19];
  assign data_o[24659] = data_o[19];
  assign data_o[24723] = data_o[19];
  assign data_o[24787] = data_o[19];
  assign data_o[24851] = data_o[19];
  assign data_o[24915] = data_o[19];
  assign data_o[24979] = data_o[19];
  assign data_o[25043] = data_o[19];
  assign data_o[25107] = data_o[19];
  assign data_o[25171] = data_o[19];
  assign data_o[25235] = data_o[19];
  assign data_o[25299] = data_o[19];
  assign data_o[25363] = data_o[19];
  assign data_o[25427] = data_o[19];
  assign data_o[25491] = data_o[19];
  assign data_o[25555] = data_o[19];
  assign data_o[25619] = data_o[19];
  assign data_o[25683] = data_o[19];
  assign data_o[25747] = data_o[19];
  assign data_o[25811] = data_o[19];
  assign data_o[25875] = data_o[19];
  assign data_o[25939] = data_o[19];
  assign data_o[26003] = data_o[19];
  assign data_o[26067] = data_o[19];
  assign data_o[26131] = data_o[19];
  assign data_o[26195] = data_o[19];
  assign data_o[26259] = data_o[19];
  assign data_o[26323] = data_o[19];
  assign data_o[26387] = data_o[19];
  assign data_o[26451] = data_o[19];
  assign data_o[26515] = data_o[19];
  assign data_o[26579] = data_o[19];
  assign data_o[26643] = data_o[19];
  assign data_o[26707] = data_o[19];
  assign data_o[26771] = data_o[19];
  assign data_o[26835] = data_o[19];
  assign data_o[26899] = data_o[19];
  assign data_o[26963] = data_o[19];
  assign data_o[27027] = data_o[19];
  assign data_o[27091] = data_o[19];
  assign data_o[27155] = data_o[19];
  assign data_o[27219] = data_o[19];
  assign data_o[27283] = data_o[19];
  assign data_o[27347] = data_o[19];
  assign data_o[27411] = data_o[19];
  assign data_o[27475] = data_o[19];
  assign data_o[27539] = data_o[19];
  assign data_o[27603] = data_o[19];
  assign data_o[27667] = data_o[19];
  assign data_o[27731] = data_o[19];
  assign data_o[27795] = data_o[19];
  assign data_o[27859] = data_o[19];
  assign data_o[27923] = data_o[19];
  assign data_o[27987] = data_o[19];
  assign data_o[28051] = data_o[19];
  assign data_o[28115] = data_o[19];
  assign data_o[28179] = data_o[19];
  assign data_o[28243] = data_o[19];
  assign data_o[28307] = data_o[19];
  assign data_o[28371] = data_o[19];
  assign data_o[28435] = data_o[19];
  assign data_o[28499] = data_o[19];
  assign data_o[28563] = data_o[19];
  assign data_o[28627] = data_o[19];
  assign data_o[28691] = data_o[19];
  assign data_o[28755] = data_o[19];
  assign data_o[28819] = data_o[19];
  assign data_o[28883] = data_o[19];
  assign data_o[28947] = data_o[19];
  assign data_o[29011] = data_o[19];
  assign data_o[29075] = data_o[19];
  assign data_o[29139] = data_o[19];
  assign data_o[29203] = data_o[19];
  assign data_o[29267] = data_o[19];
  assign data_o[29331] = data_o[19];
  assign data_o[29395] = data_o[19];
  assign data_o[29459] = data_o[19];
  assign data_o[29523] = data_o[19];
  assign data_o[29587] = data_o[19];
  assign data_o[29651] = data_o[19];
  assign data_o[29715] = data_o[19];
  assign data_o[29779] = data_o[19];
  assign data_o[29843] = data_o[19];
  assign data_o[29907] = data_o[19];
  assign data_o[29971] = data_o[19];
  assign data_o[30035] = data_o[19];
  assign data_o[30099] = data_o[19];
  assign data_o[30163] = data_o[19];
  assign data_o[30227] = data_o[19];
  assign data_o[30291] = data_o[19];
  assign data_o[30355] = data_o[19];
  assign data_o[30419] = data_o[19];
  assign data_o[30483] = data_o[19];
  assign data_o[30547] = data_o[19];
  assign data_o[30611] = data_o[19];
  assign data_o[30675] = data_o[19];
  assign data_o[30739] = data_o[19];
  assign data_o[30803] = data_o[19];
  assign data_o[30867] = data_o[19];
  assign data_o[30931] = data_o[19];
  assign data_o[30995] = data_o[19];
  assign data_o[31059] = data_o[19];
  assign data_o[31123] = data_o[19];
  assign data_o[31187] = data_o[19];
  assign data_o[31251] = data_o[19];
  assign data_o[31315] = data_o[19];
  assign data_o[31379] = data_o[19];
  assign data_o[31443] = data_o[19];
  assign data_o[31507] = data_o[19];
  assign data_o[31571] = data_o[19];
  assign data_o[31635] = data_o[19];
  assign data_o[31699] = data_o[19];
  assign data_o[31763] = data_o[19];
  assign data_o[31827] = data_o[19];
  assign data_o[31891] = data_o[19];
  assign data_o[31955] = data_o[19];
  assign data_o[82] = data_o[18];
  assign data_o[146] = data_o[18];
  assign data_o[210] = data_o[18];
  assign data_o[274] = data_o[18];
  assign data_o[338] = data_o[18];
  assign data_o[402] = data_o[18];
  assign data_o[466] = data_o[18];
  assign data_o[530] = data_o[18];
  assign data_o[594] = data_o[18];
  assign data_o[658] = data_o[18];
  assign data_o[722] = data_o[18];
  assign data_o[786] = data_o[18];
  assign data_o[850] = data_o[18];
  assign data_o[914] = data_o[18];
  assign data_o[978] = data_o[18];
  assign data_o[1042] = data_o[18];
  assign data_o[1106] = data_o[18];
  assign data_o[1170] = data_o[18];
  assign data_o[1234] = data_o[18];
  assign data_o[1298] = data_o[18];
  assign data_o[1362] = data_o[18];
  assign data_o[1426] = data_o[18];
  assign data_o[1490] = data_o[18];
  assign data_o[1554] = data_o[18];
  assign data_o[1618] = data_o[18];
  assign data_o[1682] = data_o[18];
  assign data_o[1746] = data_o[18];
  assign data_o[1810] = data_o[18];
  assign data_o[1874] = data_o[18];
  assign data_o[1938] = data_o[18];
  assign data_o[2002] = data_o[18];
  assign data_o[2066] = data_o[18];
  assign data_o[2130] = data_o[18];
  assign data_o[2194] = data_o[18];
  assign data_o[2258] = data_o[18];
  assign data_o[2322] = data_o[18];
  assign data_o[2386] = data_o[18];
  assign data_o[2450] = data_o[18];
  assign data_o[2514] = data_o[18];
  assign data_o[2578] = data_o[18];
  assign data_o[2642] = data_o[18];
  assign data_o[2706] = data_o[18];
  assign data_o[2770] = data_o[18];
  assign data_o[2834] = data_o[18];
  assign data_o[2898] = data_o[18];
  assign data_o[2962] = data_o[18];
  assign data_o[3026] = data_o[18];
  assign data_o[3090] = data_o[18];
  assign data_o[3154] = data_o[18];
  assign data_o[3218] = data_o[18];
  assign data_o[3282] = data_o[18];
  assign data_o[3346] = data_o[18];
  assign data_o[3410] = data_o[18];
  assign data_o[3474] = data_o[18];
  assign data_o[3538] = data_o[18];
  assign data_o[3602] = data_o[18];
  assign data_o[3666] = data_o[18];
  assign data_o[3730] = data_o[18];
  assign data_o[3794] = data_o[18];
  assign data_o[3858] = data_o[18];
  assign data_o[3922] = data_o[18];
  assign data_o[3986] = data_o[18];
  assign data_o[4050] = data_o[18];
  assign data_o[4114] = data_o[18];
  assign data_o[4178] = data_o[18];
  assign data_o[4242] = data_o[18];
  assign data_o[4306] = data_o[18];
  assign data_o[4370] = data_o[18];
  assign data_o[4434] = data_o[18];
  assign data_o[4498] = data_o[18];
  assign data_o[4562] = data_o[18];
  assign data_o[4626] = data_o[18];
  assign data_o[4690] = data_o[18];
  assign data_o[4754] = data_o[18];
  assign data_o[4818] = data_o[18];
  assign data_o[4882] = data_o[18];
  assign data_o[4946] = data_o[18];
  assign data_o[5010] = data_o[18];
  assign data_o[5074] = data_o[18];
  assign data_o[5138] = data_o[18];
  assign data_o[5202] = data_o[18];
  assign data_o[5266] = data_o[18];
  assign data_o[5330] = data_o[18];
  assign data_o[5394] = data_o[18];
  assign data_o[5458] = data_o[18];
  assign data_o[5522] = data_o[18];
  assign data_o[5586] = data_o[18];
  assign data_o[5650] = data_o[18];
  assign data_o[5714] = data_o[18];
  assign data_o[5778] = data_o[18];
  assign data_o[5842] = data_o[18];
  assign data_o[5906] = data_o[18];
  assign data_o[5970] = data_o[18];
  assign data_o[6034] = data_o[18];
  assign data_o[6098] = data_o[18];
  assign data_o[6162] = data_o[18];
  assign data_o[6226] = data_o[18];
  assign data_o[6290] = data_o[18];
  assign data_o[6354] = data_o[18];
  assign data_o[6418] = data_o[18];
  assign data_o[6482] = data_o[18];
  assign data_o[6546] = data_o[18];
  assign data_o[6610] = data_o[18];
  assign data_o[6674] = data_o[18];
  assign data_o[6738] = data_o[18];
  assign data_o[6802] = data_o[18];
  assign data_o[6866] = data_o[18];
  assign data_o[6930] = data_o[18];
  assign data_o[6994] = data_o[18];
  assign data_o[7058] = data_o[18];
  assign data_o[7122] = data_o[18];
  assign data_o[7186] = data_o[18];
  assign data_o[7250] = data_o[18];
  assign data_o[7314] = data_o[18];
  assign data_o[7378] = data_o[18];
  assign data_o[7442] = data_o[18];
  assign data_o[7506] = data_o[18];
  assign data_o[7570] = data_o[18];
  assign data_o[7634] = data_o[18];
  assign data_o[7698] = data_o[18];
  assign data_o[7762] = data_o[18];
  assign data_o[7826] = data_o[18];
  assign data_o[7890] = data_o[18];
  assign data_o[7954] = data_o[18];
  assign data_o[8018] = data_o[18];
  assign data_o[8082] = data_o[18];
  assign data_o[8146] = data_o[18];
  assign data_o[8210] = data_o[18];
  assign data_o[8274] = data_o[18];
  assign data_o[8338] = data_o[18];
  assign data_o[8402] = data_o[18];
  assign data_o[8466] = data_o[18];
  assign data_o[8530] = data_o[18];
  assign data_o[8594] = data_o[18];
  assign data_o[8658] = data_o[18];
  assign data_o[8722] = data_o[18];
  assign data_o[8786] = data_o[18];
  assign data_o[8850] = data_o[18];
  assign data_o[8914] = data_o[18];
  assign data_o[8978] = data_o[18];
  assign data_o[9042] = data_o[18];
  assign data_o[9106] = data_o[18];
  assign data_o[9170] = data_o[18];
  assign data_o[9234] = data_o[18];
  assign data_o[9298] = data_o[18];
  assign data_o[9362] = data_o[18];
  assign data_o[9426] = data_o[18];
  assign data_o[9490] = data_o[18];
  assign data_o[9554] = data_o[18];
  assign data_o[9618] = data_o[18];
  assign data_o[9682] = data_o[18];
  assign data_o[9746] = data_o[18];
  assign data_o[9810] = data_o[18];
  assign data_o[9874] = data_o[18];
  assign data_o[9938] = data_o[18];
  assign data_o[10002] = data_o[18];
  assign data_o[10066] = data_o[18];
  assign data_o[10130] = data_o[18];
  assign data_o[10194] = data_o[18];
  assign data_o[10258] = data_o[18];
  assign data_o[10322] = data_o[18];
  assign data_o[10386] = data_o[18];
  assign data_o[10450] = data_o[18];
  assign data_o[10514] = data_o[18];
  assign data_o[10578] = data_o[18];
  assign data_o[10642] = data_o[18];
  assign data_o[10706] = data_o[18];
  assign data_o[10770] = data_o[18];
  assign data_o[10834] = data_o[18];
  assign data_o[10898] = data_o[18];
  assign data_o[10962] = data_o[18];
  assign data_o[11026] = data_o[18];
  assign data_o[11090] = data_o[18];
  assign data_o[11154] = data_o[18];
  assign data_o[11218] = data_o[18];
  assign data_o[11282] = data_o[18];
  assign data_o[11346] = data_o[18];
  assign data_o[11410] = data_o[18];
  assign data_o[11474] = data_o[18];
  assign data_o[11538] = data_o[18];
  assign data_o[11602] = data_o[18];
  assign data_o[11666] = data_o[18];
  assign data_o[11730] = data_o[18];
  assign data_o[11794] = data_o[18];
  assign data_o[11858] = data_o[18];
  assign data_o[11922] = data_o[18];
  assign data_o[11986] = data_o[18];
  assign data_o[12050] = data_o[18];
  assign data_o[12114] = data_o[18];
  assign data_o[12178] = data_o[18];
  assign data_o[12242] = data_o[18];
  assign data_o[12306] = data_o[18];
  assign data_o[12370] = data_o[18];
  assign data_o[12434] = data_o[18];
  assign data_o[12498] = data_o[18];
  assign data_o[12562] = data_o[18];
  assign data_o[12626] = data_o[18];
  assign data_o[12690] = data_o[18];
  assign data_o[12754] = data_o[18];
  assign data_o[12818] = data_o[18];
  assign data_o[12882] = data_o[18];
  assign data_o[12946] = data_o[18];
  assign data_o[13010] = data_o[18];
  assign data_o[13074] = data_o[18];
  assign data_o[13138] = data_o[18];
  assign data_o[13202] = data_o[18];
  assign data_o[13266] = data_o[18];
  assign data_o[13330] = data_o[18];
  assign data_o[13394] = data_o[18];
  assign data_o[13458] = data_o[18];
  assign data_o[13522] = data_o[18];
  assign data_o[13586] = data_o[18];
  assign data_o[13650] = data_o[18];
  assign data_o[13714] = data_o[18];
  assign data_o[13778] = data_o[18];
  assign data_o[13842] = data_o[18];
  assign data_o[13906] = data_o[18];
  assign data_o[13970] = data_o[18];
  assign data_o[14034] = data_o[18];
  assign data_o[14098] = data_o[18];
  assign data_o[14162] = data_o[18];
  assign data_o[14226] = data_o[18];
  assign data_o[14290] = data_o[18];
  assign data_o[14354] = data_o[18];
  assign data_o[14418] = data_o[18];
  assign data_o[14482] = data_o[18];
  assign data_o[14546] = data_o[18];
  assign data_o[14610] = data_o[18];
  assign data_o[14674] = data_o[18];
  assign data_o[14738] = data_o[18];
  assign data_o[14802] = data_o[18];
  assign data_o[14866] = data_o[18];
  assign data_o[14930] = data_o[18];
  assign data_o[14994] = data_o[18];
  assign data_o[15058] = data_o[18];
  assign data_o[15122] = data_o[18];
  assign data_o[15186] = data_o[18];
  assign data_o[15250] = data_o[18];
  assign data_o[15314] = data_o[18];
  assign data_o[15378] = data_o[18];
  assign data_o[15442] = data_o[18];
  assign data_o[15506] = data_o[18];
  assign data_o[15570] = data_o[18];
  assign data_o[15634] = data_o[18];
  assign data_o[15698] = data_o[18];
  assign data_o[15762] = data_o[18];
  assign data_o[15826] = data_o[18];
  assign data_o[15890] = data_o[18];
  assign data_o[15954] = data_o[18];
  assign data_o[16018] = data_o[18];
  assign data_o[16082] = data_o[18];
  assign data_o[16146] = data_o[18];
  assign data_o[16210] = data_o[18];
  assign data_o[16274] = data_o[18];
  assign data_o[16338] = data_o[18];
  assign data_o[16402] = data_o[18];
  assign data_o[16466] = data_o[18];
  assign data_o[16530] = data_o[18];
  assign data_o[16594] = data_o[18];
  assign data_o[16658] = data_o[18];
  assign data_o[16722] = data_o[18];
  assign data_o[16786] = data_o[18];
  assign data_o[16850] = data_o[18];
  assign data_o[16914] = data_o[18];
  assign data_o[16978] = data_o[18];
  assign data_o[17042] = data_o[18];
  assign data_o[17106] = data_o[18];
  assign data_o[17170] = data_o[18];
  assign data_o[17234] = data_o[18];
  assign data_o[17298] = data_o[18];
  assign data_o[17362] = data_o[18];
  assign data_o[17426] = data_o[18];
  assign data_o[17490] = data_o[18];
  assign data_o[17554] = data_o[18];
  assign data_o[17618] = data_o[18];
  assign data_o[17682] = data_o[18];
  assign data_o[17746] = data_o[18];
  assign data_o[17810] = data_o[18];
  assign data_o[17874] = data_o[18];
  assign data_o[17938] = data_o[18];
  assign data_o[18002] = data_o[18];
  assign data_o[18066] = data_o[18];
  assign data_o[18130] = data_o[18];
  assign data_o[18194] = data_o[18];
  assign data_o[18258] = data_o[18];
  assign data_o[18322] = data_o[18];
  assign data_o[18386] = data_o[18];
  assign data_o[18450] = data_o[18];
  assign data_o[18514] = data_o[18];
  assign data_o[18578] = data_o[18];
  assign data_o[18642] = data_o[18];
  assign data_o[18706] = data_o[18];
  assign data_o[18770] = data_o[18];
  assign data_o[18834] = data_o[18];
  assign data_o[18898] = data_o[18];
  assign data_o[18962] = data_o[18];
  assign data_o[19026] = data_o[18];
  assign data_o[19090] = data_o[18];
  assign data_o[19154] = data_o[18];
  assign data_o[19218] = data_o[18];
  assign data_o[19282] = data_o[18];
  assign data_o[19346] = data_o[18];
  assign data_o[19410] = data_o[18];
  assign data_o[19474] = data_o[18];
  assign data_o[19538] = data_o[18];
  assign data_o[19602] = data_o[18];
  assign data_o[19666] = data_o[18];
  assign data_o[19730] = data_o[18];
  assign data_o[19794] = data_o[18];
  assign data_o[19858] = data_o[18];
  assign data_o[19922] = data_o[18];
  assign data_o[19986] = data_o[18];
  assign data_o[20050] = data_o[18];
  assign data_o[20114] = data_o[18];
  assign data_o[20178] = data_o[18];
  assign data_o[20242] = data_o[18];
  assign data_o[20306] = data_o[18];
  assign data_o[20370] = data_o[18];
  assign data_o[20434] = data_o[18];
  assign data_o[20498] = data_o[18];
  assign data_o[20562] = data_o[18];
  assign data_o[20626] = data_o[18];
  assign data_o[20690] = data_o[18];
  assign data_o[20754] = data_o[18];
  assign data_o[20818] = data_o[18];
  assign data_o[20882] = data_o[18];
  assign data_o[20946] = data_o[18];
  assign data_o[21010] = data_o[18];
  assign data_o[21074] = data_o[18];
  assign data_o[21138] = data_o[18];
  assign data_o[21202] = data_o[18];
  assign data_o[21266] = data_o[18];
  assign data_o[21330] = data_o[18];
  assign data_o[21394] = data_o[18];
  assign data_o[21458] = data_o[18];
  assign data_o[21522] = data_o[18];
  assign data_o[21586] = data_o[18];
  assign data_o[21650] = data_o[18];
  assign data_o[21714] = data_o[18];
  assign data_o[21778] = data_o[18];
  assign data_o[21842] = data_o[18];
  assign data_o[21906] = data_o[18];
  assign data_o[21970] = data_o[18];
  assign data_o[22034] = data_o[18];
  assign data_o[22098] = data_o[18];
  assign data_o[22162] = data_o[18];
  assign data_o[22226] = data_o[18];
  assign data_o[22290] = data_o[18];
  assign data_o[22354] = data_o[18];
  assign data_o[22418] = data_o[18];
  assign data_o[22482] = data_o[18];
  assign data_o[22546] = data_o[18];
  assign data_o[22610] = data_o[18];
  assign data_o[22674] = data_o[18];
  assign data_o[22738] = data_o[18];
  assign data_o[22802] = data_o[18];
  assign data_o[22866] = data_o[18];
  assign data_o[22930] = data_o[18];
  assign data_o[22994] = data_o[18];
  assign data_o[23058] = data_o[18];
  assign data_o[23122] = data_o[18];
  assign data_o[23186] = data_o[18];
  assign data_o[23250] = data_o[18];
  assign data_o[23314] = data_o[18];
  assign data_o[23378] = data_o[18];
  assign data_o[23442] = data_o[18];
  assign data_o[23506] = data_o[18];
  assign data_o[23570] = data_o[18];
  assign data_o[23634] = data_o[18];
  assign data_o[23698] = data_o[18];
  assign data_o[23762] = data_o[18];
  assign data_o[23826] = data_o[18];
  assign data_o[23890] = data_o[18];
  assign data_o[23954] = data_o[18];
  assign data_o[24018] = data_o[18];
  assign data_o[24082] = data_o[18];
  assign data_o[24146] = data_o[18];
  assign data_o[24210] = data_o[18];
  assign data_o[24274] = data_o[18];
  assign data_o[24338] = data_o[18];
  assign data_o[24402] = data_o[18];
  assign data_o[24466] = data_o[18];
  assign data_o[24530] = data_o[18];
  assign data_o[24594] = data_o[18];
  assign data_o[24658] = data_o[18];
  assign data_o[24722] = data_o[18];
  assign data_o[24786] = data_o[18];
  assign data_o[24850] = data_o[18];
  assign data_o[24914] = data_o[18];
  assign data_o[24978] = data_o[18];
  assign data_o[25042] = data_o[18];
  assign data_o[25106] = data_o[18];
  assign data_o[25170] = data_o[18];
  assign data_o[25234] = data_o[18];
  assign data_o[25298] = data_o[18];
  assign data_o[25362] = data_o[18];
  assign data_o[25426] = data_o[18];
  assign data_o[25490] = data_o[18];
  assign data_o[25554] = data_o[18];
  assign data_o[25618] = data_o[18];
  assign data_o[25682] = data_o[18];
  assign data_o[25746] = data_o[18];
  assign data_o[25810] = data_o[18];
  assign data_o[25874] = data_o[18];
  assign data_o[25938] = data_o[18];
  assign data_o[26002] = data_o[18];
  assign data_o[26066] = data_o[18];
  assign data_o[26130] = data_o[18];
  assign data_o[26194] = data_o[18];
  assign data_o[26258] = data_o[18];
  assign data_o[26322] = data_o[18];
  assign data_o[26386] = data_o[18];
  assign data_o[26450] = data_o[18];
  assign data_o[26514] = data_o[18];
  assign data_o[26578] = data_o[18];
  assign data_o[26642] = data_o[18];
  assign data_o[26706] = data_o[18];
  assign data_o[26770] = data_o[18];
  assign data_o[26834] = data_o[18];
  assign data_o[26898] = data_o[18];
  assign data_o[26962] = data_o[18];
  assign data_o[27026] = data_o[18];
  assign data_o[27090] = data_o[18];
  assign data_o[27154] = data_o[18];
  assign data_o[27218] = data_o[18];
  assign data_o[27282] = data_o[18];
  assign data_o[27346] = data_o[18];
  assign data_o[27410] = data_o[18];
  assign data_o[27474] = data_o[18];
  assign data_o[27538] = data_o[18];
  assign data_o[27602] = data_o[18];
  assign data_o[27666] = data_o[18];
  assign data_o[27730] = data_o[18];
  assign data_o[27794] = data_o[18];
  assign data_o[27858] = data_o[18];
  assign data_o[27922] = data_o[18];
  assign data_o[27986] = data_o[18];
  assign data_o[28050] = data_o[18];
  assign data_o[28114] = data_o[18];
  assign data_o[28178] = data_o[18];
  assign data_o[28242] = data_o[18];
  assign data_o[28306] = data_o[18];
  assign data_o[28370] = data_o[18];
  assign data_o[28434] = data_o[18];
  assign data_o[28498] = data_o[18];
  assign data_o[28562] = data_o[18];
  assign data_o[28626] = data_o[18];
  assign data_o[28690] = data_o[18];
  assign data_o[28754] = data_o[18];
  assign data_o[28818] = data_o[18];
  assign data_o[28882] = data_o[18];
  assign data_o[28946] = data_o[18];
  assign data_o[29010] = data_o[18];
  assign data_o[29074] = data_o[18];
  assign data_o[29138] = data_o[18];
  assign data_o[29202] = data_o[18];
  assign data_o[29266] = data_o[18];
  assign data_o[29330] = data_o[18];
  assign data_o[29394] = data_o[18];
  assign data_o[29458] = data_o[18];
  assign data_o[29522] = data_o[18];
  assign data_o[29586] = data_o[18];
  assign data_o[29650] = data_o[18];
  assign data_o[29714] = data_o[18];
  assign data_o[29778] = data_o[18];
  assign data_o[29842] = data_o[18];
  assign data_o[29906] = data_o[18];
  assign data_o[29970] = data_o[18];
  assign data_o[30034] = data_o[18];
  assign data_o[30098] = data_o[18];
  assign data_o[30162] = data_o[18];
  assign data_o[30226] = data_o[18];
  assign data_o[30290] = data_o[18];
  assign data_o[30354] = data_o[18];
  assign data_o[30418] = data_o[18];
  assign data_o[30482] = data_o[18];
  assign data_o[30546] = data_o[18];
  assign data_o[30610] = data_o[18];
  assign data_o[30674] = data_o[18];
  assign data_o[30738] = data_o[18];
  assign data_o[30802] = data_o[18];
  assign data_o[30866] = data_o[18];
  assign data_o[30930] = data_o[18];
  assign data_o[30994] = data_o[18];
  assign data_o[31058] = data_o[18];
  assign data_o[31122] = data_o[18];
  assign data_o[31186] = data_o[18];
  assign data_o[31250] = data_o[18];
  assign data_o[31314] = data_o[18];
  assign data_o[31378] = data_o[18];
  assign data_o[31442] = data_o[18];
  assign data_o[31506] = data_o[18];
  assign data_o[31570] = data_o[18];
  assign data_o[31634] = data_o[18];
  assign data_o[31698] = data_o[18];
  assign data_o[31762] = data_o[18];
  assign data_o[31826] = data_o[18];
  assign data_o[31890] = data_o[18];
  assign data_o[31954] = data_o[18];
  assign data_o[81] = data_o[17];
  assign data_o[145] = data_o[17];
  assign data_o[209] = data_o[17];
  assign data_o[273] = data_o[17];
  assign data_o[337] = data_o[17];
  assign data_o[401] = data_o[17];
  assign data_o[465] = data_o[17];
  assign data_o[529] = data_o[17];
  assign data_o[593] = data_o[17];
  assign data_o[657] = data_o[17];
  assign data_o[721] = data_o[17];
  assign data_o[785] = data_o[17];
  assign data_o[849] = data_o[17];
  assign data_o[913] = data_o[17];
  assign data_o[977] = data_o[17];
  assign data_o[1041] = data_o[17];
  assign data_o[1105] = data_o[17];
  assign data_o[1169] = data_o[17];
  assign data_o[1233] = data_o[17];
  assign data_o[1297] = data_o[17];
  assign data_o[1361] = data_o[17];
  assign data_o[1425] = data_o[17];
  assign data_o[1489] = data_o[17];
  assign data_o[1553] = data_o[17];
  assign data_o[1617] = data_o[17];
  assign data_o[1681] = data_o[17];
  assign data_o[1745] = data_o[17];
  assign data_o[1809] = data_o[17];
  assign data_o[1873] = data_o[17];
  assign data_o[1937] = data_o[17];
  assign data_o[2001] = data_o[17];
  assign data_o[2065] = data_o[17];
  assign data_o[2129] = data_o[17];
  assign data_o[2193] = data_o[17];
  assign data_o[2257] = data_o[17];
  assign data_o[2321] = data_o[17];
  assign data_o[2385] = data_o[17];
  assign data_o[2449] = data_o[17];
  assign data_o[2513] = data_o[17];
  assign data_o[2577] = data_o[17];
  assign data_o[2641] = data_o[17];
  assign data_o[2705] = data_o[17];
  assign data_o[2769] = data_o[17];
  assign data_o[2833] = data_o[17];
  assign data_o[2897] = data_o[17];
  assign data_o[2961] = data_o[17];
  assign data_o[3025] = data_o[17];
  assign data_o[3089] = data_o[17];
  assign data_o[3153] = data_o[17];
  assign data_o[3217] = data_o[17];
  assign data_o[3281] = data_o[17];
  assign data_o[3345] = data_o[17];
  assign data_o[3409] = data_o[17];
  assign data_o[3473] = data_o[17];
  assign data_o[3537] = data_o[17];
  assign data_o[3601] = data_o[17];
  assign data_o[3665] = data_o[17];
  assign data_o[3729] = data_o[17];
  assign data_o[3793] = data_o[17];
  assign data_o[3857] = data_o[17];
  assign data_o[3921] = data_o[17];
  assign data_o[3985] = data_o[17];
  assign data_o[4049] = data_o[17];
  assign data_o[4113] = data_o[17];
  assign data_o[4177] = data_o[17];
  assign data_o[4241] = data_o[17];
  assign data_o[4305] = data_o[17];
  assign data_o[4369] = data_o[17];
  assign data_o[4433] = data_o[17];
  assign data_o[4497] = data_o[17];
  assign data_o[4561] = data_o[17];
  assign data_o[4625] = data_o[17];
  assign data_o[4689] = data_o[17];
  assign data_o[4753] = data_o[17];
  assign data_o[4817] = data_o[17];
  assign data_o[4881] = data_o[17];
  assign data_o[4945] = data_o[17];
  assign data_o[5009] = data_o[17];
  assign data_o[5073] = data_o[17];
  assign data_o[5137] = data_o[17];
  assign data_o[5201] = data_o[17];
  assign data_o[5265] = data_o[17];
  assign data_o[5329] = data_o[17];
  assign data_o[5393] = data_o[17];
  assign data_o[5457] = data_o[17];
  assign data_o[5521] = data_o[17];
  assign data_o[5585] = data_o[17];
  assign data_o[5649] = data_o[17];
  assign data_o[5713] = data_o[17];
  assign data_o[5777] = data_o[17];
  assign data_o[5841] = data_o[17];
  assign data_o[5905] = data_o[17];
  assign data_o[5969] = data_o[17];
  assign data_o[6033] = data_o[17];
  assign data_o[6097] = data_o[17];
  assign data_o[6161] = data_o[17];
  assign data_o[6225] = data_o[17];
  assign data_o[6289] = data_o[17];
  assign data_o[6353] = data_o[17];
  assign data_o[6417] = data_o[17];
  assign data_o[6481] = data_o[17];
  assign data_o[6545] = data_o[17];
  assign data_o[6609] = data_o[17];
  assign data_o[6673] = data_o[17];
  assign data_o[6737] = data_o[17];
  assign data_o[6801] = data_o[17];
  assign data_o[6865] = data_o[17];
  assign data_o[6929] = data_o[17];
  assign data_o[6993] = data_o[17];
  assign data_o[7057] = data_o[17];
  assign data_o[7121] = data_o[17];
  assign data_o[7185] = data_o[17];
  assign data_o[7249] = data_o[17];
  assign data_o[7313] = data_o[17];
  assign data_o[7377] = data_o[17];
  assign data_o[7441] = data_o[17];
  assign data_o[7505] = data_o[17];
  assign data_o[7569] = data_o[17];
  assign data_o[7633] = data_o[17];
  assign data_o[7697] = data_o[17];
  assign data_o[7761] = data_o[17];
  assign data_o[7825] = data_o[17];
  assign data_o[7889] = data_o[17];
  assign data_o[7953] = data_o[17];
  assign data_o[8017] = data_o[17];
  assign data_o[8081] = data_o[17];
  assign data_o[8145] = data_o[17];
  assign data_o[8209] = data_o[17];
  assign data_o[8273] = data_o[17];
  assign data_o[8337] = data_o[17];
  assign data_o[8401] = data_o[17];
  assign data_o[8465] = data_o[17];
  assign data_o[8529] = data_o[17];
  assign data_o[8593] = data_o[17];
  assign data_o[8657] = data_o[17];
  assign data_o[8721] = data_o[17];
  assign data_o[8785] = data_o[17];
  assign data_o[8849] = data_o[17];
  assign data_o[8913] = data_o[17];
  assign data_o[8977] = data_o[17];
  assign data_o[9041] = data_o[17];
  assign data_o[9105] = data_o[17];
  assign data_o[9169] = data_o[17];
  assign data_o[9233] = data_o[17];
  assign data_o[9297] = data_o[17];
  assign data_o[9361] = data_o[17];
  assign data_o[9425] = data_o[17];
  assign data_o[9489] = data_o[17];
  assign data_o[9553] = data_o[17];
  assign data_o[9617] = data_o[17];
  assign data_o[9681] = data_o[17];
  assign data_o[9745] = data_o[17];
  assign data_o[9809] = data_o[17];
  assign data_o[9873] = data_o[17];
  assign data_o[9937] = data_o[17];
  assign data_o[10001] = data_o[17];
  assign data_o[10065] = data_o[17];
  assign data_o[10129] = data_o[17];
  assign data_o[10193] = data_o[17];
  assign data_o[10257] = data_o[17];
  assign data_o[10321] = data_o[17];
  assign data_o[10385] = data_o[17];
  assign data_o[10449] = data_o[17];
  assign data_o[10513] = data_o[17];
  assign data_o[10577] = data_o[17];
  assign data_o[10641] = data_o[17];
  assign data_o[10705] = data_o[17];
  assign data_o[10769] = data_o[17];
  assign data_o[10833] = data_o[17];
  assign data_o[10897] = data_o[17];
  assign data_o[10961] = data_o[17];
  assign data_o[11025] = data_o[17];
  assign data_o[11089] = data_o[17];
  assign data_o[11153] = data_o[17];
  assign data_o[11217] = data_o[17];
  assign data_o[11281] = data_o[17];
  assign data_o[11345] = data_o[17];
  assign data_o[11409] = data_o[17];
  assign data_o[11473] = data_o[17];
  assign data_o[11537] = data_o[17];
  assign data_o[11601] = data_o[17];
  assign data_o[11665] = data_o[17];
  assign data_o[11729] = data_o[17];
  assign data_o[11793] = data_o[17];
  assign data_o[11857] = data_o[17];
  assign data_o[11921] = data_o[17];
  assign data_o[11985] = data_o[17];
  assign data_o[12049] = data_o[17];
  assign data_o[12113] = data_o[17];
  assign data_o[12177] = data_o[17];
  assign data_o[12241] = data_o[17];
  assign data_o[12305] = data_o[17];
  assign data_o[12369] = data_o[17];
  assign data_o[12433] = data_o[17];
  assign data_o[12497] = data_o[17];
  assign data_o[12561] = data_o[17];
  assign data_o[12625] = data_o[17];
  assign data_o[12689] = data_o[17];
  assign data_o[12753] = data_o[17];
  assign data_o[12817] = data_o[17];
  assign data_o[12881] = data_o[17];
  assign data_o[12945] = data_o[17];
  assign data_o[13009] = data_o[17];
  assign data_o[13073] = data_o[17];
  assign data_o[13137] = data_o[17];
  assign data_o[13201] = data_o[17];
  assign data_o[13265] = data_o[17];
  assign data_o[13329] = data_o[17];
  assign data_o[13393] = data_o[17];
  assign data_o[13457] = data_o[17];
  assign data_o[13521] = data_o[17];
  assign data_o[13585] = data_o[17];
  assign data_o[13649] = data_o[17];
  assign data_o[13713] = data_o[17];
  assign data_o[13777] = data_o[17];
  assign data_o[13841] = data_o[17];
  assign data_o[13905] = data_o[17];
  assign data_o[13969] = data_o[17];
  assign data_o[14033] = data_o[17];
  assign data_o[14097] = data_o[17];
  assign data_o[14161] = data_o[17];
  assign data_o[14225] = data_o[17];
  assign data_o[14289] = data_o[17];
  assign data_o[14353] = data_o[17];
  assign data_o[14417] = data_o[17];
  assign data_o[14481] = data_o[17];
  assign data_o[14545] = data_o[17];
  assign data_o[14609] = data_o[17];
  assign data_o[14673] = data_o[17];
  assign data_o[14737] = data_o[17];
  assign data_o[14801] = data_o[17];
  assign data_o[14865] = data_o[17];
  assign data_o[14929] = data_o[17];
  assign data_o[14993] = data_o[17];
  assign data_o[15057] = data_o[17];
  assign data_o[15121] = data_o[17];
  assign data_o[15185] = data_o[17];
  assign data_o[15249] = data_o[17];
  assign data_o[15313] = data_o[17];
  assign data_o[15377] = data_o[17];
  assign data_o[15441] = data_o[17];
  assign data_o[15505] = data_o[17];
  assign data_o[15569] = data_o[17];
  assign data_o[15633] = data_o[17];
  assign data_o[15697] = data_o[17];
  assign data_o[15761] = data_o[17];
  assign data_o[15825] = data_o[17];
  assign data_o[15889] = data_o[17];
  assign data_o[15953] = data_o[17];
  assign data_o[16017] = data_o[17];
  assign data_o[16081] = data_o[17];
  assign data_o[16145] = data_o[17];
  assign data_o[16209] = data_o[17];
  assign data_o[16273] = data_o[17];
  assign data_o[16337] = data_o[17];
  assign data_o[16401] = data_o[17];
  assign data_o[16465] = data_o[17];
  assign data_o[16529] = data_o[17];
  assign data_o[16593] = data_o[17];
  assign data_o[16657] = data_o[17];
  assign data_o[16721] = data_o[17];
  assign data_o[16785] = data_o[17];
  assign data_o[16849] = data_o[17];
  assign data_o[16913] = data_o[17];
  assign data_o[16977] = data_o[17];
  assign data_o[17041] = data_o[17];
  assign data_o[17105] = data_o[17];
  assign data_o[17169] = data_o[17];
  assign data_o[17233] = data_o[17];
  assign data_o[17297] = data_o[17];
  assign data_o[17361] = data_o[17];
  assign data_o[17425] = data_o[17];
  assign data_o[17489] = data_o[17];
  assign data_o[17553] = data_o[17];
  assign data_o[17617] = data_o[17];
  assign data_o[17681] = data_o[17];
  assign data_o[17745] = data_o[17];
  assign data_o[17809] = data_o[17];
  assign data_o[17873] = data_o[17];
  assign data_o[17937] = data_o[17];
  assign data_o[18001] = data_o[17];
  assign data_o[18065] = data_o[17];
  assign data_o[18129] = data_o[17];
  assign data_o[18193] = data_o[17];
  assign data_o[18257] = data_o[17];
  assign data_o[18321] = data_o[17];
  assign data_o[18385] = data_o[17];
  assign data_o[18449] = data_o[17];
  assign data_o[18513] = data_o[17];
  assign data_o[18577] = data_o[17];
  assign data_o[18641] = data_o[17];
  assign data_o[18705] = data_o[17];
  assign data_o[18769] = data_o[17];
  assign data_o[18833] = data_o[17];
  assign data_o[18897] = data_o[17];
  assign data_o[18961] = data_o[17];
  assign data_o[19025] = data_o[17];
  assign data_o[19089] = data_o[17];
  assign data_o[19153] = data_o[17];
  assign data_o[19217] = data_o[17];
  assign data_o[19281] = data_o[17];
  assign data_o[19345] = data_o[17];
  assign data_o[19409] = data_o[17];
  assign data_o[19473] = data_o[17];
  assign data_o[19537] = data_o[17];
  assign data_o[19601] = data_o[17];
  assign data_o[19665] = data_o[17];
  assign data_o[19729] = data_o[17];
  assign data_o[19793] = data_o[17];
  assign data_o[19857] = data_o[17];
  assign data_o[19921] = data_o[17];
  assign data_o[19985] = data_o[17];
  assign data_o[20049] = data_o[17];
  assign data_o[20113] = data_o[17];
  assign data_o[20177] = data_o[17];
  assign data_o[20241] = data_o[17];
  assign data_o[20305] = data_o[17];
  assign data_o[20369] = data_o[17];
  assign data_o[20433] = data_o[17];
  assign data_o[20497] = data_o[17];
  assign data_o[20561] = data_o[17];
  assign data_o[20625] = data_o[17];
  assign data_o[20689] = data_o[17];
  assign data_o[20753] = data_o[17];
  assign data_o[20817] = data_o[17];
  assign data_o[20881] = data_o[17];
  assign data_o[20945] = data_o[17];
  assign data_o[21009] = data_o[17];
  assign data_o[21073] = data_o[17];
  assign data_o[21137] = data_o[17];
  assign data_o[21201] = data_o[17];
  assign data_o[21265] = data_o[17];
  assign data_o[21329] = data_o[17];
  assign data_o[21393] = data_o[17];
  assign data_o[21457] = data_o[17];
  assign data_o[21521] = data_o[17];
  assign data_o[21585] = data_o[17];
  assign data_o[21649] = data_o[17];
  assign data_o[21713] = data_o[17];
  assign data_o[21777] = data_o[17];
  assign data_o[21841] = data_o[17];
  assign data_o[21905] = data_o[17];
  assign data_o[21969] = data_o[17];
  assign data_o[22033] = data_o[17];
  assign data_o[22097] = data_o[17];
  assign data_o[22161] = data_o[17];
  assign data_o[22225] = data_o[17];
  assign data_o[22289] = data_o[17];
  assign data_o[22353] = data_o[17];
  assign data_o[22417] = data_o[17];
  assign data_o[22481] = data_o[17];
  assign data_o[22545] = data_o[17];
  assign data_o[22609] = data_o[17];
  assign data_o[22673] = data_o[17];
  assign data_o[22737] = data_o[17];
  assign data_o[22801] = data_o[17];
  assign data_o[22865] = data_o[17];
  assign data_o[22929] = data_o[17];
  assign data_o[22993] = data_o[17];
  assign data_o[23057] = data_o[17];
  assign data_o[23121] = data_o[17];
  assign data_o[23185] = data_o[17];
  assign data_o[23249] = data_o[17];
  assign data_o[23313] = data_o[17];
  assign data_o[23377] = data_o[17];
  assign data_o[23441] = data_o[17];
  assign data_o[23505] = data_o[17];
  assign data_o[23569] = data_o[17];
  assign data_o[23633] = data_o[17];
  assign data_o[23697] = data_o[17];
  assign data_o[23761] = data_o[17];
  assign data_o[23825] = data_o[17];
  assign data_o[23889] = data_o[17];
  assign data_o[23953] = data_o[17];
  assign data_o[24017] = data_o[17];
  assign data_o[24081] = data_o[17];
  assign data_o[24145] = data_o[17];
  assign data_o[24209] = data_o[17];
  assign data_o[24273] = data_o[17];
  assign data_o[24337] = data_o[17];
  assign data_o[24401] = data_o[17];
  assign data_o[24465] = data_o[17];
  assign data_o[24529] = data_o[17];
  assign data_o[24593] = data_o[17];
  assign data_o[24657] = data_o[17];
  assign data_o[24721] = data_o[17];
  assign data_o[24785] = data_o[17];
  assign data_o[24849] = data_o[17];
  assign data_o[24913] = data_o[17];
  assign data_o[24977] = data_o[17];
  assign data_o[25041] = data_o[17];
  assign data_o[25105] = data_o[17];
  assign data_o[25169] = data_o[17];
  assign data_o[25233] = data_o[17];
  assign data_o[25297] = data_o[17];
  assign data_o[25361] = data_o[17];
  assign data_o[25425] = data_o[17];
  assign data_o[25489] = data_o[17];
  assign data_o[25553] = data_o[17];
  assign data_o[25617] = data_o[17];
  assign data_o[25681] = data_o[17];
  assign data_o[25745] = data_o[17];
  assign data_o[25809] = data_o[17];
  assign data_o[25873] = data_o[17];
  assign data_o[25937] = data_o[17];
  assign data_o[26001] = data_o[17];
  assign data_o[26065] = data_o[17];
  assign data_o[26129] = data_o[17];
  assign data_o[26193] = data_o[17];
  assign data_o[26257] = data_o[17];
  assign data_o[26321] = data_o[17];
  assign data_o[26385] = data_o[17];
  assign data_o[26449] = data_o[17];
  assign data_o[26513] = data_o[17];
  assign data_o[26577] = data_o[17];
  assign data_o[26641] = data_o[17];
  assign data_o[26705] = data_o[17];
  assign data_o[26769] = data_o[17];
  assign data_o[26833] = data_o[17];
  assign data_o[26897] = data_o[17];
  assign data_o[26961] = data_o[17];
  assign data_o[27025] = data_o[17];
  assign data_o[27089] = data_o[17];
  assign data_o[27153] = data_o[17];
  assign data_o[27217] = data_o[17];
  assign data_o[27281] = data_o[17];
  assign data_o[27345] = data_o[17];
  assign data_o[27409] = data_o[17];
  assign data_o[27473] = data_o[17];
  assign data_o[27537] = data_o[17];
  assign data_o[27601] = data_o[17];
  assign data_o[27665] = data_o[17];
  assign data_o[27729] = data_o[17];
  assign data_o[27793] = data_o[17];
  assign data_o[27857] = data_o[17];
  assign data_o[27921] = data_o[17];
  assign data_o[27985] = data_o[17];
  assign data_o[28049] = data_o[17];
  assign data_o[28113] = data_o[17];
  assign data_o[28177] = data_o[17];
  assign data_o[28241] = data_o[17];
  assign data_o[28305] = data_o[17];
  assign data_o[28369] = data_o[17];
  assign data_o[28433] = data_o[17];
  assign data_o[28497] = data_o[17];
  assign data_o[28561] = data_o[17];
  assign data_o[28625] = data_o[17];
  assign data_o[28689] = data_o[17];
  assign data_o[28753] = data_o[17];
  assign data_o[28817] = data_o[17];
  assign data_o[28881] = data_o[17];
  assign data_o[28945] = data_o[17];
  assign data_o[29009] = data_o[17];
  assign data_o[29073] = data_o[17];
  assign data_o[29137] = data_o[17];
  assign data_o[29201] = data_o[17];
  assign data_o[29265] = data_o[17];
  assign data_o[29329] = data_o[17];
  assign data_o[29393] = data_o[17];
  assign data_o[29457] = data_o[17];
  assign data_o[29521] = data_o[17];
  assign data_o[29585] = data_o[17];
  assign data_o[29649] = data_o[17];
  assign data_o[29713] = data_o[17];
  assign data_o[29777] = data_o[17];
  assign data_o[29841] = data_o[17];
  assign data_o[29905] = data_o[17];
  assign data_o[29969] = data_o[17];
  assign data_o[30033] = data_o[17];
  assign data_o[30097] = data_o[17];
  assign data_o[30161] = data_o[17];
  assign data_o[30225] = data_o[17];
  assign data_o[30289] = data_o[17];
  assign data_o[30353] = data_o[17];
  assign data_o[30417] = data_o[17];
  assign data_o[30481] = data_o[17];
  assign data_o[30545] = data_o[17];
  assign data_o[30609] = data_o[17];
  assign data_o[30673] = data_o[17];
  assign data_o[30737] = data_o[17];
  assign data_o[30801] = data_o[17];
  assign data_o[30865] = data_o[17];
  assign data_o[30929] = data_o[17];
  assign data_o[30993] = data_o[17];
  assign data_o[31057] = data_o[17];
  assign data_o[31121] = data_o[17];
  assign data_o[31185] = data_o[17];
  assign data_o[31249] = data_o[17];
  assign data_o[31313] = data_o[17];
  assign data_o[31377] = data_o[17];
  assign data_o[31441] = data_o[17];
  assign data_o[31505] = data_o[17];
  assign data_o[31569] = data_o[17];
  assign data_o[31633] = data_o[17];
  assign data_o[31697] = data_o[17];
  assign data_o[31761] = data_o[17];
  assign data_o[31825] = data_o[17];
  assign data_o[31889] = data_o[17];
  assign data_o[31953] = data_o[17];
  assign data_o[80] = data_o[16];
  assign data_o[144] = data_o[16];
  assign data_o[208] = data_o[16];
  assign data_o[272] = data_o[16];
  assign data_o[336] = data_o[16];
  assign data_o[400] = data_o[16];
  assign data_o[464] = data_o[16];
  assign data_o[528] = data_o[16];
  assign data_o[592] = data_o[16];
  assign data_o[656] = data_o[16];
  assign data_o[720] = data_o[16];
  assign data_o[784] = data_o[16];
  assign data_o[848] = data_o[16];
  assign data_o[912] = data_o[16];
  assign data_o[976] = data_o[16];
  assign data_o[1040] = data_o[16];
  assign data_o[1104] = data_o[16];
  assign data_o[1168] = data_o[16];
  assign data_o[1232] = data_o[16];
  assign data_o[1296] = data_o[16];
  assign data_o[1360] = data_o[16];
  assign data_o[1424] = data_o[16];
  assign data_o[1488] = data_o[16];
  assign data_o[1552] = data_o[16];
  assign data_o[1616] = data_o[16];
  assign data_o[1680] = data_o[16];
  assign data_o[1744] = data_o[16];
  assign data_o[1808] = data_o[16];
  assign data_o[1872] = data_o[16];
  assign data_o[1936] = data_o[16];
  assign data_o[2000] = data_o[16];
  assign data_o[2064] = data_o[16];
  assign data_o[2128] = data_o[16];
  assign data_o[2192] = data_o[16];
  assign data_o[2256] = data_o[16];
  assign data_o[2320] = data_o[16];
  assign data_o[2384] = data_o[16];
  assign data_o[2448] = data_o[16];
  assign data_o[2512] = data_o[16];
  assign data_o[2576] = data_o[16];
  assign data_o[2640] = data_o[16];
  assign data_o[2704] = data_o[16];
  assign data_o[2768] = data_o[16];
  assign data_o[2832] = data_o[16];
  assign data_o[2896] = data_o[16];
  assign data_o[2960] = data_o[16];
  assign data_o[3024] = data_o[16];
  assign data_o[3088] = data_o[16];
  assign data_o[3152] = data_o[16];
  assign data_o[3216] = data_o[16];
  assign data_o[3280] = data_o[16];
  assign data_o[3344] = data_o[16];
  assign data_o[3408] = data_o[16];
  assign data_o[3472] = data_o[16];
  assign data_o[3536] = data_o[16];
  assign data_o[3600] = data_o[16];
  assign data_o[3664] = data_o[16];
  assign data_o[3728] = data_o[16];
  assign data_o[3792] = data_o[16];
  assign data_o[3856] = data_o[16];
  assign data_o[3920] = data_o[16];
  assign data_o[3984] = data_o[16];
  assign data_o[4048] = data_o[16];
  assign data_o[4112] = data_o[16];
  assign data_o[4176] = data_o[16];
  assign data_o[4240] = data_o[16];
  assign data_o[4304] = data_o[16];
  assign data_o[4368] = data_o[16];
  assign data_o[4432] = data_o[16];
  assign data_o[4496] = data_o[16];
  assign data_o[4560] = data_o[16];
  assign data_o[4624] = data_o[16];
  assign data_o[4688] = data_o[16];
  assign data_o[4752] = data_o[16];
  assign data_o[4816] = data_o[16];
  assign data_o[4880] = data_o[16];
  assign data_o[4944] = data_o[16];
  assign data_o[5008] = data_o[16];
  assign data_o[5072] = data_o[16];
  assign data_o[5136] = data_o[16];
  assign data_o[5200] = data_o[16];
  assign data_o[5264] = data_o[16];
  assign data_o[5328] = data_o[16];
  assign data_o[5392] = data_o[16];
  assign data_o[5456] = data_o[16];
  assign data_o[5520] = data_o[16];
  assign data_o[5584] = data_o[16];
  assign data_o[5648] = data_o[16];
  assign data_o[5712] = data_o[16];
  assign data_o[5776] = data_o[16];
  assign data_o[5840] = data_o[16];
  assign data_o[5904] = data_o[16];
  assign data_o[5968] = data_o[16];
  assign data_o[6032] = data_o[16];
  assign data_o[6096] = data_o[16];
  assign data_o[6160] = data_o[16];
  assign data_o[6224] = data_o[16];
  assign data_o[6288] = data_o[16];
  assign data_o[6352] = data_o[16];
  assign data_o[6416] = data_o[16];
  assign data_o[6480] = data_o[16];
  assign data_o[6544] = data_o[16];
  assign data_o[6608] = data_o[16];
  assign data_o[6672] = data_o[16];
  assign data_o[6736] = data_o[16];
  assign data_o[6800] = data_o[16];
  assign data_o[6864] = data_o[16];
  assign data_o[6928] = data_o[16];
  assign data_o[6992] = data_o[16];
  assign data_o[7056] = data_o[16];
  assign data_o[7120] = data_o[16];
  assign data_o[7184] = data_o[16];
  assign data_o[7248] = data_o[16];
  assign data_o[7312] = data_o[16];
  assign data_o[7376] = data_o[16];
  assign data_o[7440] = data_o[16];
  assign data_o[7504] = data_o[16];
  assign data_o[7568] = data_o[16];
  assign data_o[7632] = data_o[16];
  assign data_o[7696] = data_o[16];
  assign data_o[7760] = data_o[16];
  assign data_o[7824] = data_o[16];
  assign data_o[7888] = data_o[16];
  assign data_o[7952] = data_o[16];
  assign data_o[8016] = data_o[16];
  assign data_o[8080] = data_o[16];
  assign data_o[8144] = data_o[16];
  assign data_o[8208] = data_o[16];
  assign data_o[8272] = data_o[16];
  assign data_o[8336] = data_o[16];
  assign data_o[8400] = data_o[16];
  assign data_o[8464] = data_o[16];
  assign data_o[8528] = data_o[16];
  assign data_o[8592] = data_o[16];
  assign data_o[8656] = data_o[16];
  assign data_o[8720] = data_o[16];
  assign data_o[8784] = data_o[16];
  assign data_o[8848] = data_o[16];
  assign data_o[8912] = data_o[16];
  assign data_o[8976] = data_o[16];
  assign data_o[9040] = data_o[16];
  assign data_o[9104] = data_o[16];
  assign data_o[9168] = data_o[16];
  assign data_o[9232] = data_o[16];
  assign data_o[9296] = data_o[16];
  assign data_o[9360] = data_o[16];
  assign data_o[9424] = data_o[16];
  assign data_o[9488] = data_o[16];
  assign data_o[9552] = data_o[16];
  assign data_o[9616] = data_o[16];
  assign data_o[9680] = data_o[16];
  assign data_o[9744] = data_o[16];
  assign data_o[9808] = data_o[16];
  assign data_o[9872] = data_o[16];
  assign data_o[9936] = data_o[16];
  assign data_o[10000] = data_o[16];
  assign data_o[10064] = data_o[16];
  assign data_o[10128] = data_o[16];
  assign data_o[10192] = data_o[16];
  assign data_o[10256] = data_o[16];
  assign data_o[10320] = data_o[16];
  assign data_o[10384] = data_o[16];
  assign data_o[10448] = data_o[16];
  assign data_o[10512] = data_o[16];
  assign data_o[10576] = data_o[16];
  assign data_o[10640] = data_o[16];
  assign data_o[10704] = data_o[16];
  assign data_o[10768] = data_o[16];
  assign data_o[10832] = data_o[16];
  assign data_o[10896] = data_o[16];
  assign data_o[10960] = data_o[16];
  assign data_o[11024] = data_o[16];
  assign data_o[11088] = data_o[16];
  assign data_o[11152] = data_o[16];
  assign data_o[11216] = data_o[16];
  assign data_o[11280] = data_o[16];
  assign data_o[11344] = data_o[16];
  assign data_o[11408] = data_o[16];
  assign data_o[11472] = data_o[16];
  assign data_o[11536] = data_o[16];
  assign data_o[11600] = data_o[16];
  assign data_o[11664] = data_o[16];
  assign data_o[11728] = data_o[16];
  assign data_o[11792] = data_o[16];
  assign data_o[11856] = data_o[16];
  assign data_o[11920] = data_o[16];
  assign data_o[11984] = data_o[16];
  assign data_o[12048] = data_o[16];
  assign data_o[12112] = data_o[16];
  assign data_o[12176] = data_o[16];
  assign data_o[12240] = data_o[16];
  assign data_o[12304] = data_o[16];
  assign data_o[12368] = data_o[16];
  assign data_o[12432] = data_o[16];
  assign data_o[12496] = data_o[16];
  assign data_o[12560] = data_o[16];
  assign data_o[12624] = data_o[16];
  assign data_o[12688] = data_o[16];
  assign data_o[12752] = data_o[16];
  assign data_o[12816] = data_o[16];
  assign data_o[12880] = data_o[16];
  assign data_o[12944] = data_o[16];
  assign data_o[13008] = data_o[16];
  assign data_o[13072] = data_o[16];
  assign data_o[13136] = data_o[16];
  assign data_o[13200] = data_o[16];
  assign data_o[13264] = data_o[16];
  assign data_o[13328] = data_o[16];
  assign data_o[13392] = data_o[16];
  assign data_o[13456] = data_o[16];
  assign data_o[13520] = data_o[16];
  assign data_o[13584] = data_o[16];
  assign data_o[13648] = data_o[16];
  assign data_o[13712] = data_o[16];
  assign data_o[13776] = data_o[16];
  assign data_o[13840] = data_o[16];
  assign data_o[13904] = data_o[16];
  assign data_o[13968] = data_o[16];
  assign data_o[14032] = data_o[16];
  assign data_o[14096] = data_o[16];
  assign data_o[14160] = data_o[16];
  assign data_o[14224] = data_o[16];
  assign data_o[14288] = data_o[16];
  assign data_o[14352] = data_o[16];
  assign data_o[14416] = data_o[16];
  assign data_o[14480] = data_o[16];
  assign data_o[14544] = data_o[16];
  assign data_o[14608] = data_o[16];
  assign data_o[14672] = data_o[16];
  assign data_o[14736] = data_o[16];
  assign data_o[14800] = data_o[16];
  assign data_o[14864] = data_o[16];
  assign data_o[14928] = data_o[16];
  assign data_o[14992] = data_o[16];
  assign data_o[15056] = data_o[16];
  assign data_o[15120] = data_o[16];
  assign data_o[15184] = data_o[16];
  assign data_o[15248] = data_o[16];
  assign data_o[15312] = data_o[16];
  assign data_o[15376] = data_o[16];
  assign data_o[15440] = data_o[16];
  assign data_o[15504] = data_o[16];
  assign data_o[15568] = data_o[16];
  assign data_o[15632] = data_o[16];
  assign data_o[15696] = data_o[16];
  assign data_o[15760] = data_o[16];
  assign data_o[15824] = data_o[16];
  assign data_o[15888] = data_o[16];
  assign data_o[15952] = data_o[16];
  assign data_o[16016] = data_o[16];
  assign data_o[16080] = data_o[16];
  assign data_o[16144] = data_o[16];
  assign data_o[16208] = data_o[16];
  assign data_o[16272] = data_o[16];
  assign data_o[16336] = data_o[16];
  assign data_o[16400] = data_o[16];
  assign data_o[16464] = data_o[16];
  assign data_o[16528] = data_o[16];
  assign data_o[16592] = data_o[16];
  assign data_o[16656] = data_o[16];
  assign data_o[16720] = data_o[16];
  assign data_o[16784] = data_o[16];
  assign data_o[16848] = data_o[16];
  assign data_o[16912] = data_o[16];
  assign data_o[16976] = data_o[16];
  assign data_o[17040] = data_o[16];
  assign data_o[17104] = data_o[16];
  assign data_o[17168] = data_o[16];
  assign data_o[17232] = data_o[16];
  assign data_o[17296] = data_o[16];
  assign data_o[17360] = data_o[16];
  assign data_o[17424] = data_o[16];
  assign data_o[17488] = data_o[16];
  assign data_o[17552] = data_o[16];
  assign data_o[17616] = data_o[16];
  assign data_o[17680] = data_o[16];
  assign data_o[17744] = data_o[16];
  assign data_o[17808] = data_o[16];
  assign data_o[17872] = data_o[16];
  assign data_o[17936] = data_o[16];
  assign data_o[18000] = data_o[16];
  assign data_o[18064] = data_o[16];
  assign data_o[18128] = data_o[16];
  assign data_o[18192] = data_o[16];
  assign data_o[18256] = data_o[16];
  assign data_o[18320] = data_o[16];
  assign data_o[18384] = data_o[16];
  assign data_o[18448] = data_o[16];
  assign data_o[18512] = data_o[16];
  assign data_o[18576] = data_o[16];
  assign data_o[18640] = data_o[16];
  assign data_o[18704] = data_o[16];
  assign data_o[18768] = data_o[16];
  assign data_o[18832] = data_o[16];
  assign data_o[18896] = data_o[16];
  assign data_o[18960] = data_o[16];
  assign data_o[19024] = data_o[16];
  assign data_o[19088] = data_o[16];
  assign data_o[19152] = data_o[16];
  assign data_o[19216] = data_o[16];
  assign data_o[19280] = data_o[16];
  assign data_o[19344] = data_o[16];
  assign data_o[19408] = data_o[16];
  assign data_o[19472] = data_o[16];
  assign data_o[19536] = data_o[16];
  assign data_o[19600] = data_o[16];
  assign data_o[19664] = data_o[16];
  assign data_o[19728] = data_o[16];
  assign data_o[19792] = data_o[16];
  assign data_o[19856] = data_o[16];
  assign data_o[19920] = data_o[16];
  assign data_o[19984] = data_o[16];
  assign data_o[20048] = data_o[16];
  assign data_o[20112] = data_o[16];
  assign data_o[20176] = data_o[16];
  assign data_o[20240] = data_o[16];
  assign data_o[20304] = data_o[16];
  assign data_o[20368] = data_o[16];
  assign data_o[20432] = data_o[16];
  assign data_o[20496] = data_o[16];
  assign data_o[20560] = data_o[16];
  assign data_o[20624] = data_o[16];
  assign data_o[20688] = data_o[16];
  assign data_o[20752] = data_o[16];
  assign data_o[20816] = data_o[16];
  assign data_o[20880] = data_o[16];
  assign data_o[20944] = data_o[16];
  assign data_o[21008] = data_o[16];
  assign data_o[21072] = data_o[16];
  assign data_o[21136] = data_o[16];
  assign data_o[21200] = data_o[16];
  assign data_o[21264] = data_o[16];
  assign data_o[21328] = data_o[16];
  assign data_o[21392] = data_o[16];
  assign data_o[21456] = data_o[16];
  assign data_o[21520] = data_o[16];
  assign data_o[21584] = data_o[16];
  assign data_o[21648] = data_o[16];
  assign data_o[21712] = data_o[16];
  assign data_o[21776] = data_o[16];
  assign data_o[21840] = data_o[16];
  assign data_o[21904] = data_o[16];
  assign data_o[21968] = data_o[16];
  assign data_o[22032] = data_o[16];
  assign data_o[22096] = data_o[16];
  assign data_o[22160] = data_o[16];
  assign data_o[22224] = data_o[16];
  assign data_o[22288] = data_o[16];
  assign data_o[22352] = data_o[16];
  assign data_o[22416] = data_o[16];
  assign data_o[22480] = data_o[16];
  assign data_o[22544] = data_o[16];
  assign data_o[22608] = data_o[16];
  assign data_o[22672] = data_o[16];
  assign data_o[22736] = data_o[16];
  assign data_o[22800] = data_o[16];
  assign data_o[22864] = data_o[16];
  assign data_o[22928] = data_o[16];
  assign data_o[22992] = data_o[16];
  assign data_o[23056] = data_o[16];
  assign data_o[23120] = data_o[16];
  assign data_o[23184] = data_o[16];
  assign data_o[23248] = data_o[16];
  assign data_o[23312] = data_o[16];
  assign data_o[23376] = data_o[16];
  assign data_o[23440] = data_o[16];
  assign data_o[23504] = data_o[16];
  assign data_o[23568] = data_o[16];
  assign data_o[23632] = data_o[16];
  assign data_o[23696] = data_o[16];
  assign data_o[23760] = data_o[16];
  assign data_o[23824] = data_o[16];
  assign data_o[23888] = data_o[16];
  assign data_o[23952] = data_o[16];
  assign data_o[24016] = data_o[16];
  assign data_o[24080] = data_o[16];
  assign data_o[24144] = data_o[16];
  assign data_o[24208] = data_o[16];
  assign data_o[24272] = data_o[16];
  assign data_o[24336] = data_o[16];
  assign data_o[24400] = data_o[16];
  assign data_o[24464] = data_o[16];
  assign data_o[24528] = data_o[16];
  assign data_o[24592] = data_o[16];
  assign data_o[24656] = data_o[16];
  assign data_o[24720] = data_o[16];
  assign data_o[24784] = data_o[16];
  assign data_o[24848] = data_o[16];
  assign data_o[24912] = data_o[16];
  assign data_o[24976] = data_o[16];
  assign data_o[25040] = data_o[16];
  assign data_o[25104] = data_o[16];
  assign data_o[25168] = data_o[16];
  assign data_o[25232] = data_o[16];
  assign data_o[25296] = data_o[16];
  assign data_o[25360] = data_o[16];
  assign data_o[25424] = data_o[16];
  assign data_o[25488] = data_o[16];
  assign data_o[25552] = data_o[16];
  assign data_o[25616] = data_o[16];
  assign data_o[25680] = data_o[16];
  assign data_o[25744] = data_o[16];
  assign data_o[25808] = data_o[16];
  assign data_o[25872] = data_o[16];
  assign data_o[25936] = data_o[16];
  assign data_o[26000] = data_o[16];
  assign data_o[26064] = data_o[16];
  assign data_o[26128] = data_o[16];
  assign data_o[26192] = data_o[16];
  assign data_o[26256] = data_o[16];
  assign data_o[26320] = data_o[16];
  assign data_o[26384] = data_o[16];
  assign data_o[26448] = data_o[16];
  assign data_o[26512] = data_o[16];
  assign data_o[26576] = data_o[16];
  assign data_o[26640] = data_o[16];
  assign data_o[26704] = data_o[16];
  assign data_o[26768] = data_o[16];
  assign data_o[26832] = data_o[16];
  assign data_o[26896] = data_o[16];
  assign data_o[26960] = data_o[16];
  assign data_o[27024] = data_o[16];
  assign data_o[27088] = data_o[16];
  assign data_o[27152] = data_o[16];
  assign data_o[27216] = data_o[16];
  assign data_o[27280] = data_o[16];
  assign data_o[27344] = data_o[16];
  assign data_o[27408] = data_o[16];
  assign data_o[27472] = data_o[16];
  assign data_o[27536] = data_o[16];
  assign data_o[27600] = data_o[16];
  assign data_o[27664] = data_o[16];
  assign data_o[27728] = data_o[16];
  assign data_o[27792] = data_o[16];
  assign data_o[27856] = data_o[16];
  assign data_o[27920] = data_o[16];
  assign data_o[27984] = data_o[16];
  assign data_o[28048] = data_o[16];
  assign data_o[28112] = data_o[16];
  assign data_o[28176] = data_o[16];
  assign data_o[28240] = data_o[16];
  assign data_o[28304] = data_o[16];
  assign data_o[28368] = data_o[16];
  assign data_o[28432] = data_o[16];
  assign data_o[28496] = data_o[16];
  assign data_o[28560] = data_o[16];
  assign data_o[28624] = data_o[16];
  assign data_o[28688] = data_o[16];
  assign data_o[28752] = data_o[16];
  assign data_o[28816] = data_o[16];
  assign data_o[28880] = data_o[16];
  assign data_o[28944] = data_o[16];
  assign data_o[29008] = data_o[16];
  assign data_o[29072] = data_o[16];
  assign data_o[29136] = data_o[16];
  assign data_o[29200] = data_o[16];
  assign data_o[29264] = data_o[16];
  assign data_o[29328] = data_o[16];
  assign data_o[29392] = data_o[16];
  assign data_o[29456] = data_o[16];
  assign data_o[29520] = data_o[16];
  assign data_o[29584] = data_o[16];
  assign data_o[29648] = data_o[16];
  assign data_o[29712] = data_o[16];
  assign data_o[29776] = data_o[16];
  assign data_o[29840] = data_o[16];
  assign data_o[29904] = data_o[16];
  assign data_o[29968] = data_o[16];
  assign data_o[30032] = data_o[16];
  assign data_o[30096] = data_o[16];
  assign data_o[30160] = data_o[16];
  assign data_o[30224] = data_o[16];
  assign data_o[30288] = data_o[16];
  assign data_o[30352] = data_o[16];
  assign data_o[30416] = data_o[16];
  assign data_o[30480] = data_o[16];
  assign data_o[30544] = data_o[16];
  assign data_o[30608] = data_o[16];
  assign data_o[30672] = data_o[16];
  assign data_o[30736] = data_o[16];
  assign data_o[30800] = data_o[16];
  assign data_o[30864] = data_o[16];
  assign data_o[30928] = data_o[16];
  assign data_o[30992] = data_o[16];
  assign data_o[31056] = data_o[16];
  assign data_o[31120] = data_o[16];
  assign data_o[31184] = data_o[16];
  assign data_o[31248] = data_o[16];
  assign data_o[31312] = data_o[16];
  assign data_o[31376] = data_o[16];
  assign data_o[31440] = data_o[16];
  assign data_o[31504] = data_o[16];
  assign data_o[31568] = data_o[16];
  assign data_o[31632] = data_o[16];
  assign data_o[31696] = data_o[16];
  assign data_o[31760] = data_o[16];
  assign data_o[31824] = data_o[16];
  assign data_o[31888] = data_o[16];
  assign data_o[31952] = data_o[16];
  assign data_o[79] = data_o[15];
  assign data_o[143] = data_o[15];
  assign data_o[207] = data_o[15];
  assign data_o[271] = data_o[15];
  assign data_o[335] = data_o[15];
  assign data_o[399] = data_o[15];
  assign data_o[463] = data_o[15];
  assign data_o[527] = data_o[15];
  assign data_o[591] = data_o[15];
  assign data_o[655] = data_o[15];
  assign data_o[719] = data_o[15];
  assign data_o[783] = data_o[15];
  assign data_o[847] = data_o[15];
  assign data_o[911] = data_o[15];
  assign data_o[975] = data_o[15];
  assign data_o[1039] = data_o[15];
  assign data_o[1103] = data_o[15];
  assign data_o[1167] = data_o[15];
  assign data_o[1231] = data_o[15];
  assign data_o[1295] = data_o[15];
  assign data_o[1359] = data_o[15];
  assign data_o[1423] = data_o[15];
  assign data_o[1487] = data_o[15];
  assign data_o[1551] = data_o[15];
  assign data_o[1615] = data_o[15];
  assign data_o[1679] = data_o[15];
  assign data_o[1743] = data_o[15];
  assign data_o[1807] = data_o[15];
  assign data_o[1871] = data_o[15];
  assign data_o[1935] = data_o[15];
  assign data_o[1999] = data_o[15];
  assign data_o[2063] = data_o[15];
  assign data_o[2127] = data_o[15];
  assign data_o[2191] = data_o[15];
  assign data_o[2255] = data_o[15];
  assign data_o[2319] = data_o[15];
  assign data_o[2383] = data_o[15];
  assign data_o[2447] = data_o[15];
  assign data_o[2511] = data_o[15];
  assign data_o[2575] = data_o[15];
  assign data_o[2639] = data_o[15];
  assign data_o[2703] = data_o[15];
  assign data_o[2767] = data_o[15];
  assign data_o[2831] = data_o[15];
  assign data_o[2895] = data_o[15];
  assign data_o[2959] = data_o[15];
  assign data_o[3023] = data_o[15];
  assign data_o[3087] = data_o[15];
  assign data_o[3151] = data_o[15];
  assign data_o[3215] = data_o[15];
  assign data_o[3279] = data_o[15];
  assign data_o[3343] = data_o[15];
  assign data_o[3407] = data_o[15];
  assign data_o[3471] = data_o[15];
  assign data_o[3535] = data_o[15];
  assign data_o[3599] = data_o[15];
  assign data_o[3663] = data_o[15];
  assign data_o[3727] = data_o[15];
  assign data_o[3791] = data_o[15];
  assign data_o[3855] = data_o[15];
  assign data_o[3919] = data_o[15];
  assign data_o[3983] = data_o[15];
  assign data_o[4047] = data_o[15];
  assign data_o[4111] = data_o[15];
  assign data_o[4175] = data_o[15];
  assign data_o[4239] = data_o[15];
  assign data_o[4303] = data_o[15];
  assign data_o[4367] = data_o[15];
  assign data_o[4431] = data_o[15];
  assign data_o[4495] = data_o[15];
  assign data_o[4559] = data_o[15];
  assign data_o[4623] = data_o[15];
  assign data_o[4687] = data_o[15];
  assign data_o[4751] = data_o[15];
  assign data_o[4815] = data_o[15];
  assign data_o[4879] = data_o[15];
  assign data_o[4943] = data_o[15];
  assign data_o[5007] = data_o[15];
  assign data_o[5071] = data_o[15];
  assign data_o[5135] = data_o[15];
  assign data_o[5199] = data_o[15];
  assign data_o[5263] = data_o[15];
  assign data_o[5327] = data_o[15];
  assign data_o[5391] = data_o[15];
  assign data_o[5455] = data_o[15];
  assign data_o[5519] = data_o[15];
  assign data_o[5583] = data_o[15];
  assign data_o[5647] = data_o[15];
  assign data_o[5711] = data_o[15];
  assign data_o[5775] = data_o[15];
  assign data_o[5839] = data_o[15];
  assign data_o[5903] = data_o[15];
  assign data_o[5967] = data_o[15];
  assign data_o[6031] = data_o[15];
  assign data_o[6095] = data_o[15];
  assign data_o[6159] = data_o[15];
  assign data_o[6223] = data_o[15];
  assign data_o[6287] = data_o[15];
  assign data_o[6351] = data_o[15];
  assign data_o[6415] = data_o[15];
  assign data_o[6479] = data_o[15];
  assign data_o[6543] = data_o[15];
  assign data_o[6607] = data_o[15];
  assign data_o[6671] = data_o[15];
  assign data_o[6735] = data_o[15];
  assign data_o[6799] = data_o[15];
  assign data_o[6863] = data_o[15];
  assign data_o[6927] = data_o[15];
  assign data_o[6991] = data_o[15];
  assign data_o[7055] = data_o[15];
  assign data_o[7119] = data_o[15];
  assign data_o[7183] = data_o[15];
  assign data_o[7247] = data_o[15];
  assign data_o[7311] = data_o[15];
  assign data_o[7375] = data_o[15];
  assign data_o[7439] = data_o[15];
  assign data_o[7503] = data_o[15];
  assign data_o[7567] = data_o[15];
  assign data_o[7631] = data_o[15];
  assign data_o[7695] = data_o[15];
  assign data_o[7759] = data_o[15];
  assign data_o[7823] = data_o[15];
  assign data_o[7887] = data_o[15];
  assign data_o[7951] = data_o[15];
  assign data_o[8015] = data_o[15];
  assign data_o[8079] = data_o[15];
  assign data_o[8143] = data_o[15];
  assign data_o[8207] = data_o[15];
  assign data_o[8271] = data_o[15];
  assign data_o[8335] = data_o[15];
  assign data_o[8399] = data_o[15];
  assign data_o[8463] = data_o[15];
  assign data_o[8527] = data_o[15];
  assign data_o[8591] = data_o[15];
  assign data_o[8655] = data_o[15];
  assign data_o[8719] = data_o[15];
  assign data_o[8783] = data_o[15];
  assign data_o[8847] = data_o[15];
  assign data_o[8911] = data_o[15];
  assign data_o[8975] = data_o[15];
  assign data_o[9039] = data_o[15];
  assign data_o[9103] = data_o[15];
  assign data_o[9167] = data_o[15];
  assign data_o[9231] = data_o[15];
  assign data_o[9295] = data_o[15];
  assign data_o[9359] = data_o[15];
  assign data_o[9423] = data_o[15];
  assign data_o[9487] = data_o[15];
  assign data_o[9551] = data_o[15];
  assign data_o[9615] = data_o[15];
  assign data_o[9679] = data_o[15];
  assign data_o[9743] = data_o[15];
  assign data_o[9807] = data_o[15];
  assign data_o[9871] = data_o[15];
  assign data_o[9935] = data_o[15];
  assign data_o[9999] = data_o[15];
  assign data_o[10063] = data_o[15];
  assign data_o[10127] = data_o[15];
  assign data_o[10191] = data_o[15];
  assign data_o[10255] = data_o[15];
  assign data_o[10319] = data_o[15];
  assign data_o[10383] = data_o[15];
  assign data_o[10447] = data_o[15];
  assign data_o[10511] = data_o[15];
  assign data_o[10575] = data_o[15];
  assign data_o[10639] = data_o[15];
  assign data_o[10703] = data_o[15];
  assign data_o[10767] = data_o[15];
  assign data_o[10831] = data_o[15];
  assign data_o[10895] = data_o[15];
  assign data_o[10959] = data_o[15];
  assign data_o[11023] = data_o[15];
  assign data_o[11087] = data_o[15];
  assign data_o[11151] = data_o[15];
  assign data_o[11215] = data_o[15];
  assign data_o[11279] = data_o[15];
  assign data_o[11343] = data_o[15];
  assign data_o[11407] = data_o[15];
  assign data_o[11471] = data_o[15];
  assign data_o[11535] = data_o[15];
  assign data_o[11599] = data_o[15];
  assign data_o[11663] = data_o[15];
  assign data_o[11727] = data_o[15];
  assign data_o[11791] = data_o[15];
  assign data_o[11855] = data_o[15];
  assign data_o[11919] = data_o[15];
  assign data_o[11983] = data_o[15];
  assign data_o[12047] = data_o[15];
  assign data_o[12111] = data_o[15];
  assign data_o[12175] = data_o[15];
  assign data_o[12239] = data_o[15];
  assign data_o[12303] = data_o[15];
  assign data_o[12367] = data_o[15];
  assign data_o[12431] = data_o[15];
  assign data_o[12495] = data_o[15];
  assign data_o[12559] = data_o[15];
  assign data_o[12623] = data_o[15];
  assign data_o[12687] = data_o[15];
  assign data_o[12751] = data_o[15];
  assign data_o[12815] = data_o[15];
  assign data_o[12879] = data_o[15];
  assign data_o[12943] = data_o[15];
  assign data_o[13007] = data_o[15];
  assign data_o[13071] = data_o[15];
  assign data_o[13135] = data_o[15];
  assign data_o[13199] = data_o[15];
  assign data_o[13263] = data_o[15];
  assign data_o[13327] = data_o[15];
  assign data_o[13391] = data_o[15];
  assign data_o[13455] = data_o[15];
  assign data_o[13519] = data_o[15];
  assign data_o[13583] = data_o[15];
  assign data_o[13647] = data_o[15];
  assign data_o[13711] = data_o[15];
  assign data_o[13775] = data_o[15];
  assign data_o[13839] = data_o[15];
  assign data_o[13903] = data_o[15];
  assign data_o[13967] = data_o[15];
  assign data_o[14031] = data_o[15];
  assign data_o[14095] = data_o[15];
  assign data_o[14159] = data_o[15];
  assign data_o[14223] = data_o[15];
  assign data_o[14287] = data_o[15];
  assign data_o[14351] = data_o[15];
  assign data_o[14415] = data_o[15];
  assign data_o[14479] = data_o[15];
  assign data_o[14543] = data_o[15];
  assign data_o[14607] = data_o[15];
  assign data_o[14671] = data_o[15];
  assign data_o[14735] = data_o[15];
  assign data_o[14799] = data_o[15];
  assign data_o[14863] = data_o[15];
  assign data_o[14927] = data_o[15];
  assign data_o[14991] = data_o[15];
  assign data_o[15055] = data_o[15];
  assign data_o[15119] = data_o[15];
  assign data_o[15183] = data_o[15];
  assign data_o[15247] = data_o[15];
  assign data_o[15311] = data_o[15];
  assign data_o[15375] = data_o[15];
  assign data_o[15439] = data_o[15];
  assign data_o[15503] = data_o[15];
  assign data_o[15567] = data_o[15];
  assign data_o[15631] = data_o[15];
  assign data_o[15695] = data_o[15];
  assign data_o[15759] = data_o[15];
  assign data_o[15823] = data_o[15];
  assign data_o[15887] = data_o[15];
  assign data_o[15951] = data_o[15];
  assign data_o[16015] = data_o[15];
  assign data_o[16079] = data_o[15];
  assign data_o[16143] = data_o[15];
  assign data_o[16207] = data_o[15];
  assign data_o[16271] = data_o[15];
  assign data_o[16335] = data_o[15];
  assign data_o[16399] = data_o[15];
  assign data_o[16463] = data_o[15];
  assign data_o[16527] = data_o[15];
  assign data_o[16591] = data_o[15];
  assign data_o[16655] = data_o[15];
  assign data_o[16719] = data_o[15];
  assign data_o[16783] = data_o[15];
  assign data_o[16847] = data_o[15];
  assign data_o[16911] = data_o[15];
  assign data_o[16975] = data_o[15];
  assign data_o[17039] = data_o[15];
  assign data_o[17103] = data_o[15];
  assign data_o[17167] = data_o[15];
  assign data_o[17231] = data_o[15];
  assign data_o[17295] = data_o[15];
  assign data_o[17359] = data_o[15];
  assign data_o[17423] = data_o[15];
  assign data_o[17487] = data_o[15];
  assign data_o[17551] = data_o[15];
  assign data_o[17615] = data_o[15];
  assign data_o[17679] = data_o[15];
  assign data_o[17743] = data_o[15];
  assign data_o[17807] = data_o[15];
  assign data_o[17871] = data_o[15];
  assign data_o[17935] = data_o[15];
  assign data_o[17999] = data_o[15];
  assign data_o[18063] = data_o[15];
  assign data_o[18127] = data_o[15];
  assign data_o[18191] = data_o[15];
  assign data_o[18255] = data_o[15];
  assign data_o[18319] = data_o[15];
  assign data_o[18383] = data_o[15];
  assign data_o[18447] = data_o[15];
  assign data_o[18511] = data_o[15];
  assign data_o[18575] = data_o[15];
  assign data_o[18639] = data_o[15];
  assign data_o[18703] = data_o[15];
  assign data_o[18767] = data_o[15];
  assign data_o[18831] = data_o[15];
  assign data_o[18895] = data_o[15];
  assign data_o[18959] = data_o[15];
  assign data_o[19023] = data_o[15];
  assign data_o[19087] = data_o[15];
  assign data_o[19151] = data_o[15];
  assign data_o[19215] = data_o[15];
  assign data_o[19279] = data_o[15];
  assign data_o[19343] = data_o[15];
  assign data_o[19407] = data_o[15];
  assign data_o[19471] = data_o[15];
  assign data_o[19535] = data_o[15];
  assign data_o[19599] = data_o[15];
  assign data_o[19663] = data_o[15];
  assign data_o[19727] = data_o[15];
  assign data_o[19791] = data_o[15];
  assign data_o[19855] = data_o[15];
  assign data_o[19919] = data_o[15];
  assign data_o[19983] = data_o[15];
  assign data_o[20047] = data_o[15];
  assign data_o[20111] = data_o[15];
  assign data_o[20175] = data_o[15];
  assign data_o[20239] = data_o[15];
  assign data_o[20303] = data_o[15];
  assign data_o[20367] = data_o[15];
  assign data_o[20431] = data_o[15];
  assign data_o[20495] = data_o[15];
  assign data_o[20559] = data_o[15];
  assign data_o[20623] = data_o[15];
  assign data_o[20687] = data_o[15];
  assign data_o[20751] = data_o[15];
  assign data_o[20815] = data_o[15];
  assign data_o[20879] = data_o[15];
  assign data_o[20943] = data_o[15];
  assign data_o[21007] = data_o[15];
  assign data_o[21071] = data_o[15];
  assign data_o[21135] = data_o[15];
  assign data_o[21199] = data_o[15];
  assign data_o[21263] = data_o[15];
  assign data_o[21327] = data_o[15];
  assign data_o[21391] = data_o[15];
  assign data_o[21455] = data_o[15];
  assign data_o[21519] = data_o[15];
  assign data_o[21583] = data_o[15];
  assign data_o[21647] = data_o[15];
  assign data_o[21711] = data_o[15];
  assign data_o[21775] = data_o[15];
  assign data_o[21839] = data_o[15];
  assign data_o[21903] = data_o[15];
  assign data_o[21967] = data_o[15];
  assign data_o[22031] = data_o[15];
  assign data_o[22095] = data_o[15];
  assign data_o[22159] = data_o[15];
  assign data_o[22223] = data_o[15];
  assign data_o[22287] = data_o[15];
  assign data_o[22351] = data_o[15];
  assign data_o[22415] = data_o[15];
  assign data_o[22479] = data_o[15];
  assign data_o[22543] = data_o[15];
  assign data_o[22607] = data_o[15];
  assign data_o[22671] = data_o[15];
  assign data_o[22735] = data_o[15];
  assign data_o[22799] = data_o[15];
  assign data_o[22863] = data_o[15];
  assign data_o[22927] = data_o[15];
  assign data_o[22991] = data_o[15];
  assign data_o[23055] = data_o[15];
  assign data_o[23119] = data_o[15];
  assign data_o[23183] = data_o[15];
  assign data_o[23247] = data_o[15];
  assign data_o[23311] = data_o[15];
  assign data_o[23375] = data_o[15];
  assign data_o[23439] = data_o[15];
  assign data_o[23503] = data_o[15];
  assign data_o[23567] = data_o[15];
  assign data_o[23631] = data_o[15];
  assign data_o[23695] = data_o[15];
  assign data_o[23759] = data_o[15];
  assign data_o[23823] = data_o[15];
  assign data_o[23887] = data_o[15];
  assign data_o[23951] = data_o[15];
  assign data_o[24015] = data_o[15];
  assign data_o[24079] = data_o[15];
  assign data_o[24143] = data_o[15];
  assign data_o[24207] = data_o[15];
  assign data_o[24271] = data_o[15];
  assign data_o[24335] = data_o[15];
  assign data_o[24399] = data_o[15];
  assign data_o[24463] = data_o[15];
  assign data_o[24527] = data_o[15];
  assign data_o[24591] = data_o[15];
  assign data_o[24655] = data_o[15];
  assign data_o[24719] = data_o[15];
  assign data_o[24783] = data_o[15];
  assign data_o[24847] = data_o[15];
  assign data_o[24911] = data_o[15];
  assign data_o[24975] = data_o[15];
  assign data_o[25039] = data_o[15];
  assign data_o[25103] = data_o[15];
  assign data_o[25167] = data_o[15];
  assign data_o[25231] = data_o[15];
  assign data_o[25295] = data_o[15];
  assign data_o[25359] = data_o[15];
  assign data_o[25423] = data_o[15];
  assign data_o[25487] = data_o[15];
  assign data_o[25551] = data_o[15];
  assign data_o[25615] = data_o[15];
  assign data_o[25679] = data_o[15];
  assign data_o[25743] = data_o[15];
  assign data_o[25807] = data_o[15];
  assign data_o[25871] = data_o[15];
  assign data_o[25935] = data_o[15];
  assign data_o[25999] = data_o[15];
  assign data_o[26063] = data_o[15];
  assign data_o[26127] = data_o[15];
  assign data_o[26191] = data_o[15];
  assign data_o[26255] = data_o[15];
  assign data_o[26319] = data_o[15];
  assign data_o[26383] = data_o[15];
  assign data_o[26447] = data_o[15];
  assign data_o[26511] = data_o[15];
  assign data_o[26575] = data_o[15];
  assign data_o[26639] = data_o[15];
  assign data_o[26703] = data_o[15];
  assign data_o[26767] = data_o[15];
  assign data_o[26831] = data_o[15];
  assign data_o[26895] = data_o[15];
  assign data_o[26959] = data_o[15];
  assign data_o[27023] = data_o[15];
  assign data_o[27087] = data_o[15];
  assign data_o[27151] = data_o[15];
  assign data_o[27215] = data_o[15];
  assign data_o[27279] = data_o[15];
  assign data_o[27343] = data_o[15];
  assign data_o[27407] = data_o[15];
  assign data_o[27471] = data_o[15];
  assign data_o[27535] = data_o[15];
  assign data_o[27599] = data_o[15];
  assign data_o[27663] = data_o[15];
  assign data_o[27727] = data_o[15];
  assign data_o[27791] = data_o[15];
  assign data_o[27855] = data_o[15];
  assign data_o[27919] = data_o[15];
  assign data_o[27983] = data_o[15];
  assign data_o[28047] = data_o[15];
  assign data_o[28111] = data_o[15];
  assign data_o[28175] = data_o[15];
  assign data_o[28239] = data_o[15];
  assign data_o[28303] = data_o[15];
  assign data_o[28367] = data_o[15];
  assign data_o[28431] = data_o[15];
  assign data_o[28495] = data_o[15];
  assign data_o[28559] = data_o[15];
  assign data_o[28623] = data_o[15];
  assign data_o[28687] = data_o[15];
  assign data_o[28751] = data_o[15];
  assign data_o[28815] = data_o[15];
  assign data_o[28879] = data_o[15];
  assign data_o[28943] = data_o[15];
  assign data_o[29007] = data_o[15];
  assign data_o[29071] = data_o[15];
  assign data_o[29135] = data_o[15];
  assign data_o[29199] = data_o[15];
  assign data_o[29263] = data_o[15];
  assign data_o[29327] = data_o[15];
  assign data_o[29391] = data_o[15];
  assign data_o[29455] = data_o[15];
  assign data_o[29519] = data_o[15];
  assign data_o[29583] = data_o[15];
  assign data_o[29647] = data_o[15];
  assign data_o[29711] = data_o[15];
  assign data_o[29775] = data_o[15];
  assign data_o[29839] = data_o[15];
  assign data_o[29903] = data_o[15];
  assign data_o[29967] = data_o[15];
  assign data_o[30031] = data_o[15];
  assign data_o[30095] = data_o[15];
  assign data_o[30159] = data_o[15];
  assign data_o[30223] = data_o[15];
  assign data_o[30287] = data_o[15];
  assign data_o[30351] = data_o[15];
  assign data_o[30415] = data_o[15];
  assign data_o[30479] = data_o[15];
  assign data_o[30543] = data_o[15];
  assign data_o[30607] = data_o[15];
  assign data_o[30671] = data_o[15];
  assign data_o[30735] = data_o[15];
  assign data_o[30799] = data_o[15];
  assign data_o[30863] = data_o[15];
  assign data_o[30927] = data_o[15];
  assign data_o[30991] = data_o[15];
  assign data_o[31055] = data_o[15];
  assign data_o[31119] = data_o[15];
  assign data_o[31183] = data_o[15];
  assign data_o[31247] = data_o[15];
  assign data_o[31311] = data_o[15];
  assign data_o[31375] = data_o[15];
  assign data_o[31439] = data_o[15];
  assign data_o[31503] = data_o[15];
  assign data_o[31567] = data_o[15];
  assign data_o[31631] = data_o[15];
  assign data_o[31695] = data_o[15];
  assign data_o[31759] = data_o[15];
  assign data_o[31823] = data_o[15];
  assign data_o[31887] = data_o[15];
  assign data_o[31951] = data_o[15];
  assign data_o[78] = data_o[14];
  assign data_o[142] = data_o[14];
  assign data_o[206] = data_o[14];
  assign data_o[270] = data_o[14];
  assign data_o[334] = data_o[14];
  assign data_o[398] = data_o[14];
  assign data_o[462] = data_o[14];
  assign data_o[526] = data_o[14];
  assign data_o[590] = data_o[14];
  assign data_o[654] = data_o[14];
  assign data_o[718] = data_o[14];
  assign data_o[782] = data_o[14];
  assign data_o[846] = data_o[14];
  assign data_o[910] = data_o[14];
  assign data_o[974] = data_o[14];
  assign data_o[1038] = data_o[14];
  assign data_o[1102] = data_o[14];
  assign data_o[1166] = data_o[14];
  assign data_o[1230] = data_o[14];
  assign data_o[1294] = data_o[14];
  assign data_o[1358] = data_o[14];
  assign data_o[1422] = data_o[14];
  assign data_o[1486] = data_o[14];
  assign data_o[1550] = data_o[14];
  assign data_o[1614] = data_o[14];
  assign data_o[1678] = data_o[14];
  assign data_o[1742] = data_o[14];
  assign data_o[1806] = data_o[14];
  assign data_o[1870] = data_o[14];
  assign data_o[1934] = data_o[14];
  assign data_o[1998] = data_o[14];
  assign data_o[2062] = data_o[14];
  assign data_o[2126] = data_o[14];
  assign data_o[2190] = data_o[14];
  assign data_o[2254] = data_o[14];
  assign data_o[2318] = data_o[14];
  assign data_o[2382] = data_o[14];
  assign data_o[2446] = data_o[14];
  assign data_o[2510] = data_o[14];
  assign data_o[2574] = data_o[14];
  assign data_o[2638] = data_o[14];
  assign data_o[2702] = data_o[14];
  assign data_o[2766] = data_o[14];
  assign data_o[2830] = data_o[14];
  assign data_o[2894] = data_o[14];
  assign data_o[2958] = data_o[14];
  assign data_o[3022] = data_o[14];
  assign data_o[3086] = data_o[14];
  assign data_o[3150] = data_o[14];
  assign data_o[3214] = data_o[14];
  assign data_o[3278] = data_o[14];
  assign data_o[3342] = data_o[14];
  assign data_o[3406] = data_o[14];
  assign data_o[3470] = data_o[14];
  assign data_o[3534] = data_o[14];
  assign data_o[3598] = data_o[14];
  assign data_o[3662] = data_o[14];
  assign data_o[3726] = data_o[14];
  assign data_o[3790] = data_o[14];
  assign data_o[3854] = data_o[14];
  assign data_o[3918] = data_o[14];
  assign data_o[3982] = data_o[14];
  assign data_o[4046] = data_o[14];
  assign data_o[4110] = data_o[14];
  assign data_o[4174] = data_o[14];
  assign data_o[4238] = data_o[14];
  assign data_o[4302] = data_o[14];
  assign data_o[4366] = data_o[14];
  assign data_o[4430] = data_o[14];
  assign data_o[4494] = data_o[14];
  assign data_o[4558] = data_o[14];
  assign data_o[4622] = data_o[14];
  assign data_o[4686] = data_o[14];
  assign data_o[4750] = data_o[14];
  assign data_o[4814] = data_o[14];
  assign data_o[4878] = data_o[14];
  assign data_o[4942] = data_o[14];
  assign data_o[5006] = data_o[14];
  assign data_o[5070] = data_o[14];
  assign data_o[5134] = data_o[14];
  assign data_o[5198] = data_o[14];
  assign data_o[5262] = data_o[14];
  assign data_o[5326] = data_o[14];
  assign data_o[5390] = data_o[14];
  assign data_o[5454] = data_o[14];
  assign data_o[5518] = data_o[14];
  assign data_o[5582] = data_o[14];
  assign data_o[5646] = data_o[14];
  assign data_o[5710] = data_o[14];
  assign data_o[5774] = data_o[14];
  assign data_o[5838] = data_o[14];
  assign data_o[5902] = data_o[14];
  assign data_o[5966] = data_o[14];
  assign data_o[6030] = data_o[14];
  assign data_o[6094] = data_o[14];
  assign data_o[6158] = data_o[14];
  assign data_o[6222] = data_o[14];
  assign data_o[6286] = data_o[14];
  assign data_o[6350] = data_o[14];
  assign data_o[6414] = data_o[14];
  assign data_o[6478] = data_o[14];
  assign data_o[6542] = data_o[14];
  assign data_o[6606] = data_o[14];
  assign data_o[6670] = data_o[14];
  assign data_o[6734] = data_o[14];
  assign data_o[6798] = data_o[14];
  assign data_o[6862] = data_o[14];
  assign data_o[6926] = data_o[14];
  assign data_o[6990] = data_o[14];
  assign data_o[7054] = data_o[14];
  assign data_o[7118] = data_o[14];
  assign data_o[7182] = data_o[14];
  assign data_o[7246] = data_o[14];
  assign data_o[7310] = data_o[14];
  assign data_o[7374] = data_o[14];
  assign data_o[7438] = data_o[14];
  assign data_o[7502] = data_o[14];
  assign data_o[7566] = data_o[14];
  assign data_o[7630] = data_o[14];
  assign data_o[7694] = data_o[14];
  assign data_o[7758] = data_o[14];
  assign data_o[7822] = data_o[14];
  assign data_o[7886] = data_o[14];
  assign data_o[7950] = data_o[14];
  assign data_o[8014] = data_o[14];
  assign data_o[8078] = data_o[14];
  assign data_o[8142] = data_o[14];
  assign data_o[8206] = data_o[14];
  assign data_o[8270] = data_o[14];
  assign data_o[8334] = data_o[14];
  assign data_o[8398] = data_o[14];
  assign data_o[8462] = data_o[14];
  assign data_o[8526] = data_o[14];
  assign data_o[8590] = data_o[14];
  assign data_o[8654] = data_o[14];
  assign data_o[8718] = data_o[14];
  assign data_o[8782] = data_o[14];
  assign data_o[8846] = data_o[14];
  assign data_o[8910] = data_o[14];
  assign data_o[8974] = data_o[14];
  assign data_o[9038] = data_o[14];
  assign data_o[9102] = data_o[14];
  assign data_o[9166] = data_o[14];
  assign data_o[9230] = data_o[14];
  assign data_o[9294] = data_o[14];
  assign data_o[9358] = data_o[14];
  assign data_o[9422] = data_o[14];
  assign data_o[9486] = data_o[14];
  assign data_o[9550] = data_o[14];
  assign data_o[9614] = data_o[14];
  assign data_o[9678] = data_o[14];
  assign data_o[9742] = data_o[14];
  assign data_o[9806] = data_o[14];
  assign data_o[9870] = data_o[14];
  assign data_o[9934] = data_o[14];
  assign data_o[9998] = data_o[14];
  assign data_o[10062] = data_o[14];
  assign data_o[10126] = data_o[14];
  assign data_o[10190] = data_o[14];
  assign data_o[10254] = data_o[14];
  assign data_o[10318] = data_o[14];
  assign data_o[10382] = data_o[14];
  assign data_o[10446] = data_o[14];
  assign data_o[10510] = data_o[14];
  assign data_o[10574] = data_o[14];
  assign data_o[10638] = data_o[14];
  assign data_o[10702] = data_o[14];
  assign data_o[10766] = data_o[14];
  assign data_o[10830] = data_o[14];
  assign data_o[10894] = data_o[14];
  assign data_o[10958] = data_o[14];
  assign data_o[11022] = data_o[14];
  assign data_o[11086] = data_o[14];
  assign data_o[11150] = data_o[14];
  assign data_o[11214] = data_o[14];
  assign data_o[11278] = data_o[14];
  assign data_o[11342] = data_o[14];
  assign data_o[11406] = data_o[14];
  assign data_o[11470] = data_o[14];
  assign data_o[11534] = data_o[14];
  assign data_o[11598] = data_o[14];
  assign data_o[11662] = data_o[14];
  assign data_o[11726] = data_o[14];
  assign data_o[11790] = data_o[14];
  assign data_o[11854] = data_o[14];
  assign data_o[11918] = data_o[14];
  assign data_o[11982] = data_o[14];
  assign data_o[12046] = data_o[14];
  assign data_o[12110] = data_o[14];
  assign data_o[12174] = data_o[14];
  assign data_o[12238] = data_o[14];
  assign data_o[12302] = data_o[14];
  assign data_o[12366] = data_o[14];
  assign data_o[12430] = data_o[14];
  assign data_o[12494] = data_o[14];
  assign data_o[12558] = data_o[14];
  assign data_o[12622] = data_o[14];
  assign data_o[12686] = data_o[14];
  assign data_o[12750] = data_o[14];
  assign data_o[12814] = data_o[14];
  assign data_o[12878] = data_o[14];
  assign data_o[12942] = data_o[14];
  assign data_o[13006] = data_o[14];
  assign data_o[13070] = data_o[14];
  assign data_o[13134] = data_o[14];
  assign data_o[13198] = data_o[14];
  assign data_o[13262] = data_o[14];
  assign data_o[13326] = data_o[14];
  assign data_o[13390] = data_o[14];
  assign data_o[13454] = data_o[14];
  assign data_o[13518] = data_o[14];
  assign data_o[13582] = data_o[14];
  assign data_o[13646] = data_o[14];
  assign data_o[13710] = data_o[14];
  assign data_o[13774] = data_o[14];
  assign data_o[13838] = data_o[14];
  assign data_o[13902] = data_o[14];
  assign data_o[13966] = data_o[14];
  assign data_o[14030] = data_o[14];
  assign data_o[14094] = data_o[14];
  assign data_o[14158] = data_o[14];
  assign data_o[14222] = data_o[14];
  assign data_o[14286] = data_o[14];
  assign data_o[14350] = data_o[14];
  assign data_o[14414] = data_o[14];
  assign data_o[14478] = data_o[14];
  assign data_o[14542] = data_o[14];
  assign data_o[14606] = data_o[14];
  assign data_o[14670] = data_o[14];
  assign data_o[14734] = data_o[14];
  assign data_o[14798] = data_o[14];
  assign data_o[14862] = data_o[14];
  assign data_o[14926] = data_o[14];
  assign data_o[14990] = data_o[14];
  assign data_o[15054] = data_o[14];
  assign data_o[15118] = data_o[14];
  assign data_o[15182] = data_o[14];
  assign data_o[15246] = data_o[14];
  assign data_o[15310] = data_o[14];
  assign data_o[15374] = data_o[14];
  assign data_o[15438] = data_o[14];
  assign data_o[15502] = data_o[14];
  assign data_o[15566] = data_o[14];
  assign data_o[15630] = data_o[14];
  assign data_o[15694] = data_o[14];
  assign data_o[15758] = data_o[14];
  assign data_o[15822] = data_o[14];
  assign data_o[15886] = data_o[14];
  assign data_o[15950] = data_o[14];
  assign data_o[16014] = data_o[14];
  assign data_o[16078] = data_o[14];
  assign data_o[16142] = data_o[14];
  assign data_o[16206] = data_o[14];
  assign data_o[16270] = data_o[14];
  assign data_o[16334] = data_o[14];
  assign data_o[16398] = data_o[14];
  assign data_o[16462] = data_o[14];
  assign data_o[16526] = data_o[14];
  assign data_o[16590] = data_o[14];
  assign data_o[16654] = data_o[14];
  assign data_o[16718] = data_o[14];
  assign data_o[16782] = data_o[14];
  assign data_o[16846] = data_o[14];
  assign data_o[16910] = data_o[14];
  assign data_o[16974] = data_o[14];
  assign data_o[17038] = data_o[14];
  assign data_o[17102] = data_o[14];
  assign data_o[17166] = data_o[14];
  assign data_o[17230] = data_o[14];
  assign data_o[17294] = data_o[14];
  assign data_o[17358] = data_o[14];
  assign data_o[17422] = data_o[14];
  assign data_o[17486] = data_o[14];
  assign data_o[17550] = data_o[14];
  assign data_o[17614] = data_o[14];
  assign data_o[17678] = data_o[14];
  assign data_o[17742] = data_o[14];
  assign data_o[17806] = data_o[14];
  assign data_o[17870] = data_o[14];
  assign data_o[17934] = data_o[14];
  assign data_o[17998] = data_o[14];
  assign data_o[18062] = data_o[14];
  assign data_o[18126] = data_o[14];
  assign data_o[18190] = data_o[14];
  assign data_o[18254] = data_o[14];
  assign data_o[18318] = data_o[14];
  assign data_o[18382] = data_o[14];
  assign data_o[18446] = data_o[14];
  assign data_o[18510] = data_o[14];
  assign data_o[18574] = data_o[14];
  assign data_o[18638] = data_o[14];
  assign data_o[18702] = data_o[14];
  assign data_o[18766] = data_o[14];
  assign data_o[18830] = data_o[14];
  assign data_o[18894] = data_o[14];
  assign data_o[18958] = data_o[14];
  assign data_o[19022] = data_o[14];
  assign data_o[19086] = data_o[14];
  assign data_o[19150] = data_o[14];
  assign data_o[19214] = data_o[14];
  assign data_o[19278] = data_o[14];
  assign data_o[19342] = data_o[14];
  assign data_o[19406] = data_o[14];
  assign data_o[19470] = data_o[14];
  assign data_o[19534] = data_o[14];
  assign data_o[19598] = data_o[14];
  assign data_o[19662] = data_o[14];
  assign data_o[19726] = data_o[14];
  assign data_o[19790] = data_o[14];
  assign data_o[19854] = data_o[14];
  assign data_o[19918] = data_o[14];
  assign data_o[19982] = data_o[14];
  assign data_o[20046] = data_o[14];
  assign data_o[20110] = data_o[14];
  assign data_o[20174] = data_o[14];
  assign data_o[20238] = data_o[14];
  assign data_o[20302] = data_o[14];
  assign data_o[20366] = data_o[14];
  assign data_o[20430] = data_o[14];
  assign data_o[20494] = data_o[14];
  assign data_o[20558] = data_o[14];
  assign data_o[20622] = data_o[14];
  assign data_o[20686] = data_o[14];
  assign data_o[20750] = data_o[14];
  assign data_o[20814] = data_o[14];
  assign data_o[20878] = data_o[14];
  assign data_o[20942] = data_o[14];
  assign data_o[21006] = data_o[14];
  assign data_o[21070] = data_o[14];
  assign data_o[21134] = data_o[14];
  assign data_o[21198] = data_o[14];
  assign data_o[21262] = data_o[14];
  assign data_o[21326] = data_o[14];
  assign data_o[21390] = data_o[14];
  assign data_o[21454] = data_o[14];
  assign data_o[21518] = data_o[14];
  assign data_o[21582] = data_o[14];
  assign data_o[21646] = data_o[14];
  assign data_o[21710] = data_o[14];
  assign data_o[21774] = data_o[14];
  assign data_o[21838] = data_o[14];
  assign data_o[21902] = data_o[14];
  assign data_o[21966] = data_o[14];
  assign data_o[22030] = data_o[14];
  assign data_o[22094] = data_o[14];
  assign data_o[22158] = data_o[14];
  assign data_o[22222] = data_o[14];
  assign data_o[22286] = data_o[14];
  assign data_o[22350] = data_o[14];
  assign data_o[22414] = data_o[14];
  assign data_o[22478] = data_o[14];
  assign data_o[22542] = data_o[14];
  assign data_o[22606] = data_o[14];
  assign data_o[22670] = data_o[14];
  assign data_o[22734] = data_o[14];
  assign data_o[22798] = data_o[14];
  assign data_o[22862] = data_o[14];
  assign data_o[22926] = data_o[14];
  assign data_o[22990] = data_o[14];
  assign data_o[23054] = data_o[14];
  assign data_o[23118] = data_o[14];
  assign data_o[23182] = data_o[14];
  assign data_o[23246] = data_o[14];
  assign data_o[23310] = data_o[14];
  assign data_o[23374] = data_o[14];
  assign data_o[23438] = data_o[14];
  assign data_o[23502] = data_o[14];
  assign data_o[23566] = data_o[14];
  assign data_o[23630] = data_o[14];
  assign data_o[23694] = data_o[14];
  assign data_o[23758] = data_o[14];
  assign data_o[23822] = data_o[14];
  assign data_o[23886] = data_o[14];
  assign data_o[23950] = data_o[14];
  assign data_o[24014] = data_o[14];
  assign data_o[24078] = data_o[14];
  assign data_o[24142] = data_o[14];
  assign data_o[24206] = data_o[14];
  assign data_o[24270] = data_o[14];
  assign data_o[24334] = data_o[14];
  assign data_o[24398] = data_o[14];
  assign data_o[24462] = data_o[14];
  assign data_o[24526] = data_o[14];
  assign data_o[24590] = data_o[14];
  assign data_o[24654] = data_o[14];
  assign data_o[24718] = data_o[14];
  assign data_o[24782] = data_o[14];
  assign data_o[24846] = data_o[14];
  assign data_o[24910] = data_o[14];
  assign data_o[24974] = data_o[14];
  assign data_o[25038] = data_o[14];
  assign data_o[25102] = data_o[14];
  assign data_o[25166] = data_o[14];
  assign data_o[25230] = data_o[14];
  assign data_o[25294] = data_o[14];
  assign data_o[25358] = data_o[14];
  assign data_o[25422] = data_o[14];
  assign data_o[25486] = data_o[14];
  assign data_o[25550] = data_o[14];
  assign data_o[25614] = data_o[14];
  assign data_o[25678] = data_o[14];
  assign data_o[25742] = data_o[14];
  assign data_o[25806] = data_o[14];
  assign data_o[25870] = data_o[14];
  assign data_o[25934] = data_o[14];
  assign data_o[25998] = data_o[14];
  assign data_o[26062] = data_o[14];
  assign data_o[26126] = data_o[14];
  assign data_o[26190] = data_o[14];
  assign data_o[26254] = data_o[14];
  assign data_o[26318] = data_o[14];
  assign data_o[26382] = data_o[14];
  assign data_o[26446] = data_o[14];
  assign data_o[26510] = data_o[14];
  assign data_o[26574] = data_o[14];
  assign data_o[26638] = data_o[14];
  assign data_o[26702] = data_o[14];
  assign data_o[26766] = data_o[14];
  assign data_o[26830] = data_o[14];
  assign data_o[26894] = data_o[14];
  assign data_o[26958] = data_o[14];
  assign data_o[27022] = data_o[14];
  assign data_o[27086] = data_o[14];
  assign data_o[27150] = data_o[14];
  assign data_o[27214] = data_o[14];
  assign data_o[27278] = data_o[14];
  assign data_o[27342] = data_o[14];
  assign data_o[27406] = data_o[14];
  assign data_o[27470] = data_o[14];
  assign data_o[27534] = data_o[14];
  assign data_o[27598] = data_o[14];
  assign data_o[27662] = data_o[14];
  assign data_o[27726] = data_o[14];
  assign data_o[27790] = data_o[14];
  assign data_o[27854] = data_o[14];
  assign data_o[27918] = data_o[14];
  assign data_o[27982] = data_o[14];
  assign data_o[28046] = data_o[14];
  assign data_o[28110] = data_o[14];
  assign data_o[28174] = data_o[14];
  assign data_o[28238] = data_o[14];
  assign data_o[28302] = data_o[14];
  assign data_o[28366] = data_o[14];
  assign data_o[28430] = data_o[14];
  assign data_o[28494] = data_o[14];
  assign data_o[28558] = data_o[14];
  assign data_o[28622] = data_o[14];
  assign data_o[28686] = data_o[14];
  assign data_o[28750] = data_o[14];
  assign data_o[28814] = data_o[14];
  assign data_o[28878] = data_o[14];
  assign data_o[28942] = data_o[14];
  assign data_o[29006] = data_o[14];
  assign data_o[29070] = data_o[14];
  assign data_o[29134] = data_o[14];
  assign data_o[29198] = data_o[14];
  assign data_o[29262] = data_o[14];
  assign data_o[29326] = data_o[14];
  assign data_o[29390] = data_o[14];
  assign data_o[29454] = data_o[14];
  assign data_o[29518] = data_o[14];
  assign data_o[29582] = data_o[14];
  assign data_o[29646] = data_o[14];
  assign data_o[29710] = data_o[14];
  assign data_o[29774] = data_o[14];
  assign data_o[29838] = data_o[14];
  assign data_o[29902] = data_o[14];
  assign data_o[29966] = data_o[14];
  assign data_o[30030] = data_o[14];
  assign data_o[30094] = data_o[14];
  assign data_o[30158] = data_o[14];
  assign data_o[30222] = data_o[14];
  assign data_o[30286] = data_o[14];
  assign data_o[30350] = data_o[14];
  assign data_o[30414] = data_o[14];
  assign data_o[30478] = data_o[14];
  assign data_o[30542] = data_o[14];
  assign data_o[30606] = data_o[14];
  assign data_o[30670] = data_o[14];
  assign data_o[30734] = data_o[14];
  assign data_o[30798] = data_o[14];
  assign data_o[30862] = data_o[14];
  assign data_o[30926] = data_o[14];
  assign data_o[30990] = data_o[14];
  assign data_o[31054] = data_o[14];
  assign data_o[31118] = data_o[14];
  assign data_o[31182] = data_o[14];
  assign data_o[31246] = data_o[14];
  assign data_o[31310] = data_o[14];
  assign data_o[31374] = data_o[14];
  assign data_o[31438] = data_o[14];
  assign data_o[31502] = data_o[14];
  assign data_o[31566] = data_o[14];
  assign data_o[31630] = data_o[14];
  assign data_o[31694] = data_o[14];
  assign data_o[31758] = data_o[14];
  assign data_o[31822] = data_o[14];
  assign data_o[31886] = data_o[14];
  assign data_o[31950] = data_o[14];
  assign data_o[77] = data_o[13];
  assign data_o[141] = data_o[13];
  assign data_o[205] = data_o[13];
  assign data_o[269] = data_o[13];
  assign data_o[333] = data_o[13];
  assign data_o[397] = data_o[13];
  assign data_o[461] = data_o[13];
  assign data_o[525] = data_o[13];
  assign data_o[589] = data_o[13];
  assign data_o[653] = data_o[13];
  assign data_o[717] = data_o[13];
  assign data_o[781] = data_o[13];
  assign data_o[845] = data_o[13];
  assign data_o[909] = data_o[13];
  assign data_o[973] = data_o[13];
  assign data_o[1037] = data_o[13];
  assign data_o[1101] = data_o[13];
  assign data_o[1165] = data_o[13];
  assign data_o[1229] = data_o[13];
  assign data_o[1293] = data_o[13];
  assign data_o[1357] = data_o[13];
  assign data_o[1421] = data_o[13];
  assign data_o[1485] = data_o[13];
  assign data_o[1549] = data_o[13];
  assign data_o[1613] = data_o[13];
  assign data_o[1677] = data_o[13];
  assign data_o[1741] = data_o[13];
  assign data_o[1805] = data_o[13];
  assign data_o[1869] = data_o[13];
  assign data_o[1933] = data_o[13];
  assign data_o[1997] = data_o[13];
  assign data_o[2061] = data_o[13];
  assign data_o[2125] = data_o[13];
  assign data_o[2189] = data_o[13];
  assign data_o[2253] = data_o[13];
  assign data_o[2317] = data_o[13];
  assign data_o[2381] = data_o[13];
  assign data_o[2445] = data_o[13];
  assign data_o[2509] = data_o[13];
  assign data_o[2573] = data_o[13];
  assign data_o[2637] = data_o[13];
  assign data_o[2701] = data_o[13];
  assign data_o[2765] = data_o[13];
  assign data_o[2829] = data_o[13];
  assign data_o[2893] = data_o[13];
  assign data_o[2957] = data_o[13];
  assign data_o[3021] = data_o[13];
  assign data_o[3085] = data_o[13];
  assign data_o[3149] = data_o[13];
  assign data_o[3213] = data_o[13];
  assign data_o[3277] = data_o[13];
  assign data_o[3341] = data_o[13];
  assign data_o[3405] = data_o[13];
  assign data_o[3469] = data_o[13];
  assign data_o[3533] = data_o[13];
  assign data_o[3597] = data_o[13];
  assign data_o[3661] = data_o[13];
  assign data_o[3725] = data_o[13];
  assign data_o[3789] = data_o[13];
  assign data_o[3853] = data_o[13];
  assign data_o[3917] = data_o[13];
  assign data_o[3981] = data_o[13];
  assign data_o[4045] = data_o[13];
  assign data_o[4109] = data_o[13];
  assign data_o[4173] = data_o[13];
  assign data_o[4237] = data_o[13];
  assign data_o[4301] = data_o[13];
  assign data_o[4365] = data_o[13];
  assign data_o[4429] = data_o[13];
  assign data_o[4493] = data_o[13];
  assign data_o[4557] = data_o[13];
  assign data_o[4621] = data_o[13];
  assign data_o[4685] = data_o[13];
  assign data_o[4749] = data_o[13];
  assign data_o[4813] = data_o[13];
  assign data_o[4877] = data_o[13];
  assign data_o[4941] = data_o[13];
  assign data_o[5005] = data_o[13];
  assign data_o[5069] = data_o[13];
  assign data_o[5133] = data_o[13];
  assign data_o[5197] = data_o[13];
  assign data_o[5261] = data_o[13];
  assign data_o[5325] = data_o[13];
  assign data_o[5389] = data_o[13];
  assign data_o[5453] = data_o[13];
  assign data_o[5517] = data_o[13];
  assign data_o[5581] = data_o[13];
  assign data_o[5645] = data_o[13];
  assign data_o[5709] = data_o[13];
  assign data_o[5773] = data_o[13];
  assign data_o[5837] = data_o[13];
  assign data_o[5901] = data_o[13];
  assign data_o[5965] = data_o[13];
  assign data_o[6029] = data_o[13];
  assign data_o[6093] = data_o[13];
  assign data_o[6157] = data_o[13];
  assign data_o[6221] = data_o[13];
  assign data_o[6285] = data_o[13];
  assign data_o[6349] = data_o[13];
  assign data_o[6413] = data_o[13];
  assign data_o[6477] = data_o[13];
  assign data_o[6541] = data_o[13];
  assign data_o[6605] = data_o[13];
  assign data_o[6669] = data_o[13];
  assign data_o[6733] = data_o[13];
  assign data_o[6797] = data_o[13];
  assign data_o[6861] = data_o[13];
  assign data_o[6925] = data_o[13];
  assign data_o[6989] = data_o[13];
  assign data_o[7053] = data_o[13];
  assign data_o[7117] = data_o[13];
  assign data_o[7181] = data_o[13];
  assign data_o[7245] = data_o[13];
  assign data_o[7309] = data_o[13];
  assign data_o[7373] = data_o[13];
  assign data_o[7437] = data_o[13];
  assign data_o[7501] = data_o[13];
  assign data_o[7565] = data_o[13];
  assign data_o[7629] = data_o[13];
  assign data_o[7693] = data_o[13];
  assign data_o[7757] = data_o[13];
  assign data_o[7821] = data_o[13];
  assign data_o[7885] = data_o[13];
  assign data_o[7949] = data_o[13];
  assign data_o[8013] = data_o[13];
  assign data_o[8077] = data_o[13];
  assign data_o[8141] = data_o[13];
  assign data_o[8205] = data_o[13];
  assign data_o[8269] = data_o[13];
  assign data_o[8333] = data_o[13];
  assign data_o[8397] = data_o[13];
  assign data_o[8461] = data_o[13];
  assign data_o[8525] = data_o[13];
  assign data_o[8589] = data_o[13];
  assign data_o[8653] = data_o[13];
  assign data_o[8717] = data_o[13];
  assign data_o[8781] = data_o[13];
  assign data_o[8845] = data_o[13];
  assign data_o[8909] = data_o[13];
  assign data_o[8973] = data_o[13];
  assign data_o[9037] = data_o[13];
  assign data_o[9101] = data_o[13];
  assign data_o[9165] = data_o[13];
  assign data_o[9229] = data_o[13];
  assign data_o[9293] = data_o[13];
  assign data_o[9357] = data_o[13];
  assign data_o[9421] = data_o[13];
  assign data_o[9485] = data_o[13];
  assign data_o[9549] = data_o[13];
  assign data_o[9613] = data_o[13];
  assign data_o[9677] = data_o[13];
  assign data_o[9741] = data_o[13];
  assign data_o[9805] = data_o[13];
  assign data_o[9869] = data_o[13];
  assign data_o[9933] = data_o[13];
  assign data_o[9997] = data_o[13];
  assign data_o[10061] = data_o[13];
  assign data_o[10125] = data_o[13];
  assign data_o[10189] = data_o[13];
  assign data_o[10253] = data_o[13];
  assign data_o[10317] = data_o[13];
  assign data_o[10381] = data_o[13];
  assign data_o[10445] = data_o[13];
  assign data_o[10509] = data_o[13];
  assign data_o[10573] = data_o[13];
  assign data_o[10637] = data_o[13];
  assign data_o[10701] = data_o[13];
  assign data_o[10765] = data_o[13];
  assign data_o[10829] = data_o[13];
  assign data_o[10893] = data_o[13];
  assign data_o[10957] = data_o[13];
  assign data_o[11021] = data_o[13];
  assign data_o[11085] = data_o[13];
  assign data_o[11149] = data_o[13];
  assign data_o[11213] = data_o[13];
  assign data_o[11277] = data_o[13];
  assign data_o[11341] = data_o[13];
  assign data_o[11405] = data_o[13];
  assign data_o[11469] = data_o[13];
  assign data_o[11533] = data_o[13];
  assign data_o[11597] = data_o[13];
  assign data_o[11661] = data_o[13];
  assign data_o[11725] = data_o[13];
  assign data_o[11789] = data_o[13];
  assign data_o[11853] = data_o[13];
  assign data_o[11917] = data_o[13];
  assign data_o[11981] = data_o[13];
  assign data_o[12045] = data_o[13];
  assign data_o[12109] = data_o[13];
  assign data_o[12173] = data_o[13];
  assign data_o[12237] = data_o[13];
  assign data_o[12301] = data_o[13];
  assign data_o[12365] = data_o[13];
  assign data_o[12429] = data_o[13];
  assign data_o[12493] = data_o[13];
  assign data_o[12557] = data_o[13];
  assign data_o[12621] = data_o[13];
  assign data_o[12685] = data_o[13];
  assign data_o[12749] = data_o[13];
  assign data_o[12813] = data_o[13];
  assign data_o[12877] = data_o[13];
  assign data_o[12941] = data_o[13];
  assign data_o[13005] = data_o[13];
  assign data_o[13069] = data_o[13];
  assign data_o[13133] = data_o[13];
  assign data_o[13197] = data_o[13];
  assign data_o[13261] = data_o[13];
  assign data_o[13325] = data_o[13];
  assign data_o[13389] = data_o[13];
  assign data_o[13453] = data_o[13];
  assign data_o[13517] = data_o[13];
  assign data_o[13581] = data_o[13];
  assign data_o[13645] = data_o[13];
  assign data_o[13709] = data_o[13];
  assign data_o[13773] = data_o[13];
  assign data_o[13837] = data_o[13];
  assign data_o[13901] = data_o[13];
  assign data_o[13965] = data_o[13];
  assign data_o[14029] = data_o[13];
  assign data_o[14093] = data_o[13];
  assign data_o[14157] = data_o[13];
  assign data_o[14221] = data_o[13];
  assign data_o[14285] = data_o[13];
  assign data_o[14349] = data_o[13];
  assign data_o[14413] = data_o[13];
  assign data_o[14477] = data_o[13];
  assign data_o[14541] = data_o[13];
  assign data_o[14605] = data_o[13];
  assign data_o[14669] = data_o[13];
  assign data_o[14733] = data_o[13];
  assign data_o[14797] = data_o[13];
  assign data_o[14861] = data_o[13];
  assign data_o[14925] = data_o[13];
  assign data_o[14989] = data_o[13];
  assign data_o[15053] = data_o[13];
  assign data_o[15117] = data_o[13];
  assign data_o[15181] = data_o[13];
  assign data_o[15245] = data_o[13];
  assign data_o[15309] = data_o[13];
  assign data_o[15373] = data_o[13];
  assign data_o[15437] = data_o[13];
  assign data_o[15501] = data_o[13];
  assign data_o[15565] = data_o[13];
  assign data_o[15629] = data_o[13];
  assign data_o[15693] = data_o[13];
  assign data_o[15757] = data_o[13];
  assign data_o[15821] = data_o[13];
  assign data_o[15885] = data_o[13];
  assign data_o[15949] = data_o[13];
  assign data_o[16013] = data_o[13];
  assign data_o[16077] = data_o[13];
  assign data_o[16141] = data_o[13];
  assign data_o[16205] = data_o[13];
  assign data_o[16269] = data_o[13];
  assign data_o[16333] = data_o[13];
  assign data_o[16397] = data_o[13];
  assign data_o[16461] = data_o[13];
  assign data_o[16525] = data_o[13];
  assign data_o[16589] = data_o[13];
  assign data_o[16653] = data_o[13];
  assign data_o[16717] = data_o[13];
  assign data_o[16781] = data_o[13];
  assign data_o[16845] = data_o[13];
  assign data_o[16909] = data_o[13];
  assign data_o[16973] = data_o[13];
  assign data_o[17037] = data_o[13];
  assign data_o[17101] = data_o[13];
  assign data_o[17165] = data_o[13];
  assign data_o[17229] = data_o[13];
  assign data_o[17293] = data_o[13];
  assign data_o[17357] = data_o[13];
  assign data_o[17421] = data_o[13];
  assign data_o[17485] = data_o[13];
  assign data_o[17549] = data_o[13];
  assign data_o[17613] = data_o[13];
  assign data_o[17677] = data_o[13];
  assign data_o[17741] = data_o[13];
  assign data_o[17805] = data_o[13];
  assign data_o[17869] = data_o[13];
  assign data_o[17933] = data_o[13];
  assign data_o[17997] = data_o[13];
  assign data_o[18061] = data_o[13];
  assign data_o[18125] = data_o[13];
  assign data_o[18189] = data_o[13];
  assign data_o[18253] = data_o[13];
  assign data_o[18317] = data_o[13];
  assign data_o[18381] = data_o[13];
  assign data_o[18445] = data_o[13];
  assign data_o[18509] = data_o[13];
  assign data_o[18573] = data_o[13];
  assign data_o[18637] = data_o[13];
  assign data_o[18701] = data_o[13];
  assign data_o[18765] = data_o[13];
  assign data_o[18829] = data_o[13];
  assign data_o[18893] = data_o[13];
  assign data_o[18957] = data_o[13];
  assign data_o[19021] = data_o[13];
  assign data_o[19085] = data_o[13];
  assign data_o[19149] = data_o[13];
  assign data_o[19213] = data_o[13];
  assign data_o[19277] = data_o[13];
  assign data_o[19341] = data_o[13];
  assign data_o[19405] = data_o[13];
  assign data_o[19469] = data_o[13];
  assign data_o[19533] = data_o[13];
  assign data_o[19597] = data_o[13];
  assign data_o[19661] = data_o[13];
  assign data_o[19725] = data_o[13];
  assign data_o[19789] = data_o[13];
  assign data_o[19853] = data_o[13];
  assign data_o[19917] = data_o[13];
  assign data_o[19981] = data_o[13];
  assign data_o[20045] = data_o[13];
  assign data_o[20109] = data_o[13];
  assign data_o[20173] = data_o[13];
  assign data_o[20237] = data_o[13];
  assign data_o[20301] = data_o[13];
  assign data_o[20365] = data_o[13];
  assign data_o[20429] = data_o[13];
  assign data_o[20493] = data_o[13];
  assign data_o[20557] = data_o[13];
  assign data_o[20621] = data_o[13];
  assign data_o[20685] = data_o[13];
  assign data_o[20749] = data_o[13];
  assign data_o[20813] = data_o[13];
  assign data_o[20877] = data_o[13];
  assign data_o[20941] = data_o[13];
  assign data_o[21005] = data_o[13];
  assign data_o[21069] = data_o[13];
  assign data_o[21133] = data_o[13];
  assign data_o[21197] = data_o[13];
  assign data_o[21261] = data_o[13];
  assign data_o[21325] = data_o[13];
  assign data_o[21389] = data_o[13];
  assign data_o[21453] = data_o[13];
  assign data_o[21517] = data_o[13];
  assign data_o[21581] = data_o[13];
  assign data_o[21645] = data_o[13];
  assign data_o[21709] = data_o[13];
  assign data_o[21773] = data_o[13];
  assign data_o[21837] = data_o[13];
  assign data_o[21901] = data_o[13];
  assign data_o[21965] = data_o[13];
  assign data_o[22029] = data_o[13];
  assign data_o[22093] = data_o[13];
  assign data_o[22157] = data_o[13];
  assign data_o[22221] = data_o[13];
  assign data_o[22285] = data_o[13];
  assign data_o[22349] = data_o[13];
  assign data_o[22413] = data_o[13];
  assign data_o[22477] = data_o[13];
  assign data_o[22541] = data_o[13];
  assign data_o[22605] = data_o[13];
  assign data_o[22669] = data_o[13];
  assign data_o[22733] = data_o[13];
  assign data_o[22797] = data_o[13];
  assign data_o[22861] = data_o[13];
  assign data_o[22925] = data_o[13];
  assign data_o[22989] = data_o[13];
  assign data_o[23053] = data_o[13];
  assign data_o[23117] = data_o[13];
  assign data_o[23181] = data_o[13];
  assign data_o[23245] = data_o[13];
  assign data_o[23309] = data_o[13];
  assign data_o[23373] = data_o[13];
  assign data_o[23437] = data_o[13];
  assign data_o[23501] = data_o[13];
  assign data_o[23565] = data_o[13];
  assign data_o[23629] = data_o[13];
  assign data_o[23693] = data_o[13];
  assign data_o[23757] = data_o[13];
  assign data_o[23821] = data_o[13];
  assign data_o[23885] = data_o[13];
  assign data_o[23949] = data_o[13];
  assign data_o[24013] = data_o[13];
  assign data_o[24077] = data_o[13];
  assign data_o[24141] = data_o[13];
  assign data_o[24205] = data_o[13];
  assign data_o[24269] = data_o[13];
  assign data_o[24333] = data_o[13];
  assign data_o[24397] = data_o[13];
  assign data_o[24461] = data_o[13];
  assign data_o[24525] = data_o[13];
  assign data_o[24589] = data_o[13];
  assign data_o[24653] = data_o[13];
  assign data_o[24717] = data_o[13];
  assign data_o[24781] = data_o[13];
  assign data_o[24845] = data_o[13];
  assign data_o[24909] = data_o[13];
  assign data_o[24973] = data_o[13];
  assign data_o[25037] = data_o[13];
  assign data_o[25101] = data_o[13];
  assign data_o[25165] = data_o[13];
  assign data_o[25229] = data_o[13];
  assign data_o[25293] = data_o[13];
  assign data_o[25357] = data_o[13];
  assign data_o[25421] = data_o[13];
  assign data_o[25485] = data_o[13];
  assign data_o[25549] = data_o[13];
  assign data_o[25613] = data_o[13];
  assign data_o[25677] = data_o[13];
  assign data_o[25741] = data_o[13];
  assign data_o[25805] = data_o[13];
  assign data_o[25869] = data_o[13];
  assign data_o[25933] = data_o[13];
  assign data_o[25997] = data_o[13];
  assign data_o[26061] = data_o[13];
  assign data_o[26125] = data_o[13];
  assign data_o[26189] = data_o[13];
  assign data_o[26253] = data_o[13];
  assign data_o[26317] = data_o[13];
  assign data_o[26381] = data_o[13];
  assign data_o[26445] = data_o[13];
  assign data_o[26509] = data_o[13];
  assign data_o[26573] = data_o[13];
  assign data_o[26637] = data_o[13];
  assign data_o[26701] = data_o[13];
  assign data_o[26765] = data_o[13];
  assign data_o[26829] = data_o[13];
  assign data_o[26893] = data_o[13];
  assign data_o[26957] = data_o[13];
  assign data_o[27021] = data_o[13];
  assign data_o[27085] = data_o[13];
  assign data_o[27149] = data_o[13];
  assign data_o[27213] = data_o[13];
  assign data_o[27277] = data_o[13];
  assign data_o[27341] = data_o[13];
  assign data_o[27405] = data_o[13];
  assign data_o[27469] = data_o[13];
  assign data_o[27533] = data_o[13];
  assign data_o[27597] = data_o[13];
  assign data_o[27661] = data_o[13];
  assign data_o[27725] = data_o[13];
  assign data_o[27789] = data_o[13];
  assign data_o[27853] = data_o[13];
  assign data_o[27917] = data_o[13];
  assign data_o[27981] = data_o[13];
  assign data_o[28045] = data_o[13];
  assign data_o[28109] = data_o[13];
  assign data_o[28173] = data_o[13];
  assign data_o[28237] = data_o[13];
  assign data_o[28301] = data_o[13];
  assign data_o[28365] = data_o[13];
  assign data_o[28429] = data_o[13];
  assign data_o[28493] = data_o[13];
  assign data_o[28557] = data_o[13];
  assign data_o[28621] = data_o[13];
  assign data_o[28685] = data_o[13];
  assign data_o[28749] = data_o[13];
  assign data_o[28813] = data_o[13];
  assign data_o[28877] = data_o[13];
  assign data_o[28941] = data_o[13];
  assign data_o[29005] = data_o[13];
  assign data_o[29069] = data_o[13];
  assign data_o[29133] = data_o[13];
  assign data_o[29197] = data_o[13];
  assign data_o[29261] = data_o[13];
  assign data_o[29325] = data_o[13];
  assign data_o[29389] = data_o[13];
  assign data_o[29453] = data_o[13];
  assign data_o[29517] = data_o[13];
  assign data_o[29581] = data_o[13];
  assign data_o[29645] = data_o[13];
  assign data_o[29709] = data_o[13];
  assign data_o[29773] = data_o[13];
  assign data_o[29837] = data_o[13];
  assign data_o[29901] = data_o[13];
  assign data_o[29965] = data_o[13];
  assign data_o[30029] = data_o[13];
  assign data_o[30093] = data_o[13];
  assign data_o[30157] = data_o[13];
  assign data_o[30221] = data_o[13];
  assign data_o[30285] = data_o[13];
  assign data_o[30349] = data_o[13];
  assign data_o[30413] = data_o[13];
  assign data_o[30477] = data_o[13];
  assign data_o[30541] = data_o[13];
  assign data_o[30605] = data_o[13];
  assign data_o[30669] = data_o[13];
  assign data_o[30733] = data_o[13];
  assign data_o[30797] = data_o[13];
  assign data_o[30861] = data_o[13];
  assign data_o[30925] = data_o[13];
  assign data_o[30989] = data_o[13];
  assign data_o[31053] = data_o[13];
  assign data_o[31117] = data_o[13];
  assign data_o[31181] = data_o[13];
  assign data_o[31245] = data_o[13];
  assign data_o[31309] = data_o[13];
  assign data_o[31373] = data_o[13];
  assign data_o[31437] = data_o[13];
  assign data_o[31501] = data_o[13];
  assign data_o[31565] = data_o[13];
  assign data_o[31629] = data_o[13];
  assign data_o[31693] = data_o[13];
  assign data_o[31757] = data_o[13];
  assign data_o[31821] = data_o[13];
  assign data_o[31885] = data_o[13];
  assign data_o[31949] = data_o[13];
  assign data_o[76] = data_o[12];
  assign data_o[140] = data_o[12];
  assign data_o[204] = data_o[12];
  assign data_o[268] = data_o[12];
  assign data_o[332] = data_o[12];
  assign data_o[396] = data_o[12];
  assign data_o[460] = data_o[12];
  assign data_o[524] = data_o[12];
  assign data_o[588] = data_o[12];
  assign data_o[652] = data_o[12];
  assign data_o[716] = data_o[12];
  assign data_o[780] = data_o[12];
  assign data_o[844] = data_o[12];
  assign data_o[908] = data_o[12];
  assign data_o[972] = data_o[12];
  assign data_o[1036] = data_o[12];
  assign data_o[1100] = data_o[12];
  assign data_o[1164] = data_o[12];
  assign data_o[1228] = data_o[12];
  assign data_o[1292] = data_o[12];
  assign data_o[1356] = data_o[12];
  assign data_o[1420] = data_o[12];
  assign data_o[1484] = data_o[12];
  assign data_o[1548] = data_o[12];
  assign data_o[1612] = data_o[12];
  assign data_o[1676] = data_o[12];
  assign data_o[1740] = data_o[12];
  assign data_o[1804] = data_o[12];
  assign data_o[1868] = data_o[12];
  assign data_o[1932] = data_o[12];
  assign data_o[1996] = data_o[12];
  assign data_o[2060] = data_o[12];
  assign data_o[2124] = data_o[12];
  assign data_o[2188] = data_o[12];
  assign data_o[2252] = data_o[12];
  assign data_o[2316] = data_o[12];
  assign data_o[2380] = data_o[12];
  assign data_o[2444] = data_o[12];
  assign data_o[2508] = data_o[12];
  assign data_o[2572] = data_o[12];
  assign data_o[2636] = data_o[12];
  assign data_o[2700] = data_o[12];
  assign data_o[2764] = data_o[12];
  assign data_o[2828] = data_o[12];
  assign data_o[2892] = data_o[12];
  assign data_o[2956] = data_o[12];
  assign data_o[3020] = data_o[12];
  assign data_o[3084] = data_o[12];
  assign data_o[3148] = data_o[12];
  assign data_o[3212] = data_o[12];
  assign data_o[3276] = data_o[12];
  assign data_o[3340] = data_o[12];
  assign data_o[3404] = data_o[12];
  assign data_o[3468] = data_o[12];
  assign data_o[3532] = data_o[12];
  assign data_o[3596] = data_o[12];
  assign data_o[3660] = data_o[12];
  assign data_o[3724] = data_o[12];
  assign data_o[3788] = data_o[12];
  assign data_o[3852] = data_o[12];
  assign data_o[3916] = data_o[12];
  assign data_o[3980] = data_o[12];
  assign data_o[4044] = data_o[12];
  assign data_o[4108] = data_o[12];
  assign data_o[4172] = data_o[12];
  assign data_o[4236] = data_o[12];
  assign data_o[4300] = data_o[12];
  assign data_o[4364] = data_o[12];
  assign data_o[4428] = data_o[12];
  assign data_o[4492] = data_o[12];
  assign data_o[4556] = data_o[12];
  assign data_o[4620] = data_o[12];
  assign data_o[4684] = data_o[12];
  assign data_o[4748] = data_o[12];
  assign data_o[4812] = data_o[12];
  assign data_o[4876] = data_o[12];
  assign data_o[4940] = data_o[12];
  assign data_o[5004] = data_o[12];
  assign data_o[5068] = data_o[12];
  assign data_o[5132] = data_o[12];
  assign data_o[5196] = data_o[12];
  assign data_o[5260] = data_o[12];
  assign data_o[5324] = data_o[12];
  assign data_o[5388] = data_o[12];
  assign data_o[5452] = data_o[12];
  assign data_o[5516] = data_o[12];
  assign data_o[5580] = data_o[12];
  assign data_o[5644] = data_o[12];
  assign data_o[5708] = data_o[12];
  assign data_o[5772] = data_o[12];
  assign data_o[5836] = data_o[12];
  assign data_o[5900] = data_o[12];
  assign data_o[5964] = data_o[12];
  assign data_o[6028] = data_o[12];
  assign data_o[6092] = data_o[12];
  assign data_o[6156] = data_o[12];
  assign data_o[6220] = data_o[12];
  assign data_o[6284] = data_o[12];
  assign data_o[6348] = data_o[12];
  assign data_o[6412] = data_o[12];
  assign data_o[6476] = data_o[12];
  assign data_o[6540] = data_o[12];
  assign data_o[6604] = data_o[12];
  assign data_o[6668] = data_o[12];
  assign data_o[6732] = data_o[12];
  assign data_o[6796] = data_o[12];
  assign data_o[6860] = data_o[12];
  assign data_o[6924] = data_o[12];
  assign data_o[6988] = data_o[12];
  assign data_o[7052] = data_o[12];
  assign data_o[7116] = data_o[12];
  assign data_o[7180] = data_o[12];
  assign data_o[7244] = data_o[12];
  assign data_o[7308] = data_o[12];
  assign data_o[7372] = data_o[12];
  assign data_o[7436] = data_o[12];
  assign data_o[7500] = data_o[12];
  assign data_o[7564] = data_o[12];
  assign data_o[7628] = data_o[12];
  assign data_o[7692] = data_o[12];
  assign data_o[7756] = data_o[12];
  assign data_o[7820] = data_o[12];
  assign data_o[7884] = data_o[12];
  assign data_o[7948] = data_o[12];
  assign data_o[8012] = data_o[12];
  assign data_o[8076] = data_o[12];
  assign data_o[8140] = data_o[12];
  assign data_o[8204] = data_o[12];
  assign data_o[8268] = data_o[12];
  assign data_o[8332] = data_o[12];
  assign data_o[8396] = data_o[12];
  assign data_o[8460] = data_o[12];
  assign data_o[8524] = data_o[12];
  assign data_o[8588] = data_o[12];
  assign data_o[8652] = data_o[12];
  assign data_o[8716] = data_o[12];
  assign data_o[8780] = data_o[12];
  assign data_o[8844] = data_o[12];
  assign data_o[8908] = data_o[12];
  assign data_o[8972] = data_o[12];
  assign data_o[9036] = data_o[12];
  assign data_o[9100] = data_o[12];
  assign data_o[9164] = data_o[12];
  assign data_o[9228] = data_o[12];
  assign data_o[9292] = data_o[12];
  assign data_o[9356] = data_o[12];
  assign data_o[9420] = data_o[12];
  assign data_o[9484] = data_o[12];
  assign data_o[9548] = data_o[12];
  assign data_o[9612] = data_o[12];
  assign data_o[9676] = data_o[12];
  assign data_o[9740] = data_o[12];
  assign data_o[9804] = data_o[12];
  assign data_o[9868] = data_o[12];
  assign data_o[9932] = data_o[12];
  assign data_o[9996] = data_o[12];
  assign data_o[10060] = data_o[12];
  assign data_o[10124] = data_o[12];
  assign data_o[10188] = data_o[12];
  assign data_o[10252] = data_o[12];
  assign data_o[10316] = data_o[12];
  assign data_o[10380] = data_o[12];
  assign data_o[10444] = data_o[12];
  assign data_o[10508] = data_o[12];
  assign data_o[10572] = data_o[12];
  assign data_o[10636] = data_o[12];
  assign data_o[10700] = data_o[12];
  assign data_o[10764] = data_o[12];
  assign data_o[10828] = data_o[12];
  assign data_o[10892] = data_o[12];
  assign data_o[10956] = data_o[12];
  assign data_o[11020] = data_o[12];
  assign data_o[11084] = data_o[12];
  assign data_o[11148] = data_o[12];
  assign data_o[11212] = data_o[12];
  assign data_o[11276] = data_o[12];
  assign data_o[11340] = data_o[12];
  assign data_o[11404] = data_o[12];
  assign data_o[11468] = data_o[12];
  assign data_o[11532] = data_o[12];
  assign data_o[11596] = data_o[12];
  assign data_o[11660] = data_o[12];
  assign data_o[11724] = data_o[12];
  assign data_o[11788] = data_o[12];
  assign data_o[11852] = data_o[12];
  assign data_o[11916] = data_o[12];
  assign data_o[11980] = data_o[12];
  assign data_o[12044] = data_o[12];
  assign data_o[12108] = data_o[12];
  assign data_o[12172] = data_o[12];
  assign data_o[12236] = data_o[12];
  assign data_o[12300] = data_o[12];
  assign data_o[12364] = data_o[12];
  assign data_o[12428] = data_o[12];
  assign data_o[12492] = data_o[12];
  assign data_o[12556] = data_o[12];
  assign data_o[12620] = data_o[12];
  assign data_o[12684] = data_o[12];
  assign data_o[12748] = data_o[12];
  assign data_o[12812] = data_o[12];
  assign data_o[12876] = data_o[12];
  assign data_o[12940] = data_o[12];
  assign data_o[13004] = data_o[12];
  assign data_o[13068] = data_o[12];
  assign data_o[13132] = data_o[12];
  assign data_o[13196] = data_o[12];
  assign data_o[13260] = data_o[12];
  assign data_o[13324] = data_o[12];
  assign data_o[13388] = data_o[12];
  assign data_o[13452] = data_o[12];
  assign data_o[13516] = data_o[12];
  assign data_o[13580] = data_o[12];
  assign data_o[13644] = data_o[12];
  assign data_o[13708] = data_o[12];
  assign data_o[13772] = data_o[12];
  assign data_o[13836] = data_o[12];
  assign data_o[13900] = data_o[12];
  assign data_o[13964] = data_o[12];
  assign data_o[14028] = data_o[12];
  assign data_o[14092] = data_o[12];
  assign data_o[14156] = data_o[12];
  assign data_o[14220] = data_o[12];
  assign data_o[14284] = data_o[12];
  assign data_o[14348] = data_o[12];
  assign data_o[14412] = data_o[12];
  assign data_o[14476] = data_o[12];
  assign data_o[14540] = data_o[12];
  assign data_o[14604] = data_o[12];
  assign data_o[14668] = data_o[12];
  assign data_o[14732] = data_o[12];
  assign data_o[14796] = data_o[12];
  assign data_o[14860] = data_o[12];
  assign data_o[14924] = data_o[12];
  assign data_o[14988] = data_o[12];
  assign data_o[15052] = data_o[12];
  assign data_o[15116] = data_o[12];
  assign data_o[15180] = data_o[12];
  assign data_o[15244] = data_o[12];
  assign data_o[15308] = data_o[12];
  assign data_o[15372] = data_o[12];
  assign data_o[15436] = data_o[12];
  assign data_o[15500] = data_o[12];
  assign data_o[15564] = data_o[12];
  assign data_o[15628] = data_o[12];
  assign data_o[15692] = data_o[12];
  assign data_o[15756] = data_o[12];
  assign data_o[15820] = data_o[12];
  assign data_o[15884] = data_o[12];
  assign data_o[15948] = data_o[12];
  assign data_o[16012] = data_o[12];
  assign data_o[16076] = data_o[12];
  assign data_o[16140] = data_o[12];
  assign data_o[16204] = data_o[12];
  assign data_o[16268] = data_o[12];
  assign data_o[16332] = data_o[12];
  assign data_o[16396] = data_o[12];
  assign data_o[16460] = data_o[12];
  assign data_o[16524] = data_o[12];
  assign data_o[16588] = data_o[12];
  assign data_o[16652] = data_o[12];
  assign data_o[16716] = data_o[12];
  assign data_o[16780] = data_o[12];
  assign data_o[16844] = data_o[12];
  assign data_o[16908] = data_o[12];
  assign data_o[16972] = data_o[12];
  assign data_o[17036] = data_o[12];
  assign data_o[17100] = data_o[12];
  assign data_o[17164] = data_o[12];
  assign data_o[17228] = data_o[12];
  assign data_o[17292] = data_o[12];
  assign data_o[17356] = data_o[12];
  assign data_o[17420] = data_o[12];
  assign data_o[17484] = data_o[12];
  assign data_o[17548] = data_o[12];
  assign data_o[17612] = data_o[12];
  assign data_o[17676] = data_o[12];
  assign data_o[17740] = data_o[12];
  assign data_o[17804] = data_o[12];
  assign data_o[17868] = data_o[12];
  assign data_o[17932] = data_o[12];
  assign data_o[17996] = data_o[12];
  assign data_o[18060] = data_o[12];
  assign data_o[18124] = data_o[12];
  assign data_o[18188] = data_o[12];
  assign data_o[18252] = data_o[12];
  assign data_o[18316] = data_o[12];
  assign data_o[18380] = data_o[12];
  assign data_o[18444] = data_o[12];
  assign data_o[18508] = data_o[12];
  assign data_o[18572] = data_o[12];
  assign data_o[18636] = data_o[12];
  assign data_o[18700] = data_o[12];
  assign data_o[18764] = data_o[12];
  assign data_o[18828] = data_o[12];
  assign data_o[18892] = data_o[12];
  assign data_o[18956] = data_o[12];
  assign data_o[19020] = data_o[12];
  assign data_o[19084] = data_o[12];
  assign data_o[19148] = data_o[12];
  assign data_o[19212] = data_o[12];
  assign data_o[19276] = data_o[12];
  assign data_o[19340] = data_o[12];
  assign data_o[19404] = data_o[12];
  assign data_o[19468] = data_o[12];
  assign data_o[19532] = data_o[12];
  assign data_o[19596] = data_o[12];
  assign data_o[19660] = data_o[12];
  assign data_o[19724] = data_o[12];
  assign data_o[19788] = data_o[12];
  assign data_o[19852] = data_o[12];
  assign data_o[19916] = data_o[12];
  assign data_o[19980] = data_o[12];
  assign data_o[20044] = data_o[12];
  assign data_o[20108] = data_o[12];
  assign data_o[20172] = data_o[12];
  assign data_o[20236] = data_o[12];
  assign data_o[20300] = data_o[12];
  assign data_o[20364] = data_o[12];
  assign data_o[20428] = data_o[12];
  assign data_o[20492] = data_o[12];
  assign data_o[20556] = data_o[12];
  assign data_o[20620] = data_o[12];
  assign data_o[20684] = data_o[12];
  assign data_o[20748] = data_o[12];
  assign data_o[20812] = data_o[12];
  assign data_o[20876] = data_o[12];
  assign data_o[20940] = data_o[12];
  assign data_o[21004] = data_o[12];
  assign data_o[21068] = data_o[12];
  assign data_o[21132] = data_o[12];
  assign data_o[21196] = data_o[12];
  assign data_o[21260] = data_o[12];
  assign data_o[21324] = data_o[12];
  assign data_o[21388] = data_o[12];
  assign data_o[21452] = data_o[12];
  assign data_o[21516] = data_o[12];
  assign data_o[21580] = data_o[12];
  assign data_o[21644] = data_o[12];
  assign data_o[21708] = data_o[12];
  assign data_o[21772] = data_o[12];
  assign data_o[21836] = data_o[12];
  assign data_o[21900] = data_o[12];
  assign data_o[21964] = data_o[12];
  assign data_o[22028] = data_o[12];
  assign data_o[22092] = data_o[12];
  assign data_o[22156] = data_o[12];
  assign data_o[22220] = data_o[12];
  assign data_o[22284] = data_o[12];
  assign data_o[22348] = data_o[12];
  assign data_o[22412] = data_o[12];
  assign data_o[22476] = data_o[12];
  assign data_o[22540] = data_o[12];
  assign data_o[22604] = data_o[12];
  assign data_o[22668] = data_o[12];
  assign data_o[22732] = data_o[12];
  assign data_o[22796] = data_o[12];
  assign data_o[22860] = data_o[12];
  assign data_o[22924] = data_o[12];
  assign data_o[22988] = data_o[12];
  assign data_o[23052] = data_o[12];
  assign data_o[23116] = data_o[12];
  assign data_o[23180] = data_o[12];
  assign data_o[23244] = data_o[12];
  assign data_o[23308] = data_o[12];
  assign data_o[23372] = data_o[12];
  assign data_o[23436] = data_o[12];
  assign data_o[23500] = data_o[12];
  assign data_o[23564] = data_o[12];
  assign data_o[23628] = data_o[12];
  assign data_o[23692] = data_o[12];
  assign data_o[23756] = data_o[12];
  assign data_o[23820] = data_o[12];
  assign data_o[23884] = data_o[12];
  assign data_o[23948] = data_o[12];
  assign data_o[24012] = data_o[12];
  assign data_o[24076] = data_o[12];
  assign data_o[24140] = data_o[12];
  assign data_o[24204] = data_o[12];
  assign data_o[24268] = data_o[12];
  assign data_o[24332] = data_o[12];
  assign data_o[24396] = data_o[12];
  assign data_o[24460] = data_o[12];
  assign data_o[24524] = data_o[12];
  assign data_o[24588] = data_o[12];
  assign data_o[24652] = data_o[12];
  assign data_o[24716] = data_o[12];
  assign data_o[24780] = data_o[12];
  assign data_o[24844] = data_o[12];
  assign data_o[24908] = data_o[12];
  assign data_o[24972] = data_o[12];
  assign data_o[25036] = data_o[12];
  assign data_o[25100] = data_o[12];
  assign data_o[25164] = data_o[12];
  assign data_o[25228] = data_o[12];
  assign data_o[25292] = data_o[12];
  assign data_o[25356] = data_o[12];
  assign data_o[25420] = data_o[12];
  assign data_o[25484] = data_o[12];
  assign data_o[25548] = data_o[12];
  assign data_o[25612] = data_o[12];
  assign data_o[25676] = data_o[12];
  assign data_o[25740] = data_o[12];
  assign data_o[25804] = data_o[12];
  assign data_o[25868] = data_o[12];
  assign data_o[25932] = data_o[12];
  assign data_o[25996] = data_o[12];
  assign data_o[26060] = data_o[12];
  assign data_o[26124] = data_o[12];
  assign data_o[26188] = data_o[12];
  assign data_o[26252] = data_o[12];
  assign data_o[26316] = data_o[12];
  assign data_o[26380] = data_o[12];
  assign data_o[26444] = data_o[12];
  assign data_o[26508] = data_o[12];
  assign data_o[26572] = data_o[12];
  assign data_o[26636] = data_o[12];
  assign data_o[26700] = data_o[12];
  assign data_o[26764] = data_o[12];
  assign data_o[26828] = data_o[12];
  assign data_o[26892] = data_o[12];
  assign data_o[26956] = data_o[12];
  assign data_o[27020] = data_o[12];
  assign data_o[27084] = data_o[12];
  assign data_o[27148] = data_o[12];
  assign data_o[27212] = data_o[12];
  assign data_o[27276] = data_o[12];
  assign data_o[27340] = data_o[12];
  assign data_o[27404] = data_o[12];
  assign data_o[27468] = data_o[12];
  assign data_o[27532] = data_o[12];
  assign data_o[27596] = data_o[12];
  assign data_o[27660] = data_o[12];
  assign data_o[27724] = data_o[12];
  assign data_o[27788] = data_o[12];
  assign data_o[27852] = data_o[12];
  assign data_o[27916] = data_o[12];
  assign data_o[27980] = data_o[12];
  assign data_o[28044] = data_o[12];
  assign data_o[28108] = data_o[12];
  assign data_o[28172] = data_o[12];
  assign data_o[28236] = data_o[12];
  assign data_o[28300] = data_o[12];
  assign data_o[28364] = data_o[12];
  assign data_o[28428] = data_o[12];
  assign data_o[28492] = data_o[12];
  assign data_o[28556] = data_o[12];
  assign data_o[28620] = data_o[12];
  assign data_o[28684] = data_o[12];
  assign data_o[28748] = data_o[12];
  assign data_o[28812] = data_o[12];
  assign data_o[28876] = data_o[12];
  assign data_o[28940] = data_o[12];
  assign data_o[29004] = data_o[12];
  assign data_o[29068] = data_o[12];
  assign data_o[29132] = data_o[12];
  assign data_o[29196] = data_o[12];
  assign data_o[29260] = data_o[12];
  assign data_o[29324] = data_o[12];
  assign data_o[29388] = data_o[12];
  assign data_o[29452] = data_o[12];
  assign data_o[29516] = data_o[12];
  assign data_o[29580] = data_o[12];
  assign data_o[29644] = data_o[12];
  assign data_o[29708] = data_o[12];
  assign data_o[29772] = data_o[12];
  assign data_o[29836] = data_o[12];
  assign data_o[29900] = data_o[12];
  assign data_o[29964] = data_o[12];
  assign data_o[30028] = data_o[12];
  assign data_o[30092] = data_o[12];
  assign data_o[30156] = data_o[12];
  assign data_o[30220] = data_o[12];
  assign data_o[30284] = data_o[12];
  assign data_o[30348] = data_o[12];
  assign data_o[30412] = data_o[12];
  assign data_o[30476] = data_o[12];
  assign data_o[30540] = data_o[12];
  assign data_o[30604] = data_o[12];
  assign data_o[30668] = data_o[12];
  assign data_o[30732] = data_o[12];
  assign data_o[30796] = data_o[12];
  assign data_o[30860] = data_o[12];
  assign data_o[30924] = data_o[12];
  assign data_o[30988] = data_o[12];
  assign data_o[31052] = data_o[12];
  assign data_o[31116] = data_o[12];
  assign data_o[31180] = data_o[12];
  assign data_o[31244] = data_o[12];
  assign data_o[31308] = data_o[12];
  assign data_o[31372] = data_o[12];
  assign data_o[31436] = data_o[12];
  assign data_o[31500] = data_o[12];
  assign data_o[31564] = data_o[12];
  assign data_o[31628] = data_o[12];
  assign data_o[31692] = data_o[12];
  assign data_o[31756] = data_o[12];
  assign data_o[31820] = data_o[12];
  assign data_o[31884] = data_o[12];
  assign data_o[31948] = data_o[12];
  assign data_o[75] = data_o[11];
  assign data_o[139] = data_o[11];
  assign data_o[203] = data_o[11];
  assign data_o[267] = data_o[11];
  assign data_o[331] = data_o[11];
  assign data_o[395] = data_o[11];
  assign data_o[459] = data_o[11];
  assign data_o[523] = data_o[11];
  assign data_o[587] = data_o[11];
  assign data_o[651] = data_o[11];
  assign data_o[715] = data_o[11];
  assign data_o[779] = data_o[11];
  assign data_o[843] = data_o[11];
  assign data_o[907] = data_o[11];
  assign data_o[971] = data_o[11];
  assign data_o[1035] = data_o[11];
  assign data_o[1099] = data_o[11];
  assign data_o[1163] = data_o[11];
  assign data_o[1227] = data_o[11];
  assign data_o[1291] = data_o[11];
  assign data_o[1355] = data_o[11];
  assign data_o[1419] = data_o[11];
  assign data_o[1483] = data_o[11];
  assign data_o[1547] = data_o[11];
  assign data_o[1611] = data_o[11];
  assign data_o[1675] = data_o[11];
  assign data_o[1739] = data_o[11];
  assign data_o[1803] = data_o[11];
  assign data_o[1867] = data_o[11];
  assign data_o[1931] = data_o[11];
  assign data_o[1995] = data_o[11];
  assign data_o[2059] = data_o[11];
  assign data_o[2123] = data_o[11];
  assign data_o[2187] = data_o[11];
  assign data_o[2251] = data_o[11];
  assign data_o[2315] = data_o[11];
  assign data_o[2379] = data_o[11];
  assign data_o[2443] = data_o[11];
  assign data_o[2507] = data_o[11];
  assign data_o[2571] = data_o[11];
  assign data_o[2635] = data_o[11];
  assign data_o[2699] = data_o[11];
  assign data_o[2763] = data_o[11];
  assign data_o[2827] = data_o[11];
  assign data_o[2891] = data_o[11];
  assign data_o[2955] = data_o[11];
  assign data_o[3019] = data_o[11];
  assign data_o[3083] = data_o[11];
  assign data_o[3147] = data_o[11];
  assign data_o[3211] = data_o[11];
  assign data_o[3275] = data_o[11];
  assign data_o[3339] = data_o[11];
  assign data_o[3403] = data_o[11];
  assign data_o[3467] = data_o[11];
  assign data_o[3531] = data_o[11];
  assign data_o[3595] = data_o[11];
  assign data_o[3659] = data_o[11];
  assign data_o[3723] = data_o[11];
  assign data_o[3787] = data_o[11];
  assign data_o[3851] = data_o[11];
  assign data_o[3915] = data_o[11];
  assign data_o[3979] = data_o[11];
  assign data_o[4043] = data_o[11];
  assign data_o[4107] = data_o[11];
  assign data_o[4171] = data_o[11];
  assign data_o[4235] = data_o[11];
  assign data_o[4299] = data_o[11];
  assign data_o[4363] = data_o[11];
  assign data_o[4427] = data_o[11];
  assign data_o[4491] = data_o[11];
  assign data_o[4555] = data_o[11];
  assign data_o[4619] = data_o[11];
  assign data_o[4683] = data_o[11];
  assign data_o[4747] = data_o[11];
  assign data_o[4811] = data_o[11];
  assign data_o[4875] = data_o[11];
  assign data_o[4939] = data_o[11];
  assign data_o[5003] = data_o[11];
  assign data_o[5067] = data_o[11];
  assign data_o[5131] = data_o[11];
  assign data_o[5195] = data_o[11];
  assign data_o[5259] = data_o[11];
  assign data_o[5323] = data_o[11];
  assign data_o[5387] = data_o[11];
  assign data_o[5451] = data_o[11];
  assign data_o[5515] = data_o[11];
  assign data_o[5579] = data_o[11];
  assign data_o[5643] = data_o[11];
  assign data_o[5707] = data_o[11];
  assign data_o[5771] = data_o[11];
  assign data_o[5835] = data_o[11];
  assign data_o[5899] = data_o[11];
  assign data_o[5963] = data_o[11];
  assign data_o[6027] = data_o[11];
  assign data_o[6091] = data_o[11];
  assign data_o[6155] = data_o[11];
  assign data_o[6219] = data_o[11];
  assign data_o[6283] = data_o[11];
  assign data_o[6347] = data_o[11];
  assign data_o[6411] = data_o[11];
  assign data_o[6475] = data_o[11];
  assign data_o[6539] = data_o[11];
  assign data_o[6603] = data_o[11];
  assign data_o[6667] = data_o[11];
  assign data_o[6731] = data_o[11];
  assign data_o[6795] = data_o[11];
  assign data_o[6859] = data_o[11];
  assign data_o[6923] = data_o[11];
  assign data_o[6987] = data_o[11];
  assign data_o[7051] = data_o[11];
  assign data_o[7115] = data_o[11];
  assign data_o[7179] = data_o[11];
  assign data_o[7243] = data_o[11];
  assign data_o[7307] = data_o[11];
  assign data_o[7371] = data_o[11];
  assign data_o[7435] = data_o[11];
  assign data_o[7499] = data_o[11];
  assign data_o[7563] = data_o[11];
  assign data_o[7627] = data_o[11];
  assign data_o[7691] = data_o[11];
  assign data_o[7755] = data_o[11];
  assign data_o[7819] = data_o[11];
  assign data_o[7883] = data_o[11];
  assign data_o[7947] = data_o[11];
  assign data_o[8011] = data_o[11];
  assign data_o[8075] = data_o[11];
  assign data_o[8139] = data_o[11];
  assign data_o[8203] = data_o[11];
  assign data_o[8267] = data_o[11];
  assign data_o[8331] = data_o[11];
  assign data_o[8395] = data_o[11];
  assign data_o[8459] = data_o[11];
  assign data_o[8523] = data_o[11];
  assign data_o[8587] = data_o[11];
  assign data_o[8651] = data_o[11];
  assign data_o[8715] = data_o[11];
  assign data_o[8779] = data_o[11];
  assign data_o[8843] = data_o[11];
  assign data_o[8907] = data_o[11];
  assign data_o[8971] = data_o[11];
  assign data_o[9035] = data_o[11];
  assign data_o[9099] = data_o[11];
  assign data_o[9163] = data_o[11];
  assign data_o[9227] = data_o[11];
  assign data_o[9291] = data_o[11];
  assign data_o[9355] = data_o[11];
  assign data_o[9419] = data_o[11];
  assign data_o[9483] = data_o[11];
  assign data_o[9547] = data_o[11];
  assign data_o[9611] = data_o[11];
  assign data_o[9675] = data_o[11];
  assign data_o[9739] = data_o[11];
  assign data_o[9803] = data_o[11];
  assign data_o[9867] = data_o[11];
  assign data_o[9931] = data_o[11];
  assign data_o[9995] = data_o[11];
  assign data_o[10059] = data_o[11];
  assign data_o[10123] = data_o[11];
  assign data_o[10187] = data_o[11];
  assign data_o[10251] = data_o[11];
  assign data_o[10315] = data_o[11];
  assign data_o[10379] = data_o[11];
  assign data_o[10443] = data_o[11];
  assign data_o[10507] = data_o[11];
  assign data_o[10571] = data_o[11];
  assign data_o[10635] = data_o[11];
  assign data_o[10699] = data_o[11];
  assign data_o[10763] = data_o[11];
  assign data_o[10827] = data_o[11];
  assign data_o[10891] = data_o[11];
  assign data_o[10955] = data_o[11];
  assign data_o[11019] = data_o[11];
  assign data_o[11083] = data_o[11];
  assign data_o[11147] = data_o[11];
  assign data_o[11211] = data_o[11];
  assign data_o[11275] = data_o[11];
  assign data_o[11339] = data_o[11];
  assign data_o[11403] = data_o[11];
  assign data_o[11467] = data_o[11];
  assign data_o[11531] = data_o[11];
  assign data_o[11595] = data_o[11];
  assign data_o[11659] = data_o[11];
  assign data_o[11723] = data_o[11];
  assign data_o[11787] = data_o[11];
  assign data_o[11851] = data_o[11];
  assign data_o[11915] = data_o[11];
  assign data_o[11979] = data_o[11];
  assign data_o[12043] = data_o[11];
  assign data_o[12107] = data_o[11];
  assign data_o[12171] = data_o[11];
  assign data_o[12235] = data_o[11];
  assign data_o[12299] = data_o[11];
  assign data_o[12363] = data_o[11];
  assign data_o[12427] = data_o[11];
  assign data_o[12491] = data_o[11];
  assign data_o[12555] = data_o[11];
  assign data_o[12619] = data_o[11];
  assign data_o[12683] = data_o[11];
  assign data_o[12747] = data_o[11];
  assign data_o[12811] = data_o[11];
  assign data_o[12875] = data_o[11];
  assign data_o[12939] = data_o[11];
  assign data_o[13003] = data_o[11];
  assign data_o[13067] = data_o[11];
  assign data_o[13131] = data_o[11];
  assign data_o[13195] = data_o[11];
  assign data_o[13259] = data_o[11];
  assign data_o[13323] = data_o[11];
  assign data_o[13387] = data_o[11];
  assign data_o[13451] = data_o[11];
  assign data_o[13515] = data_o[11];
  assign data_o[13579] = data_o[11];
  assign data_o[13643] = data_o[11];
  assign data_o[13707] = data_o[11];
  assign data_o[13771] = data_o[11];
  assign data_o[13835] = data_o[11];
  assign data_o[13899] = data_o[11];
  assign data_o[13963] = data_o[11];
  assign data_o[14027] = data_o[11];
  assign data_o[14091] = data_o[11];
  assign data_o[14155] = data_o[11];
  assign data_o[14219] = data_o[11];
  assign data_o[14283] = data_o[11];
  assign data_o[14347] = data_o[11];
  assign data_o[14411] = data_o[11];
  assign data_o[14475] = data_o[11];
  assign data_o[14539] = data_o[11];
  assign data_o[14603] = data_o[11];
  assign data_o[14667] = data_o[11];
  assign data_o[14731] = data_o[11];
  assign data_o[14795] = data_o[11];
  assign data_o[14859] = data_o[11];
  assign data_o[14923] = data_o[11];
  assign data_o[14987] = data_o[11];
  assign data_o[15051] = data_o[11];
  assign data_o[15115] = data_o[11];
  assign data_o[15179] = data_o[11];
  assign data_o[15243] = data_o[11];
  assign data_o[15307] = data_o[11];
  assign data_o[15371] = data_o[11];
  assign data_o[15435] = data_o[11];
  assign data_o[15499] = data_o[11];
  assign data_o[15563] = data_o[11];
  assign data_o[15627] = data_o[11];
  assign data_o[15691] = data_o[11];
  assign data_o[15755] = data_o[11];
  assign data_o[15819] = data_o[11];
  assign data_o[15883] = data_o[11];
  assign data_o[15947] = data_o[11];
  assign data_o[16011] = data_o[11];
  assign data_o[16075] = data_o[11];
  assign data_o[16139] = data_o[11];
  assign data_o[16203] = data_o[11];
  assign data_o[16267] = data_o[11];
  assign data_o[16331] = data_o[11];
  assign data_o[16395] = data_o[11];
  assign data_o[16459] = data_o[11];
  assign data_o[16523] = data_o[11];
  assign data_o[16587] = data_o[11];
  assign data_o[16651] = data_o[11];
  assign data_o[16715] = data_o[11];
  assign data_o[16779] = data_o[11];
  assign data_o[16843] = data_o[11];
  assign data_o[16907] = data_o[11];
  assign data_o[16971] = data_o[11];
  assign data_o[17035] = data_o[11];
  assign data_o[17099] = data_o[11];
  assign data_o[17163] = data_o[11];
  assign data_o[17227] = data_o[11];
  assign data_o[17291] = data_o[11];
  assign data_o[17355] = data_o[11];
  assign data_o[17419] = data_o[11];
  assign data_o[17483] = data_o[11];
  assign data_o[17547] = data_o[11];
  assign data_o[17611] = data_o[11];
  assign data_o[17675] = data_o[11];
  assign data_o[17739] = data_o[11];
  assign data_o[17803] = data_o[11];
  assign data_o[17867] = data_o[11];
  assign data_o[17931] = data_o[11];
  assign data_o[17995] = data_o[11];
  assign data_o[18059] = data_o[11];
  assign data_o[18123] = data_o[11];
  assign data_o[18187] = data_o[11];
  assign data_o[18251] = data_o[11];
  assign data_o[18315] = data_o[11];
  assign data_o[18379] = data_o[11];
  assign data_o[18443] = data_o[11];
  assign data_o[18507] = data_o[11];
  assign data_o[18571] = data_o[11];
  assign data_o[18635] = data_o[11];
  assign data_o[18699] = data_o[11];
  assign data_o[18763] = data_o[11];
  assign data_o[18827] = data_o[11];
  assign data_o[18891] = data_o[11];
  assign data_o[18955] = data_o[11];
  assign data_o[19019] = data_o[11];
  assign data_o[19083] = data_o[11];
  assign data_o[19147] = data_o[11];
  assign data_o[19211] = data_o[11];
  assign data_o[19275] = data_o[11];
  assign data_o[19339] = data_o[11];
  assign data_o[19403] = data_o[11];
  assign data_o[19467] = data_o[11];
  assign data_o[19531] = data_o[11];
  assign data_o[19595] = data_o[11];
  assign data_o[19659] = data_o[11];
  assign data_o[19723] = data_o[11];
  assign data_o[19787] = data_o[11];
  assign data_o[19851] = data_o[11];
  assign data_o[19915] = data_o[11];
  assign data_o[19979] = data_o[11];
  assign data_o[20043] = data_o[11];
  assign data_o[20107] = data_o[11];
  assign data_o[20171] = data_o[11];
  assign data_o[20235] = data_o[11];
  assign data_o[20299] = data_o[11];
  assign data_o[20363] = data_o[11];
  assign data_o[20427] = data_o[11];
  assign data_o[20491] = data_o[11];
  assign data_o[20555] = data_o[11];
  assign data_o[20619] = data_o[11];
  assign data_o[20683] = data_o[11];
  assign data_o[20747] = data_o[11];
  assign data_o[20811] = data_o[11];
  assign data_o[20875] = data_o[11];
  assign data_o[20939] = data_o[11];
  assign data_o[21003] = data_o[11];
  assign data_o[21067] = data_o[11];
  assign data_o[21131] = data_o[11];
  assign data_o[21195] = data_o[11];
  assign data_o[21259] = data_o[11];
  assign data_o[21323] = data_o[11];
  assign data_o[21387] = data_o[11];
  assign data_o[21451] = data_o[11];
  assign data_o[21515] = data_o[11];
  assign data_o[21579] = data_o[11];
  assign data_o[21643] = data_o[11];
  assign data_o[21707] = data_o[11];
  assign data_o[21771] = data_o[11];
  assign data_o[21835] = data_o[11];
  assign data_o[21899] = data_o[11];
  assign data_o[21963] = data_o[11];
  assign data_o[22027] = data_o[11];
  assign data_o[22091] = data_o[11];
  assign data_o[22155] = data_o[11];
  assign data_o[22219] = data_o[11];
  assign data_o[22283] = data_o[11];
  assign data_o[22347] = data_o[11];
  assign data_o[22411] = data_o[11];
  assign data_o[22475] = data_o[11];
  assign data_o[22539] = data_o[11];
  assign data_o[22603] = data_o[11];
  assign data_o[22667] = data_o[11];
  assign data_o[22731] = data_o[11];
  assign data_o[22795] = data_o[11];
  assign data_o[22859] = data_o[11];
  assign data_o[22923] = data_o[11];
  assign data_o[22987] = data_o[11];
  assign data_o[23051] = data_o[11];
  assign data_o[23115] = data_o[11];
  assign data_o[23179] = data_o[11];
  assign data_o[23243] = data_o[11];
  assign data_o[23307] = data_o[11];
  assign data_o[23371] = data_o[11];
  assign data_o[23435] = data_o[11];
  assign data_o[23499] = data_o[11];
  assign data_o[23563] = data_o[11];
  assign data_o[23627] = data_o[11];
  assign data_o[23691] = data_o[11];
  assign data_o[23755] = data_o[11];
  assign data_o[23819] = data_o[11];
  assign data_o[23883] = data_o[11];
  assign data_o[23947] = data_o[11];
  assign data_o[24011] = data_o[11];
  assign data_o[24075] = data_o[11];
  assign data_o[24139] = data_o[11];
  assign data_o[24203] = data_o[11];
  assign data_o[24267] = data_o[11];
  assign data_o[24331] = data_o[11];
  assign data_o[24395] = data_o[11];
  assign data_o[24459] = data_o[11];
  assign data_o[24523] = data_o[11];
  assign data_o[24587] = data_o[11];
  assign data_o[24651] = data_o[11];
  assign data_o[24715] = data_o[11];
  assign data_o[24779] = data_o[11];
  assign data_o[24843] = data_o[11];
  assign data_o[24907] = data_o[11];
  assign data_o[24971] = data_o[11];
  assign data_o[25035] = data_o[11];
  assign data_o[25099] = data_o[11];
  assign data_o[25163] = data_o[11];
  assign data_o[25227] = data_o[11];
  assign data_o[25291] = data_o[11];
  assign data_o[25355] = data_o[11];
  assign data_o[25419] = data_o[11];
  assign data_o[25483] = data_o[11];
  assign data_o[25547] = data_o[11];
  assign data_o[25611] = data_o[11];
  assign data_o[25675] = data_o[11];
  assign data_o[25739] = data_o[11];
  assign data_o[25803] = data_o[11];
  assign data_o[25867] = data_o[11];
  assign data_o[25931] = data_o[11];
  assign data_o[25995] = data_o[11];
  assign data_o[26059] = data_o[11];
  assign data_o[26123] = data_o[11];
  assign data_o[26187] = data_o[11];
  assign data_o[26251] = data_o[11];
  assign data_o[26315] = data_o[11];
  assign data_o[26379] = data_o[11];
  assign data_o[26443] = data_o[11];
  assign data_o[26507] = data_o[11];
  assign data_o[26571] = data_o[11];
  assign data_o[26635] = data_o[11];
  assign data_o[26699] = data_o[11];
  assign data_o[26763] = data_o[11];
  assign data_o[26827] = data_o[11];
  assign data_o[26891] = data_o[11];
  assign data_o[26955] = data_o[11];
  assign data_o[27019] = data_o[11];
  assign data_o[27083] = data_o[11];
  assign data_o[27147] = data_o[11];
  assign data_o[27211] = data_o[11];
  assign data_o[27275] = data_o[11];
  assign data_o[27339] = data_o[11];
  assign data_o[27403] = data_o[11];
  assign data_o[27467] = data_o[11];
  assign data_o[27531] = data_o[11];
  assign data_o[27595] = data_o[11];
  assign data_o[27659] = data_o[11];
  assign data_o[27723] = data_o[11];
  assign data_o[27787] = data_o[11];
  assign data_o[27851] = data_o[11];
  assign data_o[27915] = data_o[11];
  assign data_o[27979] = data_o[11];
  assign data_o[28043] = data_o[11];
  assign data_o[28107] = data_o[11];
  assign data_o[28171] = data_o[11];
  assign data_o[28235] = data_o[11];
  assign data_o[28299] = data_o[11];
  assign data_o[28363] = data_o[11];
  assign data_o[28427] = data_o[11];
  assign data_o[28491] = data_o[11];
  assign data_o[28555] = data_o[11];
  assign data_o[28619] = data_o[11];
  assign data_o[28683] = data_o[11];
  assign data_o[28747] = data_o[11];
  assign data_o[28811] = data_o[11];
  assign data_o[28875] = data_o[11];
  assign data_o[28939] = data_o[11];
  assign data_o[29003] = data_o[11];
  assign data_o[29067] = data_o[11];
  assign data_o[29131] = data_o[11];
  assign data_o[29195] = data_o[11];
  assign data_o[29259] = data_o[11];
  assign data_o[29323] = data_o[11];
  assign data_o[29387] = data_o[11];
  assign data_o[29451] = data_o[11];
  assign data_o[29515] = data_o[11];
  assign data_o[29579] = data_o[11];
  assign data_o[29643] = data_o[11];
  assign data_o[29707] = data_o[11];
  assign data_o[29771] = data_o[11];
  assign data_o[29835] = data_o[11];
  assign data_o[29899] = data_o[11];
  assign data_o[29963] = data_o[11];
  assign data_o[30027] = data_o[11];
  assign data_o[30091] = data_o[11];
  assign data_o[30155] = data_o[11];
  assign data_o[30219] = data_o[11];
  assign data_o[30283] = data_o[11];
  assign data_o[30347] = data_o[11];
  assign data_o[30411] = data_o[11];
  assign data_o[30475] = data_o[11];
  assign data_o[30539] = data_o[11];
  assign data_o[30603] = data_o[11];
  assign data_o[30667] = data_o[11];
  assign data_o[30731] = data_o[11];
  assign data_o[30795] = data_o[11];
  assign data_o[30859] = data_o[11];
  assign data_o[30923] = data_o[11];
  assign data_o[30987] = data_o[11];
  assign data_o[31051] = data_o[11];
  assign data_o[31115] = data_o[11];
  assign data_o[31179] = data_o[11];
  assign data_o[31243] = data_o[11];
  assign data_o[31307] = data_o[11];
  assign data_o[31371] = data_o[11];
  assign data_o[31435] = data_o[11];
  assign data_o[31499] = data_o[11];
  assign data_o[31563] = data_o[11];
  assign data_o[31627] = data_o[11];
  assign data_o[31691] = data_o[11];
  assign data_o[31755] = data_o[11];
  assign data_o[31819] = data_o[11];
  assign data_o[31883] = data_o[11];
  assign data_o[31947] = data_o[11];
  assign data_o[74] = data_o[10];
  assign data_o[138] = data_o[10];
  assign data_o[202] = data_o[10];
  assign data_o[266] = data_o[10];
  assign data_o[330] = data_o[10];
  assign data_o[394] = data_o[10];
  assign data_o[458] = data_o[10];
  assign data_o[522] = data_o[10];
  assign data_o[586] = data_o[10];
  assign data_o[650] = data_o[10];
  assign data_o[714] = data_o[10];
  assign data_o[778] = data_o[10];
  assign data_o[842] = data_o[10];
  assign data_o[906] = data_o[10];
  assign data_o[970] = data_o[10];
  assign data_o[1034] = data_o[10];
  assign data_o[1098] = data_o[10];
  assign data_o[1162] = data_o[10];
  assign data_o[1226] = data_o[10];
  assign data_o[1290] = data_o[10];
  assign data_o[1354] = data_o[10];
  assign data_o[1418] = data_o[10];
  assign data_o[1482] = data_o[10];
  assign data_o[1546] = data_o[10];
  assign data_o[1610] = data_o[10];
  assign data_o[1674] = data_o[10];
  assign data_o[1738] = data_o[10];
  assign data_o[1802] = data_o[10];
  assign data_o[1866] = data_o[10];
  assign data_o[1930] = data_o[10];
  assign data_o[1994] = data_o[10];
  assign data_o[2058] = data_o[10];
  assign data_o[2122] = data_o[10];
  assign data_o[2186] = data_o[10];
  assign data_o[2250] = data_o[10];
  assign data_o[2314] = data_o[10];
  assign data_o[2378] = data_o[10];
  assign data_o[2442] = data_o[10];
  assign data_o[2506] = data_o[10];
  assign data_o[2570] = data_o[10];
  assign data_o[2634] = data_o[10];
  assign data_o[2698] = data_o[10];
  assign data_o[2762] = data_o[10];
  assign data_o[2826] = data_o[10];
  assign data_o[2890] = data_o[10];
  assign data_o[2954] = data_o[10];
  assign data_o[3018] = data_o[10];
  assign data_o[3082] = data_o[10];
  assign data_o[3146] = data_o[10];
  assign data_o[3210] = data_o[10];
  assign data_o[3274] = data_o[10];
  assign data_o[3338] = data_o[10];
  assign data_o[3402] = data_o[10];
  assign data_o[3466] = data_o[10];
  assign data_o[3530] = data_o[10];
  assign data_o[3594] = data_o[10];
  assign data_o[3658] = data_o[10];
  assign data_o[3722] = data_o[10];
  assign data_o[3786] = data_o[10];
  assign data_o[3850] = data_o[10];
  assign data_o[3914] = data_o[10];
  assign data_o[3978] = data_o[10];
  assign data_o[4042] = data_o[10];
  assign data_o[4106] = data_o[10];
  assign data_o[4170] = data_o[10];
  assign data_o[4234] = data_o[10];
  assign data_o[4298] = data_o[10];
  assign data_o[4362] = data_o[10];
  assign data_o[4426] = data_o[10];
  assign data_o[4490] = data_o[10];
  assign data_o[4554] = data_o[10];
  assign data_o[4618] = data_o[10];
  assign data_o[4682] = data_o[10];
  assign data_o[4746] = data_o[10];
  assign data_o[4810] = data_o[10];
  assign data_o[4874] = data_o[10];
  assign data_o[4938] = data_o[10];
  assign data_o[5002] = data_o[10];
  assign data_o[5066] = data_o[10];
  assign data_o[5130] = data_o[10];
  assign data_o[5194] = data_o[10];
  assign data_o[5258] = data_o[10];
  assign data_o[5322] = data_o[10];
  assign data_o[5386] = data_o[10];
  assign data_o[5450] = data_o[10];
  assign data_o[5514] = data_o[10];
  assign data_o[5578] = data_o[10];
  assign data_o[5642] = data_o[10];
  assign data_o[5706] = data_o[10];
  assign data_o[5770] = data_o[10];
  assign data_o[5834] = data_o[10];
  assign data_o[5898] = data_o[10];
  assign data_o[5962] = data_o[10];
  assign data_o[6026] = data_o[10];
  assign data_o[6090] = data_o[10];
  assign data_o[6154] = data_o[10];
  assign data_o[6218] = data_o[10];
  assign data_o[6282] = data_o[10];
  assign data_o[6346] = data_o[10];
  assign data_o[6410] = data_o[10];
  assign data_o[6474] = data_o[10];
  assign data_o[6538] = data_o[10];
  assign data_o[6602] = data_o[10];
  assign data_o[6666] = data_o[10];
  assign data_o[6730] = data_o[10];
  assign data_o[6794] = data_o[10];
  assign data_o[6858] = data_o[10];
  assign data_o[6922] = data_o[10];
  assign data_o[6986] = data_o[10];
  assign data_o[7050] = data_o[10];
  assign data_o[7114] = data_o[10];
  assign data_o[7178] = data_o[10];
  assign data_o[7242] = data_o[10];
  assign data_o[7306] = data_o[10];
  assign data_o[7370] = data_o[10];
  assign data_o[7434] = data_o[10];
  assign data_o[7498] = data_o[10];
  assign data_o[7562] = data_o[10];
  assign data_o[7626] = data_o[10];
  assign data_o[7690] = data_o[10];
  assign data_o[7754] = data_o[10];
  assign data_o[7818] = data_o[10];
  assign data_o[7882] = data_o[10];
  assign data_o[7946] = data_o[10];
  assign data_o[8010] = data_o[10];
  assign data_o[8074] = data_o[10];
  assign data_o[8138] = data_o[10];
  assign data_o[8202] = data_o[10];
  assign data_o[8266] = data_o[10];
  assign data_o[8330] = data_o[10];
  assign data_o[8394] = data_o[10];
  assign data_o[8458] = data_o[10];
  assign data_o[8522] = data_o[10];
  assign data_o[8586] = data_o[10];
  assign data_o[8650] = data_o[10];
  assign data_o[8714] = data_o[10];
  assign data_o[8778] = data_o[10];
  assign data_o[8842] = data_o[10];
  assign data_o[8906] = data_o[10];
  assign data_o[8970] = data_o[10];
  assign data_o[9034] = data_o[10];
  assign data_o[9098] = data_o[10];
  assign data_o[9162] = data_o[10];
  assign data_o[9226] = data_o[10];
  assign data_o[9290] = data_o[10];
  assign data_o[9354] = data_o[10];
  assign data_o[9418] = data_o[10];
  assign data_o[9482] = data_o[10];
  assign data_o[9546] = data_o[10];
  assign data_o[9610] = data_o[10];
  assign data_o[9674] = data_o[10];
  assign data_o[9738] = data_o[10];
  assign data_o[9802] = data_o[10];
  assign data_o[9866] = data_o[10];
  assign data_o[9930] = data_o[10];
  assign data_o[9994] = data_o[10];
  assign data_o[10058] = data_o[10];
  assign data_o[10122] = data_o[10];
  assign data_o[10186] = data_o[10];
  assign data_o[10250] = data_o[10];
  assign data_o[10314] = data_o[10];
  assign data_o[10378] = data_o[10];
  assign data_o[10442] = data_o[10];
  assign data_o[10506] = data_o[10];
  assign data_o[10570] = data_o[10];
  assign data_o[10634] = data_o[10];
  assign data_o[10698] = data_o[10];
  assign data_o[10762] = data_o[10];
  assign data_o[10826] = data_o[10];
  assign data_o[10890] = data_o[10];
  assign data_o[10954] = data_o[10];
  assign data_o[11018] = data_o[10];
  assign data_o[11082] = data_o[10];
  assign data_o[11146] = data_o[10];
  assign data_o[11210] = data_o[10];
  assign data_o[11274] = data_o[10];
  assign data_o[11338] = data_o[10];
  assign data_o[11402] = data_o[10];
  assign data_o[11466] = data_o[10];
  assign data_o[11530] = data_o[10];
  assign data_o[11594] = data_o[10];
  assign data_o[11658] = data_o[10];
  assign data_o[11722] = data_o[10];
  assign data_o[11786] = data_o[10];
  assign data_o[11850] = data_o[10];
  assign data_o[11914] = data_o[10];
  assign data_o[11978] = data_o[10];
  assign data_o[12042] = data_o[10];
  assign data_o[12106] = data_o[10];
  assign data_o[12170] = data_o[10];
  assign data_o[12234] = data_o[10];
  assign data_o[12298] = data_o[10];
  assign data_o[12362] = data_o[10];
  assign data_o[12426] = data_o[10];
  assign data_o[12490] = data_o[10];
  assign data_o[12554] = data_o[10];
  assign data_o[12618] = data_o[10];
  assign data_o[12682] = data_o[10];
  assign data_o[12746] = data_o[10];
  assign data_o[12810] = data_o[10];
  assign data_o[12874] = data_o[10];
  assign data_o[12938] = data_o[10];
  assign data_o[13002] = data_o[10];
  assign data_o[13066] = data_o[10];
  assign data_o[13130] = data_o[10];
  assign data_o[13194] = data_o[10];
  assign data_o[13258] = data_o[10];
  assign data_o[13322] = data_o[10];
  assign data_o[13386] = data_o[10];
  assign data_o[13450] = data_o[10];
  assign data_o[13514] = data_o[10];
  assign data_o[13578] = data_o[10];
  assign data_o[13642] = data_o[10];
  assign data_o[13706] = data_o[10];
  assign data_o[13770] = data_o[10];
  assign data_o[13834] = data_o[10];
  assign data_o[13898] = data_o[10];
  assign data_o[13962] = data_o[10];
  assign data_o[14026] = data_o[10];
  assign data_o[14090] = data_o[10];
  assign data_o[14154] = data_o[10];
  assign data_o[14218] = data_o[10];
  assign data_o[14282] = data_o[10];
  assign data_o[14346] = data_o[10];
  assign data_o[14410] = data_o[10];
  assign data_o[14474] = data_o[10];
  assign data_o[14538] = data_o[10];
  assign data_o[14602] = data_o[10];
  assign data_o[14666] = data_o[10];
  assign data_o[14730] = data_o[10];
  assign data_o[14794] = data_o[10];
  assign data_o[14858] = data_o[10];
  assign data_o[14922] = data_o[10];
  assign data_o[14986] = data_o[10];
  assign data_o[15050] = data_o[10];
  assign data_o[15114] = data_o[10];
  assign data_o[15178] = data_o[10];
  assign data_o[15242] = data_o[10];
  assign data_o[15306] = data_o[10];
  assign data_o[15370] = data_o[10];
  assign data_o[15434] = data_o[10];
  assign data_o[15498] = data_o[10];
  assign data_o[15562] = data_o[10];
  assign data_o[15626] = data_o[10];
  assign data_o[15690] = data_o[10];
  assign data_o[15754] = data_o[10];
  assign data_o[15818] = data_o[10];
  assign data_o[15882] = data_o[10];
  assign data_o[15946] = data_o[10];
  assign data_o[16010] = data_o[10];
  assign data_o[16074] = data_o[10];
  assign data_o[16138] = data_o[10];
  assign data_o[16202] = data_o[10];
  assign data_o[16266] = data_o[10];
  assign data_o[16330] = data_o[10];
  assign data_o[16394] = data_o[10];
  assign data_o[16458] = data_o[10];
  assign data_o[16522] = data_o[10];
  assign data_o[16586] = data_o[10];
  assign data_o[16650] = data_o[10];
  assign data_o[16714] = data_o[10];
  assign data_o[16778] = data_o[10];
  assign data_o[16842] = data_o[10];
  assign data_o[16906] = data_o[10];
  assign data_o[16970] = data_o[10];
  assign data_o[17034] = data_o[10];
  assign data_o[17098] = data_o[10];
  assign data_o[17162] = data_o[10];
  assign data_o[17226] = data_o[10];
  assign data_o[17290] = data_o[10];
  assign data_o[17354] = data_o[10];
  assign data_o[17418] = data_o[10];
  assign data_o[17482] = data_o[10];
  assign data_o[17546] = data_o[10];
  assign data_o[17610] = data_o[10];
  assign data_o[17674] = data_o[10];
  assign data_o[17738] = data_o[10];
  assign data_o[17802] = data_o[10];
  assign data_o[17866] = data_o[10];
  assign data_o[17930] = data_o[10];
  assign data_o[17994] = data_o[10];
  assign data_o[18058] = data_o[10];
  assign data_o[18122] = data_o[10];
  assign data_o[18186] = data_o[10];
  assign data_o[18250] = data_o[10];
  assign data_o[18314] = data_o[10];
  assign data_o[18378] = data_o[10];
  assign data_o[18442] = data_o[10];
  assign data_o[18506] = data_o[10];
  assign data_o[18570] = data_o[10];
  assign data_o[18634] = data_o[10];
  assign data_o[18698] = data_o[10];
  assign data_o[18762] = data_o[10];
  assign data_o[18826] = data_o[10];
  assign data_o[18890] = data_o[10];
  assign data_o[18954] = data_o[10];
  assign data_o[19018] = data_o[10];
  assign data_o[19082] = data_o[10];
  assign data_o[19146] = data_o[10];
  assign data_o[19210] = data_o[10];
  assign data_o[19274] = data_o[10];
  assign data_o[19338] = data_o[10];
  assign data_o[19402] = data_o[10];
  assign data_o[19466] = data_o[10];
  assign data_o[19530] = data_o[10];
  assign data_o[19594] = data_o[10];
  assign data_o[19658] = data_o[10];
  assign data_o[19722] = data_o[10];
  assign data_o[19786] = data_o[10];
  assign data_o[19850] = data_o[10];
  assign data_o[19914] = data_o[10];
  assign data_o[19978] = data_o[10];
  assign data_o[20042] = data_o[10];
  assign data_o[20106] = data_o[10];
  assign data_o[20170] = data_o[10];
  assign data_o[20234] = data_o[10];
  assign data_o[20298] = data_o[10];
  assign data_o[20362] = data_o[10];
  assign data_o[20426] = data_o[10];
  assign data_o[20490] = data_o[10];
  assign data_o[20554] = data_o[10];
  assign data_o[20618] = data_o[10];
  assign data_o[20682] = data_o[10];
  assign data_o[20746] = data_o[10];
  assign data_o[20810] = data_o[10];
  assign data_o[20874] = data_o[10];
  assign data_o[20938] = data_o[10];
  assign data_o[21002] = data_o[10];
  assign data_o[21066] = data_o[10];
  assign data_o[21130] = data_o[10];
  assign data_o[21194] = data_o[10];
  assign data_o[21258] = data_o[10];
  assign data_o[21322] = data_o[10];
  assign data_o[21386] = data_o[10];
  assign data_o[21450] = data_o[10];
  assign data_o[21514] = data_o[10];
  assign data_o[21578] = data_o[10];
  assign data_o[21642] = data_o[10];
  assign data_o[21706] = data_o[10];
  assign data_o[21770] = data_o[10];
  assign data_o[21834] = data_o[10];
  assign data_o[21898] = data_o[10];
  assign data_o[21962] = data_o[10];
  assign data_o[22026] = data_o[10];
  assign data_o[22090] = data_o[10];
  assign data_o[22154] = data_o[10];
  assign data_o[22218] = data_o[10];
  assign data_o[22282] = data_o[10];
  assign data_o[22346] = data_o[10];
  assign data_o[22410] = data_o[10];
  assign data_o[22474] = data_o[10];
  assign data_o[22538] = data_o[10];
  assign data_o[22602] = data_o[10];
  assign data_o[22666] = data_o[10];
  assign data_o[22730] = data_o[10];
  assign data_o[22794] = data_o[10];
  assign data_o[22858] = data_o[10];
  assign data_o[22922] = data_o[10];
  assign data_o[22986] = data_o[10];
  assign data_o[23050] = data_o[10];
  assign data_o[23114] = data_o[10];
  assign data_o[23178] = data_o[10];
  assign data_o[23242] = data_o[10];
  assign data_o[23306] = data_o[10];
  assign data_o[23370] = data_o[10];
  assign data_o[23434] = data_o[10];
  assign data_o[23498] = data_o[10];
  assign data_o[23562] = data_o[10];
  assign data_o[23626] = data_o[10];
  assign data_o[23690] = data_o[10];
  assign data_o[23754] = data_o[10];
  assign data_o[23818] = data_o[10];
  assign data_o[23882] = data_o[10];
  assign data_o[23946] = data_o[10];
  assign data_o[24010] = data_o[10];
  assign data_o[24074] = data_o[10];
  assign data_o[24138] = data_o[10];
  assign data_o[24202] = data_o[10];
  assign data_o[24266] = data_o[10];
  assign data_o[24330] = data_o[10];
  assign data_o[24394] = data_o[10];
  assign data_o[24458] = data_o[10];
  assign data_o[24522] = data_o[10];
  assign data_o[24586] = data_o[10];
  assign data_o[24650] = data_o[10];
  assign data_o[24714] = data_o[10];
  assign data_o[24778] = data_o[10];
  assign data_o[24842] = data_o[10];
  assign data_o[24906] = data_o[10];
  assign data_o[24970] = data_o[10];
  assign data_o[25034] = data_o[10];
  assign data_o[25098] = data_o[10];
  assign data_o[25162] = data_o[10];
  assign data_o[25226] = data_o[10];
  assign data_o[25290] = data_o[10];
  assign data_o[25354] = data_o[10];
  assign data_o[25418] = data_o[10];
  assign data_o[25482] = data_o[10];
  assign data_o[25546] = data_o[10];
  assign data_o[25610] = data_o[10];
  assign data_o[25674] = data_o[10];
  assign data_o[25738] = data_o[10];
  assign data_o[25802] = data_o[10];
  assign data_o[25866] = data_o[10];
  assign data_o[25930] = data_o[10];
  assign data_o[25994] = data_o[10];
  assign data_o[26058] = data_o[10];
  assign data_o[26122] = data_o[10];
  assign data_o[26186] = data_o[10];
  assign data_o[26250] = data_o[10];
  assign data_o[26314] = data_o[10];
  assign data_o[26378] = data_o[10];
  assign data_o[26442] = data_o[10];
  assign data_o[26506] = data_o[10];
  assign data_o[26570] = data_o[10];
  assign data_o[26634] = data_o[10];
  assign data_o[26698] = data_o[10];
  assign data_o[26762] = data_o[10];
  assign data_o[26826] = data_o[10];
  assign data_o[26890] = data_o[10];
  assign data_o[26954] = data_o[10];
  assign data_o[27018] = data_o[10];
  assign data_o[27082] = data_o[10];
  assign data_o[27146] = data_o[10];
  assign data_o[27210] = data_o[10];
  assign data_o[27274] = data_o[10];
  assign data_o[27338] = data_o[10];
  assign data_o[27402] = data_o[10];
  assign data_o[27466] = data_o[10];
  assign data_o[27530] = data_o[10];
  assign data_o[27594] = data_o[10];
  assign data_o[27658] = data_o[10];
  assign data_o[27722] = data_o[10];
  assign data_o[27786] = data_o[10];
  assign data_o[27850] = data_o[10];
  assign data_o[27914] = data_o[10];
  assign data_o[27978] = data_o[10];
  assign data_o[28042] = data_o[10];
  assign data_o[28106] = data_o[10];
  assign data_o[28170] = data_o[10];
  assign data_o[28234] = data_o[10];
  assign data_o[28298] = data_o[10];
  assign data_o[28362] = data_o[10];
  assign data_o[28426] = data_o[10];
  assign data_o[28490] = data_o[10];
  assign data_o[28554] = data_o[10];
  assign data_o[28618] = data_o[10];
  assign data_o[28682] = data_o[10];
  assign data_o[28746] = data_o[10];
  assign data_o[28810] = data_o[10];
  assign data_o[28874] = data_o[10];
  assign data_o[28938] = data_o[10];
  assign data_o[29002] = data_o[10];
  assign data_o[29066] = data_o[10];
  assign data_o[29130] = data_o[10];
  assign data_o[29194] = data_o[10];
  assign data_o[29258] = data_o[10];
  assign data_o[29322] = data_o[10];
  assign data_o[29386] = data_o[10];
  assign data_o[29450] = data_o[10];
  assign data_o[29514] = data_o[10];
  assign data_o[29578] = data_o[10];
  assign data_o[29642] = data_o[10];
  assign data_o[29706] = data_o[10];
  assign data_o[29770] = data_o[10];
  assign data_o[29834] = data_o[10];
  assign data_o[29898] = data_o[10];
  assign data_o[29962] = data_o[10];
  assign data_o[30026] = data_o[10];
  assign data_o[30090] = data_o[10];
  assign data_o[30154] = data_o[10];
  assign data_o[30218] = data_o[10];
  assign data_o[30282] = data_o[10];
  assign data_o[30346] = data_o[10];
  assign data_o[30410] = data_o[10];
  assign data_o[30474] = data_o[10];
  assign data_o[30538] = data_o[10];
  assign data_o[30602] = data_o[10];
  assign data_o[30666] = data_o[10];
  assign data_o[30730] = data_o[10];
  assign data_o[30794] = data_o[10];
  assign data_o[30858] = data_o[10];
  assign data_o[30922] = data_o[10];
  assign data_o[30986] = data_o[10];
  assign data_o[31050] = data_o[10];
  assign data_o[31114] = data_o[10];
  assign data_o[31178] = data_o[10];
  assign data_o[31242] = data_o[10];
  assign data_o[31306] = data_o[10];
  assign data_o[31370] = data_o[10];
  assign data_o[31434] = data_o[10];
  assign data_o[31498] = data_o[10];
  assign data_o[31562] = data_o[10];
  assign data_o[31626] = data_o[10];
  assign data_o[31690] = data_o[10];
  assign data_o[31754] = data_o[10];
  assign data_o[31818] = data_o[10];
  assign data_o[31882] = data_o[10];
  assign data_o[31946] = data_o[10];
  assign data_o[73] = data_o[9];
  assign data_o[137] = data_o[9];
  assign data_o[201] = data_o[9];
  assign data_o[265] = data_o[9];
  assign data_o[329] = data_o[9];
  assign data_o[393] = data_o[9];
  assign data_o[457] = data_o[9];
  assign data_o[521] = data_o[9];
  assign data_o[585] = data_o[9];
  assign data_o[649] = data_o[9];
  assign data_o[713] = data_o[9];
  assign data_o[777] = data_o[9];
  assign data_o[841] = data_o[9];
  assign data_o[905] = data_o[9];
  assign data_o[969] = data_o[9];
  assign data_o[1033] = data_o[9];
  assign data_o[1097] = data_o[9];
  assign data_o[1161] = data_o[9];
  assign data_o[1225] = data_o[9];
  assign data_o[1289] = data_o[9];
  assign data_o[1353] = data_o[9];
  assign data_o[1417] = data_o[9];
  assign data_o[1481] = data_o[9];
  assign data_o[1545] = data_o[9];
  assign data_o[1609] = data_o[9];
  assign data_o[1673] = data_o[9];
  assign data_o[1737] = data_o[9];
  assign data_o[1801] = data_o[9];
  assign data_o[1865] = data_o[9];
  assign data_o[1929] = data_o[9];
  assign data_o[1993] = data_o[9];
  assign data_o[2057] = data_o[9];
  assign data_o[2121] = data_o[9];
  assign data_o[2185] = data_o[9];
  assign data_o[2249] = data_o[9];
  assign data_o[2313] = data_o[9];
  assign data_o[2377] = data_o[9];
  assign data_o[2441] = data_o[9];
  assign data_o[2505] = data_o[9];
  assign data_o[2569] = data_o[9];
  assign data_o[2633] = data_o[9];
  assign data_o[2697] = data_o[9];
  assign data_o[2761] = data_o[9];
  assign data_o[2825] = data_o[9];
  assign data_o[2889] = data_o[9];
  assign data_o[2953] = data_o[9];
  assign data_o[3017] = data_o[9];
  assign data_o[3081] = data_o[9];
  assign data_o[3145] = data_o[9];
  assign data_o[3209] = data_o[9];
  assign data_o[3273] = data_o[9];
  assign data_o[3337] = data_o[9];
  assign data_o[3401] = data_o[9];
  assign data_o[3465] = data_o[9];
  assign data_o[3529] = data_o[9];
  assign data_o[3593] = data_o[9];
  assign data_o[3657] = data_o[9];
  assign data_o[3721] = data_o[9];
  assign data_o[3785] = data_o[9];
  assign data_o[3849] = data_o[9];
  assign data_o[3913] = data_o[9];
  assign data_o[3977] = data_o[9];
  assign data_o[4041] = data_o[9];
  assign data_o[4105] = data_o[9];
  assign data_o[4169] = data_o[9];
  assign data_o[4233] = data_o[9];
  assign data_o[4297] = data_o[9];
  assign data_o[4361] = data_o[9];
  assign data_o[4425] = data_o[9];
  assign data_o[4489] = data_o[9];
  assign data_o[4553] = data_o[9];
  assign data_o[4617] = data_o[9];
  assign data_o[4681] = data_o[9];
  assign data_o[4745] = data_o[9];
  assign data_o[4809] = data_o[9];
  assign data_o[4873] = data_o[9];
  assign data_o[4937] = data_o[9];
  assign data_o[5001] = data_o[9];
  assign data_o[5065] = data_o[9];
  assign data_o[5129] = data_o[9];
  assign data_o[5193] = data_o[9];
  assign data_o[5257] = data_o[9];
  assign data_o[5321] = data_o[9];
  assign data_o[5385] = data_o[9];
  assign data_o[5449] = data_o[9];
  assign data_o[5513] = data_o[9];
  assign data_o[5577] = data_o[9];
  assign data_o[5641] = data_o[9];
  assign data_o[5705] = data_o[9];
  assign data_o[5769] = data_o[9];
  assign data_o[5833] = data_o[9];
  assign data_o[5897] = data_o[9];
  assign data_o[5961] = data_o[9];
  assign data_o[6025] = data_o[9];
  assign data_o[6089] = data_o[9];
  assign data_o[6153] = data_o[9];
  assign data_o[6217] = data_o[9];
  assign data_o[6281] = data_o[9];
  assign data_o[6345] = data_o[9];
  assign data_o[6409] = data_o[9];
  assign data_o[6473] = data_o[9];
  assign data_o[6537] = data_o[9];
  assign data_o[6601] = data_o[9];
  assign data_o[6665] = data_o[9];
  assign data_o[6729] = data_o[9];
  assign data_o[6793] = data_o[9];
  assign data_o[6857] = data_o[9];
  assign data_o[6921] = data_o[9];
  assign data_o[6985] = data_o[9];
  assign data_o[7049] = data_o[9];
  assign data_o[7113] = data_o[9];
  assign data_o[7177] = data_o[9];
  assign data_o[7241] = data_o[9];
  assign data_o[7305] = data_o[9];
  assign data_o[7369] = data_o[9];
  assign data_o[7433] = data_o[9];
  assign data_o[7497] = data_o[9];
  assign data_o[7561] = data_o[9];
  assign data_o[7625] = data_o[9];
  assign data_o[7689] = data_o[9];
  assign data_o[7753] = data_o[9];
  assign data_o[7817] = data_o[9];
  assign data_o[7881] = data_o[9];
  assign data_o[7945] = data_o[9];
  assign data_o[8009] = data_o[9];
  assign data_o[8073] = data_o[9];
  assign data_o[8137] = data_o[9];
  assign data_o[8201] = data_o[9];
  assign data_o[8265] = data_o[9];
  assign data_o[8329] = data_o[9];
  assign data_o[8393] = data_o[9];
  assign data_o[8457] = data_o[9];
  assign data_o[8521] = data_o[9];
  assign data_o[8585] = data_o[9];
  assign data_o[8649] = data_o[9];
  assign data_o[8713] = data_o[9];
  assign data_o[8777] = data_o[9];
  assign data_o[8841] = data_o[9];
  assign data_o[8905] = data_o[9];
  assign data_o[8969] = data_o[9];
  assign data_o[9033] = data_o[9];
  assign data_o[9097] = data_o[9];
  assign data_o[9161] = data_o[9];
  assign data_o[9225] = data_o[9];
  assign data_o[9289] = data_o[9];
  assign data_o[9353] = data_o[9];
  assign data_o[9417] = data_o[9];
  assign data_o[9481] = data_o[9];
  assign data_o[9545] = data_o[9];
  assign data_o[9609] = data_o[9];
  assign data_o[9673] = data_o[9];
  assign data_o[9737] = data_o[9];
  assign data_o[9801] = data_o[9];
  assign data_o[9865] = data_o[9];
  assign data_o[9929] = data_o[9];
  assign data_o[9993] = data_o[9];
  assign data_o[10057] = data_o[9];
  assign data_o[10121] = data_o[9];
  assign data_o[10185] = data_o[9];
  assign data_o[10249] = data_o[9];
  assign data_o[10313] = data_o[9];
  assign data_o[10377] = data_o[9];
  assign data_o[10441] = data_o[9];
  assign data_o[10505] = data_o[9];
  assign data_o[10569] = data_o[9];
  assign data_o[10633] = data_o[9];
  assign data_o[10697] = data_o[9];
  assign data_o[10761] = data_o[9];
  assign data_o[10825] = data_o[9];
  assign data_o[10889] = data_o[9];
  assign data_o[10953] = data_o[9];
  assign data_o[11017] = data_o[9];
  assign data_o[11081] = data_o[9];
  assign data_o[11145] = data_o[9];
  assign data_o[11209] = data_o[9];
  assign data_o[11273] = data_o[9];
  assign data_o[11337] = data_o[9];
  assign data_o[11401] = data_o[9];
  assign data_o[11465] = data_o[9];
  assign data_o[11529] = data_o[9];
  assign data_o[11593] = data_o[9];
  assign data_o[11657] = data_o[9];
  assign data_o[11721] = data_o[9];
  assign data_o[11785] = data_o[9];
  assign data_o[11849] = data_o[9];
  assign data_o[11913] = data_o[9];
  assign data_o[11977] = data_o[9];
  assign data_o[12041] = data_o[9];
  assign data_o[12105] = data_o[9];
  assign data_o[12169] = data_o[9];
  assign data_o[12233] = data_o[9];
  assign data_o[12297] = data_o[9];
  assign data_o[12361] = data_o[9];
  assign data_o[12425] = data_o[9];
  assign data_o[12489] = data_o[9];
  assign data_o[12553] = data_o[9];
  assign data_o[12617] = data_o[9];
  assign data_o[12681] = data_o[9];
  assign data_o[12745] = data_o[9];
  assign data_o[12809] = data_o[9];
  assign data_o[12873] = data_o[9];
  assign data_o[12937] = data_o[9];
  assign data_o[13001] = data_o[9];
  assign data_o[13065] = data_o[9];
  assign data_o[13129] = data_o[9];
  assign data_o[13193] = data_o[9];
  assign data_o[13257] = data_o[9];
  assign data_o[13321] = data_o[9];
  assign data_o[13385] = data_o[9];
  assign data_o[13449] = data_o[9];
  assign data_o[13513] = data_o[9];
  assign data_o[13577] = data_o[9];
  assign data_o[13641] = data_o[9];
  assign data_o[13705] = data_o[9];
  assign data_o[13769] = data_o[9];
  assign data_o[13833] = data_o[9];
  assign data_o[13897] = data_o[9];
  assign data_o[13961] = data_o[9];
  assign data_o[14025] = data_o[9];
  assign data_o[14089] = data_o[9];
  assign data_o[14153] = data_o[9];
  assign data_o[14217] = data_o[9];
  assign data_o[14281] = data_o[9];
  assign data_o[14345] = data_o[9];
  assign data_o[14409] = data_o[9];
  assign data_o[14473] = data_o[9];
  assign data_o[14537] = data_o[9];
  assign data_o[14601] = data_o[9];
  assign data_o[14665] = data_o[9];
  assign data_o[14729] = data_o[9];
  assign data_o[14793] = data_o[9];
  assign data_o[14857] = data_o[9];
  assign data_o[14921] = data_o[9];
  assign data_o[14985] = data_o[9];
  assign data_o[15049] = data_o[9];
  assign data_o[15113] = data_o[9];
  assign data_o[15177] = data_o[9];
  assign data_o[15241] = data_o[9];
  assign data_o[15305] = data_o[9];
  assign data_o[15369] = data_o[9];
  assign data_o[15433] = data_o[9];
  assign data_o[15497] = data_o[9];
  assign data_o[15561] = data_o[9];
  assign data_o[15625] = data_o[9];
  assign data_o[15689] = data_o[9];
  assign data_o[15753] = data_o[9];
  assign data_o[15817] = data_o[9];
  assign data_o[15881] = data_o[9];
  assign data_o[15945] = data_o[9];
  assign data_o[16009] = data_o[9];
  assign data_o[16073] = data_o[9];
  assign data_o[16137] = data_o[9];
  assign data_o[16201] = data_o[9];
  assign data_o[16265] = data_o[9];
  assign data_o[16329] = data_o[9];
  assign data_o[16393] = data_o[9];
  assign data_o[16457] = data_o[9];
  assign data_o[16521] = data_o[9];
  assign data_o[16585] = data_o[9];
  assign data_o[16649] = data_o[9];
  assign data_o[16713] = data_o[9];
  assign data_o[16777] = data_o[9];
  assign data_o[16841] = data_o[9];
  assign data_o[16905] = data_o[9];
  assign data_o[16969] = data_o[9];
  assign data_o[17033] = data_o[9];
  assign data_o[17097] = data_o[9];
  assign data_o[17161] = data_o[9];
  assign data_o[17225] = data_o[9];
  assign data_o[17289] = data_o[9];
  assign data_o[17353] = data_o[9];
  assign data_o[17417] = data_o[9];
  assign data_o[17481] = data_o[9];
  assign data_o[17545] = data_o[9];
  assign data_o[17609] = data_o[9];
  assign data_o[17673] = data_o[9];
  assign data_o[17737] = data_o[9];
  assign data_o[17801] = data_o[9];
  assign data_o[17865] = data_o[9];
  assign data_o[17929] = data_o[9];
  assign data_o[17993] = data_o[9];
  assign data_o[18057] = data_o[9];
  assign data_o[18121] = data_o[9];
  assign data_o[18185] = data_o[9];
  assign data_o[18249] = data_o[9];
  assign data_o[18313] = data_o[9];
  assign data_o[18377] = data_o[9];
  assign data_o[18441] = data_o[9];
  assign data_o[18505] = data_o[9];
  assign data_o[18569] = data_o[9];
  assign data_o[18633] = data_o[9];
  assign data_o[18697] = data_o[9];
  assign data_o[18761] = data_o[9];
  assign data_o[18825] = data_o[9];
  assign data_o[18889] = data_o[9];
  assign data_o[18953] = data_o[9];
  assign data_o[19017] = data_o[9];
  assign data_o[19081] = data_o[9];
  assign data_o[19145] = data_o[9];
  assign data_o[19209] = data_o[9];
  assign data_o[19273] = data_o[9];
  assign data_o[19337] = data_o[9];
  assign data_o[19401] = data_o[9];
  assign data_o[19465] = data_o[9];
  assign data_o[19529] = data_o[9];
  assign data_o[19593] = data_o[9];
  assign data_o[19657] = data_o[9];
  assign data_o[19721] = data_o[9];
  assign data_o[19785] = data_o[9];
  assign data_o[19849] = data_o[9];
  assign data_o[19913] = data_o[9];
  assign data_o[19977] = data_o[9];
  assign data_o[20041] = data_o[9];
  assign data_o[20105] = data_o[9];
  assign data_o[20169] = data_o[9];
  assign data_o[20233] = data_o[9];
  assign data_o[20297] = data_o[9];
  assign data_o[20361] = data_o[9];
  assign data_o[20425] = data_o[9];
  assign data_o[20489] = data_o[9];
  assign data_o[20553] = data_o[9];
  assign data_o[20617] = data_o[9];
  assign data_o[20681] = data_o[9];
  assign data_o[20745] = data_o[9];
  assign data_o[20809] = data_o[9];
  assign data_o[20873] = data_o[9];
  assign data_o[20937] = data_o[9];
  assign data_o[21001] = data_o[9];
  assign data_o[21065] = data_o[9];
  assign data_o[21129] = data_o[9];
  assign data_o[21193] = data_o[9];
  assign data_o[21257] = data_o[9];
  assign data_o[21321] = data_o[9];
  assign data_o[21385] = data_o[9];
  assign data_o[21449] = data_o[9];
  assign data_o[21513] = data_o[9];
  assign data_o[21577] = data_o[9];
  assign data_o[21641] = data_o[9];
  assign data_o[21705] = data_o[9];
  assign data_o[21769] = data_o[9];
  assign data_o[21833] = data_o[9];
  assign data_o[21897] = data_o[9];
  assign data_o[21961] = data_o[9];
  assign data_o[22025] = data_o[9];
  assign data_o[22089] = data_o[9];
  assign data_o[22153] = data_o[9];
  assign data_o[22217] = data_o[9];
  assign data_o[22281] = data_o[9];
  assign data_o[22345] = data_o[9];
  assign data_o[22409] = data_o[9];
  assign data_o[22473] = data_o[9];
  assign data_o[22537] = data_o[9];
  assign data_o[22601] = data_o[9];
  assign data_o[22665] = data_o[9];
  assign data_o[22729] = data_o[9];
  assign data_o[22793] = data_o[9];
  assign data_o[22857] = data_o[9];
  assign data_o[22921] = data_o[9];
  assign data_o[22985] = data_o[9];
  assign data_o[23049] = data_o[9];
  assign data_o[23113] = data_o[9];
  assign data_o[23177] = data_o[9];
  assign data_o[23241] = data_o[9];
  assign data_o[23305] = data_o[9];
  assign data_o[23369] = data_o[9];
  assign data_o[23433] = data_o[9];
  assign data_o[23497] = data_o[9];
  assign data_o[23561] = data_o[9];
  assign data_o[23625] = data_o[9];
  assign data_o[23689] = data_o[9];
  assign data_o[23753] = data_o[9];
  assign data_o[23817] = data_o[9];
  assign data_o[23881] = data_o[9];
  assign data_o[23945] = data_o[9];
  assign data_o[24009] = data_o[9];
  assign data_o[24073] = data_o[9];
  assign data_o[24137] = data_o[9];
  assign data_o[24201] = data_o[9];
  assign data_o[24265] = data_o[9];
  assign data_o[24329] = data_o[9];
  assign data_o[24393] = data_o[9];
  assign data_o[24457] = data_o[9];
  assign data_o[24521] = data_o[9];
  assign data_o[24585] = data_o[9];
  assign data_o[24649] = data_o[9];
  assign data_o[24713] = data_o[9];
  assign data_o[24777] = data_o[9];
  assign data_o[24841] = data_o[9];
  assign data_o[24905] = data_o[9];
  assign data_o[24969] = data_o[9];
  assign data_o[25033] = data_o[9];
  assign data_o[25097] = data_o[9];
  assign data_o[25161] = data_o[9];
  assign data_o[25225] = data_o[9];
  assign data_o[25289] = data_o[9];
  assign data_o[25353] = data_o[9];
  assign data_o[25417] = data_o[9];
  assign data_o[25481] = data_o[9];
  assign data_o[25545] = data_o[9];
  assign data_o[25609] = data_o[9];
  assign data_o[25673] = data_o[9];
  assign data_o[25737] = data_o[9];
  assign data_o[25801] = data_o[9];
  assign data_o[25865] = data_o[9];
  assign data_o[25929] = data_o[9];
  assign data_o[25993] = data_o[9];
  assign data_o[26057] = data_o[9];
  assign data_o[26121] = data_o[9];
  assign data_o[26185] = data_o[9];
  assign data_o[26249] = data_o[9];
  assign data_o[26313] = data_o[9];
  assign data_o[26377] = data_o[9];
  assign data_o[26441] = data_o[9];
  assign data_o[26505] = data_o[9];
  assign data_o[26569] = data_o[9];
  assign data_o[26633] = data_o[9];
  assign data_o[26697] = data_o[9];
  assign data_o[26761] = data_o[9];
  assign data_o[26825] = data_o[9];
  assign data_o[26889] = data_o[9];
  assign data_o[26953] = data_o[9];
  assign data_o[27017] = data_o[9];
  assign data_o[27081] = data_o[9];
  assign data_o[27145] = data_o[9];
  assign data_o[27209] = data_o[9];
  assign data_o[27273] = data_o[9];
  assign data_o[27337] = data_o[9];
  assign data_o[27401] = data_o[9];
  assign data_o[27465] = data_o[9];
  assign data_o[27529] = data_o[9];
  assign data_o[27593] = data_o[9];
  assign data_o[27657] = data_o[9];
  assign data_o[27721] = data_o[9];
  assign data_o[27785] = data_o[9];
  assign data_o[27849] = data_o[9];
  assign data_o[27913] = data_o[9];
  assign data_o[27977] = data_o[9];
  assign data_o[28041] = data_o[9];
  assign data_o[28105] = data_o[9];
  assign data_o[28169] = data_o[9];
  assign data_o[28233] = data_o[9];
  assign data_o[28297] = data_o[9];
  assign data_o[28361] = data_o[9];
  assign data_o[28425] = data_o[9];
  assign data_o[28489] = data_o[9];
  assign data_o[28553] = data_o[9];
  assign data_o[28617] = data_o[9];
  assign data_o[28681] = data_o[9];
  assign data_o[28745] = data_o[9];
  assign data_o[28809] = data_o[9];
  assign data_o[28873] = data_o[9];
  assign data_o[28937] = data_o[9];
  assign data_o[29001] = data_o[9];
  assign data_o[29065] = data_o[9];
  assign data_o[29129] = data_o[9];
  assign data_o[29193] = data_o[9];
  assign data_o[29257] = data_o[9];
  assign data_o[29321] = data_o[9];
  assign data_o[29385] = data_o[9];
  assign data_o[29449] = data_o[9];
  assign data_o[29513] = data_o[9];
  assign data_o[29577] = data_o[9];
  assign data_o[29641] = data_o[9];
  assign data_o[29705] = data_o[9];
  assign data_o[29769] = data_o[9];
  assign data_o[29833] = data_o[9];
  assign data_o[29897] = data_o[9];
  assign data_o[29961] = data_o[9];
  assign data_o[30025] = data_o[9];
  assign data_o[30089] = data_o[9];
  assign data_o[30153] = data_o[9];
  assign data_o[30217] = data_o[9];
  assign data_o[30281] = data_o[9];
  assign data_o[30345] = data_o[9];
  assign data_o[30409] = data_o[9];
  assign data_o[30473] = data_o[9];
  assign data_o[30537] = data_o[9];
  assign data_o[30601] = data_o[9];
  assign data_o[30665] = data_o[9];
  assign data_o[30729] = data_o[9];
  assign data_o[30793] = data_o[9];
  assign data_o[30857] = data_o[9];
  assign data_o[30921] = data_o[9];
  assign data_o[30985] = data_o[9];
  assign data_o[31049] = data_o[9];
  assign data_o[31113] = data_o[9];
  assign data_o[31177] = data_o[9];
  assign data_o[31241] = data_o[9];
  assign data_o[31305] = data_o[9];
  assign data_o[31369] = data_o[9];
  assign data_o[31433] = data_o[9];
  assign data_o[31497] = data_o[9];
  assign data_o[31561] = data_o[9];
  assign data_o[31625] = data_o[9];
  assign data_o[31689] = data_o[9];
  assign data_o[31753] = data_o[9];
  assign data_o[31817] = data_o[9];
  assign data_o[31881] = data_o[9];
  assign data_o[31945] = data_o[9];
  assign data_o[72] = data_o[8];
  assign data_o[136] = data_o[8];
  assign data_o[200] = data_o[8];
  assign data_o[264] = data_o[8];
  assign data_o[328] = data_o[8];
  assign data_o[392] = data_o[8];
  assign data_o[456] = data_o[8];
  assign data_o[520] = data_o[8];
  assign data_o[584] = data_o[8];
  assign data_o[648] = data_o[8];
  assign data_o[712] = data_o[8];
  assign data_o[776] = data_o[8];
  assign data_o[840] = data_o[8];
  assign data_o[904] = data_o[8];
  assign data_o[968] = data_o[8];
  assign data_o[1032] = data_o[8];
  assign data_o[1096] = data_o[8];
  assign data_o[1160] = data_o[8];
  assign data_o[1224] = data_o[8];
  assign data_o[1288] = data_o[8];
  assign data_o[1352] = data_o[8];
  assign data_o[1416] = data_o[8];
  assign data_o[1480] = data_o[8];
  assign data_o[1544] = data_o[8];
  assign data_o[1608] = data_o[8];
  assign data_o[1672] = data_o[8];
  assign data_o[1736] = data_o[8];
  assign data_o[1800] = data_o[8];
  assign data_o[1864] = data_o[8];
  assign data_o[1928] = data_o[8];
  assign data_o[1992] = data_o[8];
  assign data_o[2056] = data_o[8];
  assign data_o[2120] = data_o[8];
  assign data_o[2184] = data_o[8];
  assign data_o[2248] = data_o[8];
  assign data_o[2312] = data_o[8];
  assign data_o[2376] = data_o[8];
  assign data_o[2440] = data_o[8];
  assign data_o[2504] = data_o[8];
  assign data_o[2568] = data_o[8];
  assign data_o[2632] = data_o[8];
  assign data_o[2696] = data_o[8];
  assign data_o[2760] = data_o[8];
  assign data_o[2824] = data_o[8];
  assign data_o[2888] = data_o[8];
  assign data_o[2952] = data_o[8];
  assign data_o[3016] = data_o[8];
  assign data_o[3080] = data_o[8];
  assign data_o[3144] = data_o[8];
  assign data_o[3208] = data_o[8];
  assign data_o[3272] = data_o[8];
  assign data_o[3336] = data_o[8];
  assign data_o[3400] = data_o[8];
  assign data_o[3464] = data_o[8];
  assign data_o[3528] = data_o[8];
  assign data_o[3592] = data_o[8];
  assign data_o[3656] = data_o[8];
  assign data_o[3720] = data_o[8];
  assign data_o[3784] = data_o[8];
  assign data_o[3848] = data_o[8];
  assign data_o[3912] = data_o[8];
  assign data_o[3976] = data_o[8];
  assign data_o[4040] = data_o[8];
  assign data_o[4104] = data_o[8];
  assign data_o[4168] = data_o[8];
  assign data_o[4232] = data_o[8];
  assign data_o[4296] = data_o[8];
  assign data_o[4360] = data_o[8];
  assign data_o[4424] = data_o[8];
  assign data_o[4488] = data_o[8];
  assign data_o[4552] = data_o[8];
  assign data_o[4616] = data_o[8];
  assign data_o[4680] = data_o[8];
  assign data_o[4744] = data_o[8];
  assign data_o[4808] = data_o[8];
  assign data_o[4872] = data_o[8];
  assign data_o[4936] = data_o[8];
  assign data_o[5000] = data_o[8];
  assign data_o[5064] = data_o[8];
  assign data_o[5128] = data_o[8];
  assign data_o[5192] = data_o[8];
  assign data_o[5256] = data_o[8];
  assign data_o[5320] = data_o[8];
  assign data_o[5384] = data_o[8];
  assign data_o[5448] = data_o[8];
  assign data_o[5512] = data_o[8];
  assign data_o[5576] = data_o[8];
  assign data_o[5640] = data_o[8];
  assign data_o[5704] = data_o[8];
  assign data_o[5768] = data_o[8];
  assign data_o[5832] = data_o[8];
  assign data_o[5896] = data_o[8];
  assign data_o[5960] = data_o[8];
  assign data_o[6024] = data_o[8];
  assign data_o[6088] = data_o[8];
  assign data_o[6152] = data_o[8];
  assign data_o[6216] = data_o[8];
  assign data_o[6280] = data_o[8];
  assign data_o[6344] = data_o[8];
  assign data_o[6408] = data_o[8];
  assign data_o[6472] = data_o[8];
  assign data_o[6536] = data_o[8];
  assign data_o[6600] = data_o[8];
  assign data_o[6664] = data_o[8];
  assign data_o[6728] = data_o[8];
  assign data_o[6792] = data_o[8];
  assign data_o[6856] = data_o[8];
  assign data_o[6920] = data_o[8];
  assign data_o[6984] = data_o[8];
  assign data_o[7048] = data_o[8];
  assign data_o[7112] = data_o[8];
  assign data_o[7176] = data_o[8];
  assign data_o[7240] = data_o[8];
  assign data_o[7304] = data_o[8];
  assign data_o[7368] = data_o[8];
  assign data_o[7432] = data_o[8];
  assign data_o[7496] = data_o[8];
  assign data_o[7560] = data_o[8];
  assign data_o[7624] = data_o[8];
  assign data_o[7688] = data_o[8];
  assign data_o[7752] = data_o[8];
  assign data_o[7816] = data_o[8];
  assign data_o[7880] = data_o[8];
  assign data_o[7944] = data_o[8];
  assign data_o[8008] = data_o[8];
  assign data_o[8072] = data_o[8];
  assign data_o[8136] = data_o[8];
  assign data_o[8200] = data_o[8];
  assign data_o[8264] = data_o[8];
  assign data_o[8328] = data_o[8];
  assign data_o[8392] = data_o[8];
  assign data_o[8456] = data_o[8];
  assign data_o[8520] = data_o[8];
  assign data_o[8584] = data_o[8];
  assign data_o[8648] = data_o[8];
  assign data_o[8712] = data_o[8];
  assign data_o[8776] = data_o[8];
  assign data_o[8840] = data_o[8];
  assign data_o[8904] = data_o[8];
  assign data_o[8968] = data_o[8];
  assign data_o[9032] = data_o[8];
  assign data_o[9096] = data_o[8];
  assign data_o[9160] = data_o[8];
  assign data_o[9224] = data_o[8];
  assign data_o[9288] = data_o[8];
  assign data_o[9352] = data_o[8];
  assign data_o[9416] = data_o[8];
  assign data_o[9480] = data_o[8];
  assign data_o[9544] = data_o[8];
  assign data_o[9608] = data_o[8];
  assign data_o[9672] = data_o[8];
  assign data_o[9736] = data_o[8];
  assign data_o[9800] = data_o[8];
  assign data_o[9864] = data_o[8];
  assign data_o[9928] = data_o[8];
  assign data_o[9992] = data_o[8];
  assign data_o[10056] = data_o[8];
  assign data_o[10120] = data_o[8];
  assign data_o[10184] = data_o[8];
  assign data_o[10248] = data_o[8];
  assign data_o[10312] = data_o[8];
  assign data_o[10376] = data_o[8];
  assign data_o[10440] = data_o[8];
  assign data_o[10504] = data_o[8];
  assign data_o[10568] = data_o[8];
  assign data_o[10632] = data_o[8];
  assign data_o[10696] = data_o[8];
  assign data_o[10760] = data_o[8];
  assign data_o[10824] = data_o[8];
  assign data_o[10888] = data_o[8];
  assign data_o[10952] = data_o[8];
  assign data_o[11016] = data_o[8];
  assign data_o[11080] = data_o[8];
  assign data_o[11144] = data_o[8];
  assign data_o[11208] = data_o[8];
  assign data_o[11272] = data_o[8];
  assign data_o[11336] = data_o[8];
  assign data_o[11400] = data_o[8];
  assign data_o[11464] = data_o[8];
  assign data_o[11528] = data_o[8];
  assign data_o[11592] = data_o[8];
  assign data_o[11656] = data_o[8];
  assign data_o[11720] = data_o[8];
  assign data_o[11784] = data_o[8];
  assign data_o[11848] = data_o[8];
  assign data_o[11912] = data_o[8];
  assign data_o[11976] = data_o[8];
  assign data_o[12040] = data_o[8];
  assign data_o[12104] = data_o[8];
  assign data_o[12168] = data_o[8];
  assign data_o[12232] = data_o[8];
  assign data_o[12296] = data_o[8];
  assign data_o[12360] = data_o[8];
  assign data_o[12424] = data_o[8];
  assign data_o[12488] = data_o[8];
  assign data_o[12552] = data_o[8];
  assign data_o[12616] = data_o[8];
  assign data_o[12680] = data_o[8];
  assign data_o[12744] = data_o[8];
  assign data_o[12808] = data_o[8];
  assign data_o[12872] = data_o[8];
  assign data_o[12936] = data_o[8];
  assign data_o[13000] = data_o[8];
  assign data_o[13064] = data_o[8];
  assign data_o[13128] = data_o[8];
  assign data_o[13192] = data_o[8];
  assign data_o[13256] = data_o[8];
  assign data_o[13320] = data_o[8];
  assign data_o[13384] = data_o[8];
  assign data_o[13448] = data_o[8];
  assign data_o[13512] = data_o[8];
  assign data_o[13576] = data_o[8];
  assign data_o[13640] = data_o[8];
  assign data_o[13704] = data_o[8];
  assign data_o[13768] = data_o[8];
  assign data_o[13832] = data_o[8];
  assign data_o[13896] = data_o[8];
  assign data_o[13960] = data_o[8];
  assign data_o[14024] = data_o[8];
  assign data_o[14088] = data_o[8];
  assign data_o[14152] = data_o[8];
  assign data_o[14216] = data_o[8];
  assign data_o[14280] = data_o[8];
  assign data_o[14344] = data_o[8];
  assign data_o[14408] = data_o[8];
  assign data_o[14472] = data_o[8];
  assign data_o[14536] = data_o[8];
  assign data_o[14600] = data_o[8];
  assign data_o[14664] = data_o[8];
  assign data_o[14728] = data_o[8];
  assign data_o[14792] = data_o[8];
  assign data_o[14856] = data_o[8];
  assign data_o[14920] = data_o[8];
  assign data_o[14984] = data_o[8];
  assign data_o[15048] = data_o[8];
  assign data_o[15112] = data_o[8];
  assign data_o[15176] = data_o[8];
  assign data_o[15240] = data_o[8];
  assign data_o[15304] = data_o[8];
  assign data_o[15368] = data_o[8];
  assign data_o[15432] = data_o[8];
  assign data_o[15496] = data_o[8];
  assign data_o[15560] = data_o[8];
  assign data_o[15624] = data_o[8];
  assign data_o[15688] = data_o[8];
  assign data_o[15752] = data_o[8];
  assign data_o[15816] = data_o[8];
  assign data_o[15880] = data_o[8];
  assign data_o[15944] = data_o[8];
  assign data_o[16008] = data_o[8];
  assign data_o[16072] = data_o[8];
  assign data_o[16136] = data_o[8];
  assign data_o[16200] = data_o[8];
  assign data_o[16264] = data_o[8];
  assign data_o[16328] = data_o[8];
  assign data_o[16392] = data_o[8];
  assign data_o[16456] = data_o[8];
  assign data_o[16520] = data_o[8];
  assign data_o[16584] = data_o[8];
  assign data_o[16648] = data_o[8];
  assign data_o[16712] = data_o[8];
  assign data_o[16776] = data_o[8];
  assign data_o[16840] = data_o[8];
  assign data_o[16904] = data_o[8];
  assign data_o[16968] = data_o[8];
  assign data_o[17032] = data_o[8];
  assign data_o[17096] = data_o[8];
  assign data_o[17160] = data_o[8];
  assign data_o[17224] = data_o[8];
  assign data_o[17288] = data_o[8];
  assign data_o[17352] = data_o[8];
  assign data_o[17416] = data_o[8];
  assign data_o[17480] = data_o[8];
  assign data_o[17544] = data_o[8];
  assign data_o[17608] = data_o[8];
  assign data_o[17672] = data_o[8];
  assign data_o[17736] = data_o[8];
  assign data_o[17800] = data_o[8];
  assign data_o[17864] = data_o[8];
  assign data_o[17928] = data_o[8];
  assign data_o[17992] = data_o[8];
  assign data_o[18056] = data_o[8];
  assign data_o[18120] = data_o[8];
  assign data_o[18184] = data_o[8];
  assign data_o[18248] = data_o[8];
  assign data_o[18312] = data_o[8];
  assign data_o[18376] = data_o[8];
  assign data_o[18440] = data_o[8];
  assign data_o[18504] = data_o[8];
  assign data_o[18568] = data_o[8];
  assign data_o[18632] = data_o[8];
  assign data_o[18696] = data_o[8];
  assign data_o[18760] = data_o[8];
  assign data_o[18824] = data_o[8];
  assign data_o[18888] = data_o[8];
  assign data_o[18952] = data_o[8];
  assign data_o[19016] = data_o[8];
  assign data_o[19080] = data_o[8];
  assign data_o[19144] = data_o[8];
  assign data_o[19208] = data_o[8];
  assign data_o[19272] = data_o[8];
  assign data_o[19336] = data_o[8];
  assign data_o[19400] = data_o[8];
  assign data_o[19464] = data_o[8];
  assign data_o[19528] = data_o[8];
  assign data_o[19592] = data_o[8];
  assign data_o[19656] = data_o[8];
  assign data_o[19720] = data_o[8];
  assign data_o[19784] = data_o[8];
  assign data_o[19848] = data_o[8];
  assign data_o[19912] = data_o[8];
  assign data_o[19976] = data_o[8];
  assign data_o[20040] = data_o[8];
  assign data_o[20104] = data_o[8];
  assign data_o[20168] = data_o[8];
  assign data_o[20232] = data_o[8];
  assign data_o[20296] = data_o[8];
  assign data_o[20360] = data_o[8];
  assign data_o[20424] = data_o[8];
  assign data_o[20488] = data_o[8];
  assign data_o[20552] = data_o[8];
  assign data_o[20616] = data_o[8];
  assign data_o[20680] = data_o[8];
  assign data_o[20744] = data_o[8];
  assign data_o[20808] = data_o[8];
  assign data_o[20872] = data_o[8];
  assign data_o[20936] = data_o[8];
  assign data_o[21000] = data_o[8];
  assign data_o[21064] = data_o[8];
  assign data_o[21128] = data_o[8];
  assign data_o[21192] = data_o[8];
  assign data_o[21256] = data_o[8];
  assign data_o[21320] = data_o[8];
  assign data_o[21384] = data_o[8];
  assign data_o[21448] = data_o[8];
  assign data_o[21512] = data_o[8];
  assign data_o[21576] = data_o[8];
  assign data_o[21640] = data_o[8];
  assign data_o[21704] = data_o[8];
  assign data_o[21768] = data_o[8];
  assign data_o[21832] = data_o[8];
  assign data_o[21896] = data_o[8];
  assign data_o[21960] = data_o[8];
  assign data_o[22024] = data_o[8];
  assign data_o[22088] = data_o[8];
  assign data_o[22152] = data_o[8];
  assign data_o[22216] = data_o[8];
  assign data_o[22280] = data_o[8];
  assign data_o[22344] = data_o[8];
  assign data_o[22408] = data_o[8];
  assign data_o[22472] = data_o[8];
  assign data_o[22536] = data_o[8];
  assign data_o[22600] = data_o[8];
  assign data_o[22664] = data_o[8];
  assign data_o[22728] = data_o[8];
  assign data_o[22792] = data_o[8];
  assign data_o[22856] = data_o[8];
  assign data_o[22920] = data_o[8];
  assign data_o[22984] = data_o[8];
  assign data_o[23048] = data_o[8];
  assign data_o[23112] = data_o[8];
  assign data_o[23176] = data_o[8];
  assign data_o[23240] = data_o[8];
  assign data_o[23304] = data_o[8];
  assign data_o[23368] = data_o[8];
  assign data_o[23432] = data_o[8];
  assign data_o[23496] = data_o[8];
  assign data_o[23560] = data_o[8];
  assign data_o[23624] = data_o[8];
  assign data_o[23688] = data_o[8];
  assign data_o[23752] = data_o[8];
  assign data_o[23816] = data_o[8];
  assign data_o[23880] = data_o[8];
  assign data_o[23944] = data_o[8];
  assign data_o[24008] = data_o[8];
  assign data_o[24072] = data_o[8];
  assign data_o[24136] = data_o[8];
  assign data_o[24200] = data_o[8];
  assign data_o[24264] = data_o[8];
  assign data_o[24328] = data_o[8];
  assign data_o[24392] = data_o[8];
  assign data_o[24456] = data_o[8];
  assign data_o[24520] = data_o[8];
  assign data_o[24584] = data_o[8];
  assign data_o[24648] = data_o[8];
  assign data_o[24712] = data_o[8];
  assign data_o[24776] = data_o[8];
  assign data_o[24840] = data_o[8];
  assign data_o[24904] = data_o[8];
  assign data_o[24968] = data_o[8];
  assign data_o[25032] = data_o[8];
  assign data_o[25096] = data_o[8];
  assign data_o[25160] = data_o[8];
  assign data_o[25224] = data_o[8];
  assign data_o[25288] = data_o[8];
  assign data_o[25352] = data_o[8];
  assign data_o[25416] = data_o[8];
  assign data_o[25480] = data_o[8];
  assign data_o[25544] = data_o[8];
  assign data_o[25608] = data_o[8];
  assign data_o[25672] = data_o[8];
  assign data_o[25736] = data_o[8];
  assign data_o[25800] = data_o[8];
  assign data_o[25864] = data_o[8];
  assign data_o[25928] = data_o[8];
  assign data_o[25992] = data_o[8];
  assign data_o[26056] = data_o[8];
  assign data_o[26120] = data_o[8];
  assign data_o[26184] = data_o[8];
  assign data_o[26248] = data_o[8];
  assign data_o[26312] = data_o[8];
  assign data_o[26376] = data_o[8];
  assign data_o[26440] = data_o[8];
  assign data_o[26504] = data_o[8];
  assign data_o[26568] = data_o[8];
  assign data_o[26632] = data_o[8];
  assign data_o[26696] = data_o[8];
  assign data_o[26760] = data_o[8];
  assign data_o[26824] = data_o[8];
  assign data_o[26888] = data_o[8];
  assign data_o[26952] = data_o[8];
  assign data_o[27016] = data_o[8];
  assign data_o[27080] = data_o[8];
  assign data_o[27144] = data_o[8];
  assign data_o[27208] = data_o[8];
  assign data_o[27272] = data_o[8];
  assign data_o[27336] = data_o[8];
  assign data_o[27400] = data_o[8];
  assign data_o[27464] = data_o[8];
  assign data_o[27528] = data_o[8];
  assign data_o[27592] = data_o[8];
  assign data_o[27656] = data_o[8];
  assign data_o[27720] = data_o[8];
  assign data_o[27784] = data_o[8];
  assign data_o[27848] = data_o[8];
  assign data_o[27912] = data_o[8];
  assign data_o[27976] = data_o[8];
  assign data_o[28040] = data_o[8];
  assign data_o[28104] = data_o[8];
  assign data_o[28168] = data_o[8];
  assign data_o[28232] = data_o[8];
  assign data_o[28296] = data_o[8];
  assign data_o[28360] = data_o[8];
  assign data_o[28424] = data_o[8];
  assign data_o[28488] = data_o[8];
  assign data_o[28552] = data_o[8];
  assign data_o[28616] = data_o[8];
  assign data_o[28680] = data_o[8];
  assign data_o[28744] = data_o[8];
  assign data_o[28808] = data_o[8];
  assign data_o[28872] = data_o[8];
  assign data_o[28936] = data_o[8];
  assign data_o[29000] = data_o[8];
  assign data_o[29064] = data_o[8];
  assign data_o[29128] = data_o[8];
  assign data_o[29192] = data_o[8];
  assign data_o[29256] = data_o[8];
  assign data_o[29320] = data_o[8];
  assign data_o[29384] = data_o[8];
  assign data_o[29448] = data_o[8];
  assign data_o[29512] = data_o[8];
  assign data_o[29576] = data_o[8];
  assign data_o[29640] = data_o[8];
  assign data_o[29704] = data_o[8];
  assign data_o[29768] = data_o[8];
  assign data_o[29832] = data_o[8];
  assign data_o[29896] = data_o[8];
  assign data_o[29960] = data_o[8];
  assign data_o[30024] = data_o[8];
  assign data_o[30088] = data_o[8];
  assign data_o[30152] = data_o[8];
  assign data_o[30216] = data_o[8];
  assign data_o[30280] = data_o[8];
  assign data_o[30344] = data_o[8];
  assign data_o[30408] = data_o[8];
  assign data_o[30472] = data_o[8];
  assign data_o[30536] = data_o[8];
  assign data_o[30600] = data_o[8];
  assign data_o[30664] = data_o[8];
  assign data_o[30728] = data_o[8];
  assign data_o[30792] = data_o[8];
  assign data_o[30856] = data_o[8];
  assign data_o[30920] = data_o[8];
  assign data_o[30984] = data_o[8];
  assign data_o[31048] = data_o[8];
  assign data_o[31112] = data_o[8];
  assign data_o[31176] = data_o[8];
  assign data_o[31240] = data_o[8];
  assign data_o[31304] = data_o[8];
  assign data_o[31368] = data_o[8];
  assign data_o[31432] = data_o[8];
  assign data_o[31496] = data_o[8];
  assign data_o[31560] = data_o[8];
  assign data_o[31624] = data_o[8];
  assign data_o[31688] = data_o[8];
  assign data_o[31752] = data_o[8];
  assign data_o[31816] = data_o[8];
  assign data_o[31880] = data_o[8];
  assign data_o[31944] = data_o[8];
  assign data_o[71] = data_o[7];
  assign data_o[135] = data_o[7];
  assign data_o[199] = data_o[7];
  assign data_o[263] = data_o[7];
  assign data_o[327] = data_o[7];
  assign data_o[391] = data_o[7];
  assign data_o[455] = data_o[7];
  assign data_o[519] = data_o[7];
  assign data_o[583] = data_o[7];
  assign data_o[647] = data_o[7];
  assign data_o[711] = data_o[7];
  assign data_o[775] = data_o[7];
  assign data_o[839] = data_o[7];
  assign data_o[903] = data_o[7];
  assign data_o[967] = data_o[7];
  assign data_o[1031] = data_o[7];
  assign data_o[1095] = data_o[7];
  assign data_o[1159] = data_o[7];
  assign data_o[1223] = data_o[7];
  assign data_o[1287] = data_o[7];
  assign data_o[1351] = data_o[7];
  assign data_o[1415] = data_o[7];
  assign data_o[1479] = data_o[7];
  assign data_o[1543] = data_o[7];
  assign data_o[1607] = data_o[7];
  assign data_o[1671] = data_o[7];
  assign data_o[1735] = data_o[7];
  assign data_o[1799] = data_o[7];
  assign data_o[1863] = data_o[7];
  assign data_o[1927] = data_o[7];
  assign data_o[1991] = data_o[7];
  assign data_o[2055] = data_o[7];
  assign data_o[2119] = data_o[7];
  assign data_o[2183] = data_o[7];
  assign data_o[2247] = data_o[7];
  assign data_o[2311] = data_o[7];
  assign data_o[2375] = data_o[7];
  assign data_o[2439] = data_o[7];
  assign data_o[2503] = data_o[7];
  assign data_o[2567] = data_o[7];
  assign data_o[2631] = data_o[7];
  assign data_o[2695] = data_o[7];
  assign data_o[2759] = data_o[7];
  assign data_o[2823] = data_o[7];
  assign data_o[2887] = data_o[7];
  assign data_o[2951] = data_o[7];
  assign data_o[3015] = data_o[7];
  assign data_o[3079] = data_o[7];
  assign data_o[3143] = data_o[7];
  assign data_o[3207] = data_o[7];
  assign data_o[3271] = data_o[7];
  assign data_o[3335] = data_o[7];
  assign data_o[3399] = data_o[7];
  assign data_o[3463] = data_o[7];
  assign data_o[3527] = data_o[7];
  assign data_o[3591] = data_o[7];
  assign data_o[3655] = data_o[7];
  assign data_o[3719] = data_o[7];
  assign data_o[3783] = data_o[7];
  assign data_o[3847] = data_o[7];
  assign data_o[3911] = data_o[7];
  assign data_o[3975] = data_o[7];
  assign data_o[4039] = data_o[7];
  assign data_o[4103] = data_o[7];
  assign data_o[4167] = data_o[7];
  assign data_o[4231] = data_o[7];
  assign data_o[4295] = data_o[7];
  assign data_o[4359] = data_o[7];
  assign data_o[4423] = data_o[7];
  assign data_o[4487] = data_o[7];
  assign data_o[4551] = data_o[7];
  assign data_o[4615] = data_o[7];
  assign data_o[4679] = data_o[7];
  assign data_o[4743] = data_o[7];
  assign data_o[4807] = data_o[7];
  assign data_o[4871] = data_o[7];
  assign data_o[4935] = data_o[7];
  assign data_o[4999] = data_o[7];
  assign data_o[5063] = data_o[7];
  assign data_o[5127] = data_o[7];
  assign data_o[5191] = data_o[7];
  assign data_o[5255] = data_o[7];
  assign data_o[5319] = data_o[7];
  assign data_o[5383] = data_o[7];
  assign data_o[5447] = data_o[7];
  assign data_o[5511] = data_o[7];
  assign data_o[5575] = data_o[7];
  assign data_o[5639] = data_o[7];
  assign data_o[5703] = data_o[7];
  assign data_o[5767] = data_o[7];
  assign data_o[5831] = data_o[7];
  assign data_o[5895] = data_o[7];
  assign data_o[5959] = data_o[7];
  assign data_o[6023] = data_o[7];
  assign data_o[6087] = data_o[7];
  assign data_o[6151] = data_o[7];
  assign data_o[6215] = data_o[7];
  assign data_o[6279] = data_o[7];
  assign data_o[6343] = data_o[7];
  assign data_o[6407] = data_o[7];
  assign data_o[6471] = data_o[7];
  assign data_o[6535] = data_o[7];
  assign data_o[6599] = data_o[7];
  assign data_o[6663] = data_o[7];
  assign data_o[6727] = data_o[7];
  assign data_o[6791] = data_o[7];
  assign data_o[6855] = data_o[7];
  assign data_o[6919] = data_o[7];
  assign data_o[6983] = data_o[7];
  assign data_o[7047] = data_o[7];
  assign data_o[7111] = data_o[7];
  assign data_o[7175] = data_o[7];
  assign data_o[7239] = data_o[7];
  assign data_o[7303] = data_o[7];
  assign data_o[7367] = data_o[7];
  assign data_o[7431] = data_o[7];
  assign data_o[7495] = data_o[7];
  assign data_o[7559] = data_o[7];
  assign data_o[7623] = data_o[7];
  assign data_o[7687] = data_o[7];
  assign data_o[7751] = data_o[7];
  assign data_o[7815] = data_o[7];
  assign data_o[7879] = data_o[7];
  assign data_o[7943] = data_o[7];
  assign data_o[8007] = data_o[7];
  assign data_o[8071] = data_o[7];
  assign data_o[8135] = data_o[7];
  assign data_o[8199] = data_o[7];
  assign data_o[8263] = data_o[7];
  assign data_o[8327] = data_o[7];
  assign data_o[8391] = data_o[7];
  assign data_o[8455] = data_o[7];
  assign data_o[8519] = data_o[7];
  assign data_o[8583] = data_o[7];
  assign data_o[8647] = data_o[7];
  assign data_o[8711] = data_o[7];
  assign data_o[8775] = data_o[7];
  assign data_o[8839] = data_o[7];
  assign data_o[8903] = data_o[7];
  assign data_o[8967] = data_o[7];
  assign data_o[9031] = data_o[7];
  assign data_o[9095] = data_o[7];
  assign data_o[9159] = data_o[7];
  assign data_o[9223] = data_o[7];
  assign data_o[9287] = data_o[7];
  assign data_o[9351] = data_o[7];
  assign data_o[9415] = data_o[7];
  assign data_o[9479] = data_o[7];
  assign data_o[9543] = data_o[7];
  assign data_o[9607] = data_o[7];
  assign data_o[9671] = data_o[7];
  assign data_o[9735] = data_o[7];
  assign data_o[9799] = data_o[7];
  assign data_o[9863] = data_o[7];
  assign data_o[9927] = data_o[7];
  assign data_o[9991] = data_o[7];
  assign data_o[10055] = data_o[7];
  assign data_o[10119] = data_o[7];
  assign data_o[10183] = data_o[7];
  assign data_o[10247] = data_o[7];
  assign data_o[10311] = data_o[7];
  assign data_o[10375] = data_o[7];
  assign data_o[10439] = data_o[7];
  assign data_o[10503] = data_o[7];
  assign data_o[10567] = data_o[7];
  assign data_o[10631] = data_o[7];
  assign data_o[10695] = data_o[7];
  assign data_o[10759] = data_o[7];
  assign data_o[10823] = data_o[7];
  assign data_o[10887] = data_o[7];
  assign data_o[10951] = data_o[7];
  assign data_o[11015] = data_o[7];
  assign data_o[11079] = data_o[7];
  assign data_o[11143] = data_o[7];
  assign data_o[11207] = data_o[7];
  assign data_o[11271] = data_o[7];
  assign data_o[11335] = data_o[7];
  assign data_o[11399] = data_o[7];
  assign data_o[11463] = data_o[7];
  assign data_o[11527] = data_o[7];
  assign data_o[11591] = data_o[7];
  assign data_o[11655] = data_o[7];
  assign data_o[11719] = data_o[7];
  assign data_o[11783] = data_o[7];
  assign data_o[11847] = data_o[7];
  assign data_o[11911] = data_o[7];
  assign data_o[11975] = data_o[7];
  assign data_o[12039] = data_o[7];
  assign data_o[12103] = data_o[7];
  assign data_o[12167] = data_o[7];
  assign data_o[12231] = data_o[7];
  assign data_o[12295] = data_o[7];
  assign data_o[12359] = data_o[7];
  assign data_o[12423] = data_o[7];
  assign data_o[12487] = data_o[7];
  assign data_o[12551] = data_o[7];
  assign data_o[12615] = data_o[7];
  assign data_o[12679] = data_o[7];
  assign data_o[12743] = data_o[7];
  assign data_o[12807] = data_o[7];
  assign data_o[12871] = data_o[7];
  assign data_o[12935] = data_o[7];
  assign data_o[12999] = data_o[7];
  assign data_o[13063] = data_o[7];
  assign data_o[13127] = data_o[7];
  assign data_o[13191] = data_o[7];
  assign data_o[13255] = data_o[7];
  assign data_o[13319] = data_o[7];
  assign data_o[13383] = data_o[7];
  assign data_o[13447] = data_o[7];
  assign data_o[13511] = data_o[7];
  assign data_o[13575] = data_o[7];
  assign data_o[13639] = data_o[7];
  assign data_o[13703] = data_o[7];
  assign data_o[13767] = data_o[7];
  assign data_o[13831] = data_o[7];
  assign data_o[13895] = data_o[7];
  assign data_o[13959] = data_o[7];
  assign data_o[14023] = data_o[7];
  assign data_o[14087] = data_o[7];
  assign data_o[14151] = data_o[7];
  assign data_o[14215] = data_o[7];
  assign data_o[14279] = data_o[7];
  assign data_o[14343] = data_o[7];
  assign data_o[14407] = data_o[7];
  assign data_o[14471] = data_o[7];
  assign data_o[14535] = data_o[7];
  assign data_o[14599] = data_o[7];
  assign data_o[14663] = data_o[7];
  assign data_o[14727] = data_o[7];
  assign data_o[14791] = data_o[7];
  assign data_o[14855] = data_o[7];
  assign data_o[14919] = data_o[7];
  assign data_o[14983] = data_o[7];
  assign data_o[15047] = data_o[7];
  assign data_o[15111] = data_o[7];
  assign data_o[15175] = data_o[7];
  assign data_o[15239] = data_o[7];
  assign data_o[15303] = data_o[7];
  assign data_o[15367] = data_o[7];
  assign data_o[15431] = data_o[7];
  assign data_o[15495] = data_o[7];
  assign data_o[15559] = data_o[7];
  assign data_o[15623] = data_o[7];
  assign data_o[15687] = data_o[7];
  assign data_o[15751] = data_o[7];
  assign data_o[15815] = data_o[7];
  assign data_o[15879] = data_o[7];
  assign data_o[15943] = data_o[7];
  assign data_o[16007] = data_o[7];
  assign data_o[16071] = data_o[7];
  assign data_o[16135] = data_o[7];
  assign data_o[16199] = data_o[7];
  assign data_o[16263] = data_o[7];
  assign data_o[16327] = data_o[7];
  assign data_o[16391] = data_o[7];
  assign data_o[16455] = data_o[7];
  assign data_o[16519] = data_o[7];
  assign data_o[16583] = data_o[7];
  assign data_o[16647] = data_o[7];
  assign data_o[16711] = data_o[7];
  assign data_o[16775] = data_o[7];
  assign data_o[16839] = data_o[7];
  assign data_o[16903] = data_o[7];
  assign data_o[16967] = data_o[7];
  assign data_o[17031] = data_o[7];
  assign data_o[17095] = data_o[7];
  assign data_o[17159] = data_o[7];
  assign data_o[17223] = data_o[7];
  assign data_o[17287] = data_o[7];
  assign data_o[17351] = data_o[7];
  assign data_o[17415] = data_o[7];
  assign data_o[17479] = data_o[7];
  assign data_o[17543] = data_o[7];
  assign data_o[17607] = data_o[7];
  assign data_o[17671] = data_o[7];
  assign data_o[17735] = data_o[7];
  assign data_o[17799] = data_o[7];
  assign data_o[17863] = data_o[7];
  assign data_o[17927] = data_o[7];
  assign data_o[17991] = data_o[7];
  assign data_o[18055] = data_o[7];
  assign data_o[18119] = data_o[7];
  assign data_o[18183] = data_o[7];
  assign data_o[18247] = data_o[7];
  assign data_o[18311] = data_o[7];
  assign data_o[18375] = data_o[7];
  assign data_o[18439] = data_o[7];
  assign data_o[18503] = data_o[7];
  assign data_o[18567] = data_o[7];
  assign data_o[18631] = data_o[7];
  assign data_o[18695] = data_o[7];
  assign data_o[18759] = data_o[7];
  assign data_o[18823] = data_o[7];
  assign data_o[18887] = data_o[7];
  assign data_o[18951] = data_o[7];
  assign data_o[19015] = data_o[7];
  assign data_o[19079] = data_o[7];
  assign data_o[19143] = data_o[7];
  assign data_o[19207] = data_o[7];
  assign data_o[19271] = data_o[7];
  assign data_o[19335] = data_o[7];
  assign data_o[19399] = data_o[7];
  assign data_o[19463] = data_o[7];
  assign data_o[19527] = data_o[7];
  assign data_o[19591] = data_o[7];
  assign data_o[19655] = data_o[7];
  assign data_o[19719] = data_o[7];
  assign data_o[19783] = data_o[7];
  assign data_o[19847] = data_o[7];
  assign data_o[19911] = data_o[7];
  assign data_o[19975] = data_o[7];
  assign data_o[20039] = data_o[7];
  assign data_o[20103] = data_o[7];
  assign data_o[20167] = data_o[7];
  assign data_o[20231] = data_o[7];
  assign data_o[20295] = data_o[7];
  assign data_o[20359] = data_o[7];
  assign data_o[20423] = data_o[7];
  assign data_o[20487] = data_o[7];
  assign data_o[20551] = data_o[7];
  assign data_o[20615] = data_o[7];
  assign data_o[20679] = data_o[7];
  assign data_o[20743] = data_o[7];
  assign data_o[20807] = data_o[7];
  assign data_o[20871] = data_o[7];
  assign data_o[20935] = data_o[7];
  assign data_o[20999] = data_o[7];
  assign data_o[21063] = data_o[7];
  assign data_o[21127] = data_o[7];
  assign data_o[21191] = data_o[7];
  assign data_o[21255] = data_o[7];
  assign data_o[21319] = data_o[7];
  assign data_o[21383] = data_o[7];
  assign data_o[21447] = data_o[7];
  assign data_o[21511] = data_o[7];
  assign data_o[21575] = data_o[7];
  assign data_o[21639] = data_o[7];
  assign data_o[21703] = data_o[7];
  assign data_o[21767] = data_o[7];
  assign data_o[21831] = data_o[7];
  assign data_o[21895] = data_o[7];
  assign data_o[21959] = data_o[7];
  assign data_o[22023] = data_o[7];
  assign data_o[22087] = data_o[7];
  assign data_o[22151] = data_o[7];
  assign data_o[22215] = data_o[7];
  assign data_o[22279] = data_o[7];
  assign data_o[22343] = data_o[7];
  assign data_o[22407] = data_o[7];
  assign data_o[22471] = data_o[7];
  assign data_o[22535] = data_o[7];
  assign data_o[22599] = data_o[7];
  assign data_o[22663] = data_o[7];
  assign data_o[22727] = data_o[7];
  assign data_o[22791] = data_o[7];
  assign data_o[22855] = data_o[7];
  assign data_o[22919] = data_o[7];
  assign data_o[22983] = data_o[7];
  assign data_o[23047] = data_o[7];
  assign data_o[23111] = data_o[7];
  assign data_o[23175] = data_o[7];
  assign data_o[23239] = data_o[7];
  assign data_o[23303] = data_o[7];
  assign data_o[23367] = data_o[7];
  assign data_o[23431] = data_o[7];
  assign data_o[23495] = data_o[7];
  assign data_o[23559] = data_o[7];
  assign data_o[23623] = data_o[7];
  assign data_o[23687] = data_o[7];
  assign data_o[23751] = data_o[7];
  assign data_o[23815] = data_o[7];
  assign data_o[23879] = data_o[7];
  assign data_o[23943] = data_o[7];
  assign data_o[24007] = data_o[7];
  assign data_o[24071] = data_o[7];
  assign data_o[24135] = data_o[7];
  assign data_o[24199] = data_o[7];
  assign data_o[24263] = data_o[7];
  assign data_o[24327] = data_o[7];
  assign data_o[24391] = data_o[7];
  assign data_o[24455] = data_o[7];
  assign data_o[24519] = data_o[7];
  assign data_o[24583] = data_o[7];
  assign data_o[24647] = data_o[7];
  assign data_o[24711] = data_o[7];
  assign data_o[24775] = data_o[7];
  assign data_o[24839] = data_o[7];
  assign data_o[24903] = data_o[7];
  assign data_o[24967] = data_o[7];
  assign data_o[25031] = data_o[7];
  assign data_o[25095] = data_o[7];
  assign data_o[25159] = data_o[7];
  assign data_o[25223] = data_o[7];
  assign data_o[25287] = data_o[7];
  assign data_o[25351] = data_o[7];
  assign data_o[25415] = data_o[7];
  assign data_o[25479] = data_o[7];
  assign data_o[25543] = data_o[7];
  assign data_o[25607] = data_o[7];
  assign data_o[25671] = data_o[7];
  assign data_o[25735] = data_o[7];
  assign data_o[25799] = data_o[7];
  assign data_o[25863] = data_o[7];
  assign data_o[25927] = data_o[7];
  assign data_o[25991] = data_o[7];
  assign data_o[26055] = data_o[7];
  assign data_o[26119] = data_o[7];
  assign data_o[26183] = data_o[7];
  assign data_o[26247] = data_o[7];
  assign data_o[26311] = data_o[7];
  assign data_o[26375] = data_o[7];
  assign data_o[26439] = data_o[7];
  assign data_o[26503] = data_o[7];
  assign data_o[26567] = data_o[7];
  assign data_o[26631] = data_o[7];
  assign data_o[26695] = data_o[7];
  assign data_o[26759] = data_o[7];
  assign data_o[26823] = data_o[7];
  assign data_o[26887] = data_o[7];
  assign data_o[26951] = data_o[7];
  assign data_o[27015] = data_o[7];
  assign data_o[27079] = data_o[7];
  assign data_o[27143] = data_o[7];
  assign data_o[27207] = data_o[7];
  assign data_o[27271] = data_o[7];
  assign data_o[27335] = data_o[7];
  assign data_o[27399] = data_o[7];
  assign data_o[27463] = data_o[7];
  assign data_o[27527] = data_o[7];
  assign data_o[27591] = data_o[7];
  assign data_o[27655] = data_o[7];
  assign data_o[27719] = data_o[7];
  assign data_o[27783] = data_o[7];
  assign data_o[27847] = data_o[7];
  assign data_o[27911] = data_o[7];
  assign data_o[27975] = data_o[7];
  assign data_o[28039] = data_o[7];
  assign data_o[28103] = data_o[7];
  assign data_o[28167] = data_o[7];
  assign data_o[28231] = data_o[7];
  assign data_o[28295] = data_o[7];
  assign data_o[28359] = data_o[7];
  assign data_o[28423] = data_o[7];
  assign data_o[28487] = data_o[7];
  assign data_o[28551] = data_o[7];
  assign data_o[28615] = data_o[7];
  assign data_o[28679] = data_o[7];
  assign data_o[28743] = data_o[7];
  assign data_o[28807] = data_o[7];
  assign data_o[28871] = data_o[7];
  assign data_o[28935] = data_o[7];
  assign data_o[28999] = data_o[7];
  assign data_o[29063] = data_o[7];
  assign data_o[29127] = data_o[7];
  assign data_o[29191] = data_o[7];
  assign data_o[29255] = data_o[7];
  assign data_o[29319] = data_o[7];
  assign data_o[29383] = data_o[7];
  assign data_o[29447] = data_o[7];
  assign data_o[29511] = data_o[7];
  assign data_o[29575] = data_o[7];
  assign data_o[29639] = data_o[7];
  assign data_o[29703] = data_o[7];
  assign data_o[29767] = data_o[7];
  assign data_o[29831] = data_o[7];
  assign data_o[29895] = data_o[7];
  assign data_o[29959] = data_o[7];
  assign data_o[30023] = data_o[7];
  assign data_o[30087] = data_o[7];
  assign data_o[30151] = data_o[7];
  assign data_o[30215] = data_o[7];
  assign data_o[30279] = data_o[7];
  assign data_o[30343] = data_o[7];
  assign data_o[30407] = data_o[7];
  assign data_o[30471] = data_o[7];
  assign data_o[30535] = data_o[7];
  assign data_o[30599] = data_o[7];
  assign data_o[30663] = data_o[7];
  assign data_o[30727] = data_o[7];
  assign data_o[30791] = data_o[7];
  assign data_o[30855] = data_o[7];
  assign data_o[30919] = data_o[7];
  assign data_o[30983] = data_o[7];
  assign data_o[31047] = data_o[7];
  assign data_o[31111] = data_o[7];
  assign data_o[31175] = data_o[7];
  assign data_o[31239] = data_o[7];
  assign data_o[31303] = data_o[7];
  assign data_o[31367] = data_o[7];
  assign data_o[31431] = data_o[7];
  assign data_o[31495] = data_o[7];
  assign data_o[31559] = data_o[7];
  assign data_o[31623] = data_o[7];
  assign data_o[31687] = data_o[7];
  assign data_o[31751] = data_o[7];
  assign data_o[31815] = data_o[7];
  assign data_o[31879] = data_o[7];
  assign data_o[31943] = data_o[7];
  assign data_o[70] = data_o[6];
  assign data_o[134] = data_o[6];
  assign data_o[198] = data_o[6];
  assign data_o[262] = data_o[6];
  assign data_o[326] = data_o[6];
  assign data_o[390] = data_o[6];
  assign data_o[454] = data_o[6];
  assign data_o[518] = data_o[6];
  assign data_o[582] = data_o[6];
  assign data_o[646] = data_o[6];
  assign data_o[710] = data_o[6];
  assign data_o[774] = data_o[6];
  assign data_o[838] = data_o[6];
  assign data_o[902] = data_o[6];
  assign data_o[966] = data_o[6];
  assign data_o[1030] = data_o[6];
  assign data_o[1094] = data_o[6];
  assign data_o[1158] = data_o[6];
  assign data_o[1222] = data_o[6];
  assign data_o[1286] = data_o[6];
  assign data_o[1350] = data_o[6];
  assign data_o[1414] = data_o[6];
  assign data_o[1478] = data_o[6];
  assign data_o[1542] = data_o[6];
  assign data_o[1606] = data_o[6];
  assign data_o[1670] = data_o[6];
  assign data_o[1734] = data_o[6];
  assign data_o[1798] = data_o[6];
  assign data_o[1862] = data_o[6];
  assign data_o[1926] = data_o[6];
  assign data_o[1990] = data_o[6];
  assign data_o[2054] = data_o[6];
  assign data_o[2118] = data_o[6];
  assign data_o[2182] = data_o[6];
  assign data_o[2246] = data_o[6];
  assign data_o[2310] = data_o[6];
  assign data_o[2374] = data_o[6];
  assign data_o[2438] = data_o[6];
  assign data_o[2502] = data_o[6];
  assign data_o[2566] = data_o[6];
  assign data_o[2630] = data_o[6];
  assign data_o[2694] = data_o[6];
  assign data_o[2758] = data_o[6];
  assign data_o[2822] = data_o[6];
  assign data_o[2886] = data_o[6];
  assign data_o[2950] = data_o[6];
  assign data_o[3014] = data_o[6];
  assign data_o[3078] = data_o[6];
  assign data_o[3142] = data_o[6];
  assign data_o[3206] = data_o[6];
  assign data_o[3270] = data_o[6];
  assign data_o[3334] = data_o[6];
  assign data_o[3398] = data_o[6];
  assign data_o[3462] = data_o[6];
  assign data_o[3526] = data_o[6];
  assign data_o[3590] = data_o[6];
  assign data_o[3654] = data_o[6];
  assign data_o[3718] = data_o[6];
  assign data_o[3782] = data_o[6];
  assign data_o[3846] = data_o[6];
  assign data_o[3910] = data_o[6];
  assign data_o[3974] = data_o[6];
  assign data_o[4038] = data_o[6];
  assign data_o[4102] = data_o[6];
  assign data_o[4166] = data_o[6];
  assign data_o[4230] = data_o[6];
  assign data_o[4294] = data_o[6];
  assign data_o[4358] = data_o[6];
  assign data_o[4422] = data_o[6];
  assign data_o[4486] = data_o[6];
  assign data_o[4550] = data_o[6];
  assign data_o[4614] = data_o[6];
  assign data_o[4678] = data_o[6];
  assign data_o[4742] = data_o[6];
  assign data_o[4806] = data_o[6];
  assign data_o[4870] = data_o[6];
  assign data_o[4934] = data_o[6];
  assign data_o[4998] = data_o[6];
  assign data_o[5062] = data_o[6];
  assign data_o[5126] = data_o[6];
  assign data_o[5190] = data_o[6];
  assign data_o[5254] = data_o[6];
  assign data_o[5318] = data_o[6];
  assign data_o[5382] = data_o[6];
  assign data_o[5446] = data_o[6];
  assign data_o[5510] = data_o[6];
  assign data_o[5574] = data_o[6];
  assign data_o[5638] = data_o[6];
  assign data_o[5702] = data_o[6];
  assign data_o[5766] = data_o[6];
  assign data_o[5830] = data_o[6];
  assign data_o[5894] = data_o[6];
  assign data_o[5958] = data_o[6];
  assign data_o[6022] = data_o[6];
  assign data_o[6086] = data_o[6];
  assign data_o[6150] = data_o[6];
  assign data_o[6214] = data_o[6];
  assign data_o[6278] = data_o[6];
  assign data_o[6342] = data_o[6];
  assign data_o[6406] = data_o[6];
  assign data_o[6470] = data_o[6];
  assign data_o[6534] = data_o[6];
  assign data_o[6598] = data_o[6];
  assign data_o[6662] = data_o[6];
  assign data_o[6726] = data_o[6];
  assign data_o[6790] = data_o[6];
  assign data_o[6854] = data_o[6];
  assign data_o[6918] = data_o[6];
  assign data_o[6982] = data_o[6];
  assign data_o[7046] = data_o[6];
  assign data_o[7110] = data_o[6];
  assign data_o[7174] = data_o[6];
  assign data_o[7238] = data_o[6];
  assign data_o[7302] = data_o[6];
  assign data_o[7366] = data_o[6];
  assign data_o[7430] = data_o[6];
  assign data_o[7494] = data_o[6];
  assign data_o[7558] = data_o[6];
  assign data_o[7622] = data_o[6];
  assign data_o[7686] = data_o[6];
  assign data_o[7750] = data_o[6];
  assign data_o[7814] = data_o[6];
  assign data_o[7878] = data_o[6];
  assign data_o[7942] = data_o[6];
  assign data_o[8006] = data_o[6];
  assign data_o[8070] = data_o[6];
  assign data_o[8134] = data_o[6];
  assign data_o[8198] = data_o[6];
  assign data_o[8262] = data_o[6];
  assign data_o[8326] = data_o[6];
  assign data_o[8390] = data_o[6];
  assign data_o[8454] = data_o[6];
  assign data_o[8518] = data_o[6];
  assign data_o[8582] = data_o[6];
  assign data_o[8646] = data_o[6];
  assign data_o[8710] = data_o[6];
  assign data_o[8774] = data_o[6];
  assign data_o[8838] = data_o[6];
  assign data_o[8902] = data_o[6];
  assign data_o[8966] = data_o[6];
  assign data_o[9030] = data_o[6];
  assign data_o[9094] = data_o[6];
  assign data_o[9158] = data_o[6];
  assign data_o[9222] = data_o[6];
  assign data_o[9286] = data_o[6];
  assign data_o[9350] = data_o[6];
  assign data_o[9414] = data_o[6];
  assign data_o[9478] = data_o[6];
  assign data_o[9542] = data_o[6];
  assign data_o[9606] = data_o[6];
  assign data_o[9670] = data_o[6];
  assign data_o[9734] = data_o[6];
  assign data_o[9798] = data_o[6];
  assign data_o[9862] = data_o[6];
  assign data_o[9926] = data_o[6];
  assign data_o[9990] = data_o[6];
  assign data_o[10054] = data_o[6];
  assign data_o[10118] = data_o[6];
  assign data_o[10182] = data_o[6];
  assign data_o[10246] = data_o[6];
  assign data_o[10310] = data_o[6];
  assign data_o[10374] = data_o[6];
  assign data_o[10438] = data_o[6];
  assign data_o[10502] = data_o[6];
  assign data_o[10566] = data_o[6];
  assign data_o[10630] = data_o[6];
  assign data_o[10694] = data_o[6];
  assign data_o[10758] = data_o[6];
  assign data_o[10822] = data_o[6];
  assign data_o[10886] = data_o[6];
  assign data_o[10950] = data_o[6];
  assign data_o[11014] = data_o[6];
  assign data_o[11078] = data_o[6];
  assign data_o[11142] = data_o[6];
  assign data_o[11206] = data_o[6];
  assign data_o[11270] = data_o[6];
  assign data_o[11334] = data_o[6];
  assign data_o[11398] = data_o[6];
  assign data_o[11462] = data_o[6];
  assign data_o[11526] = data_o[6];
  assign data_o[11590] = data_o[6];
  assign data_o[11654] = data_o[6];
  assign data_o[11718] = data_o[6];
  assign data_o[11782] = data_o[6];
  assign data_o[11846] = data_o[6];
  assign data_o[11910] = data_o[6];
  assign data_o[11974] = data_o[6];
  assign data_o[12038] = data_o[6];
  assign data_o[12102] = data_o[6];
  assign data_o[12166] = data_o[6];
  assign data_o[12230] = data_o[6];
  assign data_o[12294] = data_o[6];
  assign data_o[12358] = data_o[6];
  assign data_o[12422] = data_o[6];
  assign data_o[12486] = data_o[6];
  assign data_o[12550] = data_o[6];
  assign data_o[12614] = data_o[6];
  assign data_o[12678] = data_o[6];
  assign data_o[12742] = data_o[6];
  assign data_o[12806] = data_o[6];
  assign data_o[12870] = data_o[6];
  assign data_o[12934] = data_o[6];
  assign data_o[12998] = data_o[6];
  assign data_o[13062] = data_o[6];
  assign data_o[13126] = data_o[6];
  assign data_o[13190] = data_o[6];
  assign data_o[13254] = data_o[6];
  assign data_o[13318] = data_o[6];
  assign data_o[13382] = data_o[6];
  assign data_o[13446] = data_o[6];
  assign data_o[13510] = data_o[6];
  assign data_o[13574] = data_o[6];
  assign data_o[13638] = data_o[6];
  assign data_o[13702] = data_o[6];
  assign data_o[13766] = data_o[6];
  assign data_o[13830] = data_o[6];
  assign data_o[13894] = data_o[6];
  assign data_o[13958] = data_o[6];
  assign data_o[14022] = data_o[6];
  assign data_o[14086] = data_o[6];
  assign data_o[14150] = data_o[6];
  assign data_o[14214] = data_o[6];
  assign data_o[14278] = data_o[6];
  assign data_o[14342] = data_o[6];
  assign data_o[14406] = data_o[6];
  assign data_o[14470] = data_o[6];
  assign data_o[14534] = data_o[6];
  assign data_o[14598] = data_o[6];
  assign data_o[14662] = data_o[6];
  assign data_o[14726] = data_o[6];
  assign data_o[14790] = data_o[6];
  assign data_o[14854] = data_o[6];
  assign data_o[14918] = data_o[6];
  assign data_o[14982] = data_o[6];
  assign data_o[15046] = data_o[6];
  assign data_o[15110] = data_o[6];
  assign data_o[15174] = data_o[6];
  assign data_o[15238] = data_o[6];
  assign data_o[15302] = data_o[6];
  assign data_o[15366] = data_o[6];
  assign data_o[15430] = data_o[6];
  assign data_o[15494] = data_o[6];
  assign data_o[15558] = data_o[6];
  assign data_o[15622] = data_o[6];
  assign data_o[15686] = data_o[6];
  assign data_o[15750] = data_o[6];
  assign data_o[15814] = data_o[6];
  assign data_o[15878] = data_o[6];
  assign data_o[15942] = data_o[6];
  assign data_o[16006] = data_o[6];
  assign data_o[16070] = data_o[6];
  assign data_o[16134] = data_o[6];
  assign data_o[16198] = data_o[6];
  assign data_o[16262] = data_o[6];
  assign data_o[16326] = data_o[6];
  assign data_o[16390] = data_o[6];
  assign data_o[16454] = data_o[6];
  assign data_o[16518] = data_o[6];
  assign data_o[16582] = data_o[6];
  assign data_o[16646] = data_o[6];
  assign data_o[16710] = data_o[6];
  assign data_o[16774] = data_o[6];
  assign data_o[16838] = data_o[6];
  assign data_o[16902] = data_o[6];
  assign data_o[16966] = data_o[6];
  assign data_o[17030] = data_o[6];
  assign data_o[17094] = data_o[6];
  assign data_o[17158] = data_o[6];
  assign data_o[17222] = data_o[6];
  assign data_o[17286] = data_o[6];
  assign data_o[17350] = data_o[6];
  assign data_o[17414] = data_o[6];
  assign data_o[17478] = data_o[6];
  assign data_o[17542] = data_o[6];
  assign data_o[17606] = data_o[6];
  assign data_o[17670] = data_o[6];
  assign data_o[17734] = data_o[6];
  assign data_o[17798] = data_o[6];
  assign data_o[17862] = data_o[6];
  assign data_o[17926] = data_o[6];
  assign data_o[17990] = data_o[6];
  assign data_o[18054] = data_o[6];
  assign data_o[18118] = data_o[6];
  assign data_o[18182] = data_o[6];
  assign data_o[18246] = data_o[6];
  assign data_o[18310] = data_o[6];
  assign data_o[18374] = data_o[6];
  assign data_o[18438] = data_o[6];
  assign data_o[18502] = data_o[6];
  assign data_o[18566] = data_o[6];
  assign data_o[18630] = data_o[6];
  assign data_o[18694] = data_o[6];
  assign data_o[18758] = data_o[6];
  assign data_o[18822] = data_o[6];
  assign data_o[18886] = data_o[6];
  assign data_o[18950] = data_o[6];
  assign data_o[19014] = data_o[6];
  assign data_o[19078] = data_o[6];
  assign data_o[19142] = data_o[6];
  assign data_o[19206] = data_o[6];
  assign data_o[19270] = data_o[6];
  assign data_o[19334] = data_o[6];
  assign data_o[19398] = data_o[6];
  assign data_o[19462] = data_o[6];
  assign data_o[19526] = data_o[6];
  assign data_o[19590] = data_o[6];
  assign data_o[19654] = data_o[6];
  assign data_o[19718] = data_o[6];
  assign data_o[19782] = data_o[6];
  assign data_o[19846] = data_o[6];
  assign data_o[19910] = data_o[6];
  assign data_o[19974] = data_o[6];
  assign data_o[20038] = data_o[6];
  assign data_o[20102] = data_o[6];
  assign data_o[20166] = data_o[6];
  assign data_o[20230] = data_o[6];
  assign data_o[20294] = data_o[6];
  assign data_o[20358] = data_o[6];
  assign data_o[20422] = data_o[6];
  assign data_o[20486] = data_o[6];
  assign data_o[20550] = data_o[6];
  assign data_o[20614] = data_o[6];
  assign data_o[20678] = data_o[6];
  assign data_o[20742] = data_o[6];
  assign data_o[20806] = data_o[6];
  assign data_o[20870] = data_o[6];
  assign data_o[20934] = data_o[6];
  assign data_o[20998] = data_o[6];
  assign data_o[21062] = data_o[6];
  assign data_o[21126] = data_o[6];
  assign data_o[21190] = data_o[6];
  assign data_o[21254] = data_o[6];
  assign data_o[21318] = data_o[6];
  assign data_o[21382] = data_o[6];
  assign data_o[21446] = data_o[6];
  assign data_o[21510] = data_o[6];
  assign data_o[21574] = data_o[6];
  assign data_o[21638] = data_o[6];
  assign data_o[21702] = data_o[6];
  assign data_o[21766] = data_o[6];
  assign data_o[21830] = data_o[6];
  assign data_o[21894] = data_o[6];
  assign data_o[21958] = data_o[6];
  assign data_o[22022] = data_o[6];
  assign data_o[22086] = data_o[6];
  assign data_o[22150] = data_o[6];
  assign data_o[22214] = data_o[6];
  assign data_o[22278] = data_o[6];
  assign data_o[22342] = data_o[6];
  assign data_o[22406] = data_o[6];
  assign data_o[22470] = data_o[6];
  assign data_o[22534] = data_o[6];
  assign data_o[22598] = data_o[6];
  assign data_o[22662] = data_o[6];
  assign data_o[22726] = data_o[6];
  assign data_o[22790] = data_o[6];
  assign data_o[22854] = data_o[6];
  assign data_o[22918] = data_o[6];
  assign data_o[22982] = data_o[6];
  assign data_o[23046] = data_o[6];
  assign data_o[23110] = data_o[6];
  assign data_o[23174] = data_o[6];
  assign data_o[23238] = data_o[6];
  assign data_o[23302] = data_o[6];
  assign data_o[23366] = data_o[6];
  assign data_o[23430] = data_o[6];
  assign data_o[23494] = data_o[6];
  assign data_o[23558] = data_o[6];
  assign data_o[23622] = data_o[6];
  assign data_o[23686] = data_o[6];
  assign data_o[23750] = data_o[6];
  assign data_o[23814] = data_o[6];
  assign data_o[23878] = data_o[6];
  assign data_o[23942] = data_o[6];
  assign data_o[24006] = data_o[6];
  assign data_o[24070] = data_o[6];
  assign data_o[24134] = data_o[6];
  assign data_o[24198] = data_o[6];
  assign data_o[24262] = data_o[6];
  assign data_o[24326] = data_o[6];
  assign data_o[24390] = data_o[6];
  assign data_o[24454] = data_o[6];
  assign data_o[24518] = data_o[6];
  assign data_o[24582] = data_o[6];
  assign data_o[24646] = data_o[6];
  assign data_o[24710] = data_o[6];
  assign data_o[24774] = data_o[6];
  assign data_o[24838] = data_o[6];
  assign data_o[24902] = data_o[6];
  assign data_o[24966] = data_o[6];
  assign data_o[25030] = data_o[6];
  assign data_o[25094] = data_o[6];
  assign data_o[25158] = data_o[6];
  assign data_o[25222] = data_o[6];
  assign data_o[25286] = data_o[6];
  assign data_o[25350] = data_o[6];
  assign data_o[25414] = data_o[6];
  assign data_o[25478] = data_o[6];
  assign data_o[25542] = data_o[6];
  assign data_o[25606] = data_o[6];
  assign data_o[25670] = data_o[6];
  assign data_o[25734] = data_o[6];
  assign data_o[25798] = data_o[6];
  assign data_o[25862] = data_o[6];
  assign data_o[25926] = data_o[6];
  assign data_o[25990] = data_o[6];
  assign data_o[26054] = data_o[6];
  assign data_o[26118] = data_o[6];
  assign data_o[26182] = data_o[6];
  assign data_o[26246] = data_o[6];
  assign data_o[26310] = data_o[6];
  assign data_o[26374] = data_o[6];
  assign data_o[26438] = data_o[6];
  assign data_o[26502] = data_o[6];
  assign data_o[26566] = data_o[6];
  assign data_o[26630] = data_o[6];
  assign data_o[26694] = data_o[6];
  assign data_o[26758] = data_o[6];
  assign data_o[26822] = data_o[6];
  assign data_o[26886] = data_o[6];
  assign data_o[26950] = data_o[6];
  assign data_o[27014] = data_o[6];
  assign data_o[27078] = data_o[6];
  assign data_o[27142] = data_o[6];
  assign data_o[27206] = data_o[6];
  assign data_o[27270] = data_o[6];
  assign data_o[27334] = data_o[6];
  assign data_o[27398] = data_o[6];
  assign data_o[27462] = data_o[6];
  assign data_o[27526] = data_o[6];
  assign data_o[27590] = data_o[6];
  assign data_o[27654] = data_o[6];
  assign data_o[27718] = data_o[6];
  assign data_o[27782] = data_o[6];
  assign data_o[27846] = data_o[6];
  assign data_o[27910] = data_o[6];
  assign data_o[27974] = data_o[6];
  assign data_o[28038] = data_o[6];
  assign data_o[28102] = data_o[6];
  assign data_o[28166] = data_o[6];
  assign data_o[28230] = data_o[6];
  assign data_o[28294] = data_o[6];
  assign data_o[28358] = data_o[6];
  assign data_o[28422] = data_o[6];
  assign data_o[28486] = data_o[6];
  assign data_o[28550] = data_o[6];
  assign data_o[28614] = data_o[6];
  assign data_o[28678] = data_o[6];
  assign data_o[28742] = data_o[6];
  assign data_o[28806] = data_o[6];
  assign data_o[28870] = data_o[6];
  assign data_o[28934] = data_o[6];
  assign data_o[28998] = data_o[6];
  assign data_o[29062] = data_o[6];
  assign data_o[29126] = data_o[6];
  assign data_o[29190] = data_o[6];
  assign data_o[29254] = data_o[6];
  assign data_o[29318] = data_o[6];
  assign data_o[29382] = data_o[6];
  assign data_o[29446] = data_o[6];
  assign data_o[29510] = data_o[6];
  assign data_o[29574] = data_o[6];
  assign data_o[29638] = data_o[6];
  assign data_o[29702] = data_o[6];
  assign data_o[29766] = data_o[6];
  assign data_o[29830] = data_o[6];
  assign data_o[29894] = data_o[6];
  assign data_o[29958] = data_o[6];
  assign data_o[30022] = data_o[6];
  assign data_o[30086] = data_o[6];
  assign data_o[30150] = data_o[6];
  assign data_o[30214] = data_o[6];
  assign data_o[30278] = data_o[6];
  assign data_o[30342] = data_o[6];
  assign data_o[30406] = data_o[6];
  assign data_o[30470] = data_o[6];
  assign data_o[30534] = data_o[6];
  assign data_o[30598] = data_o[6];
  assign data_o[30662] = data_o[6];
  assign data_o[30726] = data_o[6];
  assign data_o[30790] = data_o[6];
  assign data_o[30854] = data_o[6];
  assign data_o[30918] = data_o[6];
  assign data_o[30982] = data_o[6];
  assign data_o[31046] = data_o[6];
  assign data_o[31110] = data_o[6];
  assign data_o[31174] = data_o[6];
  assign data_o[31238] = data_o[6];
  assign data_o[31302] = data_o[6];
  assign data_o[31366] = data_o[6];
  assign data_o[31430] = data_o[6];
  assign data_o[31494] = data_o[6];
  assign data_o[31558] = data_o[6];
  assign data_o[31622] = data_o[6];
  assign data_o[31686] = data_o[6];
  assign data_o[31750] = data_o[6];
  assign data_o[31814] = data_o[6];
  assign data_o[31878] = data_o[6];
  assign data_o[31942] = data_o[6];
  assign data_o[69] = data_o[5];
  assign data_o[133] = data_o[5];
  assign data_o[197] = data_o[5];
  assign data_o[261] = data_o[5];
  assign data_o[325] = data_o[5];
  assign data_o[389] = data_o[5];
  assign data_o[453] = data_o[5];
  assign data_o[517] = data_o[5];
  assign data_o[581] = data_o[5];
  assign data_o[645] = data_o[5];
  assign data_o[709] = data_o[5];
  assign data_o[773] = data_o[5];
  assign data_o[837] = data_o[5];
  assign data_o[901] = data_o[5];
  assign data_o[965] = data_o[5];
  assign data_o[1029] = data_o[5];
  assign data_o[1093] = data_o[5];
  assign data_o[1157] = data_o[5];
  assign data_o[1221] = data_o[5];
  assign data_o[1285] = data_o[5];
  assign data_o[1349] = data_o[5];
  assign data_o[1413] = data_o[5];
  assign data_o[1477] = data_o[5];
  assign data_o[1541] = data_o[5];
  assign data_o[1605] = data_o[5];
  assign data_o[1669] = data_o[5];
  assign data_o[1733] = data_o[5];
  assign data_o[1797] = data_o[5];
  assign data_o[1861] = data_o[5];
  assign data_o[1925] = data_o[5];
  assign data_o[1989] = data_o[5];
  assign data_o[2053] = data_o[5];
  assign data_o[2117] = data_o[5];
  assign data_o[2181] = data_o[5];
  assign data_o[2245] = data_o[5];
  assign data_o[2309] = data_o[5];
  assign data_o[2373] = data_o[5];
  assign data_o[2437] = data_o[5];
  assign data_o[2501] = data_o[5];
  assign data_o[2565] = data_o[5];
  assign data_o[2629] = data_o[5];
  assign data_o[2693] = data_o[5];
  assign data_o[2757] = data_o[5];
  assign data_o[2821] = data_o[5];
  assign data_o[2885] = data_o[5];
  assign data_o[2949] = data_o[5];
  assign data_o[3013] = data_o[5];
  assign data_o[3077] = data_o[5];
  assign data_o[3141] = data_o[5];
  assign data_o[3205] = data_o[5];
  assign data_o[3269] = data_o[5];
  assign data_o[3333] = data_o[5];
  assign data_o[3397] = data_o[5];
  assign data_o[3461] = data_o[5];
  assign data_o[3525] = data_o[5];
  assign data_o[3589] = data_o[5];
  assign data_o[3653] = data_o[5];
  assign data_o[3717] = data_o[5];
  assign data_o[3781] = data_o[5];
  assign data_o[3845] = data_o[5];
  assign data_o[3909] = data_o[5];
  assign data_o[3973] = data_o[5];
  assign data_o[4037] = data_o[5];
  assign data_o[4101] = data_o[5];
  assign data_o[4165] = data_o[5];
  assign data_o[4229] = data_o[5];
  assign data_o[4293] = data_o[5];
  assign data_o[4357] = data_o[5];
  assign data_o[4421] = data_o[5];
  assign data_o[4485] = data_o[5];
  assign data_o[4549] = data_o[5];
  assign data_o[4613] = data_o[5];
  assign data_o[4677] = data_o[5];
  assign data_o[4741] = data_o[5];
  assign data_o[4805] = data_o[5];
  assign data_o[4869] = data_o[5];
  assign data_o[4933] = data_o[5];
  assign data_o[4997] = data_o[5];
  assign data_o[5061] = data_o[5];
  assign data_o[5125] = data_o[5];
  assign data_o[5189] = data_o[5];
  assign data_o[5253] = data_o[5];
  assign data_o[5317] = data_o[5];
  assign data_o[5381] = data_o[5];
  assign data_o[5445] = data_o[5];
  assign data_o[5509] = data_o[5];
  assign data_o[5573] = data_o[5];
  assign data_o[5637] = data_o[5];
  assign data_o[5701] = data_o[5];
  assign data_o[5765] = data_o[5];
  assign data_o[5829] = data_o[5];
  assign data_o[5893] = data_o[5];
  assign data_o[5957] = data_o[5];
  assign data_o[6021] = data_o[5];
  assign data_o[6085] = data_o[5];
  assign data_o[6149] = data_o[5];
  assign data_o[6213] = data_o[5];
  assign data_o[6277] = data_o[5];
  assign data_o[6341] = data_o[5];
  assign data_o[6405] = data_o[5];
  assign data_o[6469] = data_o[5];
  assign data_o[6533] = data_o[5];
  assign data_o[6597] = data_o[5];
  assign data_o[6661] = data_o[5];
  assign data_o[6725] = data_o[5];
  assign data_o[6789] = data_o[5];
  assign data_o[6853] = data_o[5];
  assign data_o[6917] = data_o[5];
  assign data_o[6981] = data_o[5];
  assign data_o[7045] = data_o[5];
  assign data_o[7109] = data_o[5];
  assign data_o[7173] = data_o[5];
  assign data_o[7237] = data_o[5];
  assign data_o[7301] = data_o[5];
  assign data_o[7365] = data_o[5];
  assign data_o[7429] = data_o[5];
  assign data_o[7493] = data_o[5];
  assign data_o[7557] = data_o[5];
  assign data_o[7621] = data_o[5];
  assign data_o[7685] = data_o[5];
  assign data_o[7749] = data_o[5];
  assign data_o[7813] = data_o[5];
  assign data_o[7877] = data_o[5];
  assign data_o[7941] = data_o[5];
  assign data_o[8005] = data_o[5];
  assign data_o[8069] = data_o[5];
  assign data_o[8133] = data_o[5];
  assign data_o[8197] = data_o[5];
  assign data_o[8261] = data_o[5];
  assign data_o[8325] = data_o[5];
  assign data_o[8389] = data_o[5];
  assign data_o[8453] = data_o[5];
  assign data_o[8517] = data_o[5];
  assign data_o[8581] = data_o[5];
  assign data_o[8645] = data_o[5];
  assign data_o[8709] = data_o[5];
  assign data_o[8773] = data_o[5];
  assign data_o[8837] = data_o[5];
  assign data_o[8901] = data_o[5];
  assign data_o[8965] = data_o[5];
  assign data_o[9029] = data_o[5];
  assign data_o[9093] = data_o[5];
  assign data_o[9157] = data_o[5];
  assign data_o[9221] = data_o[5];
  assign data_o[9285] = data_o[5];
  assign data_o[9349] = data_o[5];
  assign data_o[9413] = data_o[5];
  assign data_o[9477] = data_o[5];
  assign data_o[9541] = data_o[5];
  assign data_o[9605] = data_o[5];
  assign data_o[9669] = data_o[5];
  assign data_o[9733] = data_o[5];
  assign data_o[9797] = data_o[5];
  assign data_o[9861] = data_o[5];
  assign data_o[9925] = data_o[5];
  assign data_o[9989] = data_o[5];
  assign data_o[10053] = data_o[5];
  assign data_o[10117] = data_o[5];
  assign data_o[10181] = data_o[5];
  assign data_o[10245] = data_o[5];
  assign data_o[10309] = data_o[5];
  assign data_o[10373] = data_o[5];
  assign data_o[10437] = data_o[5];
  assign data_o[10501] = data_o[5];
  assign data_o[10565] = data_o[5];
  assign data_o[10629] = data_o[5];
  assign data_o[10693] = data_o[5];
  assign data_o[10757] = data_o[5];
  assign data_o[10821] = data_o[5];
  assign data_o[10885] = data_o[5];
  assign data_o[10949] = data_o[5];
  assign data_o[11013] = data_o[5];
  assign data_o[11077] = data_o[5];
  assign data_o[11141] = data_o[5];
  assign data_o[11205] = data_o[5];
  assign data_o[11269] = data_o[5];
  assign data_o[11333] = data_o[5];
  assign data_o[11397] = data_o[5];
  assign data_o[11461] = data_o[5];
  assign data_o[11525] = data_o[5];
  assign data_o[11589] = data_o[5];
  assign data_o[11653] = data_o[5];
  assign data_o[11717] = data_o[5];
  assign data_o[11781] = data_o[5];
  assign data_o[11845] = data_o[5];
  assign data_o[11909] = data_o[5];
  assign data_o[11973] = data_o[5];
  assign data_o[12037] = data_o[5];
  assign data_o[12101] = data_o[5];
  assign data_o[12165] = data_o[5];
  assign data_o[12229] = data_o[5];
  assign data_o[12293] = data_o[5];
  assign data_o[12357] = data_o[5];
  assign data_o[12421] = data_o[5];
  assign data_o[12485] = data_o[5];
  assign data_o[12549] = data_o[5];
  assign data_o[12613] = data_o[5];
  assign data_o[12677] = data_o[5];
  assign data_o[12741] = data_o[5];
  assign data_o[12805] = data_o[5];
  assign data_o[12869] = data_o[5];
  assign data_o[12933] = data_o[5];
  assign data_o[12997] = data_o[5];
  assign data_o[13061] = data_o[5];
  assign data_o[13125] = data_o[5];
  assign data_o[13189] = data_o[5];
  assign data_o[13253] = data_o[5];
  assign data_o[13317] = data_o[5];
  assign data_o[13381] = data_o[5];
  assign data_o[13445] = data_o[5];
  assign data_o[13509] = data_o[5];
  assign data_o[13573] = data_o[5];
  assign data_o[13637] = data_o[5];
  assign data_o[13701] = data_o[5];
  assign data_o[13765] = data_o[5];
  assign data_o[13829] = data_o[5];
  assign data_o[13893] = data_o[5];
  assign data_o[13957] = data_o[5];
  assign data_o[14021] = data_o[5];
  assign data_o[14085] = data_o[5];
  assign data_o[14149] = data_o[5];
  assign data_o[14213] = data_o[5];
  assign data_o[14277] = data_o[5];
  assign data_o[14341] = data_o[5];
  assign data_o[14405] = data_o[5];
  assign data_o[14469] = data_o[5];
  assign data_o[14533] = data_o[5];
  assign data_o[14597] = data_o[5];
  assign data_o[14661] = data_o[5];
  assign data_o[14725] = data_o[5];
  assign data_o[14789] = data_o[5];
  assign data_o[14853] = data_o[5];
  assign data_o[14917] = data_o[5];
  assign data_o[14981] = data_o[5];
  assign data_o[15045] = data_o[5];
  assign data_o[15109] = data_o[5];
  assign data_o[15173] = data_o[5];
  assign data_o[15237] = data_o[5];
  assign data_o[15301] = data_o[5];
  assign data_o[15365] = data_o[5];
  assign data_o[15429] = data_o[5];
  assign data_o[15493] = data_o[5];
  assign data_o[15557] = data_o[5];
  assign data_o[15621] = data_o[5];
  assign data_o[15685] = data_o[5];
  assign data_o[15749] = data_o[5];
  assign data_o[15813] = data_o[5];
  assign data_o[15877] = data_o[5];
  assign data_o[15941] = data_o[5];
  assign data_o[16005] = data_o[5];
  assign data_o[16069] = data_o[5];
  assign data_o[16133] = data_o[5];
  assign data_o[16197] = data_o[5];
  assign data_o[16261] = data_o[5];
  assign data_o[16325] = data_o[5];
  assign data_o[16389] = data_o[5];
  assign data_o[16453] = data_o[5];
  assign data_o[16517] = data_o[5];
  assign data_o[16581] = data_o[5];
  assign data_o[16645] = data_o[5];
  assign data_o[16709] = data_o[5];
  assign data_o[16773] = data_o[5];
  assign data_o[16837] = data_o[5];
  assign data_o[16901] = data_o[5];
  assign data_o[16965] = data_o[5];
  assign data_o[17029] = data_o[5];
  assign data_o[17093] = data_o[5];
  assign data_o[17157] = data_o[5];
  assign data_o[17221] = data_o[5];
  assign data_o[17285] = data_o[5];
  assign data_o[17349] = data_o[5];
  assign data_o[17413] = data_o[5];
  assign data_o[17477] = data_o[5];
  assign data_o[17541] = data_o[5];
  assign data_o[17605] = data_o[5];
  assign data_o[17669] = data_o[5];
  assign data_o[17733] = data_o[5];
  assign data_o[17797] = data_o[5];
  assign data_o[17861] = data_o[5];
  assign data_o[17925] = data_o[5];
  assign data_o[17989] = data_o[5];
  assign data_o[18053] = data_o[5];
  assign data_o[18117] = data_o[5];
  assign data_o[18181] = data_o[5];
  assign data_o[18245] = data_o[5];
  assign data_o[18309] = data_o[5];
  assign data_o[18373] = data_o[5];
  assign data_o[18437] = data_o[5];
  assign data_o[18501] = data_o[5];
  assign data_o[18565] = data_o[5];
  assign data_o[18629] = data_o[5];
  assign data_o[18693] = data_o[5];
  assign data_o[18757] = data_o[5];
  assign data_o[18821] = data_o[5];
  assign data_o[18885] = data_o[5];
  assign data_o[18949] = data_o[5];
  assign data_o[19013] = data_o[5];
  assign data_o[19077] = data_o[5];
  assign data_o[19141] = data_o[5];
  assign data_o[19205] = data_o[5];
  assign data_o[19269] = data_o[5];
  assign data_o[19333] = data_o[5];
  assign data_o[19397] = data_o[5];
  assign data_o[19461] = data_o[5];
  assign data_o[19525] = data_o[5];
  assign data_o[19589] = data_o[5];
  assign data_o[19653] = data_o[5];
  assign data_o[19717] = data_o[5];
  assign data_o[19781] = data_o[5];
  assign data_o[19845] = data_o[5];
  assign data_o[19909] = data_o[5];
  assign data_o[19973] = data_o[5];
  assign data_o[20037] = data_o[5];
  assign data_o[20101] = data_o[5];
  assign data_o[20165] = data_o[5];
  assign data_o[20229] = data_o[5];
  assign data_o[20293] = data_o[5];
  assign data_o[20357] = data_o[5];
  assign data_o[20421] = data_o[5];
  assign data_o[20485] = data_o[5];
  assign data_o[20549] = data_o[5];
  assign data_o[20613] = data_o[5];
  assign data_o[20677] = data_o[5];
  assign data_o[20741] = data_o[5];
  assign data_o[20805] = data_o[5];
  assign data_o[20869] = data_o[5];
  assign data_o[20933] = data_o[5];
  assign data_o[20997] = data_o[5];
  assign data_o[21061] = data_o[5];
  assign data_o[21125] = data_o[5];
  assign data_o[21189] = data_o[5];
  assign data_o[21253] = data_o[5];
  assign data_o[21317] = data_o[5];
  assign data_o[21381] = data_o[5];
  assign data_o[21445] = data_o[5];
  assign data_o[21509] = data_o[5];
  assign data_o[21573] = data_o[5];
  assign data_o[21637] = data_o[5];
  assign data_o[21701] = data_o[5];
  assign data_o[21765] = data_o[5];
  assign data_o[21829] = data_o[5];
  assign data_o[21893] = data_o[5];
  assign data_o[21957] = data_o[5];
  assign data_o[22021] = data_o[5];
  assign data_o[22085] = data_o[5];
  assign data_o[22149] = data_o[5];
  assign data_o[22213] = data_o[5];
  assign data_o[22277] = data_o[5];
  assign data_o[22341] = data_o[5];
  assign data_o[22405] = data_o[5];
  assign data_o[22469] = data_o[5];
  assign data_o[22533] = data_o[5];
  assign data_o[22597] = data_o[5];
  assign data_o[22661] = data_o[5];
  assign data_o[22725] = data_o[5];
  assign data_o[22789] = data_o[5];
  assign data_o[22853] = data_o[5];
  assign data_o[22917] = data_o[5];
  assign data_o[22981] = data_o[5];
  assign data_o[23045] = data_o[5];
  assign data_o[23109] = data_o[5];
  assign data_o[23173] = data_o[5];
  assign data_o[23237] = data_o[5];
  assign data_o[23301] = data_o[5];
  assign data_o[23365] = data_o[5];
  assign data_o[23429] = data_o[5];
  assign data_o[23493] = data_o[5];
  assign data_o[23557] = data_o[5];
  assign data_o[23621] = data_o[5];
  assign data_o[23685] = data_o[5];
  assign data_o[23749] = data_o[5];
  assign data_o[23813] = data_o[5];
  assign data_o[23877] = data_o[5];
  assign data_o[23941] = data_o[5];
  assign data_o[24005] = data_o[5];
  assign data_o[24069] = data_o[5];
  assign data_o[24133] = data_o[5];
  assign data_o[24197] = data_o[5];
  assign data_o[24261] = data_o[5];
  assign data_o[24325] = data_o[5];
  assign data_o[24389] = data_o[5];
  assign data_o[24453] = data_o[5];
  assign data_o[24517] = data_o[5];
  assign data_o[24581] = data_o[5];
  assign data_o[24645] = data_o[5];
  assign data_o[24709] = data_o[5];
  assign data_o[24773] = data_o[5];
  assign data_o[24837] = data_o[5];
  assign data_o[24901] = data_o[5];
  assign data_o[24965] = data_o[5];
  assign data_o[25029] = data_o[5];
  assign data_o[25093] = data_o[5];
  assign data_o[25157] = data_o[5];
  assign data_o[25221] = data_o[5];
  assign data_o[25285] = data_o[5];
  assign data_o[25349] = data_o[5];
  assign data_o[25413] = data_o[5];
  assign data_o[25477] = data_o[5];
  assign data_o[25541] = data_o[5];
  assign data_o[25605] = data_o[5];
  assign data_o[25669] = data_o[5];
  assign data_o[25733] = data_o[5];
  assign data_o[25797] = data_o[5];
  assign data_o[25861] = data_o[5];
  assign data_o[25925] = data_o[5];
  assign data_o[25989] = data_o[5];
  assign data_o[26053] = data_o[5];
  assign data_o[26117] = data_o[5];
  assign data_o[26181] = data_o[5];
  assign data_o[26245] = data_o[5];
  assign data_o[26309] = data_o[5];
  assign data_o[26373] = data_o[5];
  assign data_o[26437] = data_o[5];
  assign data_o[26501] = data_o[5];
  assign data_o[26565] = data_o[5];
  assign data_o[26629] = data_o[5];
  assign data_o[26693] = data_o[5];
  assign data_o[26757] = data_o[5];
  assign data_o[26821] = data_o[5];
  assign data_o[26885] = data_o[5];
  assign data_o[26949] = data_o[5];
  assign data_o[27013] = data_o[5];
  assign data_o[27077] = data_o[5];
  assign data_o[27141] = data_o[5];
  assign data_o[27205] = data_o[5];
  assign data_o[27269] = data_o[5];
  assign data_o[27333] = data_o[5];
  assign data_o[27397] = data_o[5];
  assign data_o[27461] = data_o[5];
  assign data_o[27525] = data_o[5];
  assign data_o[27589] = data_o[5];
  assign data_o[27653] = data_o[5];
  assign data_o[27717] = data_o[5];
  assign data_o[27781] = data_o[5];
  assign data_o[27845] = data_o[5];
  assign data_o[27909] = data_o[5];
  assign data_o[27973] = data_o[5];
  assign data_o[28037] = data_o[5];
  assign data_o[28101] = data_o[5];
  assign data_o[28165] = data_o[5];
  assign data_o[28229] = data_o[5];
  assign data_o[28293] = data_o[5];
  assign data_o[28357] = data_o[5];
  assign data_o[28421] = data_o[5];
  assign data_o[28485] = data_o[5];
  assign data_o[28549] = data_o[5];
  assign data_o[28613] = data_o[5];
  assign data_o[28677] = data_o[5];
  assign data_o[28741] = data_o[5];
  assign data_o[28805] = data_o[5];
  assign data_o[28869] = data_o[5];
  assign data_o[28933] = data_o[5];
  assign data_o[28997] = data_o[5];
  assign data_o[29061] = data_o[5];
  assign data_o[29125] = data_o[5];
  assign data_o[29189] = data_o[5];
  assign data_o[29253] = data_o[5];
  assign data_o[29317] = data_o[5];
  assign data_o[29381] = data_o[5];
  assign data_o[29445] = data_o[5];
  assign data_o[29509] = data_o[5];
  assign data_o[29573] = data_o[5];
  assign data_o[29637] = data_o[5];
  assign data_o[29701] = data_o[5];
  assign data_o[29765] = data_o[5];
  assign data_o[29829] = data_o[5];
  assign data_o[29893] = data_o[5];
  assign data_o[29957] = data_o[5];
  assign data_o[30021] = data_o[5];
  assign data_o[30085] = data_o[5];
  assign data_o[30149] = data_o[5];
  assign data_o[30213] = data_o[5];
  assign data_o[30277] = data_o[5];
  assign data_o[30341] = data_o[5];
  assign data_o[30405] = data_o[5];
  assign data_o[30469] = data_o[5];
  assign data_o[30533] = data_o[5];
  assign data_o[30597] = data_o[5];
  assign data_o[30661] = data_o[5];
  assign data_o[30725] = data_o[5];
  assign data_o[30789] = data_o[5];
  assign data_o[30853] = data_o[5];
  assign data_o[30917] = data_o[5];
  assign data_o[30981] = data_o[5];
  assign data_o[31045] = data_o[5];
  assign data_o[31109] = data_o[5];
  assign data_o[31173] = data_o[5];
  assign data_o[31237] = data_o[5];
  assign data_o[31301] = data_o[5];
  assign data_o[31365] = data_o[5];
  assign data_o[31429] = data_o[5];
  assign data_o[31493] = data_o[5];
  assign data_o[31557] = data_o[5];
  assign data_o[31621] = data_o[5];
  assign data_o[31685] = data_o[5];
  assign data_o[31749] = data_o[5];
  assign data_o[31813] = data_o[5];
  assign data_o[31877] = data_o[5];
  assign data_o[31941] = data_o[5];
  assign data_o[68] = data_o[4];
  assign data_o[132] = data_o[4];
  assign data_o[196] = data_o[4];
  assign data_o[260] = data_o[4];
  assign data_o[324] = data_o[4];
  assign data_o[388] = data_o[4];
  assign data_o[452] = data_o[4];
  assign data_o[516] = data_o[4];
  assign data_o[580] = data_o[4];
  assign data_o[644] = data_o[4];
  assign data_o[708] = data_o[4];
  assign data_o[772] = data_o[4];
  assign data_o[836] = data_o[4];
  assign data_o[900] = data_o[4];
  assign data_o[964] = data_o[4];
  assign data_o[1028] = data_o[4];
  assign data_o[1092] = data_o[4];
  assign data_o[1156] = data_o[4];
  assign data_o[1220] = data_o[4];
  assign data_o[1284] = data_o[4];
  assign data_o[1348] = data_o[4];
  assign data_o[1412] = data_o[4];
  assign data_o[1476] = data_o[4];
  assign data_o[1540] = data_o[4];
  assign data_o[1604] = data_o[4];
  assign data_o[1668] = data_o[4];
  assign data_o[1732] = data_o[4];
  assign data_o[1796] = data_o[4];
  assign data_o[1860] = data_o[4];
  assign data_o[1924] = data_o[4];
  assign data_o[1988] = data_o[4];
  assign data_o[2052] = data_o[4];
  assign data_o[2116] = data_o[4];
  assign data_o[2180] = data_o[4];
  assign data_o[2244] = data_o[4];
  assign data_o[2308] = data_o[4];
  assign data_o[2372] = data_o[4];
  assign data_o[2436] = data_o[4];
  assign data_o[2500] = data_o[4];
  assign data_o[2564] = data_o[4];
  assign data_o[2628] = data_o[4];
  assign data_o[2692] = data_o[4];
  assign data_o[2756] = data_o[4];
  assign data_o[2820] = data_o[4];
  assign data_o[2884] = data_o[4];
  assign data_o[2948] = data_o[4];
  assign data_o[3012] = data_o[4];
  assign data_o[3076] = data_o[4];
  assign data_o[3140] = data_o[4];
  assign data_o[3204] = data_o[4];
  assign data_o[3268] = data_o[4];
  assign data_o[3332] = data_o[4];
  assign data_o[3396] = data_o[4];
  assign data_o[3460] = data_o[4];
  assign data_o[3524] = data_o[4];
  assign data_o[3588] = data_o[4];
  assign data_o[3652] = data_o[4];
  assign data_o[3716] = data_o[4];
  assign data_o[3780] = data_o[4];
  assign data_o[3844] = data_o[4];
  assign data_o[3908] = data_o[4];
  assign data_o[3972] = data_o[4];
  assign data_o[4036] = data_o[4];
  assign data_o[4100] = data_o[4];
  assign data_o[4164] = data_o[4];
  assign data_o[4228] = data_o[4];
  assign data_o[4292] = data_o[4];
  assign data_o[4356] = data_o[4];
  assign data_o[4420] = data_o[4];
  assign data_o[4484] = data_o[4];
  assign data_o[4548] = data_o[4];
  assign data_o[4612] = data_o[4];
  assign data_o[4676] = data_o[4];
  assign data_o[4740] = data_o[4];
  assign data_o[4804] = data_o[4];
  assign data_o[4868] = data_o[4];
  assign data_o[4932] = data_o[4];
  assign data_o[4996] = data_o[4];
  assign data_o[5060] = data_o[4];
  assign data_o[5124] = data_o[4];
  assign data_o[5188] = data_o[4];
  assign data_o[5252] = data_o[4];
  assign data_o[5316] = data_o[4];
  assign data_o[5380] = data_o[4];
  assign data_o[5444] = data_o[4];
  assign data_o[5508] = data_o[4];
  assign data_o[5572] = data_o[4];
  assign data_o[5636] = data_o[4];
  assign data_o[5700] = data_o[4];
  assign data_o[5764] = data_o[4];
  assign data_o[5828] = data_o[4];
  assign data_o[5892] = data_o[4];
  assign data_o[5956] = data_o[4];
  assign data_o[6020] = data_o[4];
  assign data_o[6084] = data_o[4];
  assign data_o[6148] = data_o[4];
  assign data_o[6212] = data_o[4];
  assign data_o[6276] = data_o[4];
  assign data_o[6340] = data_o[4];
  assign data_o[6404] = data_o[4];
  assign data_o[6468] = data_o[4];
  assign data_o[6532] = data_o[4];
  assign data_o[6596] = data_o[4];
  assign data_o[6660] = data_o[4];
  assign data_o[6724] = data_o[4];
  assign data_o[6788] = data_o[4];
  assign data_o[6852] = data_o[4];
  assign data_o[6916] = data_o[4];
  assign data_o[6980] = data_o[4];
  assign data_o[7044] = data_o[4];
  assign data_o[7108] = data_o[4];
  assign data_o[7172] = data_o[4];
  assign data_o[7236] = data_o[4];
  assign data_o[7300] = data_o[4];
  assign data_o[7364] = data_o[4];
  assign data_o[7428] = data_o[4];
  assign data_o[7492] = data_o[4];
  assign data_o[7556] = data_o[4];
  assign data_o[7620] = data_o[4];
  assign data_o[7684] = data_o[4];
  assign data_o[7748] = data_o[4];
  assign data_o[7812] = data_o[4];
  assign data_o[7876] = data_o[4];
  assign data_o[7940] = data_o[4];
  assign data_o[8004] = data_o[4];
  assign data_o[8068] = data_o[4];
  assign data_o[8132] = data_o[4];
  assign data_o[8196] = data_o[4];
  assign data_o[8260] = data_o[4];
  assign data_o[8324] = data_o[4];
  assign data_o[8388] = data_o[4];
  assign data_o[8452] = data_o[4];
  assign data_o[8516] = data_o[4];
  assign data_o[8580] = data_o[4];
  assign data_o[8644] = data_o[4];
  assign data_o[8708] = data_o[4];
  assign data_o[8772] = data_o[4];
  assign data_o[8836] = data_o[4];
  assign data_o[8900] = data_o[4];
  assign data_o[8964] = data_o[4];
  assign data_o[9028] = data_o[4];
  assign data_o[9092] = data_o[4];
  assign data_o[9156] = data_o[4];
  assign data_o[9220] = data_o[4];
  assign data_o[9284] = data_o[4];
  assign data_o[9348] = data_o[4];
  assign data_o[9412] = data_o[4];
  assign data_o[9476] = data_o[4];
  assign data_o[9540] = data_o[4];
  assign data_o[9604] = data_o[4];
  assign data_o[9668] = data_o[4];
  assign data_o[9732] = data_o[4];
  assign data_o[9796] = data_o[4];
  assign data_o[9860] = data_o[4];
  assign data_o[9924] = data_o[4];
  assign data_o[9988] = data_o[4];
  assign data_o[10052] = data_o[4];
  assign data_o[10116] = data_o[4];
  assign data_o[10180] = data_o[4];
  assign data_o[10244] = data_o[4];
  assign data_o[10308] = data_o[4];
  assign data_o[10372] = data_o[4];
  assign data_o[10436] = data_o[4];
  assign data_o[10500] = data_o[4];
  assign data_o[10564] = data_o[4];
  assign data_o[10628] = data_o[4];
  assign data_o[10692] = data_o[4];
  assign data_o[10756] = data_o[4];
  assign data_o[10820] = data_o[4];
  assign data_o[10884] = data_o[4];
  assign data_o[10948] = data_o[4];
  assign data_o[11012] = data_o[4];
  assign data_o[11076] = data_o[4];
  assign data_o[11140] = data_o[4];
  assign data_o[11204] = data_o[4];
  assign data_o[11268] = data_o[4];
  assign data_o[11332] = data_o[4];
  assign data_o[11396] = data_o[4];
  assign data_o[11460] = data_o[4];
  assign data_o[11524] = data_o[4];
  assign data_o[11588] = data_o[4];
  assign data_o[11652] = data_o[4];
  assign data_o[11716] = data_o[4];
  assign data_o[11780] = data_o[4];
  assign data_o[11844] = data_o[4];
  assign data_o[11908] = data_o[4];
  assign data_o[11972] = data_o[4];
  assign data_o[12036] = data_o[4];
  assign data_o[12100] = data_o[4];
  assign data_o[12164] = data_o[4];
  assign data_o[12228] = data_o[4];
  assign data_o[12292] = data_o[4];
  assign data_o[12356] = data_o[4];
  assign data_o[12420] = data_o[4];
  assign data_o[12484] = data_o[4];
  assign data_o[12548] = data_o[4];
  assign data_o[12612] = data_o[4];
  assign data_o[12676] = data_o[4];
  assign data_o[12740] = data_o[4];
  assign data_o[12804] = data_o[4];
  assign data_o[12868] = data_o[4];
  assign data_o[12932] = data_o[4];
  assign data_o[12996] = data_o[4];
  assign data_o[13060] = data_o[4];
  assign data_o[13124] = data_o[4];
  assign data_o[13188] = data_o[4];
  assign data_o[13252] = data_o[4];
  assign data_o[13316] = data_o[4];
  assign data_o[13380] = data_o[4];
  assign data_o[13444] = data_o[4];
  assign data_o[13508] = data_o[4];
  assign data_o[13572] = data_o[4];
  assign data_o[13636] = data_o[4];
  assign data_o[13700] = data_o[4];
  assign data_o[13764] = data_o[4];
  assign data_o[13828] = data_o[4];
  assign data_o[13892] = data_o[4];
  assign data_o[13956] = data_o[4];
  assign data_o[14020] = data_o[4];
  assign data_o[14084] = data_o[4];
  assign data_o[14148] = data_o[4];
  assign data_o[14212] = data_o[4];
  assign data_o[14276] = data_o[4];
  assign data_o[14340] = data_o[4];
  assign data_o[14404] = data_o[4];
  assign data_o[14468] = data_o[4];
  assign data_o[14532] = data_o[4];
  assign data_o[14596] = data_o[4];
  assign data_o[14660] = data_o[4];
  assign data_o[14724] = data_o[4];
  assign data_o[14788] = data_o[4];
  assign data_o[14852] = data_o[4];
  assign data_o[14916] = data_o[4];
  assign data_o[14980] = data_o[4];
  assign data_o[15044] = data_o[4];
  assign data_o[15108] = data_o[4];
  assign data_o[15172] = data_o[4];
  assign data_o[15236] = data_o[4];
  assign data_o[15300] = data_o[4];
  assign data_o[15364] = data_o[4];
  assign data_o[15428] = data_o[4];
  assign data_o[15492] = data_o[4];
  assign data_o[15556] = data_o[4];
  assign data_o[15620] = data_o[4];
  assign data_o[15684] = data_o[4];
  assign data_o[15748] = data_o[4];
  assign data_o[15812] = data_o[4];
  assign data_o[15876] = data_o[4];
  assign data_o[15940] = data_o[4];
  assign data_o[16004] = data_o[4];
  assign data_o[16068] = data_o[4];
  assign data_o[16132] = data_o[4];
  assign data_o[16196] = data_o[4];
  assign data_o[16260] = data_o[4];
  assign data_o[16324] = data_o[4];
  assign data_o[16388] = data_o[4];
  assign data_o[16452] = data_o[4];
  assign data_o[16516] = data_o[4];
  assign data_o[16580] = data_o[4];
  assign data_o[16644] = data_o[4];
  assign data_o[16708] = data_o[4];
  assign data_o[16772] = data_o[4];
  assign data_o[16836] = data_o[4];
  assign data_o[16900] = data_o[4];
  assign data_o[16964] = data_o[4];
  assign data_o[17028] = data_o[4];
  assign data_o[17092] = data_o[4];
  assign data_o[17156] = data_o[4];
  assign data_o[17220] = data_o[4];
  assign data_o[17284] = data_o[4];
  assign data_o[17348] = data_o[4];
  assign data_o[17412] = data_o[4];
  assign data_o[17476] = data_o[4];
  assign data_o[17540] = data_o[4];
  assign data_o[17604] = data_o[4];
  assign data_o[17668] = data_o[4];
  assign data_o[17732] = data_o[4];
  assign data_o[17796] = data_o[4];
  assign data_o[17860] = data_o[4];
  assign data_o[17924] = data_o[4];
  assign data_o[17988] = data_o[4];
  assign data_o[18052] = data_o[4];
  assign data_o[18116] = data_o[4];
  assign data_o[18180] = data_o[4];
  assign data_o[18244] = data_o[4];
  assign data_o[18308] = data_o[4];
  assign data_o[18372] = data_o[4];
  assign data_o[18436] = data_o[4];
  assign data_o[18500] = data_o[4];
  assign data_o[18564] = data_o[4];
  assign data_o[18628] = data_o[4];
  assign data_o[18692] = data_o[4];
  assign data_o[18756] = data_o[4];
  assign data_o[18820] = data_o[4];
  assign data_o[18884] = data_o[4];
  assign data_o[18948] = data_o[4];
  assign data_o[19012] = data_o[4];
  assign data_o[19076] = data_o[4];
  assign data_o[19140] = data_o[4];
  assign data_o[19204] = data_o[4];
  assign data_o[19268] = data_o[4];
  assign data_o[19332] = data_o[4];
  assign data_o[19396] = data_o[4];
  assign data_o[19460] = data_o[4];
  assign data_o[19524] = data_o[4];
  assign data_o[19588] = data_o[4];
  assign data_o[19652] = data_o[4];
  assign data_o[19716] = data_o[4];
  assign data_o[19780] = data_o[4];
  assign data_o[19844] = data_o[4];
  assign data_o[19908] = data_o[4];
  assign data_o[19972] = data_o[4];
  assign data_o[20036] = data_o[4];
  assign data_o[20100] = data_o[4];
  assign data_o[20164] = data_o[4];
  assign data_o[20228] = data_o[4];
  assign data_o[20292] = data_o[4];
  assign data_o[20356] = data_o[4];
  assign data_o[20420] = data_o[4];
  assign data_o[20484] = data_o[4];
  assign data_o[20548] = data_o[4];
  assign data_o[20612] = data_o[4];
  assign data_o[20676] = data_o[4];
  assign data_o[20740] = data_o[4];
  assign data_o[20804] = data_o[4];
  assign data_o[20868] = data_o[4];
  assign data_o[20932] = data_o[4];
  assign data_o[20996] = data_o[4];
  assign data_o[21060] = data_o[4];
  assign data_o[21124] = data_o[4];
  assign data_o[21188] = data_o[4];
  assign data_o[21252] = data_o[4];
  assign data_o[21316] = data_o[4];
  assign data_o[21380] = data_o[4];
  assign data_o[21444] = data_o[4];
  assign data_o[21508] = data_o[4];
  assign data_o[21572] = data_o[4];
  assign data_o[21636] = data_o[4];
  assign data_o[21700] = data_o[4];
  assign data_o[21764] = data_o[4];
  assign data_o[21828] = data_o[4];
  assign data_o[21892] = data_o[4];
  assign data_o[21956] = data_o[4];
  assign data_o[22020] = data_o[4];
  assign data_o[22084] = data_o[4];
  assign data_o[22148] = data_o[4];
  assign data_o[22212] = data_o[4];
  assign data_o[22276] = data_o[4];
  assign data_o[22340] = data_o[4];
  assign data_o[22404] = data_o[4];
  assign data_o[22468] = data_o[4];
  assign data_o[22532] = data_o[4];
  assign data_o[22596] = data_o[4];
  assign data_o[22660] = data_o[4];
  assign data_o[22724] = data_o[4];
  assign data_o[22788] = data_o[4];
  assign data_o[22852] = data_o[4];
  assign data_o[22916] = data_o[4];
  assign data_o[22980] = data_o[4];
  assign data_o[23044] = data_o[4];
  assign data_o[23108] = data_o[4];
  assign data_o[23172] = data_o[4];
  assign data_o[23236] = data_o[4];
  assign data_o[23300] = data_o[4];
  assign data_o[23364] = data_o[4];
  assign data_o[23428] = data_o[4];
  assign data_o[23492] = data_o[4];
  assign data_o[23556] = data_o[4];
  assign data_o[23620] = data_o[4];
  assign data_o[23684] = data_o[4];
  assign data_o[23748] = data_o[4];
  assign data_o[23812] = data_o[4];
  assign data_o[23876] = data_o[4];
  assign data_o[23940] = data_o[4];
  assign data_o[24004] = data_o[4];
  assign data_o[24068] = data_o[4];
  assign data_o[24132] = data_o[4];
  assign data_o[24196] = data_o[4];
  assign data_o[24260] = data_o[4];
  assign data_o[24324] = data_o[4];
  assign data_o[24388] = data_o[4];
  assign data_o[24452] = data_o[4];
  assign data_o[24516] = data_o[4];
  assign data_o[24580] = data_o[4];
  assign data_o[24644] = data_o[4];
  assign data_o[24708] = data_o[4];
  assign data_o[24772] = data_o[4];
  assign data_o[24836] = data_o[4];
  assign data_o[24900] = data_o[4];
  assign data_o[24964] = data_o[4];
  assign data_o[25028] = data_o[4];
  assign data_o[25092] = data_o[4];
  assign data_o[25156] = data_o[4];
  assign data_o[25220] = data_o[4];
  assign data_o[25284] = data_o[4];
  assign data_o[25348] = data_o[4];
  assign data_o[25412] = data_o[4];
  assign data_o[25476] = data_o[4];
  assign data_o[25540] = data_o[4];
  assign data_o[25604] = data_o[4];
  assign data_o[25668] = data_o[4];
  assign data_o[25732] = data_o[4];
  assign data_o[25796] = data_o[4];
  assign data_o[25860] = data_o[4];
  assign data_o[25924] = data_o[4];
  assign data_o[25988] = data_o[4];
  assign data_o[26052] = data_o[4];
  assign data_o[26116] = data_o[4];
  assign data_o[26180] = data_o[4];
  assign data_o[26244] = data_o[4];
  assign data_o[26308] = data_o[4];
  assign data_o[26372] = data_o[4];
  assign data_o[26436] = data_o[4];
  assign data_o[26500] = data_o[4];
  assign data_o[26564] = data_o[4];
  assign data_o[26628] = data_o[4];
  assign data_o[26692] = data_o[4];
  assign data_o[26756] = data_o[4];
  assign data_o[26820] = data_o[4];
  assign data_o[26884] = data_o[4];
  assign data_o[26948] = data_o[4];
  assign data_o[27012] = data_o[4];
  assign data_o[27076] = data_o[4];
  assign data_o[27140] = data_o[4];
  assign data_o[27204] = data_o[4];
  assign data_o[27268] = data_o[4];
  assign data_o[27332] = data_o[4];
  assign data_o[27396] = data_o[4];
  assign data_o[27460] = data_o[4];
  assign data_o[27524] = data_o[4];
  assign data_o[27588] = data_o[4];
  assign data_o[27652] = data_o[4];
  assign data_o[27716] = data_o[4];
  assign data_o[27780] = data_o[4];
  assign data_o[27844] = data_o[4];
  assign data_o[27908] = data_o[4];
  assign data_o[27972] = data_o[4];
  assign data_o[28036] = data_o[4];
  assign data_o[28100] = data_o[4];
  assign data_o[28164] = data_o[4];
  assign data_o[28228] = data_o[4];
  assign data_o[28292] = data_o[4];
  assign data_o[28356] = data_o[4];
  assign data_o[28420] = data_o[4];
  assign data_o[28484] = data_o[4];
  assign data_o[28548] = data_o[4];
  assign data_o[28612] = data_o[4];
  assign data_o[28676] = data_o[4];
  assign data_o[28740] = data_o[4];
  assign data_o[28804] = data_o[4];
  assign data_o[28868] = data_o[4];
  assign data_o[28932] = data_o[4];
  assign data_o[28996] = data_o[4];
  assign data_o[29060] = data_o[4];
  assign data_o[29124] = data_o[4];
  assign data_o[29188] = data_o[4];
  assign data_o[29252] = data_o[4];
  assign data_o[29316] = data_o[4];
  assign data_o[29380] = data_o[4];
  assign data_o[29444] = data_o[4];
  assign data_o[29508] = data_o[4];
  assign data_o[29572] = data_o[4];
  assign data_o[29636] = data_o[4];
  assign data_o[29700] = data_o[4];
  assign data_o[29764] = data_o[4];
  assign data_o[29828] = data_o[4];
  assign data_o[29892] = data_o[4];
  assign data_o[29956] = data_o[4];
  assign data_o[30020] = data_o[4];
  assign data_o[30084] = data_o[4];
  assign data_o[30148] = data_o[4];
  assign data_o[30212] = data_o[4];
  assign data_o[30276] = data_o[4];
  assign data_o[30340] = data_o[4];
  assign data_o[30404] = data_o[4];
  assign data_o[30468] = data_o[4];
  assign data_o[30532] = data_o[4];
  assign data_o[30596] = data_o[4];
  assign data_o[30660] = data_o[4];
  assign data_o[30724] = data_o[4];
  assign data_o[30788] = data_o[4];
  assign data_o[30852] = data_o[4];
  assign data_o[30916] = data_o[4];
  assign data_o[30980] = data_o[4];
  assign data_o[31044] = data_o[4];
  assign data_o[31108] = data_o[4];
  assign data_o[31172] = data_o[4];
  assign data_o[31236] = data_o[4];
  assign data_o[31300] = data_o[4];
  assign data_o[31364] = data_o[4];
  assign data_o[31428] = data_o[4];
  assign data_o[31492] = data_o[4];
  assign data_o[31556] = data_o[4];
  assign data_o[31620] = data_o[4];
  assign data_o[31684] = data_o[4];
  assign data_o[31748] = data_o[4];
  assign data_o[31812] = data_o[4];
  assign data_o[31876] = data_o[4];
  assign data_o[31940] = data_o[4];
  assign data_o[67] = data_o[3];
  assign data_o[131] = data_o[3];
  assign data_o[195] = data_o[3];
  assign data_o[259] = data_o[3];
  assign data_o[323] = data_o[3];
  assign data_o[387] = data_o[3];
  assign data_o[451] = data_o[3];
  assign data_o[515] = data_o[3];
  assign data_o[579] = data_o[3];
  assign data_o[643] = data_o[3];
  assign data_o[707] = data_o[3];
  assign data_o[771] = data_o[3];
  assign data_o[835] = data_o[3];
  assign data_o[899] = data_o[3];
  assign data_o[963] = data_o[3];
  assign data_o[1027] = data_o[3];
  assign data_o[1091] = data_o[3];
  assign data_o[1155] = data_o[3];
  assign data_o[1219] = data_o[3];
  assign data_o[1283] = data_o[3];
  assign data_o[1347] = data_o[3];
  assign data_o[1411] = data_o[3];
  assign data_o[1475] = data_o[3];
  assign data_o[1539] = data_o[3];
  assign data_o[1603] = data_o[3];
  assign data_o[1667] = data_o[3];
  assign data_o[1731] = data_o[3];
  assign data_o[1795] = data_o[3];
  assign data_o[1859] = data_o[3];
  assign data_o[1923] = data_o[3];
  assign data_o[1987] = data_o[3];
  assign data_o[2051] = data_o[3];
  assign data_o[2115] = data_o[3];
  assign data_o[2179] = data_o[3];
  assign data_o[2243] = data_o[3];
  assign data_o[2307] = data_o[3];
  assign data_o[2371] = data_o[3];
  assign data_o[2435] = data_o[3];
  assign data_o[2499] = data_o[3];
  assign data_o[2563] = data_o[3];
  assign data_o[2627] = data_o[3];
  assign data_o[2691] = data_o[3];
  assign data_o[2755] = data_o[3];
  assign data_o[2819] = data_o[3];
  assign data_o[2883] = data_o[3];
  assign data_o[2947] = data_o[3];
  assign data_o[3011] = data_o[3];
  assign data_o[3075] = data_o[3];
  assign data_o[3139] = data_o[3];
  assign data_o[3203] = data_o[3];
  assign data_o[3267] = data_o[3];
  assign data_o[3331] = data_o[3];
  assign data_o[3395] = data_o[3];
  assign data_o[3459] = data_o[3];
  assign data_o[3523] = data_o[3];
  assign data_o[3587] = data_o[3];
  assign data_o[3651] = data_o[3];
  assign data_o[3715] = data_o[3];
  assign data_o[3779] = data_o[3];
  assign data_o[3843] = data_o[3];
  assign data_o[3907] = data_o[3];
  assign data_o[3971] = data_o[3];
  assign data_o[4035] = data_o[3];
  assign data_o[4099] = data_o[3];
  assign data_o[4163] = data_o[3];
  assign data_o[4227] = data_o[3];
  assign data_o[4291] = data_o[3];
  assign data_o[4355] = data_o[3];
  assign data_o[4419] = data_o[3];
  assign data_o[4483] = data_o[3];
  assign data_o[4547] = data_o[3];
  assign data_o[4611] = data_o[3];
  assign data_o[4675] = data_o[3];
  assign data_o[4739] = data_o[3];
  assign data_o[4803] = data_o[3];
  assign data_o[4867] = data_o[3];
  assign data_o[4931] = data_o[3];
  assign data_o[4995] = data_o[3];
  assign data_o[5059] = data_o[3];
  assign data_o[5123] = data_o[3];
  assign data_o[5187] = data_o[3];
  assign data_o[5251] = data_o[3];
  assign data_o[5315] = data_o[3];
  assign data_o[5379] = data_o[3];
  assign data_o[5443] = data_o[3];
  assign data_o[5507] = data_o[3];
  assign data_o[5571] = data_o[3];
  assign data_o[5635] = data_o[3];
  assign data_o[5699] = data_o[3];
  assign data_o[5763] = data_o[3];
  assign data_o[5827] = data_o[3];
  assign data_o[5891] = data_o[3];
  assign data_o[5955] = data_o[3];
  assign data_o[6019] = data_o[3];
  assign data_o[6083] = data_o[3];
  assign data_o[6147] = data_o[3];
  assign data_o[6211] = data_o[3];
  assign data_o[6275] = data_o[3];
  assign data_o[6339] = data_o[3];
  assign data_o[6403] = data_o[3];
  assign data_o[6467] = data_o[3];
  assign data_o[6531] = data_o[3];
  assign data_o[6595] = data_o[3];
  assign data_o[6659] = data_o[3];
  assign data_o[6723] = data_o[3];
  assign data_o[6787] = data_o[3];
  assign data_o[6851] = data_o[3];
  assign data_o[6915] = data_o[3];
  assign data_o[6979] = data_o[3];
  assign data_o[7043] = data_o[3];
  assign data_o[7107] = data_o[3];
  assign data_o[7171] = data_o[3];
  assign data_o[7235] = data_o[3];
  assign data_o[7299] = data_o[3];
  assign data_o[7363] = data_o[3];
  assign data_o[7427] = data_o[3];
  assign data_o[7491] = data_o[3];
  assign data_o[7555] = data_o[3];
  assign data_o[7619] = data_o[3];
  assign data_o[7683] = data_o[3];
  assign data_o[7747] = data_o[3];
  assign data_o[7811] = data_o[3];
  assign data_o[7875] = data_o[3];
  assign data_o[7939] = data_o[3];
  assign data_o[8003] = data_o[3];
  assign data_o[8067] = data_o[3];
  assign data_o[8131] = data_o[3];
  assign data_o[8195] = data_o[3];
  assign data_o[8259] = data_o[3];
  assign data_o[8323] = data_o[3];
  assign data_o[8387] = data_o[3];
  assign data_o[8451] = data_o[3];
  assign data_o[8515] = data_o[3];
  assign data_o[8579] = data_o[3];
  assign data_o[8643] = data_o[3];
  assign data_o[8707] = data_o[3];
  assign data_o[8771] = data_o[3];
  assign data_o[8835] = data_o[3];
  assign data_o[8899] = data_o[3];
  assign data_o[8963] = data_o[3];
  assign data_o[9027] = data_o[3];
  assign data_o[9091] = data_o[3];
  assign data_o[9155] = data_o[3];
  assign data_o[9219] = data_o[3];
  assign data_o[9283] = data_o[3];
  assign data_o[9347] = data_o[3];
  assign data_o[9411] = data_o[3];
  assign data_o[9475] = data_o[3];
  assign data_o[9539] = data_o[3];
  assign data_o[9603] = data_o[3];
  assign data_o[9667] = data_o[3];
  assign data_o[9731] = data_o[3];
  assign data_o[9795] = data_o[3];
  assign data_o[9859] = data_o[3];
  assign data_o[9923] = data_o[3];
  assign data_o[9987] = data_o[3];
  assign data_o[10051] = data_o[3];
  assign data_o[10115] = data_o[3];
  assign data_o[10179] = data_o[3];
  assign data_o[10243] = data_o[3];
  assign data_o[10307] = data_o[3];
  assign data_o[10371] = data_o[3];
  assign data_o[10435] = data_o[3];
  assign data_o[10499] = data_o[3];
  assign data_o[10563] = data_o[3];
  assign data_o[10627] = data_o[3];
  assign data_o[10691] = data_o[3];
  assign data_o[10755] = data_o[3];
  assign data_o[10819] = data_o[3];
  assign data_o[10883] = data_o[3];
  assign data_o[10947] = data_o[3];
  assign data_o[11011] = data_o[3];
  assign data_o[11075] = data_o[3];
  assign data_o[11139] = data_o[3];
  assign data_o[11203] = data_o[3];
  assign data_o[11267] = data_o[3];
  assign data_o[11331] = data_o[3];
  assign data_o[11395] = data_o[3];
  assign data_o[11459] = data_o[3];
  assign data_o[11523] = data_o[3];
  assign data_o[11587] = data_o[3];
  assign data_o[11651] = data_o[3];
  assign data_o[11715] = data_o[3];
  assign data_o[11779] = data_o[3];
  assign data_o[11843] = data_o[3];
  assign data_o[11907] = data_o[3];
  assign data_o[11971] = data_o[3];
  assign data_o[12035] = data_o[3];
  assign data_o[12099] = data_o[3];
  assign data_o[12163] = data_o[3];
  assign data_o[12227] = data_o[3];
  assign data_o[12291] = data_o[3];
  assign data_o[12355] = data_o[3];
  assign data_o[12419] = data_o[3];
  assign data_o[12483] = data_o[3];
  assign data_o[12547] = data_o[3];
  assign data_o[12611] = data_o[3];
  assign data_o[12675] = data_o[3];
  assign data_o[12739] = data_o[3];
  assign data_o[12803] = data_o[3];
  assign data_o[12867] = data_o[3];
  assign data_o[12931] = data_o[3];
  assign data_o[12995] = data_o[3];
  assign data_o[13059] = data_o[3];
  assign data_o[13123] = data_o[3];
  assign data_o[13187] = data_o[3];
  assign data_o[13251] = data_o[3];
  assign data_o[13315] = data_o[3];
  assign data_o[13379] = data_o[3];
  assign data_o[13443] = data_o[3];
  assign data_o[13507] = data_o[3];
  assign data_o[13571] = data_o[3];
  assign data_o[13635] = data_o[3];
  assign data_o[13699] = data_o[3];
  assign data_o[13763] = data_o[3];
  assign data_o[13827] = data_o[3];
  assign data_o[13891] = data_o[3];
  assign data_o[13955] = data_o[3];
  assign data_o[14019] = data_o[3];
  assign data_o[14083] = data_o[3];
  assign data_o[14147] = data_o[3];
  assign data_o[14211] = data_o[3];
  assign data_o[14275] = data_o[3];
  assign data_o[14339] = data_o[3];
  assign data_o[14403] = data_o[3];
  assign data_o[14467] = data_o[3];
  assign data_o[14531] = data_o[3];
  assign data_o[14595] = data_o[3];
  assign data_o[14659] = data_o[3];
  assign data_o[14723] = data_o[3];
  assign data_o[14787] = data_o[3];
  assign data_o[14851] = data_o[3];
  assign data_o[14915] = data_o[3];
  assign data_o[14979] = data_o[3];
  assign data_o[15043] = data_o[3];
  assign data_o[15107] = data_o[3];
  assign data_o[15171] = data_o[3];
  assign data_o[15235] = data_o[3];
  assign data_o[15299] = data_o[3];
  assign data_o[15363] = data_o[3];
  assign data_o[15427] = data_o[3];
  assign data_o[15491] = data_o[3];
  assign data_o[15555] = data_o[3];
  assign data_o[15619] = data_o[3];
  assign data_o[15683] = data_o[3];
  assign data_o[15747] = data_o[3];
  assign data_o[15811] = data_o[3];
  assign data_o[15875] = data_o[3];
  assign data_o[15939] = data_o[3];
  assign data_o[16003] = data_o[3];
  assign data_o[16067] = data_o[3];
  assign data_o[16131] = data_o[3];
  assign data_o[16195] = data_o[3];
  assign data_o[16259] = data_o[3];
  assign data_o[16323] = data_o[3];
  assign data_o[16387] = data_o[3];
  assign data_o[16451] = data_o[3];
  assign data_o[16515] = data_o[3];
  assign data_o[16579] = data_o[3];
  assign data_o[16643] = data_o[3];
  assign data_o[16707] = data_o[3];
  assign data_o[16771] = data_o[3];
  assign data_o[16835] = data_o[3];
  assign data_o[16899] = data_o[3];
  assign data_o[16963] = data_o[3];
  assign data_o[17027] = data_o[3];
  assign data_o[17091] = data_o[3];
  assign data_o[17155] = data_o[3];
  assign data_o[17219] = data_o[3];
  assign data_o[17283] = data_o[3];
  assign data_o[17347] = data_o[3];
  assign data_o[17411] = data_o[3];
  assign data_o[17475] = data_o[3];
  assign data_o[17539] = data_o[3];
  assign data_o[17603] = data_o[3];
  assign data_o[17667] = data_o[3];
  assign data_o[17731] = data_o[3];
  assign data_o[17795] = data_o[3];
  assign data_o[17859] = data_o[3];
  assign data_o[17923] = data_o[3];
  assign data_o[17987] = data_o[3];
  assign data_o[18051] = data_o[3];
  assign data_o[18115] = data_o[3];
  assign data_o[18179] = data_o[3];
  assign data_o[18243] = data_o[3];
  assign data_o[18307] = data_o[3];
  assign data_o[18371] = data_o[3];
  assign data_o[18435] = data_o[3];
  assign data_o[18499] = data_o[3];
  assign data_o[18563] = data_o[3];
  assign data_o[18627] = data_o[3];
  assign data_o[18691] = data_o[3];
  assign data_o[18755] = data_o[3];
  assign data_o[18819] = data_o[3];
  assign data_o[18883] = data_o[3];
  assign data_o[18947] = data_o[3];
  assign data_o[19011] = data_o[3];
  assign data_o[19075] = data_o[3];
  assign data_o[19139] = data_o[3];
  assign data_o[19203] = data_o[3];
  assign data_o[19267] = data_o[3];
  assign data_o[19331] = data_o[3];
  assign data_o[19395] = data_o[3];
  assign data_o[19459] = data_o[3];
  assign data_o[19523] = data_o[3];
  assign data_o[19587] = data_o[3];
  assign data_o[19651] = data_o[3];
  assign data_o[19715] = data_o[3];
  assign data_o[19779] = data_o[3];
  assign data_o[19843] = data_o[3];
  assign data_o[19907] = data_o[3];
  assign data_o[19971] = data_o[3];
  assign data_o[20035] = data_o[3];
  assign data_o[20099] = data_o[3];
  assign data_o[20163] = data_o[3];
  assign data_o[20227] = data_o[3];
  assign data_o[20291] = data_o[3];
  assign data_o[20355] = data_o[3];
  assign data_o[20419] = data_o[3];
  assign data_o[20483] = data_o[3];
  assign data_o[20547] = data_o[3];
  assign data_o[20611] = data_o[3];
  assign data_o[20675] = data_o[3];
  assign data_o[20739] = data_o[3];
  assign data_o[20803] = data_o[3];
  assign data_o[20867] = data_o[3];
  assign data_o[20931] = data_o[3];
  assign data_o[20995] = data_o[3];
  assign data_o[21059] = data_o[3];
  assign data_o[21123] = data_o[3];
  assign data_o[21187] = data_o[3];
  assign data_o[21251] = data_o[3];
  assign data_o[21315] = data_o[3];
  assign data_o[21379] = data_o[3];
  assign data_o[21443] = data_o[3];
  assign data_o[21507] = data_o[3];
  assign data_o[21571] = data_o[3];
  assign data_o[21635] = data_o[3];
  assign data_o[21699] = data_o[3];
  assign data_o[21763] = data_o[3];
  assign data_o[21827] = data_o[3];
  assign data_o[21891] = data_o[3];
  assign data_o[21955] = data_o[3];
  assign data_o[22019] = data_o[3];
  assign data_o[22083] = data_o[3];
  assign data_o[22147] = data_o[3];
  assign data_o[22211] = data_o[3];
  assign data_o[22275] = data_o[3];
  assign data_o[22339] = data_o[3];
  assign data_o[22403] = data_o[3];
  assign data_o[22467] = data_o[3];
  assign data_o[22531] = data_o[3];
  assign data_o[22595] = data_o[3];
  assign data_o[22659] = data_o[3];
  assign data_o[22723] = data_o[3];
  assign data_o[22787] = data_o[3];
  assign data_o[22851] = data_o[3];
  assign data_o[22915] = data_o[3];
  assign data_o[22979] = data_o[3];
  assign data_o[23043] = data_o[3];
  assign data_o[23107] = data_o[3];
  assign data_o[23171] = data_o[3];
  assign data_o[23235] = data_o[3];
  assign data_o[23299] = data_o[3];
  assign data_o[23363] = data_o[3];
  assign data_o[23427] = data_o[3];
  assign data_o[23491] = data_o[3];
  assign data_o[23555] = data_o[3];
  assign data_o[23619] = data_o[3];
  assign data_o[23683] = data_o[3];
  assign data_o[23747] = data_o[3];
  assign data_o[23811] = data_o[3];
  assign data_o[23875] = data_o[3];
  assign data_o[23939] = data_o[3];
  assign data_o[24003] = data_o[3];
  assign data_o[24067] = data_o[3];
  assign data_o[24131] = data_o[3];
  assign data_o[24195] = data_o[3];
  assign data_o[24259] = data_o[3];
  assign data_o[24323] = data_o[3];
  assign data_o[24387] = data_o[3];
  assign data_o[24451] = data_o[3];
  assign data_o[24515] = data_o[3];
  assign data_o[24579] = data_o[3];
  assign data_o[24643] = data_o[3];
  assign data_o[24707] = data_o[3];
  assign data_o[24771] = data_o[3];
  assign data_o[24835] = data_o[3];
  assign data_o[24899] = data_o[3];
  assign data_o[24963] = data_o[3];
  assign data_o[25027] = data_o[3];
  assign data_o[25091] = data_o[3];
  assign data_o[25155] = data_o[3];
  assign data_o[25219] = data_o[3];
  assign data_o[25283] = data_o[3];
  assign data_o[25347] = data_o[3];
  assign data_o[25411] = data_o[3];
  assign data_o[25475] = data_o[3];
  assign data_o[25539] = data_o[3];
  assign data_o[25603] = data_o[3];
  assign data_o[25667] = data_o[3];
  assign data_o[25731] = data_o[3];
  assign data_o[25795] = data_o[3];
  assign data_o[25859] = data_o[3];
  assign data_o[25923] = data_o[3];
  assign data_o[25987] = data_o[3];
  assign data_o[26051] = data_o[3];
  assign data_o[26115] = data_o[3];
  assign data_o[26179] = data_o[3];
  assign data_o[26243] = data_o[3];
  assign data_o[26307] = data_o[3];
  assign data_o[26371] = data_o[3];
  assign data_o[26435] = data_o[3];
  assign data_o[26499] = data_o[3];
  assign data_o[26563] = data_o[3];
  assign data_o[26627] = data_o[3];
  assign data_o[26691] = data_o[3];
  assign data_o[26755] = data_o[3];
  assign data_o[26819] = data_o[3];
  assign data_o[26883] = data_o[3];
  assign data_o[26947] = data_o[3];
  assign data_o[27011] = data_o[3];
  assign data_o[27075] = data_o[3];
  assign data_o[27139] = data_o[3];
  assign data_o[27203] = data_o[3];
  assign data_o[27267] = data_o[3];
  assign data_o[27331] = data_o[3];
  assign data_o[27395] = data_o[3];
  assign data_o[27459] = data_o[3];
  assign data_o[27523] = data_o[3];
  assign data_o[27587] = data_o[3];
  assign data_o[27651] = data_o[3];
  assign data_o[27715] = data_o[3];
  assign data_o[27779] = data_o[3];
  assign data_o[27843] = data_o[3];
  assign data_o[27907] = data_o[3];
  assign data_o[27971] = data_o[3];
  assign data_o[28035] = data_o[3];
  assign data_o[28099] = data_o[3];
  assign data_o[28163] = data_o[3];
  assign data_o[28227] = data_o[3];
  assign data_o[28291] = data_o[3];
  assign data_o[28355] = data_o[3];
  assign data_o[28419] = data_o[3];
  assign data_o[28483] = data_o[3];
  assign data_o[28547] = data_o[3];
  assign data_o[28611] = data_o[3];
  assign data_o[28675] = data_o[3];
  assign data_o[28739] = data_o[3];
  assign data_o[28803] = data_o[3];
  assign data_o[28867] = data_o[3];
  assign data_o[28931] = data_o[3];
  assign data_o[28995] = data_o[3];
  assign data_o[29059] = data_o[3];
  assign data_o[29123] = data_o[3];
  assign data_o[29187] = data_o[3];
  assign data_o[29251] = data_o[3];
  assign data_o[29315] = data_o[3];
  assign data_o[29379] = data_o[3];
  assign data_o[29443] = data_o[3];
  assign data_o[29507] = data_o[3];
  assign data_o[29571] = data_o[3];
  assign data_o[29635] = data_o[3];
  assign data_o[29699] = data_o[3];
  assign data_o[29763] = data_o[3];
  assign data_o[29827] = data_o[3];
  assign data_o[29891] = data_o[3];
  assign data_o[29955] = data_o[3];
  assign data_o[30019] = data_o[3];
  assign data_o[30083] = data_o[3];
  assign data_o[30147] = data_o[3];
  assign data_o[30211] = data_o[3];
  assign data_o[30275] = data_o[3];
  assign data_o[30339] = data_o[3];
  assign data_o[30403] = data_o[3];
  assign data_o[30467] = data_o[3];
  assign data_o[30531] = data_o[3];
  assign data_o[30595] = data_o[3];
  assign data_o[30659] = data_o[3];
  assign data_o[30723] = data_o[3];
  assign data_o[30787] = data_o[3];
  assign data_o[30851] = data_o[3];
  assign data_o[30915] = data_o[3];
  assign data_o[30979] = data_o[3];
  assign data_o[31043] = data_o[3];
  assign data_o[31107] = data_o[3];
  assign data_o[31171] = data_o[3];
  assign data_o[31235] = data_o[3];
  assign data_o[31299] = data_o[3];
  assign data_o[31363] = data_o[3];
  assign data_o[31427] = data_o[3];
  assign data_o[31491] = data_o[3];
  assign data_o[31555] = data_o[3];
  assign data_o[31619] = data_o[3];
  assign data_o[31683] = data_o[3];
  assign data_o[31747] = data_o[3];
  assign data_o[31811] = data_o[3];
  assign data_o[31875] = data_o[3];
  assign data_o[31939] = data_o[3];
  assign data_o[66] = data_o[2];
  assign data_o[130] = data_o[2];
  assign data_o[194] = data_o[2];
  assign data_o[258] = data_o[2];
  assign data_o[322] = data_o[2];
  assign data_o[386] = data_o[2];
  assign data_o[450] = data_o[2];
  assign data_o[514] = data_o[2];
  assign data_o[578] = data_o[2];
  assign data_o[642] = data_o[2];
  assign data_o[706] = data_o[2];
  assign data_o[770] = data_o[2];
  assign data_o[834] = data_o[2];
  assign data_o[898] = data_o[2];
  assign data_o[962] = data_o[2];
  assign data_o[1026] = data_o[2];
  assign data_o[1090] = data_o[2];
  assign data_o[1154] = data_o[2];
  assign data_o[1218] = data_o[2];
  assign data_o[1282] = data_o[2];
  assign data_o[1346] = data_o[2];
  assign data_o[1410] = data_o[2];
  assign data_o[1474] = data_o[2];
  assign data_o[1538] = data_o[2];
  assign data_o[1602] = data_o[2];
  assign data_o[1666] = data_o[2];
  assign data_o[1730] = data_o[2];
  assign data_o[1794] = data_o[2];
  assign data_o[1858] = data_o[2];
  assign data_o[1922] = data_o[2];
  assign data_o[1986] = data_o[2];
  assign data_o[2050] = data_o[2];
  assign data_o[2114] = data_o[2];
  assign data_o[2178] = data_o[2];
  assign data_o[2242] = data_o[2];
  assign data_o[2306] = data_o[2];
  assign data_o[2370] = data_o[2];
  assign data_o[2434] = data_o[2];
  assign data_o[2498] = data_o[2];
  assign data_o[2562] = data_o[2];
  assign data_o[2626] = data_o[2];
  assign data_o[2690] = data_o[2];
  assign data_o[2754] = data_o[2];
  assign data_o[2818] = data_o[2];
  assign data_o[2882] = data_o[2];
  assign data_o[2946] = data_o[2];
  assign data_o[3010] = data_o[2];
  assign data_o[3074] = data_o[2];
  assign data_o[3138] = data_o[2];
  assign data_o[3202] = data_o[2];
  assign data_o[3266] = data_o[2];
  assign data_o[3330] = data_o[2];
  assign data_o[3394] = data_o[2];
  assign data_o[3458] = data_o[2];
  assign data_o[3522] = data_o[2];
  assign data_o[3586] = data_o[2];
  assign data_o[3650] = data_o[2];
  assign data_o[3714] = data_o[2];
  assign data_o[3778] = data_o[2];
  assign data_o[3842] = data_o[2];
  assign data_o[3906] = data_o[2];
  assign data_o[3970] = data_o[2];
  assign data_o[4034] = data_o[2];
  assign data_o[4098] = data_o[2];
  assign data_o[4162] = data_o[2];
  assign data_o[4226] = data_o[2];
  assign data_o[4290] = data_o[2];
  assign data_o[4354] = data_o[2];
  assign data_o[4418] = data_o[2];
  assign data_o[4482] = data_o[2];
  assign data_o[4546] = data_o[2];
  assign data_o[4610] = data_o[2];
  assign data_o[4674] = data_o[2];
  assign data_o[4738] = data_o[2];
  assign data_o[4802] = data_o[2];
  assign data_o[4866] = data_o[2];
  assign data_o[4930] = data_o[2];
  assign data_o[4994] = data_o[2];
  assign data_o[5058] = data_o[2];
  assign data_o[5122] = data_o[2];
  assign data_o[5186] = data_o[2];
  assign data_o[5250] = data_o[2];
  assign data_o[5314] = data_o[2];
  assign data_o[5378] = data_o[2];
  assign data_o[5442] = data_o[2];
  assign data_o[5506] = data_o[2];
  assign data_o[5570] = data_o[2];
  assign data_o[5634] = data_o[2];
  assign data_o[5698] = data_o[2];
  assign data_o[5762] = data_o[2];
  assign data_o[5826] = data_o[2];
  assign data_o[5890] = data_o[2];
  assign data_o[5954] = data_o[2];
  assign data_o[6018] = data_o[2];
  assign data_o[6082] = data_o[2];
  assign data_o[6146] = data_o[2];
  assign data_o[6210] = data_o[2];
  assign data_o[6274] = data_o[2];
  assign data_o[6338] = data_o[2];
  assign data_o[6402] = data_o[2];
  assign data_o[6466] = data_o[2];
  assign data_o[6530] = data_o[2];
  assign data_o[6594] = data_o[2];
  assign data_o[6658] = data_o[2];
  assign data_o[6722] = data_o[2];
  assign data_o[6786] = data_o[2];
  assign data_o[6850] = data_o[2];
  assign data_o[6914] = data_o[2];
  assign data_o[6978] = data_o[2];
  assign data_o[7042] = data_o[2];
  assign data_o[7106] = data_o[2];
  assign data_o[7170] = data_o[2];
  assign data_o[7234] = data_o[2];
  assign data_o[7298] = data_o[2];
  assign data_o[7362] = data_o[2];
  assign data_o[7426] = data_o[2];
  assign data_o[7490] = data_o[2];
  assign data_o[7554] = data_o[2];
  assign data_o[7618] = data_o[2];
  assign data_o[7682] = data_o[2];
  assign data_o[7746] = data_o[2];
  assign data_o[7810] = data_o[2];
  assign data_o[7874] = data_o[2];
  assign data_o[7938] = data_o[2];
  assign data_o[8002] = data_o[2];
  assign data_o[8066] = data_o[2];
  assign data_o[8130] = data_o[2];
  assign data_o[8194] = data_o[2];
  assign data_o[8258] = data_o[2];
  assign data_o[8322] = data_o[2];
  assign data_o[8386] = data_o[2];
  assign data_o[8450] = data_o[2];
  assign data_o[8514] = data_o[2];
  assign data_o[8578] = data_o[2];
  assign data_o[8642] = data_o[2];
  assign data_o[8706] = data_o[2];
  assign data_o[8770] = data_o[2];
  assign data_o[8834] = data_o[2];
  assign data_o[8898] = data_o[2];
  assign data_o[8962] = data_o[2];
  assign data_o[9026] = data_o[2];
  assign data_o[9090] = data_o[2];
  assign data_o[9154] = data_o[2];
  assign data_o[9218] = data_o[2];
  assign data_o[9282] = data_o[2];
  assign data_o[9346] = data_o[2];
  assign data_o[9410] = data_o[2];
  assign data_o[9474] = data_o[2];
  assign data_o[9538] = data_o[2];
  assign data_o[9602] = data_o[2];
  assign data_o[9666] = data_o[2];
  assign data_o[9730] = data_o[2];
  assign data_o[9794] = data_o[2];
  assign data_o[9858] = data_o[2];
  assign data_o[9922] = data_o[2];
  assign data_o[9986] = data_o[2];
  assign data_o[10050] = data_o[2];
  assign data_o[10114] = data_o[2];
  assign data_o[10178] = data_o[2];
  assign data_o[10242] = data_o[2];
  assign data_o[10306] = data_o[2];
  assign data_o[10370] = data_o[2];
  assign data_o[10434] = data_o[2];
  assign data_o[10498] = data_o[2];
  assign data_o[10562] = data_o[2];
  assign data_o[10626] = data_o[2];
  assign data_o[10690] = data_o[2];
  assign data_o[10754] = data_o[2];
  assign data_o[10818] = data_o[2];
  assign data_o[10882] = data_o[2];
  assign data_o[10946] = data_o[2];
  assign data_o[11010] = data_o[2];
  assign data_o[11074] = data_o[2];
  assign data_o[11138] = data_o[2];
  assign data_o[11202] = data_o[2];
  assign data_o[11266] = data_o[2];
  assign data_o[11330] = data_o[2];
  assign data_o[11394] = data_o[2];
  assign data_o[11458] = data_o[2];
  assign data_o[11522] = data_o[2];
  assign data_o[11586] = data_o[2];
  assign data_o[11650] = data_o[2];
  assign data_o[11714] = data_o[2];
  assign data_o[11778] = data_o[2];
  assign data_o[11842] = data_o[2];
  assign data_o[11906] = data_o[2];
  assign data_o[11970] = data_o[2];
  assign data_o[12034] = data_o[2];
  assign data_o[12098] = data_o[2];
  assign data_o[12162] = data_o[2];
  assign data_o[12226] = data_o[2];
  assign data_o[12290] = data_o[2];
  assign data_o[12354] = data_o[2];
  assign data_o[12418] = data_o[2];
  assign data_o[12482] = data_o[2];
  assign data_o[12546] = data_o[2];
  assign data_o[12610] = data_o[2];
  assign data_o[12674] = data_o[2];
  assign data_o[12738] = data_o[2];
  assign data_o[12802] = data_o[2];
  assign data_o[12866] = data_o[2];
  assign data_o[12930] = data_o[2];
  assign data_o[12994] = data_o[2];
  assign data_o[13058] = data_o[2];
  assign data_o[13122] = data_o[2];
  assign data_o[13186] = data_o[2];
  assign data_o[13250] = data_o[2];
  assign data_o[13314] = data_o[2];
  assign data_o[13378] = data_o[2];
  assign data_o[13442] = data_o[2];
  assign data_o[13506] = data_o[2];
  assign data_o[13570] = data_o[2];
  assign data_o[13634] = data_o[2];
  assign data_o[13698] = data_o[2];
  assign data_o[13762] = data_o[2];
  assign data_o[13826] = data_o[2];
  assign data_o[13890] = data_o[2];
  assign data_o[13954] = data_o[2];
  assign data_o[14018] = data_o[2];
  assign data_o[14082] = data_o[2];
  assign data_o[14146] = data_o[2];
  assign data_o[14210] = data_o[2];
  assign data_o[14274] = data_o[2];
  assign data_o[14338] = data_o[2];
  assign data_o[14402] = data_o[2];
  assign data_o[14466] = data_o[2];
  assign data_o[14530] = data_o[2];
  assign data_o[14594] = data_o[2];
  assign data_o[14658] = data_o[2];
  assign data_o[14722] = data_o[2];
  assign data_o[14786] = data_o[2];
  assign data_o[14850] = data_o[2];
  assign data_o[14914] = data_o[2];
  assign data_o[14978] = data_o[2];
  assign data_o[15042] = data_o[2];
  assign data_o[15106] = data_o[2];
  assign data_o[15170] = data_o[2];
  assign data_o[15234] = data_o[2];
  assign data_o[15298] = data_o[2];
  assign data_o[15362] = data_o[2];
  assign data_o[15426] = data_o[2];
  assign data_o[15490] = data_o[2];
  assign data_o[15554] = data_o[2];
  assign data_o[15618] = data_o[2];
  assign data_o[15682] = data_o[2];
  assign data_o[15746] = data_o[2];
  assign data_o[15810] = data_o[2];
  assign data_o[15874] = data_o[2];
  assign data_o[15938] = data_o[2];
  assign data_o[16002] = data_o[2];
  assign data_o[16066] = data_o[2];
  assign data_o[16130] = data_o[2];
  assign data_o[16194] = data_o[2];
  assign data_o[16258] = data_o[2];
  assign data_o[16322] = data_o[2];
  assign data_o[16386] = data_o[2];
  assign data_o[16450] = data_o[2];
  assign data_o[16514] = data_o[2];
  assign data_o[16578] = data_o[2];
  assign data_o[16642] = data_o[2];
  assign data_o[16706] = data_o[2];
  assign data_o[16770] = data_o[2];
  assign data_o[16834] = data_o[2];
  assign data_o[16898] = data_o[2];
  assign data_o[16962] = data_o[2];
  assign data_o[17026] = data_o[2];
  assign data_o[17090] = data_o[2];
  assign data_o[17154] = data_o[2];
  assign data_o[17218] = data_o[2];
  assign data_o[17282] = data_o[2];
  assign data_o[17346] = data_o[2];
  assign data_o[17410] = data_o[2];
  assign data_o[17474] = data_o[2];
  assign data_o[17538] = data_o[2];
  assign data_o[17602] = data_o[2];
  assign data_o[17666] = data_o[2];
  assign data_o[17730] = data_o[2];
  assign data_o[17794] = data_o[2];
  assign data_o[17858] = data_o[2];
  assign data_o[17922] = data_o[2];
  assign data_o[17986] = data_o[2];
  assign data_o[18050] = data_o[2];
  assign data_o[18114] = data_o[2];
  assign data_o[18178] = data_o[2];
  assign data_o[18242] = data_o[2];
  assign data_o[18306] = data_o[2];
  assign data_o[18370] = data_o[2];
  assign data_o[18434] = data_o[2];
  assign data_o[18498] = data_o[2];
  assign data_o[18562] = data_o[2];
  assign data_o[18626] = data_o[2];
  assign data_o[18690] = data_o[2];
  assign data_o[18754] = data_o[2];
  assign data_o[18818] = data_o[2];
  assign data_o[18882] = data_o[2];
  assign data_o[18946] = data_o[2];
  assign data_o[19010] = data_o[2];
  assign data_o[19074] = data_o[2];
  assign data_o[19138] = data_o[2];
  assign data_o[19202] = data_o[2];
  assign data_o[19266] = data_o[2];
  assign data_o[19330] = data_o[2];
  assign data_o[19394] = data_o[2];
  assign data_o[19458] = data_o[2];
  assign data_o[19522] = data_o[2];
  assign data_o[19586] = data_o[2];
  assign data_o[19650] = data_o[2];
  assign data_o[19714] = data_o[2];
  assign data_o[19778] = data_o[2];
  assign data_o[19842] = data_o[2];
  assign data_o[19906] = data_o[2];
  assign data_o[19970] = data_o[2];
  assign data_o[20034] = data_o[2];
  assign data_o[20098] = data_o[2];
  assign data_o[20162] = data_o[2];
  assign data_o[20226] = data_o[2];
  assign data_o[20290] = data_o[2];
  assign data_o[20354] = data_o[2];
  assign data_o[20418] = data_o[2];
  assign data_o[20482] = data_o[2];
  assign data_o[20546] = data_o[2];
  assign data_o[20610] = data_o[2];
  assign data_o[20674] = data_o[2];
  assign data_o[20738] = data_o[2];
  assign data_o[20802] = data_o[2];
  assign data_o[20866] = data_o[2];
  assign data_o[20930] = data_o[2];
  assign data_o[20994] = data_o[2];
  assign data_o[21058] = data_o[2];
  assign data_o[21122] = data_o[2];
  assign data_o[21186] = data_o[2];
  assign data_o[21250] = data_o[2];
  assign data_o[21314] = data_o[2];
  assign data_o[21378] = data_o[2];
  assign data_o[21442] = data_o[2];
  assign data_o[21506] = data_o[2];
  assign data_o[21570] = data_o[2];
  assign data_o[21634] = data_o[2];
  assign data_o[21698] = data_o[2];
  assign data_o[21762] = data_o[2];
  assign data_o[21826] = data_o[2];
  assign data_o[21890] = data_o[2];
  assign data_o[21954] = data_o[2];
  assign data_o[22018] = data_o[2];
  assign data_o[22082] = data_o[2];
  assign data_o[22146] = data_o[2];
  assign data_o[22210] = data_o[2];
  assign data_o[22274] = data_o[2];
  assign data_o[22338] = data_o[2];
  assign data_o[22402] = data_o[2];
  assign data_o[22466] = data_o[2];
  assign data_o[22530] = data_o[2];
  assign data_o[22594] = data_o[2];
  assign data_o[22658] = data_o[2];
  assign data_o[22722] = data_o[2];
  assign data_o[22786] = data_o[2];
  assign data_o[22850] = data_o[2];
  assign data_o[22914] = data_o[2];
  assign data_o[22978] = data_o[2];
  assign data_o[23042] = data_o[2];
  assign data_o[23106] = data_o[2];
  assign data_o[23170] = data_o[2];
  assign data_o[23234] = data_o[2];
  assign data_o[23298] = data_o[2];
  assign data_o[23362] = data_o[2];
  assign data_o[23426] = data_o[2];
  assign data_o[23490] = data_o[2];
  assign data_o[23554] = data_o[2];
  assign data_o[23618] = data_o[2];
  assign data_o[23682] = data_o[2];
  assign data_o[23746] = data_o[2];
  assign data_o[23810] = data_o[2];
  assign data_o[23874] = data_o[2];
  assign data_o[23938] = data_o[2];
  assign data_o[24002] = data_o[2];
  assign data_o[24066] = data_o[2];
  assign data_o[24130] = data_o[2];
  assign data_o[24194] = data_o[2];
  assign data_o[24258] = data_o[2];
  assign data_o[24322] = data_o[2];
  assign data_o[24386] = data_o[2];
  assign data_o[24450] = data_o[2];
  assign data_o[24514] = data_o[2];
  assign data_o[24578] = data_o[2];
  assign data_o[24642] = data_o[2];
  assign data_o[24706] = data_o[2];
  assign data_o[24770] = data_o[2];
  assign data_o[24834] = data_o[2];
  assign data_o[24898] = data_o[2];
  assign data_o[24962] = data_o[2];
  assign data_o[25026] = data_o[2];
  assign data_o[25090] = data_o[2];
  assign data_o[25154] = data_o[2];
  assign data_o[25218] = data_o[2];
  assign data_o[25282] = data_o[2];
  assign data_o[25346] = data_o[2];
  assign data_o[25410] = data_o[2];
  assign data_o[25474] = data_o[2];
  assign data_o[25538] = data_o[2];
  assign data_o[25602] = data_o[2];
  assign data_o[25666] = data_o[2];
  assign data_o[25730] = data_o[2];
  assign data_o[25794] = data_o[2];
  assign data_o[25858] = data_o[2];
  assign data_o[25922] = data_o[2];
  assign data_o[25986] = data_o[2];
  assign data_o[26050] = data_o[2];
  assign data_o[26114] = data_o[2];
  assign data_o[26178] = data_o[2];
  assign data_o[26242] = data_o[2];
  assign data_o[26306] = data_o[2];
  assign data_o[26370] = data_o[2];
  assign data_o[26434] = data_o[2];
  assign data_o[26498] = data_o[2];
  assign data_o[26562] = data_o[2];
  assign data_o[26626] = data_o[2];
  assign data_o[26690] = data_o[2];
  assign data_o[26754] = data_o[2];
  assign data_o[26818] = data_o[2];
  assign data_o[26882] = data_o[2];
  assign data_o[26946] = data_o[2];
  assign data_o[27010] = data_o[2];
  assign data_o[27074] = data_o[2];
  assign data_o[27138] = data_o[2];
  assign data_o[27202] = data_o[2];
  assign data_o[27266] = data_o[2];
  assign data_o[27330] = data_o[2];
  assign data_o[27394] = data_o[2];
  assign data_o[27458] = data_o[2];
  assign data_o[27522] = data_o[2];
  assign data_o[27586] = data_o[2];
  assign data_o[27650] = data_o[2];
  assign data_o[27714] = data_o[2];
  assign data_o[27778] = data_o[2];
  assign data_o[27842] = data_o[2];
  assign data_o[27906] = data_o[2];
  assign data_o[27970] = data_o[2];
  assign data_o[28034] = data_o[2];
  assign data_o[28098] = data_o[2];
  assign data_o[28162] = data_o[2];
  assign data_o[28226] = data_o[2];
  assign data_o[28290] = data_o[2];
  assign data_o[28354] = data_o[2];
  assign data_o[28418] = data_o[2];
  assign data_o[28482] = data_o[2];
  assign data_o[28546] = data_o[2];
  assign data_o[28610] = data_o[2];
  assign data_o[28674] = data_o[2];
  assign data_o[28738] = data_o[2];
  assign data_o[28802] = data_o[2];
  assign data_o[28866] = data_o[2];
  assign data_o[28930] = data_o[2];
  assign data_o[28994] = data_o[2];
  assign data_o[29058] = data_o[2];
  assign data_o[29122] = data_o[2];
  assign data_o[29186] = data_o[2];
  assign data_o[29250] = data_o[2];
  assign data_o[29314] = data_o[2];
  assign data_o[29378] = data_o[2];
  assign data_o[29442] = data_o[2];
  assign data_o[29506] = data_o[2];
  assign data_o[29570] = data_o[2];
  assign data_o[29634] = data_o[2];
  assign data_o[29698] = data_o[2];
  assign data_o[29762] = data_o[2];
  assign data_o[29826] = data_o[2];
  assign data_o[29890] = data_o[2];
  assign data_o[29954] = data_o[2];
  assign data_o[30018] = data_o[2];
  assign data_o[30082] = data_o[2];
  assign data_o[30146] = data_o[2];
  assign data_o[30210] = data_o[2];
  assign data_o[30274] = data_o[2];
  assign data_o[30338] = data_o[2];
  assign data_o[30402] = data_o[2];
  assign data_o[30466] = data_o[2];
  assign data_o[30530] = data_o[2];
  assign data_o[30594] = data_o[2];
  assign data_o[30658] = data_o[2];
  assign data_o[30722] = data_o[2];
  assign data_o[30786] = data_o[2];
  assign data_o[30850] = data_o[2];
  assign data_o[30914] = data_o[2];
  assign data_o[30978] = data_o[2];
  assign data_o[31042] = data_o[2];
  assign data_o[31106] = data_o[2];
  assign data_o[31170] = data_o[2];
  assign data_o[31234] = data_o[2];
  assign data_o[31298] = data_o[2];
  assign data_o[31362] = data_o[2];
  assign data_o[31426] = data_o[2];
  assign data_o[31490] = data_o[2];
  assign data_o[31554] = data_o[2];
  assign data_o[31618] = data_o[2];
  assign data_o[31682] = data_o[2];
  assign data_o[31746] = data_o[2];
  assign data_o[31810] = data_o[2];
  assign data_o[31874] = data_o[2];
  assign data_o[31938] = data_o[2];
  assign data_o[65] = data_o[1];
  assign data_o[129] = data_o[1];
  assign data_o[193] = data_o[1];
  assign data_o[257] = data_o[1];
  assign data_o[321] = data_o[1];
  assign data_o[385] = data_o[1];
  assign data_o[449] = data_o[1];
  assign data_o[513] = data_o[1];
  assign data_o[577] = data_o[1];
  assign data_o[641] = data_o[1];
  assign data_o[705] = data_o[1];
  assign data_o[769] = data_o[1];
  assign data_o[833] = data_o[1];
  assign data_o[897] = data_o[1];
  assign data_o[961] = data_o[1];
  assign data_o[1025] = data_o[1];
  assign data_o[1089] = data_o[1];
  assign data_o[1153] = data_o[1];
  assign data_o[1217] = data_o[1];
  assign data_o[1281] = data_o[1];
  assign data_o[1345] = data_o[1];
  assign data_o[1409] = data_o[1];
  assign data_o[1473] = data_o[1];
  assign data_o[1537] = data_o[1];
  assign data_o[1601] = data_o[1];
  assign data_o[1665] = data_o[1];
  assign data_o[1729] = data_o[1];
  assign data_o[1793] = data_o[1];
  assign data_o[1857] = data_o[1];
  assign data_o[1921] = data_o[1];
  assign data_o[1985] = data_o[1];
  assign data_o[2049] = data_o[1];
  assign data_o[2113] = data_o[1];
  assign data_o[2177] = data_o[1];
  assign data_o[2241] = data_o[1];
  assign data_o[2305] = data_o[1];
  assign data_o[2369] = data_o[1];
  assign data_o[2433] = data_o[1];
  assign data_o[2497] = data_o[1];
  assign data_o[2561] = data_o[1];
  assign data_o[2625] = data_o[1];
  assign data_o[2689] = data_o[1];
  assign data_o[2753] = data_o[1];
  assign data_o[2817] = data_o[1];
  assign data_o[2881] = data_o[1];
  assign data_o[2945] = data_o[1];
  assign data_o[3009] = data_o[1];
  assign data_o[3073] = data_o[1];
  assign data_o[3137] = data_o[1];
  assign data_o[3201] = data_o[1];
  assign data_o[3265] = data_o[1];
  assign data_o[3329] = data_o[1];
  assign data_o[3393] = data_o[1];
  assign data_o[3457] = data_o[1];
  assign data_o[3521] = data_o[1];
  assign data_o[3585] = data_o[1];
  assign data_o[3649] = data_o[1];
  assign data_o[3713] = data_o[1];
  assign data_o[3777] = data_o[1];
  assign data_o[3841] = data_o[1];
  assign data_o[3905] = data_o[1];
  assign data_o[3969] = data_o[1];
  assign data_o[4033] = data_o[1];
  assign data_o[4097] = data_o[1];
  assign data_o[4161] = data_o[1];
  assign data_o[4225] = data_o[1];
  assign data_o[4289] = data_o[1];
  assign data_o[4353] = data_o[1];
  assign data_o[4417] = data_o[1];
  assign data_o[4481] = data_o[1];
  assign data_o[4545] = data_o[1];
  assign data_o[4609] = data_o[1];
  assign data_o[4673] = data_o[1];
  assign data_o[4737] = data_o[1];
  assign data_o[4801] = data_o[1];
  assign data_o[4865] = data_o[1];
  assign data_o[4929] = data_o[1];
  assign data_o[4993] = data_o[1];
  assign data_o[5057] = data_o[1];
  assign data_o[5121] = data_o[1];
  assign data_o[5185] = data_o[1];
  assign data_o[5249] = data_o[1];
  assign data_o[5313] = data_o[1];
  assign data_o[5377] = data_o[1];
  assign data_o[5441] = data_o[1];
  assign data_o[5505] = data_o[1];
  assign data_o[5569] = data_o[1];
  assign data_o[5633] = data_o[1];
  assign data_o[5697] = data_o[1];
  assign data_o[5761] = data_o[1];
  assign data_o[5825] = data_o[1];
  assign data_o[5889] = data_o[1];
  assign data_o[5953] = data_o[1];
  assign data_o[6017] = data_o[1];
  assign data_o[6081] = data_o[1];
  assign data_o[6145] = data_o[1];
  assign data_o[6209] = data_o[1];
  assign data_o[6273] = data_o[1];
  assign data_o[6337] = data_o[1];
  assign data_o[6401] = data_o[1];
  assign data_o[6465] = data_o[1];
  assign data_o[6529] = data_o[1];
  assign data_o[6593] = data_o[1];
  assign data_o[6657] = data_o[1];
  assign data_o[6721] = data_o[1];
  assign data_o[6785] = data_o[1];
  assign data_o[6849] = data_o[1];
  assign data_o[6913] = data_o[1];
  assign data_o[6977] = data_o[1];
  assign data_o[7041] = data_o[1];
  assign data_o[7105] = data_o[1];
  assign data_o[7169] = data_o[1];
  assign data_o[7233] = data_o[1];
  assign data_o[7297] = data_o[1];
  assign data_o[7361] = data_o[1];
  assign data_o[7425] = data_o[1];
  assign data_o[7489] = data_o[1];
  assign data_o[7553] = data_o[1];
  assign data_o[7617] = data_o[1];
  assign data_o[7681] = data_o[1];
  assign data_o[7745] = data_o[1];
  assign data_o[7809] = data_o[1];
  assign data_o[7873] = data_o[1];
  assign data_o[7937] = data_o[1];
  assign data_o[8001] = data_o[1];
  assign data_o[8065] = data_o[1];
  assign data_o[8129] = data_o[1];
  assign data_o[8193] = data_o[1];
  assign data_o[8257] = data_o[1];
  assign data_o[8321] = data_o[1];
  assign data_o[8385] = data_o[1];
  assign data_o[8449] = data_o[1];
  assign data_o[8513] = data_o[1];
  assign data_o[8577] = data_o[1];
  assign data_o[8641] = data_o[1];
  assign data_o[8705] = data_o[1];
  assign data_o[8769] = data_o[1];
  assign data_o[8833] = data_o[1];
  assign data_o[8897] = data_o[1];
  assign data_o[8961] = data_o[1];
  assign data_o[9025] = data_o[1];
  assign data_o[9089] = data_o[1];
  assign data_o[9153] = data_o[1];
  assign data_o[9217] = data_o[1];
  assign data_o[9281] = data_o[1];
  assign data_o[9345] = data_o[1];
  assign data_o[9409] = data_o[1];
  assign data_o[9473] = data_o[1];
  assign data_o[9537] = data_o[1];
  assign data_o[9601] = data_o[1];
  assign data_o[9665] = data_o[1];
  assign data_o[9729] = data_o[1];
  assign data_o[9793] = data_o[1];
  assign data_o[9857] = data_o[1];
  assign data_o[9921] = data_o[1];
  assign data_o[9985] = data_o[1];
  assign data_o[10049] = data_o[1];
  assign data_o[10113] = data_o[1];
  assign data_o[10177] = data_o[1];
  assign data_o[10241] = data_o[1];
  assign data_o[10305] = data_o[1];
  assign data_o[10369] = data_o[1];
  assign data_o[10433] = data_o[1];
  assign data_o[10497] = data_o[1];
  assign data_o[10561] = data_o[1];
  assign data_o[10625] = data_o[1];
  assign data_o[10689] = data_o[1];
  assign data_o[10753] = data_o[1];
  assign data_o[10817] = data_o[1];
  assign data_o[10881] = data_o[1];
  assign data_o[10945] = data_o[1];
  assign data_o[11009] = data_o[1];
  assign data_o[11073] = data_o[1];
  assign data_o[11137] = data_o[1];
  assign data_o[11201] = data_o[1];
  assign data_o[11265] = data_o[1];
  assign data_o[11329] = data_o[1];
  assign data_o[11393] = data_o[1];
  assign data_o[11457] = data_o[1];
  assign data_o[11521] = data_o[1];
  assign data_o[11585] = data_o[1];
  assign data_o[11649] = data_o[1];
  assign data_o[11713] = data_o[1];
  assign data_o[11777] = data_o[1];
  assign data_o[11841] = data_o[1];
  assign data_o[11905] = data_o[1];
  assign data_o[11969] = data_o[1];
  assign data_o[12033] = data_o[1];
  assign data_o[12097] = data_o[1];
  assign data_o[12161] = data_o[1];
  assign data_o[12225] = data_o[1];
  assign data_o[12289] = data_o[1];
  assign data_o[12353] = data_o[1];
  assign data_o[12417] = data_o[1];
  assign data_o[12481] = data_o[1];
  assign data_o[12545] = data_o[1];
  assign data_o[12609] = data_o[1];
  assign data_o[12673] = data_o[1];
  assign data_o[12737] = data_o[1];
  assign data_o[12801] = data_o[1];
  assign data_o[12865] = data_o[1];
  assign data_o[12929] = data_o[1];
  assign data_o[12993] = data_o[1];
  assign data_o[13057] = data_o[1];
  assign data_o[13121] = data_o[1];
  assign data_o[13185] = data_o[1];
  assign data_o[13249] = data_o[1];
  assign data_o[13313] = data_o[1];
  assign data_o[13377] = data_o[1];
  assign data_o[13441] = data_o[1];
  assign data_o[13505] = data_o[1];
  assign data_o[13569] = data_o[1];
  assign data_o[13633] = data_o[1];
  assign data_o[13697] = data_o[1];
  assign data_o[13761] = data_o[1];
  assign data_o[13825] = data_o[1];
  assign data_o[13889] = data_o[1];
  assign data_o[13953] = data_o[1];
  assign data_o[14017] = data_o[1];
  assign data_o[14081] = data_o[1];
  assign data_o[14145] = data_o[1];
  assign data_o[14209] = data_o[1];
  assign data_o[14273] = data_o[1];
  assign data_o[14337] = data_o[1];
  assign data_o[14401] = data_o[1];
  assign data_o[14465] = data_o[1];
  assign data_o[14529] = data_o[1];
  assign data_o[14593] = data_o[1];
  assign data_o[14657] = data_o[1];
  assign data_o[14721] = data_o[1];
  assign data_o[14785] = data_o[1];
  assign data_o[14849] = data_o[1];
  assign data_o[14913] = data_o[1];
  assign data_o[14977] = data_o[1];
  assign data_o[15041] = data_o[1];
  assign data_o[15105] = data_o[1];
  assign data_o[15169] = data_o[1];
  assign data_o[15233] = data_o[1];
  assign data_o[15297] = data_o[1];
  assign data_o[15361] = data_o[1];
  assign data_o[15425] = data_o[1];
  assign data_o[15489] = data_o[1];
  assign data_o[15553] = data_o[1];
  assign data_o[15617] = data_o[1];
  assign data_o[15681] = data_o[1];
  assign data_o[15745] = data_o[1];
  assign data_o[15809] = data_o[1];
  assign data_o[15873] = data_o[1];
  assign data_o[15937] = data_o[1];
  assign data_o[16001] = data_o[1];
  assign data_o[16065] = data_o[1];
  assign data_o[16129] = data_o[1];
  assign data_o[16193] = data_o[1];
  assign data_o[16257] = data_o[1];
  assign data_o[16321] = data_o[1];
  assign data_o[16385] = data_o[1];
  assign data_o[16449] = data_o[1];
  assign data_o[16513] = data_o[1];
  assign data_o[16577] = data_o[1];
  assign data_o[16641] = data_o[1];
  assign data_o[16705] = data_o[1];
  assign data_o[16769] = data_o[1];
  assign data_o[16833] = data_o[1];
  assign data_o[16897] = data_o[1];
  assign data_o[16961] = data_o[1];
  assign data_o[17025] = data_o[1];
  assign data_o[17089] = data_o[1];
  assign data_o[17153] = data_o[1];
  assign data_o[17217] = data_o[1];
  assign data_o[17281] = data_o[1];
  assign data_o[17345] = data_o[1];
  assign data_o[17409] = data_o[1];
  assign data_o[17473] = data_o[1];
  assign data_o[17537] = data_o[1];
  assign data_o[17601] = data_o[1];
  assign data_o[17665] = data_o[1];
  assign data_o[17729] = data_o[1];
  assign data_o[17793] = data_o[1];
  assign data_o[17857] = data_o[1];
  assign data_o[17921] = data_o[1];
  assign data_o[17985] = data_o[1];
  assign data_o[18049] = data_o[1];
  assign data_o[18113] = data_o[1];
  assign data_o[18177] = data_o[1];
  assign data_o[18241] = data_o[1];
  assign data_o[18305] = data_o[1];
  assign data_o[18369] = data_o[1];
  assign data_o[18433] = data_o[1];
  assign data_o[18497] = data_o[1];
  assign data_o[18561] = data_o[1];
  assign data_o[18625] = data_o[1];
  assign data_o[18689] = data_o[1];
  assign data_o[18753] = data_o[1];
  assign data_o[18817] = data_o[1];
  assign data_o[18881] = data_o[1];
  assign data_o[18945] = data_o[1];
  assign data_o[19009] = data_o[1];
  assign data_o[19073] = data_o[1];
  assign data_o[19137] = data_o[1];
  assign data_o[19201] = data_o[1];
  assign data_o[19265] = data_o[1];
  assign data_o[19329] = data_o[1];
  assign data_o[19393] = data_o[1];
  assign data_o[19457] = data_o[1];
  assign data_o[19521] = data_o[1];
  assign data_o[19585] = data_o[1];
  assign data_o[19649] = data_o[1];
  assign data_o[19713] = data_o[1];
  assign data_o[19777] = data_o[1];
  assign data_o[19841] = data_o[1];
  assign data_o[19905] = data_o[1];
  assign data_o[19969] = data_o[1];
  assign data_o[20033] = data_o[1];
  assign data_o[20097] = data_o[1];
  assign data_o[20161] = data_o[1];
  assign data_o[20225] = data_o[1];
  assign data_o[20289] = data_o[1];
  assign data_o[20353] = data_o[1];
  assign data_o[20417] = data_o[1];
  assign data_o[20481] = data_o[1];
  assign data_o[20545] = data_o[1];
  assign data_o[20609] = data_o[1];
  assign data_o[20673] = data_o[1];
  assign data_o[20737] = data_o[1];
  assign data_o[20801] = data_o[1];
  assign data_o[20865] = data_o[1];
  assign data_o[20929] = data_o[1];
  assign data_o[20993] = data_o[1];
  assign data_o[21057] = data_o[1];
  assign data_o[21121] = data_o[1];
  assign data_o[21185] = data_o[1];
  assign data_o[21249] = data_o[1];
  assign data_o[21313] = data_o[1];
  assign data_o[21377] = data_o[1];
  assign data_o[21441] = data_o[1];
  assign data_o[21505] = data_o[1];
  assign data_o[21569] = data_o[1];
  assign data_o[21633] = data_o[1];
  assign data_o[21697] = data_o[1];
  assign data_o[21761] = data_o[1];
  assign data_o[21825] = data_o[1];
  assign data_o[21889] = data_o[1];
  assign data_o[21953] = data_o[1];
  assign data_o[22017] = data_o[1];
  assign data_o[22081] = data_o[1];
  assign data_o[22145] = data_o[1];
  assign data_o[22209] = data_o[1];
  assign data_o[22273] = data_o[1];
  assign data_o[22337] = data_o[1];
  assign data_o[22401] = data_o[1];
  assign data_o[22465] = data_o[1];
  assign data_o[22529] = data_o[1];
  assign data_o[22593] = data_o[1];
  assign data_o[22657] = data_o[1];
  assign data_o[22721] = data_o[1];
  assign data_o[22785] = data_o[1];
  assign data_o[22849] = data_o[1];
  assign data_o[22913] = data_o[1];
  assign data_o[22977] = data_o[1];
  assign data_o[23041] = data_o[1];
  assign data_o[23105] = data_o[1];
  assign data_o[23169] = data_o[1];
  assign data_o[23233] = data_o[1];
  assign data_o[23297] = data_o[1];
  assign data_o[23361] = data_o[1];
  assign data_o[23425] = data_o[1];
  assign data_o[23489] = data_o[1];
  assign data_o[23553] = data_o[1];
  assign data_o[23617] = data_o[1];
  assign data_o[23681] = data_o[1];
  assign data_o[23745] = data_o[1];
  assign data_o[23809] = data_o[1];
  assign data_o[23873] = data_o[1];
  assign data_o[23937] = data_o[1];
  assign data_o[24001] = data_o[1];
  assign data_o[24065] = data_o[1];
  assign data_o[24129] = data_o[1];
  assign data_o[24193] = data_o[1];
  assign data_o[24257] = data_o[1];
  assign data_o[24321] = data_o[1];
  assign data_o[24385] = data_o[1];
  assign data_o[24449] = data_o[1];
  assign data_o[24513] = data_o[1];
  assign data_o[24577] = data_o[1];
  assign data_o[24641] = data_o[1];
  assign data_o[24705] = data_o[1];
  assign data_o[24769] = data_o[1];
  assign data_o[24833] = data_o[1];
  assign data_o[24897] = data_o[1];
  assign data_o[24961] = data_o[1];
  assign data_o[25025] = data_o[1];
  assign data_o[25089] = data_o[1];
  assign data_o[25153] = data_o[1];
  assign data_o[25217] = data_o[1];
  assign data_o[25281] = data_o[1];
  assign data_o[25345] = data_o[1];
  assign data_o[25409] = data_o[1];
  assign data_o[25473] = data_o[1];
  assign data_o[25537] = data_o[1];
  assign data_o[25601] = data_o[1];
  assign data_o[25665] = data_o[1];
  assign data_o[25729] = data_o[1];
  assign data_o[25793] = data_o[1];
  assign data_o[25857] = data_o[1];
  assign data_o[25921] = data_o[1];
  assign data_o[25985] = data_o[1];
  assign data_o[26049] = data_o[1];
  assign data_o[26113] = data_o[1];
  assign data_o[26177] = data_o[1];
  assign data_o[26241] = data_o[1];
  assign data_o[26305] = data_o[1];
  assign data_o[26369] = data_o[1];
  assign data_o[26433] = data_o[1];
  assign data_o[26497] = data_o[1];
  assign data_o[26561] = data_o[1];
  assign data_o[26625] = data_o[1];
  assign data_o[26689] = data_o[1];
  assign data_o[26753] = data_o[1];
  assign data_o[26817] = data_o[1];
  assign data_o[26881] = data_o[1];
  assign data_o[26945] = data_o[1];
  assign data_o[27009] = data_o[1];
  assign data_o[27073] = data_o[1];
  assign data_o[27137] = data_o[1];
  assign data_o[27201] = data_o[1];
  assign data_o[27265] = data_o[1];
  assign data_o[27329] = data_o[1];
  assign data_o[27393] = data_o[1];
  assign data_o[27457] = data_o[1];
  assign data_o[27521] = data_o[1];
  assign data_o[27585] = data_o[1];
  assign data_o[27649] = data_o[1];
  assign data_o[27713] = data_o[1];
  assign data_o[27777] = data_o[1];
  assign data_o[27841] = data_o[1];
  assign data_o[27905] = data_o[1];
  assign data_o[27969] = data_o[1];
  assign data_o[28033] = data_o[1];
  assign data_o[28097] = data_o[1];
  assign data_o[28161] = data_o[1];
  assign data_o[28225] = data_o[1];
  assign data_o[28289] = data_o[1];
  assign data_o[28353] = data_o[1];
  assign data_o[28417] = data_o[1];
  assign data_o[28481] = data_o[1];
  assign data_o[28545] = data_o[1];
  assign data_o[28609] = data_o[1];
  assign data_o[28673] = data_o[1];
  assign data_o[28737] = data_o[1];
  assign data_o[28801] = data_o[1];
  assign data_o[28865] = data_o[1];
  assign data_o[28929] = data_o[1];
  assign data_o[28993] = data_o[1];
  assign data_o[29057] = data_o[1];
  assign data_o[29121] = data_o[1];
  assign data_o[29185] = data_o[1];
  assign data_o[29249] = data_o[1];
  assign data_o[29313] = data_o[1];
  assign data_o[29377] = data_o[1];
  assign data_o[29441] = data_o[1];
  assign data_o[29505] = data_o[1];
  assign data_o[29569] = data_o[1];
  assign data_o[29633] = data_o[1];
  assign data_o[29697] = data_o[1];
  assign data_o[29761] = data_o[1];
  assign data_o[29825] = data_o[1];
  assign data_o[29889] = data_o[1];
  assign data_o[29953] = data_o[1];
  assign data_o[30017] = data_o[1];
  assign data_o[30081] = data_o[1];
  assign data_o[30145] = data_o[1];
  assign data_o[30209] = data_o[1];
  assign data_o[30273] = data_o[1];
  assign data_o[30337] = data_o[1];
  assign data_o[30401] = data_o[1];
  assign data_o[30465] = data_o[1];
  assign data_o[30529] = data_o[1];
  assign data_o[30593] = data_o[1];
  assign data_o[30657] = data_o[1];
  assign data_o[30721] = data_o[1];
  assign data_o[30785] = data_o[1];
  assign data_o[30849] = data_o[1];
  assign data_o[30913] = data_o[1];
  assign data_o[30977] = data_o[1];
  assign data_o[31041] = data_o[1];
  assign data_o[31105] = data_o[1];
  assign data_o[31169] = data_o[1];
  assign data_o[31233] = data_o[1];
  assign data_o[31297] = data_o[1];
  assign data_o[31361] = data_o[1];
  assign data_o[31425] = data_o[1];
  assign data_o[31489] = data_o[1];
  assign data_o[31553] = data_o[1];
  assign data_o[31617] = data_o[1];
  assign data_o[31681] = data_o[1];
  assign data_o[31745] = data_o[1];
  assign data_o[31809] = data_o[1];
  assign data_o[31873] = data_o[1];
  assign data_o[31937] = data_o[1];
  assign data_o[64] = data_o[0];
  assign data_o[128] = data_o[0];
  assign data_o[192] = data_o[0];
  assign data_o[256] = data_o[0];
  assign data_o[320] = data_o[0];
  assign data_o[384] = data_o[0];
  assign data_o[448] = data_o[0];
  assign data_o[512] = data_o[0];
  assign data_o[576] = data_o[0];
  assign data_o[640] = data_o[0];
  assign data_o[704] = data_o[0];
  assign data_o[768] = data_o[0];
  assign data_o[832] = data_o[0];
  assign data_o[896] = data_o[0];
  assign data_o[960] = data_o[0];
  assign data_o[1024] = data_o[0];
  assign data_o[1088] = data_o[0];
  assign data_o[1152] = data_o[0];
  assign data_o[1216] = data_o[0];
  assign data_o[1280] = data_o[0];
  assign data_o[1344] = data_o[0];
  assign data_o[1408] = data_o[0];
  assign data_o[1472] = data_o[0];
  assign data_o[1536] = data_o[0];
  assign data_o[1600] = data_o[0];
  assign data_o[1664] = data_o[0];
  assign data_o[1728] = data_o[0];
  assign data_o[1792] = data_o[0];
  assign data_o[1856] = data_o[0];
  assign data_o[1920] = data_o[0];
  assign data_o[1984] = data_o[0];
  assign data_o[2048] = data_o[0];
  assign data_o[2112] = data_o[0];
  assign data_o[2176] = data_o[0];
  assign data_o[2240] = data_o[0];
  assign data_o[2304] = data_o[0];
  assign data_o[2368] = data_o[0];
  assign data_o[2432] = data_o[0];
  assign data_o[2496] = data_o[0];
  assign data_o[2560] = data_o[0];
  assign data_o[2624] = data_o[0];
  assign data_o[2688] = data_o[0];
  assign data_o[2752] = data_o[0];
  assign data_o[2816] = data_o[0];
  assign data_o[2880] = data_o[0];
  assign data_o[2944] = data_o[0];
  assign data_o[3008] = data_o[0];
  assign data_o[3072] = data_o[0];
  assign data_o[3136] = data_o[0];
  assign data_o[3200] = data_o[0];
  assign data_o[3264] = data_o[0];
  assign data_o[3328] = data_o[0];
  assign data_o[3392] = data_o[0];
  assign data_o[3456] = data_o[0];
  assign data_o[3520] = data_o[0];
  assign data_o[3584] = data_o[0];
  assign data_o[3648] = data_o[0];
  assign data_o[3712] = data_o[0];
  assign data_o[3776] = data_o[0];
  assign data_o[3840] = data_o[0];
  assign data_o[3904] = data_o[0];
  assign data_o[3968] = data_o[0];
  assign data_o[4032] = data_o[0];
  assign data_o[4096] = data_o[0];
  assign data_o[4160] = data_o[0];
  assign data_o[4224] = data_o[0];
  assign data_o[4288] = data_o[0];
  assign data_o[4352] = data_o[0];
  assign data_o[4416] = data_o[0];
  assign data_o[4480] = data_o[0];
  assign data_o[4544] = data_o[0];
  assign data_o[4608] = data_o[0];
  assign data_o[4672] = data_o[0];
  assign data_o[4736] = data_o[0];
  assign data_o[4800] = data_o[0];
  assign data_o[4864] = data_o[0];
  assign data_o[4928] = data_o[0];
  assign data_o[4992] = data_o[0];
  assign data_o[5056] = data_o[0];
  assign data_o[5120] = data_o[0];
  assign data_o[5184] = data_o[0];
  assign data_o[5248] = data_o[0];
  assign data_o[5312] = data_o[0];
  assign data_o[5376] = data_o[0];
  assign data_o[5440] = data_o[0];
  assign data_o[5504] = data_o[0];
  assign data_o[5568] = data_o[0];
  assign data_o[5632] = data_o[0];
  assign data_o[5696] = data_o[0];
  assign data_o[5760] = data_o[0];
  assign data_o[5824] = data_o[0];
  assign data_o[5888] = data_o[0];
  assign data_o[5952] = data_o[0];
  assign data_o[6016] = data_o[0];
  assign data_o[6080] = data_o[0];
  assign data_o[6144] = data_o[0];
  assign data_o[6208] = data_o[0];
  assign data_o[6272] = data_o[0];
  assign data_o[6336] = data_o[0];
  assign data_o[6400] = data_o[0];
  assign data_o[6464] = data_o[0];
  assign data_o[6528] = data_o[0];
  assign data_o[6592] = data_o[0];
  assign data_o[6656] = data_o[0];
  assign data_o[6720] = data_o[0];
  assign data_o[6784] = data_o[0];
  assign data_o[6848] = data_o[0];
  assign data_o[6912] = data_o[0];
  assign data_o[6976] = data_o[0];
  assign data_o[7040] = data_o[0];
  assign data_o[7104] = data_o[0];
  assign data_o[7168] = data_o[0];
  assign data_o[7232] = data_o[0];
  assign data_o[7296] = data_o[0];
  assign data_o[7360] = data_o[0];
  assign data_o[7424] = data_o[0];
  assign data_o[7488] = data_o[0];
  assign data_o[7552] = data_o[0];
  assign data_o[7616] = data_o[0];
  assign data_o[7680] = data_o[0];
  assign data_o[7744] = data_o[0];
  assign data_o[7808] = data_o[0];
  assign data_o[7872] = data_o[0];
  assign data_o[7936] = data_o[0];
  assign data_o[8000] = data_o[0];
  assign data_o[8064] = data_o[0];
  assign data_o[8128] = data_o[0];
  assign data_o[8192] = data_o[0];
  assign data_o[8256] = data_o[0];
  assign data_o[8320] = data_o[0];
  assign data_o[8384] = data_o[0];
  assign data_o[8448] = data_o[0];
  assign data_o[8512] = data_o[0];
  assign data_o[8576] = data_o[0];
  assign data_o[8640] = data_o[0];
  assign data_o[8704] = data_o[0];
  assign data_o[8768] = data_o[0];
  assign data_o[8832] = data_o[0];
  assign data_o[8896] = data_o[0];
  assign data_o[8960] = data_o[0];
  assign data_o[9024] = data_o[0];
  assign data_o[9088] = data_o[0];
  assign data_o[9152] = data_o[0];
  assign data_o[9216] = data_o[0];
  assign data_o[9280] = data_o[0];
  assign data_o[9344] = data_o[0];
  assign data_o[9408] = data_o[0];
  assign data_o[9472] = data_o[0];
  assign data_o[9536] = data_o[0];
  assign data_o[9600] = data_o[0];
  assign data_o[9664] = data_o[0];
  assign data_o[9728] = data_o[0];
  assign data_o[9792] = data_o[0];
  assign data_o[9856] = data_o[0];
  assign data_o[9920] = data_o[0];
  assign data_o[9984] = data_o[0];
  assign data_o[10048] = data_o[0];
  assign data_o[10112] = data_o[0];
  assign data_o[10176] = data_o[0];
  assign data_o[10240] = data_o[0];
  assign data_o[10304] = data_o[0];
  assign data_o[10368] = data_o[0];
  assign data_o[10432] = data_o[0];
  assign data_o[10496] = data_o[0];
  assign data_o[10560] = data_o[0];
  assign data_o[10624] = data_o[0];
  assign data_o[10688] = data_o[0];
  assign data_o[10752] = data_o[0];
  assign data_o[10816] = data_o[0];
  assign data_o[10880] = data_o[0];
  assign data_o[10944] = data_o[0];
  assign data_o[11008] = data_o[0];
  assign data_o[11072] = data_o[0];
  assign data_o[11136] = data_o[0];
  assign data_o[11200] = data_o[0];
  assign data_o[11264] = data_o[0];
  assign data_o[11328] = data_o[0];
  assign data_o[11392] = data_o[0];
  assign data_o[11456] = data_o[0];
  assign data_o[11520] = data_o[0];
  assign data_o[11584] = data_o[0];
  assign data_o[11648] = data_o[0];
  assign data_o[11712] = data_o[0];
  assign data_o[11776] = data_o[0];
  assign data_o[11840] = data_o[0];
  assign data_o[11904] = data_o[0];
  assign data_o[11968] = data_o[0];
  assign data_o[12032] = data_o[0];
  assign data_o[12096] = data_o[0];
  assign data_o[12160] = data_o[0];
  assign data_o[12224] = data_o[0];
  assign data_o[12288] = data_o[0];
  assign data_o[12352] = data_o[0];
  assign data_o[12416] = data_o[0];
  assign data_o[12480] = data_o[0];
  assign data_o[12544] = data_o[0];
  assign data_o[12608] = data_o[0];
  assign data_o[12672] = data_o[0];
  assign data_o[12736] = data_o[0];
  assign data_o[12800] = data_o[0];
  assign data_o[12864] = data_o[0];
  assign data_o[12928] = data_o[0];
  assign data_o[12992] = data_o[0];
  assign data_o[13056] = data_o[0];
  assign data_o[13120] = data_o[0];
  assign data_o[13184] = data_o[0];
  assign data_o[13248] = data_o[0];
  assign data_o[13312] = data_o[0];
  assign data_o[13376] = data_o[0];
  assign data_o[13440] = data_o[0];
  assign data_o[13504] = data_o[0];
  assign data_o[13568] = data_o[0];
  assign data_o[13632] = data_o[0];
  assign data_o[13696] = data_o[0];
  assign data_o[13760] = data_o[0];
  assign data_o[13824] = data_o[0];
  assign data_o[13888] = data_o[0];
  assign data_o[13952] = data_o[0];
  assign data_o[14016] = data_o[0];
  assign data_o[14080] = data_o[0];
  assign data_o[14144] = data_o[0];
  assign data_o[14208] = data_o[0];
  assign data_o[14272] = data_o[0];
  assign data_o[14336] = data_o[0];
  assign data_o[14400] = data_o[0];
  assign data_o[14464] = data_o[0];
  assign data_o[14528] = data_o[0];
  assign data_o[14592] = data_o[0];
  assign data_o[14656] = data_o[0];
  assign data_o[14720] = data_o[0];
  assign data_o[14784] = data_o[0];
  assign data_o[14848] = data_o[0];
  assign data_o[14912] = data_o[0];
  assign data_o[14976] = data_o[0];
  assign data_o[15040] = data_o[0];
  assign data_o[15104] = data_o[0];
  assign data_o[15168] = data_o[0];
  assign data_o[15232] = data_o[0];
  assign data_o[15296] = data_o[0];
  assign data_o[15360] = data_o[0];
  assign data_o[15424] = data_o[0];
  assign data_o[15488] = data_o[0];
  assign data_o[15552] = data_o[0];
  assign data_o[15616] = data_o[0];
  assign data_o[15680] = data_o[0];
  assign data_o[15744] = data_o[0];
  assign data_o[15808] = data_o[0];
  assign data_o[15872] = data_o[0];
  assign data_o[15936] = data_o[0];
  assign data_o[16000] = data_o[0];
  assign data_o[16064] = data_o[0];
  assign data_o[16128] = data_o[0];
  assign data_o[16192] = data_o[0];
  assign data_o[16256] = data_o[0];
  assign data_o[16320] = data_o[0];
  assign data_o[16384] = data_o[0];
  assign data_o[16448] = data_o[0];
  assign data_o[16512] = data_o[0];
  assign data_o[16576] = data_o[0];
  assign data_o[16640] = data_o[0];
  assign data_o[16704] = data_o[0];
  assign data_o[16768] = data_o[0];
  assign data_o[16832] = data_o[0];
  assign data_o[16896] = data_o[0];
  assign data_o[16960] = data_o[0];
  assign data_o[17024] = data_o[0];
  assign data_o[17088] = data_o[0];
  assign data_o[17152] = data_o[0];
  assign data_o[17216] = data_o[0];
  assign data_o[17280] = data_o[0];
  assign data_o[17344] = data_o[0];
  assign data_o[17408] = data_o[0];
  assign data_o[17472] = data_o[0];
  assign data_o[17536] = data_o[0];
  assign data_o[17600] = data_o[0];
  assign data_o[17664] = data_o[0];
  assign data_o[17728] = data_o[0];
  assign data_o[17792] = data_o[0];
  assign data_o[17856] = data_o[0];
  assign data_o[17920] = data_o[0];
  assign data_o[17984] = data_o[0];
  assign data_o[18048] = data_o[0];
  assign data_o[18112] = data_o[0];
  assign data_o[18176] = data_o[0];
  assign data_o[18240] = data_o[0];
  assign data_o[18304] = data_o[0];
  assign data_o[18368] = data_o[0];
  assign data_o[18432] = data_o[0];
  assign data_o[18496] = data_o[0];
  assign data_o[18560] = data_o[0];
  assign data_o[18624] = data_o[0];
  assign data_o[18688] = data_o[0];
  assign data_o[18752] = data_o[0];
  assign data_o[18816] = data_o[0];
  assign data_o[18880] = data_o[0];
  assign data_o[18944] = data_o[0];
  assign data_o[19008] = data_o[0];
  assign data_o[19072] = data_o[0];
  assign data_o[19136] = data_o[0];
  assign data_o[19200] = data_o[0];
  assign data_o[19264] = data_o[0];
  assign data_o[19328] = data_o[0];
  assign data_o[19392] = data_o[0];
  assign data_o[19456] = data_o[0];
  assign data_o[19520] = data_o[0];
  assign data_o[19584] = data_o[0];
  assign data_o[19648] = data_o[0];
  assign data_o[19712] = data_o[0];
  assign data_o[19776] = data_o[0];
  assign data_o[19840] = data_o[0];
  assign data_o[19904] = data_o[0];
  assign data_o[19968] = data_o[0];
  assign data_o[20032] = data_o[0];
  assign data_o[20096] = data_o[0];
  assign data_o[20160] = data_o[0];
  assign data_o[20224] = data_o[0];
  assign data_o[20288] = data_o[0];
  assign data_o[20352] = data_o[0];
  assign data_o[20416] = data_o[0];
  assign data_o[20480] = data_o[0];
  assign data_o[20544] = data_o[0];
  assign data_o[20608] = data_o[0];
  assign data_o[20672] = data_o[0];
  assign data_o[20736] = data_o[0];
  assign data_o[20800] = data_o[0];
  assign data_o[20864] = data_o[0];
  assign data_o[20928] = data_o[0];
  assign data_o[20992] = data_o[0];
  assign data_o[21056] = data_o[0];
  assign data_o[21120] = data_o[0];
  assign data_o[21184] = data_o[0];
  assign data_o[21248] = data_o[0];
  assign data_o[21312] = data_o[0];
  assign data_o[21376] = data_o[0];
  assign data_o[21440] = data_o[0];
  assign data_o[21504] = data_o[0];
  assign data_o[21568] = data_o[0];
  assign data_o[21632] = data_o[0];
  assign data_o[21696] = data_o[0];
  assign data_o[21760] = data_o[0];
  assign data_o[21824] = data_o[0];
  assign data_o[21888] = data_o[0];
  assign data_o[21952] = data_o[0];
  assign data_o[22016] = data_o[0];
  assign data_o[22080] = data_o[0];
  assign data_o[22144] = data_o[0];
  assign data_o[22208] = data_o[0];
  assign data_o[22272] = data_o[0];
  assign data_o[22336] = data_o[0];
  assign data_o[22400] = data_o[0];
  assign data_o[22464] = data_o[0];
  assign data_o[22528] = data_o[0];
  assign data_o[22592] = data_o[0];
  assign data_o[22656] = data_o[0];
  assign data_o[22720] = data_o[0];
  assign data_o[22784] = data_o[0];
  assign data_o[22848] = data_o[0];
  assign data_o[22912] = data_o[0];
  assign data_o[22976] = data_o[0];
  assign data_o[23040] = data_o[0];
  assign data_o[23104] = data_o[0];
  assign data_o[23168] = data_o[0];
  assign data_o[23232] = data_o[0];
  assign data_o[23296] = data_o[0];
  assign data_o[23360] = data_o[0];
  assign data_o[23424] = data_o[0];
  assign data_o[23488] = data_o[0];
  assign data_o[23552] = data_o[0];
  assign data_o[23616] = data_o[0];
  assign data_o[23680] = data_o[0];
  assign data_o[23744] = data_o[0];
  assign data_o[23808] = data_o[0];
  assign data_o[23872] = data_o[0];
  assign data_o[23936] = data_o[0];
  assign data_o[24000] = data_o[0];
  assign data_o[24064] = data_o[0];
  assign data_o[24128] = data_o[0];
  assign data_o[24192] = data_o[0];
  assign data_o[24256] = data_o[0];
  assign data_o[24320] = data_o[0];
  assign data_o[24384] = data_o[0];
  assign data_o[24448] = data_o[0];
  assign data_o[24512] = data_o[0];
  assign data_o[24576] = data_o[0];
  assign data_o[24640] = data_o[0];
  assign data_o[24704] = data_o[0];
  assign data_o[24768] = data_o[0];
  assign data_o[24832] = data_o[0];
  assign data_o[24896] = data_o[0];
  assign data_o[24960] = data_o[0];
  assign data_o[25024] = data_o[0];
  assign data_o[25088] = data_o[0];
  assign data_o[25152] = data_o[0];
  assign data_o[25216] = data_o[0];
  assign data_o[25280] = data_o[0];
  assign data_o[25344] = data_o[0];
  assign data_o[25408] = data_o[0];
  assign data_o[25472] = data_o[0];
  assign data_o[25536] = data_o[0];
  assign data_o[25600] = data_o[0];
  assign data_o[25664] = data_o[0];
  assign data_o[25728] = data_o[0];
  assign data_o[25792] = data_o[0];
  assign data_o[25856] = data_o[0];
  assign data_o[25920] = data_o[0];
  assign data_o[25984] = data_o[0];
  assign data_o[26048] = data_o[0];
  assign data_o[26112] = data_o[0];
  assign data_o[26176] = data_o[0];
  assign data_o[26240] = data_o[0];
  assign data_o[26304] = data_o[0];
  assign data_o[26368] = data_o[0];
  assign data_o[26432] = data_o[0];
  assign data_o[26496] = data_o[0];
  assign data_o[26560] = data_o[0];
  assign data_o[26624] = data_o[0];
  assign data_o[26688] = data_o[0];
  assign data_o[26752] = data_o[0];
  assign data_o[26816] = data_o[0];
  assign data_o[26880] = data_o[0];
  assign data_o[26944] = data_o[0];
  assign data_o[27008] = data_o[0];
  assign data_o[27072] = data_o[0];
  assign data_o[27136] = data_o[0];
  assign data_o[27200] = data_o[0];
  assign data_o[27264] = data_o[0];
  assign data_o[27328] = data_o[0];
  assign data_o[27392] = data_o[0];
  assign data_o[27456] = data_o[0];
  assign data_o[27520] = data_o[0];
  assign data_o[27584] = data_o[0];
  assign data_o[27648] = data_o[0];
  assign data_o[27712] = data_o[0];
  assign data_o[27776] = data_o[0];
  assign data_o[27840] = data_o[0];
  assign data_o[27904] = data_o[0];
  assign data_o[27968] = data_o[0];
  assign data_o[28032] = data_o[0];
  assign data_o[28096] = data_o[0];
  assign data_o[28160] = data_o[0];
  assign data_o[28224] = data_o[0];
  assign data_o[28288] = data_o[0];
  assign data_o[28352] = data_o[0];
  assign data_o[28416] = data_o[0];
  assign data_o[28480] = data_o[0];
  assign data_o[28544] = data_o[0];
  assign data_o[28608] = data_o[0];
  assign data_o[28672] = data_o[0];
  assign data_o[28736] = data_o[0];
  assign data_o[28800] = data_o[0];
  assign data_o[28864] = data_o[0];
  assign data_o[28928] = data_o[0];
  assign data_o[28992] = data_o[0];
  assign data_o[29056] = data_o[0];
  assign data_o[29120] = data_o[0];
  assign data_o[29184] = data_o[0];
  assign data_o[29248] = data_o[0];
  assign data_o[29312] = data_o[0];
  assign data_o[29376] = data_o[0];
  assign data_o[29440] = data_o[0];
  assign data_o[29504] = data_o[0];
  assign data_o[29568] = data_o[0];
  assign data_o[29632] = data_o[0];
  assign data_o[29696] = data_o[0];
  assign data_o[29760] = data_o[0];
  assign data_o[29824] = data_o[0];
  assign data_o[29888] = data_o[0];
  assign data_o[29952] = data_o[0];
  assign data_o[30016] = data_o[0];
  assign data_o[30080] = data_o[0];
  assign data_o[30144] = data_o[0];
  assign data_o[30208] = data_o[0];
  assign data_o[30272] = data_o[0];
  assign data_o[30336] = data_o[0];
  assign data_o[30400] = data_o[0];
  assign data_o[30464] = data_o[0];
  assign data_o[30528] = data_o[0];
  assign data_o[30592] = data_o[0];
  assign data_o[30656] = data_o[0];
  assign data_o[30720] = data_o[0];
  assign data_o[30784] = data_o[0];
  assign data_o[30848] = data_o[0];
  assign data_o[30912] = data_o[0];
  assign data_o[30976] = data_o[0];
  assign data_o[31040] = data_o[0];
  assign data_o[31104] = data_o[0];
  assign data_o[31168] = data_o[0];
  assign data_o[31232] = data_o[0];
  assign data_o[31296] = data_o[0];
  assign data_o[31360] = data_o[0];
  assign data_o[31424] = data_o[0];
  assign data_o[31488] = data_o[0];
  assign data_o[31552] = data_o[0];
  assign data_o[31616] = data_o[0];
  assign data_o[31680] = data_o[0];
  assign data_o[31744] = data_o[0];
  assign data_o[31808] = data_o[0];
  assign data_o[31872] = data_o[0];
  assign data_o[31936] = data_o[0];

  bsg_two_fifo_width_p64
  fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_i(v_i),
    .v_o(fifo_v),
    .data_o(data_o[63:0]),
    .yumi_i(fifo_yumi)
  );

  assign N1503 = (N0)? 1'b0 : 
                 (N1)? N1502 : 1'b0;
  assign N0 = N1501;
  assign N1 = N1500;
  assign sent_n[0] = (N2)? 1'b1 : 
                     (N1505)? sent_r[0] : 1'b0;
  assign N2 = N1504;
  assign N1509 = (N3)? 1'b0 : 
                 (N4)? N1508 : 1'b0;
  assign N3 = N1507;
  assign N4 = N1506;
  assign sent_n[1] = (N5)? 1'b1 : 
                     (N1511)? sent_r[1] : 1'b0;
  assign N5 = N1510;
  assign N1515 = (N6)? 1'b0 : 
                 (N7)? N1514 : 1'b0;
  assign N6 = N1513;
  assign N7 = N1512;
  assign sent_n[2] = (N8)? 1'b1 : 
                     (N1517)? sent_r[2] : 1'b0;
  assign N8 = N1516;
  assign N1521 = (N9)? 1'b0 : 
                 (N10)? N1520 : 1'b0;
  assign N9 = N1519;
  assign N10 = N1518;
  assign sent_n[3] = (N11)? 1'b1 : 
                     (N1523)? sent_r[3] : 1'b0;
  assign N11 = N1522;
  assign N1527 = (N12)? 1'b0 : 
                 (N13)? N1526 : 1'b0;
  assign N12 = N1525;
  assign N13 = N1524;
  assign sent_n[4] = (N14)? 1'b1 : 
                     (N1529)? sent_r[4] : 1'b0;
  assign N14 = N1528;
  assign N1533 = (N15)? 1'b0 : 
                 (N16)? N1532 : 1'b0;
  assign N15 = N1531;
  assign N16 = N1530;
  assign sent_n[5] = (N17)? 1'b1 : 
                     (N1535)? sent_r[5] : 1'b0;
  assign N17 = N1534;
  assign N1539 = (N18)? 1'b0 : 
                 (N19)? N1538 : 1'b0;
  assign N18 = N1537;
  assign N19 = N1536;
  assign sent_n[6] = (N20)? 1'b1 : 
                     (N1541)? sent_r[6] : 1'b0;
  assign N20 = N1540;
  assign N1545 = (N21)? 1'b0 : 
                 (N22)? N1544 : 1'b0;
  assign N21 = N1543;
  assign N22 = N1542;
  assign sent_n[7] = (N23)? 1'b1 : 
                     (N1547)? sent_r[7] : 1'b0;
  assign N23 = N1546;
  assign N1551 = (N24)? 1'b0 : 
                 (N25)? N1550 : 1'b0;
  assign N24 = N1549;
  assign N25 = N1548;
  assign sent_n[8] = (N26)? 1'b1 : 
                     (N1553)? sent_r[8] : 1'b0;
  assign N26 = N1552;
  assign N1557 = (N27)? 1'b0 : 
                 (N28)? N1556 : 1'b0;
  assign N27 = N1555;
  assign N28 = N1554;
  assign sent_n[9] = (N29)? 1'b1 : 
                     (N1559)? sent_r[9] : 1'b0;
  assign N29 = N1558;
  assign N1563 = (N30)? 1'b0 : 
                 (N31)? N1562 : 1'b0;
  assign N30 = N1561;
  assign N31 = N1560;
  assign sent_n[10] = (N32)? 1'b1 : 
                      (N1565)? sent_r[10] : 1'b0;
  assign N32 = N1564;
  assign N1569 = (N33)? 1'b0 : 
                 (N34)? N1568 : 1'b0;
  assign N33 = N1567;
  assign N34 = N1566;
  assign sent_n[11] = (N35)? 1'b1 : 
                      (N1571)? sent_r[11] : 1'b0;
  assign N35 = N1570;
  assign N1575 = (N36)? 1'b0 : 
                 (N37)? N1574 : 1'b0;
  assign N36 = N1573;
  assign N37 = N1572;
  assign sent_n[12] = (N38)? 1'b1 : 
                      (N1577)? sent_r[12] : 1'b0;
  assign N38 = N1576;
  assign N1581 = (N39)? 1'b0 : 
                 (N40)? N1580 : 1'b0;
  assign N39 = N1579;
  assign N40 = N1578;
  assign sent_n[13] = (N41)? 1'b1 : 
                      (N1583)? sent_r[13] : 1'b0;
  assign N41 = N1582;
  assign N1587 = (N42)? 1'b0 : 
                 (N43)? N1586 : 1'b0;
  assign N42 = N1585;
  assign N43 = N1584;
  assign sent_n[14] = (N44)? 1'b1 : 
                      (N1589)? sent_r[14] : 1'b0;
  assign N44 = N1588;
  assign N1593 = (N45)? 1'b0 : 
                 (N46)? N1592 : 1'b0;
  assign N45 = N1591;
  assign N46 = N1590;
  assign sent_n[15] = (N47)? 1'b1 : 
                      (N1595)? sent_r[15] : 1'b0;
  assign N47 = N1594;
  assign N1599 = (N48)? 1'b0 : 
                 (N49)? N1598 : 1'b0;
  assign N48 = N1597;
  assign N49 = N1596;
  assign sent_n[16] = (N50)? 1'b1 : 
                      (N1601)? sent_r[16] : 1'b0;
  assign N50 = N1600;
  assign N1605 = (N51)? 1'b0 : 
                 (N52)? N1604 : 1'b0;
  assign N51 = N1603;
  assign N52 = N1602;
  assign sent_n[17] = (N53)? 1'b1 : 
                      (N1607)? sent_r[17] : 1'b0;
  assign N53 = N1606;
  assign N1611 = (N54)? 1'b0 : 
                 (N55)? N1610 : 1'b0;
  assign N54 = N1609;
  assign N55 = N1608;
  assign sent_n[18] = (N56)? 1'b1 : 
                      (N1613)? sent_r[18] : 1'b0;
  assign N56 = N1612;
  assign N1617 = (N57)? 1'b0 : 
                 (N58)? N1616 : 1'b0;
  assign N57 = N1615;
  assign N58 = N1614;
  assign sent_n[19] = (N59)? 1'b1 : 
                      (N1619)? sent_r[19] : 1'b0;
  assign N59 = N1618;
  assign N1623 = (N60)? 1'b0 : 
                 (N61)? N1622 : 1'b0;
  assign N60 = N1621;
  assign N61 = N1620;
  assign sent_n[20] = (N62)? 1'b1 : 
                      (N1625)? sent_r[20] : 1'b0;
  assign N62 = N1624;
  assign N1629 = (N63)? 1'b0 : 
                 (N64)? N1628 : 1'b0;
  assign N63 = N1627;
  assign N64 = N1626;
  assign sent_n[21] = (N65)? 1'b1 : 
                      (N1631)? sent_r[21] : 1'b0;
  assign N65 = N1630;
  assign N1635 = (N66)? 1'b0 : 
                 (N67)? N1634 : 1'b0;
  assign N66 = N1633;
  assign N67 = N1632;
  assign sent_n[22] = (N68)? 1'b1 : 
                      (N1637)? sent_r[22] : 1'b0;
  assign N68 = N1636;
  assign N1641 = (N69)? 1'b0 : 
                 (N70)? N1640 : 1'b0;
  assign N69 = N1639;
  assign N70 = N1638;
  assign sent_n[23] = (N71)? 1'b1 : 
                      (N1643)? sent_r[23] : 1'b0;
  assign N71 = N1642;
  assign N1647 = (N72)? 1'b0 : 
                 (N73)? N1646 : 1'b0;
  assign N72 = N1645;
  assign N73 = N1644;
  assign sent_n[24] = (N74)? 1'b1 : 
                      (N1649)? sent_r[24] : 1'b0;
  assign N74 = N1648;
  assign N1653 = (N75)? 1'b0 : 
                 (N76)? N1652 : 1'b0;
  assign N75 = N1651;
  assign N76 = N1650;
  assign sent_n[25] = (N77)? 1'b1 : 
                      (N1655)? sent_r[25] : 1'b0;
  assign N77 = N1654;
  assign N1659 = (N78)? 1'b0 : 
                 (N79)? N1658 : 1'b0;
  assign N78 = N1657;
  assign N79 = N1656;
  assign sent_n[26] = (N80)? 1'b1 : 
                      (N1661)? sent_r[26] : 1'b0;
  assign N80 = N1660;
  assign N1665 = (N81)? 1'b0 : 
                 (N82)? N1664 : 1'b0;
  assign N81 = N1663;
  assign N82 = N1662;
  assign sent_n[27] = (N83)? 1'b1 : 
                      (N1667)? sent_r[27] : 1'b0;
  assign N83 = N1666;
  assign N1671 = (N84)? 1'b0 : 
                 (N85)? N1670 : 1'b0;
  assign N84 = N1669;
  assign N85 = N1668;
  assign sent_n[28] = (N86)? 1'b1 : 
                      (N1673)? sent_r[28] : 1'b0;
  assign N86 = N1672;
  assign N1677 = (N87)? 1'b0 : 
                 (N88)? N1676 : 1'b0;
  assign N87 = N1675;
  assign N88 = N1674;
  assign sent_n[29] = (N89)? 1'b1 : 
                      (N1679)? sent_r[29] : 1'b0;
  assign N89 = N1678;
  assign N1683 = (N90)? 1'b0 : 
                 (N91)? N1682 : 1'b0;
  assign N90 = N1681;
  assign N91 = N1680;
  assign sent_n[30] = (N92)? 1'b1 : 
                      (N1685)? sent_r[30] : 1'b0;
  assign N92 = N1684;
  assign N1689 = (N93)? 1'b0 : 
                 (N94)? N1688 : 1'b0;
  assign N93 = N1687;
  assign N94 = N1686;
  assign sent_n[31] = (N95)? 1'b1 : 
                      (N1691)? sent_r[31] : 1'b0;
  assign N95 = N1690;
  assign N1695 = (N96)? 1'b0 : 
                 (N97)? N1694 : 1'b0;
  assign N96 = N1693;
  assign N97 = N1692;
  assign sent_n[32] = (N98)? 1'b1 : 
                      (N1697)? sent_r[32] : 1'b0;
  assign N98 = N1696;
  assign N1701 = (N99)? 1'b0 : 
                 (N100)? N1700 : 1'b0;
  assign N99 = N1699;
  assign N100 = N1698;
  assign sent_n[33] = (N101)? 1'b1 : 
                      (N1703)? sent_r[33] : 1'b0;
  assign N101 = N1702;
  assign N1707 = (N102)? 1'b0 : 
                 (N103)? N1706 : 1'b0;
  assign N102 = N1705;
  assign N103 = N1704;
  assign sent_n[34] = (N104)? 1'b1 : 
                      (N1709)? sent_r[34] : 1'b0;
  assign N104 = N1708;
  assign N1713 = (N105)? 1'b0 : 
                 (N106)? N1712 : 1'b0;
  assign N105 = N1711;
  assign N106 = N1710;
  assign sent_n[35] = (N107)? 1'b1 : 
                      (N1715)? sent_r[35] : 1'b0;
  assign N107 = N1714;
  assign N1719 = (N108)? 1'b0 : 
                 (N109)? N1718 : 1'b0;
  assign N108 = N1717;
  assign N109 = N1716;
  assign sent_n[36] = (N110)? 1'b1 : 
                      (N1721)? sent_r[36] : 1'b0;
  assign N110 = N1720;
  assign N1725 = (N111)? 1'b0 : 
                 (N112)? N1724 : 1'b0;
  assign N111 = N1723;
  assign N112 = N1722;
  assign sent_n[37] = (N113)? 1'b1 : 
                      (N1727)? sent_r[37] : 1'b0;
  assign N113 = N1726;
  assign N1731 = (N114)? 1'b0 : 
                 (N115)? N1730 : 1'b0;
  assign N114 = N1729;
  assign N115 = N1728;
  assign sent_n[38] = (N116)? 1'b1 : 
                      (N1733)? sent_r[38] : 1'b0;
  assign N116 = N1732;
  assign N1737 = (N117)? 1'b0 : 
                 (N118)? N1736 : 1'b0;
  assign N117 = N1735;
  assign N118 = N1734;
  assign sent_n[39] = (N119)? 1'b1 : 
                      (N1739)? sent_r[39] : 1'b0;
  assign N119 = N1738;
  assign N1743 = (N120)? 1'b0 : 
                 (N121)? N1742 : 1'b0;
  assign N120 = N1741;
  assign N121 = N1740;
  assign sent_n[40] = (N122)? 1'b1 : 
                      (N1745)? sent_r[40] : 1'b0;
  assign N122 = N1744;
  assign N1749 = (N123)? 1'b0 : 
                 (N124)? N1748 : 1'b0;
  assign N123 = N1747;
  assign N124 = N1746;
  assign sent_n[41] = (N125)? 1'b1 : 
                      (N1751)? sent_r[41] : 1'b0;
  assign N125 = N1750;
  assign N1755 = (N126)? 1'b0 : 
                 (N127)? N1754 : 1'b0;
  assign N126 = N1753;
  assign N127 = N1752;
  assign sent_n[42] = (N128)? 1'b1 : 
                      (N1757)? sent_r[42] : 1'b0;
  assign N128 = N1756;
  assign N1761 = (N129)? 1'b0 : 
                 (N130)? N1760 : 1'b0;
  assign N129 = N1759;
  assign N130 = N1758;
  assign sent_n[43] = (N131)? 1'b1 : 
                      (N1763)? sent_r[43] : 1'b0;
  assign N131 = N1762;
  assign N1767 = (N132)? 1'b0 : 
                 (N133)? N1766 : 1'b0;
  assign N132 = N1765;
  assign N133 = N1764;
  assign sent_n[44] = (N134)? 1'b1 : 
                      (N1769)? sent_r[44] : 1'b0;
  assign N134 = N1768;
  assign N1773 = (N135)? 1'b0 : 
                 (N136)? N1772 : 1'b0;
  assign N135 = N1771;
  assign N136 = N1770;
  assign sent_n[45] = (N137)? 1'b1 : 
                      (N1775)? sent_r[45] : 1'b0;
  assign N137 = N1774;
  assign N1779 = (N138)? 1'b0 : 
                 (N139)? N1778 : 1'b0;
  assign N138 = N1777;
  assign N139 = N1776;
  assign sent_n[46] = (N140)? 1'b1 : 
                      (N1781)? sent_r[46] : 1'b0;
  assign N140 = N1780;
  assign N1785 = (N141)? 1'b0 : 
                 (N142)? N1784 : 1'b0;
  assign N141 = N1783;
  assign N142 = N1782;
  assign sent_n[47] = (N143)? 1'b1 : 
                      (N1787)? sent_r[47] : 1'b0;
  assign N143 = N1786;
  assign N1791 = (N144)? 1'b0 : 
                 (N145)? N1790 : 1'b0;
  assign N144 = N1789;
  assign N145 = N1788;
  assign sent_n[48] = (N146)? 1'b1 : 
                      (N1793)? sent_r[48] : 1'b0;
  assign N146 = N1792;
  assign N1797 = (N147)? 1'b0 : 
                 (N148)? N1796 : 1'b0;
  assign N147 = N1795;
  assign N148 = N1794;
  assign sent_n[49] = (N149)? 1'b1 : 
                      (N1799)? sent_r[49] : 1'b0;
  assign N149 = N1798;
  assign N1803 = (N150)? 1'b0 : 
                 (N151)? N1802 : 1'b0;
  assign N150 = N1801;
  assign N151 = N1800;
  assign sent_n[50] = (N152)? 1'b1 : 
                      (N1805)? sent_r[50] : 1'b0;
  assign N152 = N1804;
  assign N1809 = (N153)? 1'b0 : 
                 (N154)? N1808 : 1'b0;
  assign N153 = N1807;
  assign N154 = N1806;
  assign sent_n[51] = (N155)? 1'b1 : 
                      (N1811)? sent_r[51] : 1'b0;
  assign N155 = N1810;
  assign N1815 = (N156)? 1'b0 : 
                 (N157)? N1814 : 1'b0;
  assign N156 = N1813;
  assign N157 = N1812;
  assign sent_n[52] = (N158)? 1'b1 : 
                      (N1817)? sent_r[52] : 1'b0;
  assign N158 = N1816;
  assign N1821 = (N159)? 1'b0 : 
                 (N160)? N1820 : 1'b0;
  assign N159 = N1819;
  assign N160 = N1818;
  assign sent_n[53] = (N161)? 1'b1 : 
                      (N1823)? sent_r[53] : 1'b0;
  assign N161 = N1822;
  assign N1827 = (N162)? 1'b0 : 
                 (N163)? N1826 : 1'b0;
  assign N162 = N1825;
  assign N163 = N1824;
  assign sent_n[54] = (N164)? 1'b1 : 
                      (N1829)? sent_r[54] : 1'b0;
  assign N164 = N1828;
  assign N1833 = (N165)? 1'b0 : 
                 (N166)? N1832 : 1'b0;
  assign N165 = N1831;
  assign N166 = N1830;
  assign sent_n[55] = (N167)? 1'b1 : 
                      (N1835)? sent_r[55] : 1'b0;
  assign N167 = N1834;
  assign N1839 = (N168)? 1'b0 : 
                 (N169)? N1838 : 1'b0;
  assign N168 = N1837;
  assign N169 = N1836;
  assign sent_n[56] = (N170)? 1'b1 : 
                      (N1841)? sent_r[56] : 1'b0;
  assign N170 = N1840;
  assign N1845 = (N171)? 1'b0 : 
                 (N172)? N1844 : 1'b0;
  assign N171 = N1843;
  assign N172 = N1842;
  assign sent_n[57] = (N173)? 1'b1 : 
                      (N1847)? sent_r[57] : 1'b0;
  assign N173 = N1846;
  assign N1851 = (N174)? 1'b0 : 
                 (N175)? N1850 : 1'b0;
  assign N174 = N1849;
  assign N175 = N1848;
  assign sent_n[58] = (N176)? 1'b1 : 
                      (N1853)? sent_r[58] : 1'b0;
  assign N176 = N1852;
  assign N1857 = (N177)? 1'b0 : 
                 (N178)? N1856 : 1'b0;
  assign N177 = N1855;
  assign N178 = N1854;
  assign sent_n[59] = (N179)? 1'b1 : 
                      (N1859)? sent_r[59] : 1'b0;
  assign N179 = N1858;
  assign N1863 = (N180)? 1'b0 : 
                 (N181)? N1862 : 1'b0;
  assign N180 = N1861;
  assign N181 = N1860;
  assign sent_n[60] = (N182)? 1'b1 : 
                      (N1865)? sent_r[60] : 1'b0;
  assign N182 = N1864;
  assign N1869 = (N183)? 1'b0 : 
                 (N184)? N1868 : 1'b0;
  assign N183 = N1867;
  assign N184 = N1866;
  assign sent_n[61] = (N185)? 1'b1 : 
                      (N1871)? sent_r[61] : 1'b0;
  assign N185 = N1870;
  assign N1875 = (N186)? 1'b0 : 
                 (N187)? N1874 : 1'b0;
  assign N186 = N1873;
  assign N187 = N1872;
  assign sent_n[62] = (N188)? 1'b1 : 
                      (N1877)? sent_r[62] : 1'b0;
  assign N188 = N1876;
  assign N1881 = (N189)? 1'b0 : 
                 (N190)? N1880 : 1'b0;
  assign N189 = N1879;
  assign N190 = N1878;
  assign sent_n[63] = (N191)? 1'b1 : 
                      (N1883)? sent_r[63] : 1'b0;
  assign N191 = N1882;
  assign N1887 = (N192)? 1'b0 : 
                 (N193)? N1886 : 1'b0;
  assign N192 = N1885;
  assign N193 = N1884;
  assign sent_n[64] = (N194)? 1'b1 : 
                      (N1889)? sent_r[64] : 1'b0;
  assign N194 = N1888;
  assign N1893 = (N195)? 1'b0 : 
                 (N196)? N1892 : 1'b0;
  assign N195 = N1891;
  assign N196 = N1890;
  assign sent_n[65] = (N197)? 1'b1 : 
                      (N1895)? sent_r[65] : 1'b0;
  assign N197 = N1894;
  assign N1899 = (N198)? 1'b0 : 
                 (N199)? N1898 : 1'b0;
  assign N198 = N1897;
  assign N199 = N1896;
  assign sent_n[66] = (N200)? 1'b1 : 
                      (N1901)? sent_r[66] : 1'b0;
  assign N200 = N1900;
  assign N1905 = (N201)? 1'b0 : 
                 (N202)? N1904 : 1'b0;
  assign N201 = N1903;
  assign N202 = N1902;
  assign sent_n[67] = (N203)? 1'b1 : 
                      (N1907)? sent_r[67] : 1'b0;
  assign N203 = N1906;
  assign N1911 = (N204)? 1'b0 : 
                 (N205)? N1910 : 1'b0;
  assign N204 = N1909;
  assign N205 = N1908;
  assign sent_n[68] = (N206)? 1'b1 : 
                      (N1913)? sent_r[68] : 1'b0;
  assign N206 = N1912;
  assign N1917 = (N207)? 1'b0 : 
                 (N208)? N1916 : 1'b0;
  assign N207 = N1915;
  assign N208 = N1914;
  assign sent_n[69] = (N209)? 1'b1 : 
                      (N1919)? sent_r[69] : 1'b0;
  assign N209 = N1918;
  assign N1923 = (N210)? 1'b0 : 
                 (N211)? N1922 : 1'b0;
  assign N210 = N1921;
  assign N211 = N1920;
  assign sent_n[70] = (N212)? 1'b1 : 
                      (N1925)? sent_r[70] : 1'b0;
  assign N212 = N1924;
  assign N1929 = (N213)? 1'b0 : 
                 (N214)? N1928 : 1'b0;
  assign N213 = N1927;
  assign N214 = N1926;
  assign sent_n[71] = (N215)? 1'b1 : 
                      (N1931)? sent_r[71] : 1'b0;
  assign N215 = N1930;
  assign N1935 = (N216)? 1'b0 : 
                 (N217)? N1934 : 1'b0;
  assign N216 = N1933;
  assign N217 = N1932;
  assign sent_n[72] = (N218)? 1'b1 : 
                      (N1937)? sent_r[72] : 1'b0;
  assign N218 = N1936;
  assign N1941 = (N219)? 1'b0 : 
                 (N220)? N1940 : 1'b0;
  assign N219 = N1939;
  assign N220 = N1938;
  assign sent_n[73] = (N221)? 1'b1 : 
                      (N1943)? sent_r[73] : 1'b0;
  assign N221 = N1942;
  assign N1947 = (N222)? 1'b0 : 
                 (N223)? N1946 : 1'b0;
  assign N222 = N1945;
  assign N223 = N1944;
  assign sent_n[74] = (N224)? 1'b1 : 
                      (N1949)? sent_r[74] : 1'b0;
  assign N224 = N1948;
  assign N1953 = (N225)? 1'b0 : 
                 (N226)? N1952 : 1'b0;
  assign N225 = N1951;
  assign N226 = N1950;
  assign sent_n[75] = (N227)? 1'b1 : 
                      (N1955)? sent_r[75] : 1'b0;
  assign N227 = N1954;
  assign N1959 = (N228)? 1'b0 : 
                 (N229)? N1958 : 1'b0;
  assign N228 = N1957;
  assign N229 = N1956;
  assign sent_n[76] = (N230)? 1'b1 : 
                      (N1961)? sent_r[76] : 1'b0;
  assign N230 = N1960;
  assign N1965 = (N231)? 1'b0 : 
                 (N232)? N1964 : 1'b0;
  assign N231 = N1963;
  assign N232 = N1962;
  assign sent_n[77] = (N233)? 1'b1 : 
                      (N1967)? sent_r[77] : 1'b0;
  assign N233 = N1966;
  assign N1971 = (N234)? 1'b0 : 
                 (N235)? N1970 : 1'b0;
  assign N234 = N1969;
  assign N235 = N1968;
  assign sent_n[78] = (N236)? 1'b1 : 
                      (N1973)? sent_r[78] : 1'b0;
  assign N236 = N1972;
  assign N1977 = (N237)? 1'b0 : 
                 (N238)? N1976 : 1'b0;
  assign N237 = N1975;
  assign N238 = N1974;
  assign sent_n[79] = (N239)? 1'b1 : 
                      (N1979)? sent_r[79] : 1'b0;
  assign N239 = N1978;
  assign N1983 = (N240)? 1'b0 : 
                 (N241)? N1982 : 1'b0;
  assign N240 = N1981;
  assign N241 = N1980;
  assign sent_n[80] = (N242)? 1'b1 : 
                      (N1985)? sent_r[80] : 1'b0;
  assign N242 = N1984;
  assign N1989 = (N243)? 1'b0 : 
                 (N244)? N1988 : 1'b0;
  assign N243 = N1987;
  assign N244 = N1986;
  assign sent_n[81] = (N245)? 1'b1 : 
                      (N1991)? sent_r[81] : 1'b0;
  assign N245 = N1990;
  assign N1995 = (N246)? 1'b0 : 
                 (N247)? N1994 : 1'b0;
  assign N246 = N1993;
  assign N247 = N1992;
  assign sent_n[82] = (N248)? 1'b1 : 
                      (N1997)? sent_r[82] : 1'b0;
  assign N248 = N1996;
  assign N2001 = (N249)? 1'b0 : 
                 (N250)? N2000 : 1'b0;
  assign N249 = N1999;
  assign N250 = N1998;
  assign sent_n[83] = (N251)? 1'b1 : 
                      (N2003)? sent_r[83] : 1'b0;
  assign N251 = N2002;
  assign N2007 = (N252)? 1'b0 : 
                 (N253)? N2006 : 1'b0;
  assign N252 = N2005;
  assign N253 = N2004;
  assign sent_n[84] = (N254)? 1'b1 : 
                      (N2009)? sent_r[84] : 1'b0;
  assign N254 = N2008;
  assign N2013 = (N255)? 1'b0 : 
                 (N256)? N2012 : 1'b0;
  assign N255 = N2011;
  assign N256 = N2010;
  assign sent_n[85] = (N257)? 1'b1 : 
                      (N2015)? sent_r[85] : 1'b0;
  assign N257 = N2014;
  assign N2019 = (N258)? 1'b0 : 
                 (N259)? N2018 : 1'b0;
  assign N258 = N2017;
  assign N259 = N2016;
  assign sent_n[86] = (N260)? 1'b1 : 
                      (N2021)? sent_r[86] : 1'b0;
  assign N260 = N2020;
  assign N2025 = (N261)? 1'b0 : 
                 (N262)? N2024 : 1'b0;
  assign N261 = N2023;
  assign N262 = N2022;
  assign sent_n[87] = (N263)? 1'b1 : 
                      (N2027)? sent_r[87] : 1'b0;
  assign N263 = N2026;
  assign N2031 = (N264)? 1'b0 : 
                 (N265)? N2030 : 1'b0;
  assign N264 = N2029;
  assign N265 = N2028;
  assign sent_n[88] = (N266)? 1'b1 : 
                      (N2033)? sent_r[88] : 1'b0;
  assign N266 = N2032;
  assign N2037 = (N267)? 1'b0 : 
                 (N268)? N2036 : 1'b0;
  assign N267 = N2035;
  assign N268 = N2034;
  assign sent_n[89] = (N269)? 1'b1 : 
                      (N2039)? sent_r[89] : 1'b0;
  assign N269 = N2038;
  assign N2043 = (N270)? 1'b0 : 
                 (N271)? N2042 : 1'b0;
  assign N270 = N2041;
  assign N271 = N2040;
  assign sent_n[90] = (N272)? 1'b1 : 
                      (N2045)? sent_r[90] : 1'b0;
  assign N272 = N2044;
  assign N2049 = (N273)? 1'b0 : 
                 (N274)? N2048 : 1'b0;
  assign N273 = N2047;
  assign N274 = N2046;
  assign sent_n[91] = (N275)? 1'b1 : 
                      (N2051)? sent_r[91] : 1'b0;
  assign N275 = N2050;
  assign N2055 = (N276)? 1'b0 : 
                 (N277)? N2054 : 1'b0;
  assign N276 = N2053;
  assign N277 = N2052;
  assign sent_n[92] = (N278)? 1'b1 : 
                      (N2057)? sent_r[92] : 1'b0;
  assign N278 = N2056;
  assign N2061 = (N279)? 1'b0 : 
                 (N280)? N2060 : 1'b0;
  assign N279 = N2059;
  assign N280 = N2058;
  assign sent_n[93] = (N281)? 1'b1 : 
                      (N2063)? sent_r[93] : 1'b0;
  assign N281 = N2062;
  assign N2067 = (N282)? 1'b0 : 
                 (N283)? N2066 : 1'b0;
  assign N282 = N2065;
  assign N283 = N2064;
  assign sent_n[94] = (N284)? 1'b1 : 
                      (N2069)? sent_r[94] : 1'b0;
  assign N284 = N2068;
  assign N2073 = (N285)? 1'b0 : 
                 (N286)? N2072 : 1'b0;
  assign N285 = N2071;
  assign N286 = N2070;
  assign sent_n[95] = (N287)? 1'b1 : 
                      (N2075)? sent_r[95] : 1'b0;
  assign N287 = N2074;
  assign N2079 = (N288)? 1'b0 : 
                 (N289)? N2078 : 1'b0;
  assign N288 = N2077;
  assign N289 = N2076;
  assign sent_n[96] = (N290)? 1'b1 : 
                      (N2081)? sent_r[96] : 1'b0;
  assign N290 = N2080;
  assign N2085 = (N291)? 1'b0 : 
                 (N292)? N2084 : 1'b0;
  assign N291 = N2083;
  assign N292 = N2082;
  assign sent_n[97] = (N293)? 1'b1 : 
                      (N2087)? sent_r[97] : 1'b0;
  assign N293 = N2086;
  assign N2091 = (N294)? 1'b0 : 
                 (N295)? N2090 : 1'b0;
  assign N294 = N2089;
  assign N295 = N2088;
  assign sent_n[98] = (N296)? 1'b1 : 
                      (N2093)? sent_r[98] : 1'b0;
  assign N296 = N2092;
  assign N2097 = (N297)? 1'b0 : 
                 (N298)? N2096 : 1'b0;
  assign N297 = N2095;
  assign N298 = N2094;
  assign sent_n[99] = (N299)? 1'b1 : 
                      (N2099)? sent_r[99] : 1'b0;
  assign N299 = N2098;
  assign N2103 = (N300)? 1'b0 : 
                 (N301)? N2102 : 1'b0;
  assign N300 = N2101;
  assign N301 = N2100;
  assign sent_n[100] = (N302)? 1'b1 : 
                       (N2105)? sent_r[100] : 1'b0;
  assign N302 = N2104;
  assign N2109 = (N303)? 1'b0 : 
                 (N304)? N2108 : 1'b0;
  assign N303 = N2107;
  assign N304 = N2106;
  assign sent_n[101] = (N305)? 1'b1 : 
                       (N2111)? sent_r[101] : 1'b0;
  assign N305 = N2110;
  assign N2115 = (N306)? 1'b0 : 
                 (N307)? N2114 : 1'b0;
  assign N306 = N2113;
  assign N307 = N2112;
  assign sent_n[102] = (N308)? 1'b1 : 
                       (N2117)? sent_r[102] : 1'b0;
  assign N308 = N2116;
  assign N2121 = (N309)? 1'b0 : 
                 (N310)? N2120 : 1'b0;
  assign N309 = N2119;
  assign N310 = N2118;
  assign sent_n[103] = (N311)? 1'b1 : 
                       (N2123)? sent_r[103] : 1'b0;
  assign N311 = N2122;
  assign N2127 = (N312)? 1'b0 : 
                 (N313)? N2126 : 1'b0;
  assign N312 = N2125;
  assign N313 = N2124;
  assign sent_n[104] = (N314)? 1'b1 : 
                       (N2129)? sent_r[104] : 1'b0;
  assign N314 = N2128;
  assign N2133 = (N315)? 1'b0 : 
                 (N316)? N2132 : 1'b0;
  assign N315 = N2131;
  assign N316 = N2130;
  assign sent_n[105] = (N317)? 1'b1 : 
                       (N2135)? sent_r[105] : 1'b0;
  assign N317 = N2134;
  assign N2139 = (N318)? 1'b0 : 
                 (N319)? N2138 : 1'b0;
  assign N318 = N2137;
  assign N319 = N2136;
  assign sent_n[106] = (N320)? 1'b1 : 
                       (N2141)? sent_r[106] : 1'b0;
  assign N320 = N2140;
  assign N2145 = (N321)? 1'b0 : 
                 (N322)? N2144 : 1'b0;
  assign N321 = N2143;
  assign N322 = N2142;
  assign sent_n[107] = (N323)? 1'b1 : 
                       (N2147)? sent_r[107] : 1'b0;
  assign N323 = N2146;
  assign N2151 = (N324)? 1'b0 : 
                 (N325)? N2150 : 1'b0;
  assign N324 = N2149;
  assign N325 = N2148;
  assign sent_n[108] = (N326)? 1'b1 : 
                       (N2153)? sent_r[108] : 1'b0;
  assign N326 = N2152;
  assign N2157 = (N327)? 1'b0 : 
                 (N328)? N2156 : 1'b0;
  assign N327 = N2155;
  assign N328 = N2154;
  assign sent_n[109] = (N329)? 1'b1 : 
                       (N2159)? sent_r[109] : 1'b0;
  assign N329 = N2158;
  assign N2163 = (N330)? 1'b0 : 
                 (N331)? N2162 : 1'b0;
  assign N330 = N2161;
  assign N331 = N2160;
  assign sent_n[110] = (N332)? 1'b1 : 
                       (N2165)? sent_r[110] : 1'b0;
  assign N332 = N2164;
  assign N2169 = (N333)? 1'b0 : 
                 (N334)? N2168 : 1'b0;
  assign N333 = N2167;
  assign N334 = N2166;
  assign sent_n[111] = (N335)? 1'b1 : 
                       (N2171)? sent_r[111] : 1'b0;
  assign N335 = N2170;
  assign N2175 = (N336)? 1'b0 : 
                 (N337)? N2174 : 1'b0;
  assign N336 = N2173;
  assign N337 = N2172;
  assign sent_n[112] = (N338)? 1'b1 : 
                       (N2177)? sent_r[112] : 1'b0;
  assign N338 = N2176;
  assign N2181 = (N339)? 1'b0 : 
                 (N340)? N2180 : 1'b0;
  assign N339 = N2179;
  assign N340 = N2178;
  assign sent_n[113] = (N341)? 1'b1 : 
                       (N2183)? sent_r[113] : 1'b0;
  assign N341 = N2182;
  assign N2187 = (N342)? 1'b0 : 
                 (N343)? N2186 : 1'b0;
  assign N342 = N2185;
  assign N343 = N2184;
  assign sent_n[114] = (N344)? 1'b1 : 
                       (N2189)? sent_r[114] : 1'b0;
  assign N344 = N2188;
  assign N2193 = (N345)? 1'b0 : 
                 (N346)? N2192 : 1'b0;
  assign N345 = N2191;
  assign N346 = N2190;
  assign sent_n[115] = (N347)? 1'b1 : 
                       (N2195)? sent_r[115] : 1'b0;
  assign N347 = N2194;
  assign N2199 = (N348)? 1'b0 : 
                 (N349)? N2198 : 1'b0;
  assign N348 = N2197;
  assign N349 = N2196;
  assign sent_n[116] = (N350)? 1'b1 : 
                       (N2201)? sent_r[116] : 1'b0;
  assign N350 = N2200;
  assign N2205 = (N351)? 1'b0 : 
                 (N352)? N2204 : 1'b0;
  assign N351 = N2203;
  assign N352 = N2202;
  assign sent_n[117] = (N353)? 1'b1 : 
                       (N2207)? sent_r[117] : 1'b0;
  assign N353 = N2206;
  assign N2211 = (N354)? 1'b0 : 
                 (N355)? N2210 : 1'b0;
  assign N354 = N2209;
  assign N355 = N2208;
  assign sent_n[118] = (N356)? 1'b1 : 
                       (N2213)? sent_r[118] : 1'b0;
  assign N356 = N2212;
  assign N2217 = (N357)? 1'b0 : 
                 (N358)? N2216 : 1'b0;
  assign N357 = N2215;
  assign N358 = N2214;
  assign sent_n[119] = (N359)? 1'b1 : 
                       (N2219)? sent_r[119] : 1'b0;
  assign N359 = N2218;
  assign N2223 = (N360)? 1'b0 : 
                 (N361)? N2222 : 1'b0;
  assign N360 = N2221;
  assign N361 = N2220;
  assign sent_n[120] = (N362)? 1'b1 : 
                       (N2225)? sent_r[120] : 1'b0;
  assign N362 = N2224;
  assign N2229 = (N363)? 1'b0 : 
                 (N364)? N2228 : 1'b0;
  assign N363 = N2227;
  assign N364 = N2226;
  assign sent_n[121] = (N365)? 1'b1 : 
                       (N2231)? sent_r[121] : 1'b0;
  assign N365 = N2230;
  assign N2235 = (N366)? 1'b0 : 
                 (N367)? N2234 : 1'b0;
  assign N366 = N2233;
  assign N367 = N2232;
  assign sent_n[122] = (N368)? 1'b1 : 
                       (N2237)? sent_r[122] : 1'b0;
  assign N368 = N2236;
  assign N2241 = (N369)? 1'b0 : 
                 (N370)? N2240 : 1'b0;
  assign N369 = N2239;
  assign N370 = N2238;
  assign sent_n[123] = (N371)? 1'b1 : 
                       (N2243)? sent_r[123] : 1'b0;
  assign N371 = N2242;
  assign N2247 = (N372)? 1'b0 : 
                 (N373)? N2246 : 1'b0;
  assign N372 = N2245;
  assign N373 = N2244;
  assign sent_n[124] = (N374)? 1'b1 : 
                       (N2249)? sent_r[124] : 1'b0;
  assign N374 = N2248;
  assign N2253 = (N375)? 1'b0 : 
                 (N376)? N2252 : 1'b0;
  assign N375 = N2251;
  assign N376 = N2250;
  assign sent_n[125] = (N377)? 1'b1 : 
                       (N2255)? sent_r[125] : 1'b0;
  assign N377 = N2254;
  assign N2259 = (N378)? 1'b0 : 
                 (N379)? N2258 : 1'b0;
  assign N378 = N2257;
  assign N379 = N2256;
  assign sent_n[126] = (N380)? 1'b1 : 
                       (N2261)? sent_r[126] : 1'b0;
  assign N380 = N2260;
  assign N2265 = (N381)? 1'b0 : 
                 (N382)? N2264 : 1'b0;
  assign N381 = N2263;
  assign N382 = N2262;
  assign sent_n[127] = (N383)? 1'b1 : 
                       (N2267)? sent_r[127] : 1'b0;
  assign N383 = N2266;
  assign N2271 = (N384)? 1'b0 : 
                 (N385)? N2270 : 1'b0;
  assign N384 = N2269;
  assign N385 = N2268;
  assign sent_n[128] = (N386)? 1'b1 : 
                       (N2273)? sent_r[128] : 1'b0;
  assign N386 = N2272;
  assign N2277 = (N387)? 1'b0 : 
                 (N388)? N2276 : 1'b0;
  assign N387 = N2275;
  assign N388 = N2274;
  assign sent_n[129] = (N389)? 1'b1 : 
                       (N2279)? sent_r[129] : 1'b0;
  assign N389 = N2278;
  assign N2283 = (N390)? 1'b0 : 
                 (N391)? N2282 : 1'b0;
  assign N390 = N2281;
  assign N391 = N2280;
  assign sent_n[130] = (N392)? 1'b1 : 
                       (N2285)? sent_r[130] : 1'b0;
  assign N392 = N2284;
  assign N2289 = (N393)? 1'b0 : 
                 (N394)? N2288 : 1'b0;
  assign N393 = N2287;
  assign N394 = N2286;
  assign sent_n[131] = (N395)? 1'b1 : 
                       (N2291)? sent_r[131] : 1'b0;
  assign N395 = N2290;
  assign N2295 = (N396)? 1'b0 : 
                 (N397)? N2294 : 1'b0;
  assign N396 = N2293;
  assign N397 = N2292;
  assign sent_n[132] = (N398)? 1'b1 : 
                       (N2297)? sent_r[132] : 1'b0;
  assign N398 = N2296;
  assign N2301 = (N399)? 1'b0 : 
                 (N400)? N2300 : 1'b0;
  assign N399 = N2299;
  assign N400 = N2298;
  assign sent_n[133] = (N401)? 1'b1 : 
                       (N2303)? sent_r[133] : 1'b0;
  assign N401 = N2302;
  assign N2307 = (N402)? 1'b0 : 
                 (N403)? N2306 : 1'b0;
  assign N402 = N2305;
  assign N403 = N2304;
  assign sent_n[134] = (N404)? 1'b1 : 
                       (N2309)? sent_r[134] : 1'b0;
  assign N404 = N2308;
  assign N2313 = (N405)? 1'b0 : 
                 (N406)? N2312 : 1'b0;
  assign N405 = N2311;
  assign N406 = N2310;
  assign sent_n[135] = (N407)? 1'b1 : 
                       (N2315)? sent_r[135] : 1'b0;
  assign N407 = N2314;
  assign N2319 = (N408)? 1'b0 : 
                 (N409)? N2318 : 1'b0;
  assign N408 = N2317;
  assign N409 = N2316;
  assign sent_n[136] = (N410)? 1'b1 : 
                       (N2321)? sent_r[136] : 1'b0;
  assign N410 = N2320;
  assign N2325 = (N411)? 1'b0 : 
                 (N412)? N2324 : 1'b0;
  assign N411 = N2323;
  assign N412 = N2322;
  assign sent_n[137] = (N413)? 1'b1 : 
                       (N2327)? sent_r[137] : 1'b0;
  assign N413 = N2326;
  assign N2331 = (N414)? 1'b0 : 
                 (N415)? N2330 : 1'b0;
  assign N414 = N2329;
  assign N415 = N2328;
  assign sent_n[138] = (N416)? 1'b1 : 
                       (N2333)? sent_r[138] : 1'b0;
  assign N416 = N2332;
  assign N2337 = (N417)? 1'b0 : 
                 (N418)? N2336 : 1'b0;
  assign N417 = N2335;
  assign N418 = N2334;
  assign sent_n[139] = (N419)? 1'b1 : 
                       (N2339)? sent_r[139] : 1'b0;
  assign N419 = N2338;
  assign N2343 = (N420)? 1'b0 : 
                 (N421)? N2342 : 1'b0;
  assign N420 = N2341;
  assign N421 = N2340;
  assign sent_n[140] = (N422)? 1'b1 : 
                       (N2345)? sent_r[140] : 1'b0;
  assign N422 = N2344;
  assign N2349 = (N423)? 1'b0 : 
                 (N424)? N2348 : 1'b0;
  assign N423 = N2347;
  assign N424 = N2346;
  assign sent_n[141] = (N425)? 1'b1 : 
                       (N2351)? sent_r[141] : 1'b0;
  assign N425 = N2350;
  assign N2355 = (N426)? 1'b0 : 
                 (N427)? N2354 : 1'b0;
  assign N426 = N2353;
  assign N427 = N2352;
  assign sent_n[142] = (N428)? 1'b1 : 
                       (N2357)? sent_r[142] : 1'b0;
  assign N428 = N2356;
  assign N2361 = (N429)? 1'b0 : 
                 (N430)? N2360 : 1'b0;
  assign N429 = N2359;
  assign N430 = N2358;
  assign sent_n[143] = (N431)? 1'b1 : 
                       (N2363)? sent_r[143] : 1'b0;
  assign N431 = N2362;
  assign N2367 = (N432)? 1'b0 : 
                 (N433)? N2366 : 1'b0;
  assign N432 = N2365;
  assign N433 = N2364;
  assign sent_n[144] = (N434)? 1'b1 : 
                       (N2369)? sent_r[144] : 1'b0;
  assign N434 = N2368;
  assign N2373 = (N435)? 1'b0 : 
                 (N436)? N2372 : 1'b0;
  assign N435 = N2371;
  assign N436 = N2370;
  assign sent_n[145] = (N437)? 1'b1 : 
                       (N2375)? sent_r[145] : 1'b0;
  assign N437 = N2374;
  assign N2379 = (N438)? 1'b0 : 
                 (N439)? N2378 : 1'b0;
  assign N438 = N2377;
  assign N439 = N2376;
  assign sent_n[146] = (N440)? 1'b1 : 
                       (N2381)? sent_r[146] : 1'b0;
  assign N440 = N2380;
  assign N2385 = (N441)? 1'b0 : 
                 (N442)? N2384 : 1'b0;
  assign N441 = N2383;
  assign N442 = N2382;
  assign sent_n[147] = (N443)? 1'b1 : 
                       (N2387)? sent_r[147] : 1'b0;
  assign N443 = N2386;
  assign N2391 = (N444)? 1'b0 : 
                 (N445)? N2390 : 1'b0;
  assign N444 = N2389;
  assign N445 = N2388;
  assign sent_n[148] = (N446)? 1'b1 : 
                       (N2393)? sent_r[148] : 1'b0;
  assign N446 = N2392;
  assign N2397 = (N447)? 1'b0 : 
                 (N448)? N2396 : 1'b0;
  assign N447 = N2395;
  assign N448 = N2394;
  assign sent_n[149] = (N449)? 1'b1 : 
                       (N2399)? sent_r[149] : 1'b0;
  assign N449 = N2398;
  assign N2403 = (N450)? 1'b0 : 
                 (N451)? N2402 : 1'b0;
  assign N450 = N2401;
  assign N451 = N2400;
  assign sent_n[150] = (N452)? 1'b1 : 
                       (N2405)? sent_r[150] : 1'b0;
  assign N452 = N2404;
  assign N2409 = (N453)? 1'b0 : 
                 (N454)? N2408 : 1'b0;
  assign N453 = N2407;
  assign N454 = N2406;
  assign sent_n[151] = (N455)? 1'b1 : 
                       (N2411)? sent_r[151] : 1'b0;
  assign N455 = N2410;
  assign N2415 = (N456)? 1'b0 : 
                 (N457)? N2414 : 1'b0;
  assign N456 = N2413;
  assign N457 = N2412;
  assign sent_n[152] = (N458)? 1'b1 : 
                       (N2417)? sent_r[152] : 1'b0;
  assign N458 = N2416;
  assign N2421 = (N459)? 1'b0 : 
                 (N460)? N2420 : 1'b0;
  assign N459 = N2419;
  assign N460 = N2418;
  assign sent_n[153] = (N461)? 1'b1 : 
                       (N2423)? sent_r[153] : 1'b0;
  assign N461 = N2422;
  assign N2427 = (N462)? 1'b0 : 
                 (N463)? N2426 : 1'b0;
  assign N462 = N2425;
  assign N463 = N2424;
  assign sent_n[154] = (N464)? 1'b1 : 
                       (N2429)? sent_r[154] : 1'b0;
  assign N464 = N2428;
  assign N2433 = (N465)? 1'b0 : 
                 (N466)? N2432 : 1'b0;
  assign N465 = N2431;
  assign N466 = N2430;
  assign sent_n[155] = (N467)? 1'b1 : 
                       (N2435)? sent_r[155] : 1'b0;
  assign N467 = N2434;
  assign N2439 = (N468)? 1'b0 : 
                 (N469)? N2438 : 1'b0;
  assign N468 = N2437;
  assign N469 = N2436;
  assign sent_n[156] = (N470)? 1'b1 : 
                       (N2441)? sent_r[156] : 1'b0;
  assign N470 = N2440;
  assign N2445 = (N471)? 1'b0 : 
                 (N472)? N2444 : 1'b0;
  assign N471 = N2443;
  assign N472 = N2442;
  assign sent_n[157] = (N473)? 1'b1 : 
                       (N2447)? sent_r[157] : 1'b0;
  assign N473 = N2446;
  assign N2451 = (N474)? 1'b0 : 
                 (N475)? N2450 : 1'b0;
  assign N474 = N2449;
  assign N475 = N2448;
  assign sent_n[158] = (N476)? 1'b1 : 
                       (N2453)? sent_r[158] : 1'b0;
  assign N476 = N2452;
  assign N2457 = (N477)? 1'b0 : 
                 (N478)? N2456 : 1'b0;
  assign N477 = N2455;
  assign N478 = N2454;
  assign sent_n[159] = (N479)? 1'b1 : 
                       (N2459)? sent_r[159] : 1'b0;
  assign N479 = N2458;
  assign N2463 = (N480)? 1'b0 : 
                 (N481)? N2462 : 1'b0;
  assign N480 = N2461;
  assign N481 = N2460;
  assign sent_n[160] = (N482)? 1'b1 : 
                       (N2465)? sent_r[160] : 1'b0;
  assign N482 = N2464;
  assign N2469 = (N483)? 1'b0 : 
                 (N484)? N2468 : 1'b0;
  assign N483 = N2467;
  assign N484 = N2466;
  assign sent_n[161] = (N485)? 1'b1 : 
                       (N2471)? sent_r[161] : 1'b0;
  assign N485 = N2470;
  assign N2475 = (N486)? 1'b0 : 
                 (N487)? N2474 : 1'b0;
  assign N486 = N2473;
  assign N487 = N2472;
  assign sent_n[162] = (N488)? 1'b1 : 
                       (N2477)? sent_r[162] : 1'b0;
  assign N488 = N2476;
  assign N2481 = (N489)? 1'b0 : 
                 (N490)? N2480 : 1'b0;
  assign N489 = N2479;
  assign N490 = N2478;
  assign sent_n[163] = (N491)? 1'b1 : 
                       (N2483)? sent_r[163] : 1'b0;
  assign N491 = N2482;
  assign N2487 = (N492)? 1'b0 : 
                 (N493)? N2486 : 1'b0;
  assign N492 = N2485;
  assign N493 = N2484;
  assign sent_n[164] = (N494)? 1'b1 : 
                       (N2489)? sent_r[164] : 1'b0;
  assign N494 = N2488;
  assign N2493 = (N495)? 1'b0 : 
                 (N496)? N2492 : 1'b0;
  assign N495 = N2491;
  assign N496 = N2490;
  assign sent_n[165] = (N497)? 1'b1 : 
                       (N2495)? sent_r[165] : 1'b0;
  assign N497 = N2494;
  assign N2499 = (N498)? 1'b0 : 
                 (N499)? N2498 : 1'b0;
  assign N498 = N2497;
  assign N499 = N2496;
  assign sent_n[166] = (N500)? 1'b1 : 
                       (N2501)? sent_r[166] : 1'b0;
  assign N500 = N2500;
  assign N2505 = (N501)? 1'b0 : 
                 (N502)? N2504 : 1'b0;
  assign N501 = N2503;
  assign N502 = N2502;
  assign sent_n[167] = (N503)? 1'b1 : 
                       (N2507)? sent_r[167] : 1'b0;
  assign N503 = N2506;
  assign N2511 = (N504)? 1'b0 : 
                 (N505)? N2510 : 1'b0;
  assign N504 = N2509;
  assign N505 = N2508;
  assign sent_n[168] = (N506)? 1'b1 : 
                       (N2513)? sent_r[168] : 1'b0;
  assign N506 = N2512;
  assign N2517 = (N507)? 1'b0 : 
                 (N508)? N2516 : 1'b0;
  assign N507 = N2515;
  assign N508 = N2514;
  assign sent_n[169] = (N509)? 1'b1 : 
                       (N2519)? sent_r[169] : 1'b0;
  assign N509 = N2518;
  assign N2523 = (N510)? 1'b0 : 
                 (N511)? N2522 : 1'b0;
  assign N510 = N2521;
  assign N511 = N2520;
  assign sent_n[170] = (N512)? 1'b1 : 
                       (N2525)? sent_r[170] : 1'b0;
  assign N512 = N2524;
  assign N2529 = (N513)? 1'b0 : 
                 (N514)? N2528 : 1'b0;
  assign N513 = N2527;
  assign N514 = N2526;
  assign sent_n[171] = (N515)? 1'b1 : 
                       (N2531)? sent_r[171] : 1'b0;
  assign N515 = N2530;
  assign N2535 = (N516)? 1'b0 : 
                 (N517)? N2534 : 1'b0;
  assign N516 = N2533;
  assign N517 = N2532;
  assign sent_n[172] = (N518)? 1'b1 : 
                       (N2537)? sent_r[172] : 1'b0;
  assign N518 = N2536;
  assign N2541 = (N519)? 1'b0 : 
                 (N520)? N2540 : 1'b0;
  assign N519 = N2539;
  assign N520 = N2538;
  assign sent_n[173] = (N521)? 1'b1 : 
                       (N2543)? sent_r[173] : 1'b0;
  assign N521 = N2542;
  assign N2547 = (N522)? 1'b0 : 
                 (N523)? N2546 : 1'b0;
  assign N522 = N2545;
  assign N523 = N2544;
  assign sent_n[174] = (N524)? 1'b1 : 
                       (N2549)? sent_r[174] : 1'b0;
  assign N524 = N2548;
  assign N2553 = (N525)? 1'b0 : 
                 (N526)? N2552 : 1'b0;
  assign N525 = N2551;
  assign N526 = N2550;
  assign sent_n[175] = (N527)? 1'b1 : 
                       (N2555)? sent_r[175] : 1'b0;
  assign N527 = N2554;
  assign N2559 = (N528)? 1'b0 : 
                 (N529)? N2558 : 1'b0;
  assign N528 = N2557;
  assign N529 = N2556;
  assign sent_n[176] = (N530)? 1'b1 : 
                       (N2561)? sent_r[176] : 1'b0;
  assign N530 = N2560;
  assign N2565 = (N531)? 1'b0 : 
                 (N532)? N2564 : 1'b0;
  assign N531 = N2563;
  assign N532 = N2562;
  assign sent_n[177] = (N533)? 1'b1 : 
                       (N2567)? sent_r[177] : 1'b0;
  assign N533 = N2566;
  assign N2571 = (N534)? 1'b0 : 
                 (N535)? N2570 : 1'b0;
  assign N534 = N2569;
  assign N535 = N2568;
  assign sent_n[178] = (N536)? 1'b1 : 
                       (N2573)? sent_r[178] : 1'b0;
  assign N536 = N2572;
  assign N2577 = (N537)? 1'b0 : 
                 (N538)? N2576 : 1'b0;
  assign N537 = N2575;
  assign N538 = N2574;
  assign sent_n[179] = (N539)? 1'b1 : 
                       (N2579)? sent_r[179] : 1'b0;
  assign N539 = N2578;
  assign N2583 = (N540)? 1'b0 : 
                 (N541)? N2582 : 1'b0;
  assign N540 = N2581;
  assign N541 = N2580;
  assign sent_n[180] = (N542)? 1'b1 : 
                       (N2585)? sent_r[180] : 1'b0;
  assign N542 = N2584;
  assign N2589 = (N543)? 1'b0 : 
                 (N544)? N2588 : 1'b0;
  assign N543 = N2587;
  assign N544 = N2586;
  assign sent_n[181] = (N545)? 1'b1 : 
                       (N2591)? sent_r[181] : 1'b0;
  assign N545 = N2590;
  assign N2595 = (N546)? 1'b0 : 
                 (N547)? N2594 : 1'b0;
  assign N546 = N2593;
  assign N547 = N2592;
  assign sent_n[182] = (N548)? 1'b1 : 
                       (N2597)? sent_r[182] : 1'b0;
  assign N548 = N2596;
  assign N2601 = (N549)? 1'b0 : 
                 (N550)? N2600 : 1'b0;
  assign N549 = N2599;
  assign N550 = N2598;
  assign sent_n[183] = (N551)? 1'b1 : 
                       (N2603)? sent_r[183] : 1'b0;
  assign N551 = N2602;
  assign N2607 = (N552)? 1'b0 : 
                 (N553)? N2606 : 1'b0;
  assign N552 = N2605;
  assign N553 = N2604;
  assign sent_n[184] = (N554)? 1'b1 : 
                       (N2609)? sent_r[184] : 1'b0;
  assign N554 = N2608;
  assign N2613 = (N555)? 1'b0 : 
                 (N556)? N2612 : 1'b0;
  assign N555 = N2611;
  assign N556 = N2610;
  assign sent_n[185] = (N557)? 1'b1 : 
                       (N2615)? sent_r[185] : 1'b0;
  assign N557 = N2614;
  assign N2619 = (N558)? 1'b0 : 
                 (N559)? N2618 : 1'b0;
  assign N558 = N2617;
  assign N559 = N2616;
  assign sent_n[186] = (N560)? 1'b1 : 
                       (N2621)? sent_r[186] : 1'b0;
  assign N560 = N2620;
  assign N2625 = (N561)? 1'b0 : 
                 (N562)? N2624 : 1'b0;
  assign N561 = N2623;
  assign N562 = N2622;
  assign sent_n[187] = (N563)? 1'b1 : 
                       (N2627)? sent_r[187] : 1'b0;
  assign N563 = N2626;
  assign N2631 = (N564)? 1'b0 : 
                 (N565)? N2630 : 1'b0;
  assign N564 = N2629;
  assign N565 = N2628;
  assign sent_n[188] = (N566)? 1'b1 : 
                       (N2633)? sent_r[188] : 1'b0;
  assign N566 = N2632;
  assign N2637 = (N567)? 1'b0 : 
                 (N568)? N2636 : 1'b0;
  assign N567 = N2635;
  assign N568 = N2634;
  assign sent_n[189] = (N569)? 1'b1 : 
                       (N2639)? sent_r[189] : 1'b0;
  assign N569 = N2638;
  assign N2643 = (N570)? 1'b0 : 
                 (N571)? N2642 : 1'b0;
  assign N570 = N2641;
  assign N571 = N2640;
  assign sent_n[190] = (N572)? 1'b1 : 
                       (N2645)? sent_r[190] : 1'b0;
  assign N572 = N2644;
  assign N2649 = (N573)? 1'b0 : 
                 (N574)? N2648 : 1'b0;
  assign N573 = N2647;
  assign N574 = N2646;
  assign sent_n[191] = (N575)? 1'b1 : 
                       (N2651)? sent_r[191] : 1'b0;
  assign N575 = N2650;
  assign N2655 = (N576)? 1'b0 : 
                 (N577)? N2654 : 1'b0;
  assign N576 = N2653;
  assign N577 = N2652;
  assign sent_n[192] = (N578)? 1'b1 : 
                       (N2657)? sent_r[192] : 1'b0;
  assign N578 = N2656;
  assign N2661 = (N579)? 1'b0 : 
                 (N580)? N2660 : 1'b0;
  assign N579 = N2659;
  assign N580 = N2658;
  assign sent_n[193] = (N581)? 1'b1 : 
                       (N2663)? sent_r[193] : 1'b0;
  assign N581 = N2662;
  assign N2667 = (N582)? 1'b0 : 
                 (N583)? N2666 : 1'b0;
  assign N582 = N2665;
  assign N583 = N2664;
  assign sent_n[194] = (N584)? 1'b1 : 
                       (N2669)? sent_r[194] : 1'b0;
  assign N584 = N2668;
  assign N2673 = (N585)? 1'b0 : 
                 (N586)? N2672 : 1'b0;
  assign N585 = N2671;
  assign N586 = N2670;
  assign sent_n[195] = (N587)? 1'b1 : 
                       (N2675)? sent_r[195] : 1'b0;
  assign N587 = N2674;
  assign N2679 = (N588)? 1'b0 : 
                 (N589)? N2678 : 1'b0;
  assign N588 = N2677;
  assign N589 = N2676;
  assign sent_n[196] = (N590)? 1'b1 : 
                       (N2681)? sent_r[196] : 1'b0;
  assign N590 = N2680;
  assign N2685 = (N591)? 1'b0 : 
                 (N592)? N2684 : 1'b0;
  assign N591 = N2683;
  assign N592 = N2682;
  assign sent_n[197] = (N593)? 1'b1 : 
                       (N2687)? sent_r[197] : 1'b0;
  assign N593 = N2686;
  assign N2691 = (N594)? 1'b0 : 
                 (N595)? N2690 : 1'b0;
  assign N594 = N2689;
  assign N595 = N2688;
  assign sent_n[198] = (N596)? 1'b1 : 
                       (N2693)? sent_r[198] : 1'b0;
  assign N596 = N2692;
  assign N2697 = (N597)? 1'b0 : 
                 (N598)? N2696 : 1'b0;
  assign N597 = N2695;
  assign N598 = N2694;
  assign sent_n[199] = (N599)? 1'b1 : 
                       (N2699)? sent_r[199] : 1'b0;
  assign N599 = N2698;
  assign N2703 = (N600)? 1'b0 : 
                 (N601)? N2702 : 1'b0;
  assign N600 = N2701;
  assign N601 = N2700;
  assign sent_n[200] = (N602)? 1'b1 : 
                       (N2705)? sent_r[200] : 1'b0;
  assign N602 = N2704;
  assign N2709 = (N603)? 1'b0 : 
                 (N604)? N2708 : 1'b0;
  assign N603 = N2707;
  assign N604 = N2706;
  assign sent_n[201] = (N605)? 1'b1 : 
                       (N2711)? sent_r[201] : 1'b0;
  assign N605 = N2710;
  assign N2715 = (N606)? 1'b0 : 
                 (N607)? N2714 : 1'b0;
  assign N606 = N2713;
  assign N607 = N2712;
  assign sent_n[202] = (N608)? 1'b1 : 
                       (N2717)? sent_r[202] : 1'b0;
  assign N608 = N2716;
  assign N2721 = (N609)? 1'b0 : 
                 (N610)? N2720 : 1'b0;
  assign N609 = N2719;
  assign N610 = N2718;
  assign sent_n[203] = (N611)? 1'b1 : 
                       (N2723)? sent_r[203] : 1'b0;
  assign N611 = N2722;
  assign N2727 = (N612)? 1'b0 : 
                 (N613)? N2726 : 1'b0;
  assign N612 = N2725;
  assign N613 = N2724;
  assign sent_n[204] = (N614)? 1'b1 : 
                       (N2729)? sent_r[204] : 1'b0;
  assign N614 = N2728;
  assign N2733 = (N615)? 1'b0 : 
                 (N616)? N2732 : 1'b0;
  assign N615 = N2731;
  assign N616 = N2730;
  assign sent_n[205] = (N617)? 1'b1 : 
                       (N2735)? sent_r[205] : 1'b0;
  assign N617 = N2734;
  assign N2739 = (N618)? 1'b0 : 
                 (N619)? N2738 : 1'b0;
  assign N618 = N2737;
  assign N619 = N2736;
  assign sent_n[206] = (N620)? 1'b1 : 
                       (N2741)? sent_r[206] : 1'b0;
  assign N620 = N2740;
  assign N2745 = (N621)? 1'b0 : 
                 (N622)? N2744 : 1'b0;
  assign N621 = N2743;
  assign N622 = N2742;
  assign sent_n[207] = (N623)? 1'b1 : 
                       (N2747)? sent_r[207] : 1'b0;
  assign N623 = N2746;
  assign N2751 = (N624)? 1'b0 : 
                 (N625)? N2750 : 1'b0;
  assign N624 = N2749;
  assign N625 = N2748;
  assign sent_n[208] = (N626)? 1'b1 : 
                       (N2753)? sent_r[208] : 1'b0;
  assign N626 = N2752;
  assign N2757 = (N627)? 1'b0 : 
                 (N628)? N2756 : 1'b0;
  assign N627 = N2755;
  assign N628 = N2754;
  assign sent_n[209] = (N629)? 1'b1 : 
                       (N2759)? sent_r[209] : 1'b0;
  assign N629 = N2758;
  assign N2763 = (N630)? 1'b0 : 
                 (N631)? N2762 : 1'b0;
  assign N630 = N2761;
  assign N631 = N2760;
  assign sent_n[210] = (N632)? 1'b1 : 
                       (N2765)? sent_r[210] : 1'b0;
  assign N632 = N2764;
  assign N2769 = (N633)? 1'b0 : 
                 (N634)? N2768 : 1'b0;
  assign N633 = N2767;
  assign N634 = N2766;
  assign sent_n[211] = (N635)? 1'b1 : 
                       (N2771)? sent_r[211] : 1'b0;
  assign N635 = N2770;
  assign N2775 = (N636)? 1'b0 : 
                 (N637)? N2774 : 1'b0;
  assign N636 = N2773;
  assign N637 = N2772;
  assign sent_n[212] = (N638)? 1'b1 : 
                       (N2777)? sent_r[212] : 1'b0;
  assign N638 = N2776;
  assign N2781 = (N639)? 1'b0 : 
                 (N640)? N2780 : 1'b0;
  assign N639 = N2779;
  assign N640 = N2778;
  assign sent_n[213] = (N641)? 1'b1 : 
                       (N2783)? sent_r[213] : 1'b0;
  assign N641 = N2782;
  assign N2787 = (N642)? 1'b0 : 
                 (N643)? N2786 : 1'b0;
  assign N642 = N2785;
  assign N643 = N2784;
  assign sent_n[214] = (N644)? 1'b1 : 
                       (N2789)? sent_r[214] : 1'b0;
  assign N644 = N2788;
  assign N2793 = (N645)? 1'b0 : 
                 (N646)? N2792 : 1'b0;
  assign N645 = N2791;
  assign N646 = N2790;
  assign sent_n[215] = (N647)? 1'b1 : 
                       (N2795)? sent_r[215] : 1'b0;
  assign N647 = N2794;
  assign N2799 = (N648)? 1'b0 : 
                 (N649)? N2798 : 1'b0;
  assign N648 = N2797;
  assign N649 = N2796;
  assign sent_n[216] = (N650)? 1'b1 : 
                       (N2801)? sent_r[216] : 1'b0;
  assign N650 = N2800;
  assign N2805 = (N651)? 1'b0 : 
                 (N652)? N2804 : 1'b0;
  assign N651 = N2803;
  assign N652 = N2802;
  assign sent_n[217] = (N653)? 1'b1 : 
                       (N2807)? sent_r[217] : 1'b0;
  assign N653 = N2806;
  assign N2811 = (N654)? 1'b0 : 
                 (N655)? N2810 : 1'b0;
  assign N654 = N2809;
  assign N655 = N2808;
  assign sent_n[218] = (N656)? 1'b1 : 
                       (N2813)? sent_r[218] : 1'b0;
  assign N656 = N2812;
  assign N2817 = (N657)? 1'b0 : 
                 (N658)? N2816 : 1'b0;
  assign N657 = N2815;
  assign N658 = N2814;
  assign sent_n[219] = (N659)? 1'b1 : 
                       (N2819)? sent_r[219] : 1'b0;
  assign N659 = N2818;
  assign N2823 = (N660)? 1'b0 : 
                 (N661)? N2822 : 1'b0;
  assign N660 = N2821;
  assign N661 = N2820;
  assign sent_n[220] = (N662)? 1'b1 : 
                       (N2825)? sent_r[220] : 1'b0;
  assign N662 = N2824;
  assign N2829 = (N663)? 1'b0 : 
                 (N664)? N2828 : 1'b0;
  assign N663 = N2827;
  assign N664 = N2826;
  assign sent_n[221] = (N665)? 1'b1 : 
                       (N2831)? sent_r[221] : 1'b0;
  assign N665 = N2830;
  assign N2835 = (N666)? 1'b0 : 
                 (N667)? N2834 : 1'b0;
  assign N666 = N2833;
  assign N667 = N2832;
  assign sent_n[222] = (N668)? 1'b1 : 
                       (N2837)? sent_r[222] : 1'b0;
  assign N668 = N2836;
  assign N2841 = (N669)? 1'b0 : 
                 (N670)? N2840 : 1'b0;
  assign N669 = N2839;
  assign N670 = N2838;
  assign sent_n[223] = (N671)? 1'b1 : 
                       (N2843)? sent_r[223] : 1'b0;
  assign N671 = N2842;
  assign N2847 = (N672)? 1'b0 : 
                 (N673)? N2846 : 1'b0;
  assign N672 = N2845;
  assign N673 = N2844;
  assign sent_n[224] = (N674)? 1'b1 : 
                       (N2849)? sent_r[224] : 1'b0;
  assign N674 = N2848;
  assign N2853 = (N675)? 1'b0 : 
                 (N676)? N2852 : 1'b0;
  assign N675 = N2851;
  assign N676 = N2850;
  assign sent_n[225] = (N677)? 1'b1 : 
                       (N2855)? sent_r[225] : 1'b0;
  assign N677 = N2854;
  assign N2859 = (N678)? 1'b0 : 
                 (N679)? N2858 : 1'b0;
  assign N678 = N2857;
  assign N679 = N2856;
  assign sent_n[226] = (N680)? 1'b1 : 
                       (N2861)? sent_r[226] : 1'b0;
  assign N680 = N2860;
  assign N2865 = (N681)? 1'b0 : 
                 (N682)? N2864 : 1'b0;
  assign N681 = N2863;
  assign N682 = N2862;
  assign sent_n[227] = (N683)? 1'b1 : 
                       (N2867)? sent_r[227] : 1'b0;
  assign N683 = N2866;
  assign N2871 = (N684)? 1'b0 : 
                 (N685)? N2870 : 1'b0;
  assign N684 = N2869;
  assign N685 = N2868;
  assign sent_n[228] = (N686)? 1'b1 : 
                       (N2873)? sent_r[228] : 1'b0;
  assign N686 = N2872;
  assign N2877 = (N687)? 1'b0 : 
                 (N688)? N2876 : 1'b0;
  assign N687 = N2875;
  assign N688 = N2874;
  assign sent_n[229] = (N689)? 1'b1 : 
                       (N2879)? sent_r[229] : 1'b0;
  assign N689 = N2878;
  assign N2883 = (N690)? 1'b0 : 
                 (N691)? N2882 : 1'b0;
  assign N690 = N2881;
  assign N691 = N2880;
  assign sent_n[230] = (N692)? 1'b1 : 
                       (N2885)? sent_r[230] : 1'b0;
  assign N692 = N2884;
  assign N2889 = (N693)? 1'b0 : 
                 (N694)? N2888 : 1'b0;
  assign N693 = N2887;
  assign N694 = N2886;
  assign sent_n[231] = (N695)? 1'b1 : 
                       (N2891)? sent_r[231] : 1'b0;
  assign N695 = N2890;
  assign N2895 = (N696)? 1'b0 : 
                 (N697)? N2894 : 1'b0;
  assign N696 = N2893;
  assign N697 = N2892;
  assign sent_n[232] = (N698)? 1'b1 : 
                       (N2897)? sent_r[232] : 1'b0;
  assign N698 = N2896;
  assign N2901 = (N699)? 1'b0 : 
                 (N700)? N2900 : 1'b0;
  assign N699 = N2899;
  assign N700 = N2898;
  assign sent_n[233] = (N701)? 1'b1 : 
                       (N2903)? sent_r[233] : 1'b0;
  assign N701 = N2902;
  assign N2907 = (N702)? 1'b0 : 
                 (N703)? N2906 : 1'b0;
  assign N702 = N2905;
  assign N703 = N2904;
  assign sent_n[234] = (N704)? 1'b1 : 
                       (N2909)? sent_r[234] : 1'b0;
  assign N704 = N2908;
  assign N2913 = (N705)? 1'b0 : 
                 (N706)? N2912 : 1'b0;
  assign N705 = N2911;
  assign N706 = N2910;
  assign sent_n[235] = (N707)? 1'b1 : 
                       (N2915)? sent_r[235] : 1'b0;
  assign N707 = N2914;
  assign N2919 = (N708)? 1'b0 : 
                 (N709)? N2918 : 1'b0;
  assign N708 = N2917;
  assign N709 = N2916;
  assign sent_n[236] = (N710)? 1'b1 : 
                       (N2921)? sent_r[236] : 1'b0;
  assign N710 = N2920;
  assign N2925 = (N711)? 1'b0 : 
                 (N712)? N2924 : 1'b0;
  assign N711 = N2923;
  assign N712 = N2922;
  assign sent_n[237] = (N713)? 1'b1 : 
                       (N2927)? sent_r[237] : 1'b0;
  assign N713 = N2926;
  assign N2931 = (N714)? 1'b0 : 
                 (N715)? N2930 : 1'b0;
  assign N714 = N2929;
  assign N715 = N2928;
  assign sent_n[238] = (N716)? 1'b1 : 
                       (N2933)? sent_r[238] : 1'b0;
  assign N716 = N2932;
  assign N2937 = (N717)? 1'b0 : 
                 (N718)? N2936 : 1'b0;
  assign N717 = N2935;
  assign N718 = N2934;
  assign sent_n[239] = (N719)? 1'b1 : 
                       (N2939)? sent_r[239] : 1'b0;
  assign N719 = N2938;
  assign N2943 = (N720)? 1'b0 : 
                 (N721)? N2942 : 1'b0;
  assign N720 = N2941;
  assign N721 = N2940;
  assign sent_n[240] = (N722)? 1'b1 : 
                       (N2945)? sent_r[240] : 1'b0;
  assign N722 = N2944;
  assign N2949 = (N723)? 1'b0 : 
                 (N724)? N2948 : 1'b0;
  assign N723 = N2947;
  assign N724 = N2946;
  assign sent_n[241] = (N725)? 1'b1 : 
                       (N2951)? sent_r[241] : 1'b0;
  assign N725 = N2950;
  assign N2955 = (N726)? 1'b0 : 
                 (N727)? N2954 : 1'b0;
  assign N726 = N2953;
  assign N727 = N2952;
  assign sent_n[242] = (N728)? 1'b1 : 
                       (N2957)? sent_r[242] : 1'b0;
  assign N728 = N2956;
  assign N2961 = (N729)? 1'b0 : 
                 (N730)? N2960 : 1'b0;
  assign N729 = N2959;
  assign N730 = N2958;
  assign sent_n[243] = (N731)? 1'b1 : 
                       (N2963)? sent_r[243] : 1'b0;
  assign N731 = N2962;
  assign N2967 = (N732)? 1'b0 : 
                 (N733)? N2966 : 1'b0;
  assign N732 = N2965;
  assign N733 = N2964;
  assign sent_n[244] = (N734)? 1'b1 : 
                       (N2969)? sent_r[244] : 1'b0;
  assign N734 = N2968;
  assign N2973 = (N735)? 1'b0 : 
                 (N736)? N2972 : 1'b0;
  assign N735 = N2971;
  assign N736 = N2970;
  assign sent_n[245] = (N737)? 1'b1 : 
                       (N2975)? sent_r[245] : 1'b0;
  assign N737 = N2974;
  assign N2979 = (N738)? 1'b0 : 
                 (N739)? N2978 : 1'b0;
  assign N738 = N2977;
  assign N739 = N2976;
  assign sent_n[246] = (N740)? 1'b1 : 
                       (N2981)? sent_r[246] : 1'b0;
  assign N740 = N2980;
  assign N2985 = (N741)? 1'b0 : 
                 (N742)? N2984 : 1'b0;
  assign N741 = N2983;
  assign N742 = N2982;
  assign sent_n[247] = (N743)? 1'b1 : 
                       (N2987)? sent_r[247] : 1'b0;
  assign N743 = N2986;
  assign N2991 = (N744)? 1'b0 : 
                 (N745)? N2990 : 1'b0;
  assign N744 = N2989;
  assign N745 = N2988;
  assign sent_n[248] = (N746)? 1'b1 : 
                       (N2993)? sent_r[248] : 1'b0;
  assign N746 = N2992;
  assign N2997 = (N747)? 1'b0 : 
                 (N748)? N2996 : 1'b0;
  assign N747 = N2995;
  assign N748 = N2994;
  assign sent_n[249] = (N749)? 1'b1 : 
                       (N2999)? sent_r[249] : 1'b0;
  assign N749 = N2998;
  assign N3003 = (N750)? 1'b0 : 
                 (N751)? N3002 : 1'b0;
  assign N750 = N3001;
  assign N751 = N3000;
  assign sent_n[250] = (N752)? 1'b1 : 
                       (N3005)? sent_r[250] : 1'b0;
  assign N752 = N3004;
  assign N3009 = (N753)? 1'b0 : 
                 (N754)? N3008 : 1'b0;
  assign N753 = N3007;
  assign N754 = N3006;
  assign sent_n[251] = (N755)? 1'b1 : 
                       (N3011)? sent_r[251] : 1'b0;
  assign N755 = N3010;
  assign N3015 = (N756)? 1'b0 : 
                 (N757)? N3014 : 1'b0;
  assign N756 = N3013;
  assign N757 = N3012;
  assign sent_n[252] = (N758)? 1'b1 : 
                       (N3017)? sent_r[252] : 1'b0;
  assign N758 = N3016;
  assign N3021 = (N759)? 1'b0 : 
                 (N760)? N3020 : 1'b0;
  assign N759 = N3019;
  assign N760 = N3018;
  assign sent_n[253] = (N761)? 1'b1 : 
                       (N3023)? sent_r[253] : 1'b0;
  assign N761 = N3022;
  assign N3027 = (N762)? 1'b0 : 
                 (N763)? N3026 : 1'b0;
  assign N762 = N3025;
  assign N763 = N3024;
  assign sent_n[254] = (N764)? 1'b1 : 
                       (N3029)? sent_r[254] : 1'b0;
  assign N764 = N3028;
  assign N3033 = (N765)? 1'b0 : 
                 (N766)? N3032 : 1'b0;
  assign N765 = N3031;
  assign N766 = N3030;
  assign sent_n[255] = (N767)? 1'b1 : 
                       (N3035)? sent_r[255] : 1'b0;
  assign N767 = N3034;
  assign N3039 = (N768)? 1'b0 : 
                 (N769)? N3038 : 1'b0;
  assign N768 = N3037;
  assign N769 = N3036;
  assign sent_n[256] = (N770)? 1'b1 : 
                       (N3041)? sent_r[256] : 1'b0;
  assign N770 = N3040;
  assign N3045 = (N771)? 1'b0 : 
                 (N772)? N3044 : 1'b0;
  assign N771 = N3043;
  assign N772 = N3042;
  assign sent_n[257] = (N773)? 1'b1 : 
                       (N3047)? sent_r[257] : 1'b0;
  assign N773 = N3046;
  assign N3051 = (N774)? 1'b0 : 
                 (N775)? N3050 : 1'b0;
  assign N774 = N3049;
  assign N775 = N3048;
  assign sent_n[258] = (N776)? 1'b1 : 
                       (N3053)? sent_r[258] : 1'b0;
  assign N776 = N3052;
  assign N3057 = (N777)? 1'b0 : 
                 (N778)? N3056 : 1'b0;
  assign N777 = N3055;
  assign N778 = N3054;
  assign sent_n[259] = (N779)? 1'b1 : 
                       (N3059)? sent_r[259] : 1'b0;
  assign N779 = N3058;
  assign N3063 = (N780)? 1'b0 : 
                 (N781)? N3062 : 1'b0;
  assign N780 = N3061;
  assign N781 = N3060;
  assign sent_n[260] = (N782)? 1'b1 : 
                       (N3065)? sent_r[260] : 1'b0;
  assign N782 = N3064;
  assign N3069 = (N783)? 1'b0 : 
                 (N784)? N3068 : 1'b0;
  assign N783 = N3067;
  assign N784 = N3066;
  assign sent_n[261] = (N785)? 1'b1 : 
                       (N3071)? sent_r[261] : 1'b0;
  assign N785 = N3070;
  assign N3075 = (N786)? 1'b0 : 
                 (N787)? N3074 : 1'b0;
  assign N786 = N3073;
  assign N787 = N3072;
  assign sent_n[262] = (N788)? 1'b1 : 
                       (N3077)? sent_r[262] : 1'b0;
  assign N788 = N3076;
  assign N3081 = (N789)? 1'b0 : 
                 (N790)? N3080 : 1'b0;
  assign N789 = N3079;
  assign N790 = N3078;
  assign sent_n[263] = (N791)? 1'b1 : 
                       (N3083)? sent_r[263] : 1'b0;
  assign N791 = N3082;
  assign N3087 = (N792)? 1'b0 : 
                 (N793)? N3086 : 1'b0;
  assign N792 = N3085;
  assign N793 = N3084;
  assign sent_n[264] = (N794)? 1'b1 : 
                       (N3089)? sent_r[264] : 1'b0;
  assign N794 = N3088;
  assign N3093 = (N795)? 1'b0 : 
                 (N796)? N3092 : 1'b0;
  assign N795 = N3091;
  assign N796 = N3090;
  assign sent_n[265] = (N797)? 1'b1 : 
                       (N3095)? sent_r[265] : 1'b0;
  assign N797 = N3094;
  assign N3099 = (N798)? 1'b0 : 
                 (N799)? N3098 : 1'b0;
  assign N798 = N3097;
  assign N799 = N3096;
  assign sent_n[266] = (N800)? 1'b1 : 
                       (N3101)? sent_r[266] : 1'b0;
  assign N800 = N3100;
  assign N3105 = (N801)? 1'b0 : 
                 (N802)? N3104 : 1'b0;
  assign N801 = N3103;
  assign N802 = N3102;
  assign sent_n[267] = (N803)? 1'b1 : 
                       (N3107)? sent_r[267] : 1'b0;
  assign N803 = N3106;
  assign N3111 = (N804)? 1'b0 : 
                 (N805)? N3110 : 1'b0;
  assign N804 = N3109;
  assign N805 = N3108;
  assign sent_n[268] = (N806)? 1'b1 : 
                       (N3113)? sent_r[268] : 1'b0;
  assign N806 = N3112;
  assign N3117 = (N807)? 1'b0 : 
                 (N808)? N3116 : 1'b0;
  assign N807 = N3115;
  assign N808 = N3114;
  assign sent_n[269] = (N809)? 1'b1 : 
                       (N3119)? sent_r[269] : 1'b0;
  assign N809 = N3118;
  assign N3123 = (N810)? 1'b0 : 
                 (N811)? N3122 : 1'b0;
  assign N810 = N3121;
  assign N811 = N3120;
  assign sent_n[270] = (N812)? 1'b1 : 
                       (N3125)? sent_r[270] : 1'b0;
  assign N812 = N3124;
  assign N3129 = (N813)? 1'b0 : 
                 (N814)? N3128 : 1'b0;
  assign N813 = N3127;
  assign N814 = N3126;
  assign sent_n[271] = (N815)? 1'b1 : 
                       (N3131)? sent_r[271] : 1'b0;
  assign N815 = N3130;
  assign N3135 = (N816)? 1'b0 : 
                 (N817)? N3134 : 1'b0;
  assign N816 = N3133;
  assign N817 = N3132;
  assign sent_n[272] = (N818)? 1'b1 : 
                       (N3137)? sent_r[272] : 1'b0;
  assign N818 = N3136;
  assign N3141 = (N819)? 1'b0 : 
                 (N820)? N3140 : 1'b0;
  assign N819 = N3139;
  assign N820 = N3138;
  assign sent_n[273] = (N821)? 1'b1 : 
                       (N3143)? sent_r[273] : 1'b0;
  assign N821 = N3142;
  assign N3147 = (N822)? 1'b0 : 
                 (N823)? N3146 : 1'b0;
  assign N822 = N3145;
  assign N823 = N3144;
  assign sent_n[274] = (N824)? 1'b1 : 
                       (N3149)? sent_r[274] : 1'b0;
  assign N824 = N3148;
  assign N3153 = (N825)? 1'b0 : 
                 (N826)? N3152 : 1'b0;
  assign N825 = N3151;
  assign N826 = N3150;
  assign sent_n[275] = (N827)? 1'b1 : 
                       (N3155)? sent_r[275] : 1'b0;
  assign N827 = N3154;
  assign N3159 = (N828)? 1'b0 : 
                 (N829)? N3158 : 1'b0;
  assign N828 = N3157;
  assign N829 = N3156;
  assign sent_n[276] = (N830)? 1'b1 : 
                       (N3161)? sent_r[276] : 1'b0;
  assign N830 = N3160;
  assign N3165 = (N831)? 1'b0 : 
                 (N832)? N3164 : 1'b0;
  assign N831 = N3163;
  assign N832 = N3162;
  assign sent_n[277] = (N833)? 1'b1 : 
                       (N3167)? sent_r[277] : 1'b0;
  assign N833 = N3166;
  assign N3171 = (N834)? 1'b0 : 
                 (N835)? N3170 : 1'b0;
  assign N834 = N3169;
  assign N835 = N3168;
  assign sent_n[278] = (N836)? 1'b1 : 
                       (N3173)? sent_r[278] : 1'b0;
  assign N836 = N3172;
  assign N3177 = (N837)? 1'b0 : 
                 (N838)? N3176 : 1'b0;
  assign N837 = N3175;
  assign N838 = N3174;
  assign sent_n[279] = (N839)? 1'b1 : 
                       (N3179)? sent_r[279] : 1'b0;
  assign N839 = N3178;
  assign N3183 = (N840)? 1'b0 : 
                 (N841)? N3182 : 1'b0;
  assign N840 = N3181;
  assign N841 = N3180;
  assign sent_n[280] = (N842)? 1'b1 : 
                       (N3185)? sent_r[280] : 1'b0;
  assign N842 = N3184;
  assign N3189 = (N843)? 1'b0 : 
                 (N844)? N3188 : 1'b0;
  assign N843 = N3187;
  assign N844 = N3186;
  assign sent_n[281] = (N845)? 1'b1 : 
                       (N3191)? sent_r[281] : 1'b0;
  assign N845 = N3190;
  assign N3195 = (N846)? 1'b0 : 
                 (N847)? N3194 : 1'b0;
  assign N846 = N3193;
  assign N847 = N3192;
  assign sent_n[282] = (N848)? 1'b1 : 
                       (N3197)? sent_r[282] : 1'b0;
  assign N848 = N3196;
  assign N3201 = (N849)? 1'b0 : 
                 (N850)? N3200 : 1'b0;
  assign N849 = N3199;
  assign N850 = N3198;
  assign sent_n[283] = (N851)? 1'b1 : 
                       (N3203)? sent_r[283] : 1'b0;
  assign N851 = N3202;
  assign N3207 = (N852)? 1'b0 : 
                 (N853)? N3206 : 1'b0;
  assign N852 = N3205;
  assign N853 = N3204;
  assign sent_n[284] = (N854)? 1'b1 : 
                       (N3209)? sent_r[284] : 1'b0;
  assign N854 = N3208;
  assign N3213 = (N855)? 1'b0 : 
                 (N856)? N3212 : 1'b0;
  assign N855 = N3211;
  assign N856 = N3210;
  assign sent_n[285] = (N857)? 1'b1 : 
                       (N3215)? sent_r[285] : 1'b0;
  assign N857 = N3214;
  assign N3219 = (N858)? 1'b0 : 
                 (N859)? N3218 : 1'b0;
  assign N858 = N3217;
  assign N859 = N3216;
  assign sent_n[286] = (N860)? 1'b1 : 
                       (N3221)? sent_r[286] : 1'b0;
  assign N860 = N3220;
  assign N3225 = (N861)? 1'b0 : 
                 (N862)? N3224 : 1'b0;
  assign N861 = N3223;
  assign N862 = N3222;
  assign sent_n[287] = (N863)? 1'b1 : 
                       (N3227)? sent_r[287] : 1'b0;
  assign N863 = N3226;
  assign N3231 = (N864)? 1'b0 : 
                 (N865)? N3230 : 1'b0;
  assign N864 = N3229;
  assign N865 = N3228;
  assign sent_n[288] = (N866)? 1'b1 : 
                       (N3233)? sent_r[288] : 1'b0;
  assign N866 = N3232;
  assign N3237 = (N867)? 1'b0 : 
                 (N868)? N3236 : 1'b0;
  assign N867 = N3235;
  assign N868 = N3234;
  assign sent_n[289] = (N869)? 1'b1 : 
                       (N3239)? sent_r[289] : 1'b0;
  assign N869 = N3238;
  assign N3243 = (N870)? 1'b0 : 
                 (N871)? N3242 : 1'b0;
  assign N870 = N3241;
  assign N871 = N3240;
  assign sent_n[290] = (N872)? 1'b1 : 
                       (N3245)? sent_r[290] : 1'b0;
  assign N872 = N3244;
  assign N3249 = (N873)? 1'b0 : 
                 (N874)? N3248 : 1'b0;
  assign N873 = N3247;
  assign N874 = N3246;
  assign sent_n[291] = (N875)? 1'b1 : 
                       (N3251)? sent_r[291] : 1'b0;
  assign N875 = N3250;
  assign N3255 = (N876)? 1'b0 : 
                 (N877)? N3254 : 1'b0;
  assign N876 = N3253;
  assign N877 = N3252;
  assign sent_n[292] = (N878)? 1'b1 : 
                       (N3257)? sent_r[292] : 1'b0;
  assign N878 = N3256;
  assign N3261 = (N879)? 1'b0 : 
                 (N880)? N3260 : 1'b0;
  assign N879 = N3259;
  assign N880 = N3258;
  assign sent_n[293] = (N881)? 1'b1 : 
                       (N3263)? sent_r[293] : 1'b0;
  assign N881 = N3262;
  assign N3267 = (N882)? 1'b0 : 
                 (N883)? N3266 : 1'b0;
  assign N882 = N3265;
  assign N883 = N3264;
  assign sent_n[294] = (N884)? 1'b1 : 
                       (N3269)? sent_r[294] : 1'b0;
  assign N884 = N3268;
  assign N3273 = (N885)? 1'b0 : 
                 (N886)? N3272 : 1'b0;
  assign N885 = N3271;
  assign N886 = N3270;
  assign sent_n[295] = (N887)? 1'b1 : 
                       (N3275)? sent_r[295] : 1'b0;
  assign N887 = N3274;
  assign N3279 = (N888)? 1'b0 : 
                 (N889)? N3278 : 1'b0;
  assign N888 = N3277;
  assign N889 = N3276;
  assign sent_n[296] = (N890)? 1'b1 : 
                       (N3281)? sent_r[296] : 1'b0;
  assign N890 = N3280;
  assign N3285 = (N891)? 1'b0 : 
                 (N892)? N3284 : 1'b0;
  assign N891 = N3283;
  assign N892 = N3282;
  assign sent_n[297] = (N893)? 1'b1 : 
                       (N3287)? sent_r[297] : 1'b0;
  assign N893 = N3286;
  assign N3291 = (N894)? 1'b0 : 
                 (N895)? N3290 : 1'b0;
  assign N894 = N3289;
  assign N895 = N3288;
  assign sent_n[298] = (N896)? 1'b1 : 
                       (N3293)? sent_r[298] : 1'b0;
  assign N896 = N3292;
  assign N3297 = (N897)? 1'b0 : 
                 (N898)? N3296 : 1'b0;
  assign N897 = N3295;
  assign N898 = N3294;
  assign sent_n[299] = (N899)? 1'b1 : 
                       (N3299)? sent_r[299] : 1'b0;
  assign N899 = N3298;
  assign N3303 = (N900)? 1'b0 : 
                 (N901)? N3302 : 1'b0;
  assign N900 = N3301;
  assign N901 = N3300;
  assign sent_n[300] = (N902)? 1'b1 : 
                       (N3305)? sent_r[300] : 1'b0;
  assign N902 = N3304;
  assign N3309 = (N903)? 1'b0 : 
                 (N904)? N3308 : 1'b0;
  assign N903 = N3307;
  assign N904 = N3306;
  assign sent_n[301] = (N905)? 1'b1 : 
                       (N3311)? sent_r[301] : 1'b0;
  assign N905 = N3310;
  assign N3315 = (N906)? 1'b0 : 
                 (N907)? N3314 : 1'b0;
  assign N906 = N3313;
  assign N907 = N3312;
  assign sent_n[302] = (N908)? 1'b1 : 
                       (N3317)? sent_r[302] : 1'b0;
  assign N908 = N3316;
  assign N3321 = (N909)? 1'b0 : 
                 (N910)? N3320 : 1'b0;
  assign N909 = N3319;
  assign N910 = N3318;
  assign sent_n[303] = (N911)? 1'b1 : 
                       (N3323)? sent_r[303] : 1'b0;
  assign N911 = N3322;
  assign N3327 = (N912)? 1'b0 : 
                 (N913)? N3326 : 1'b0;
  assign N912 = N3325;
  assign N913 = N3324;
  assign sent_n[304] = (N914)? 1'b1 : 
                       (N3329)? sent_r[304] : 1'b0;
  assign N914 = N3328;
  assign N3333 = (N915)? 1'b0 : 
                 (N916)? N3332 : 1'b0;
  assign N915 = N3331;
  assign N916 = N3330;
  assign sent_n[305] = (N917)? 1'b1 : 
                       (N3335)? sent_r[305] : 1'b0;
  assign N917 = N3334;
  assign N3339 = (N918)? 1'b0 : 
                 (N919)? N3338 : 1'b0;
  assign N918 = N3337;
  assign N919 = N3336;
  assign sent_n[306] = (N920)? 1'b1 : 
                       (N3341)? sent_r[306] : 1'b0;
  assign N920 = N3340;
  assign N3345 = (N921)? 1'b0 : 
                 (N922)? N3344 : 1'b0;
  assign N921 = N3343;
  assign N922 = N3342;
  assign sent_n[307] = (N923)? 1'b1 : 
                       (N3347)? sent_r[307] : 1'b0;
  assign N923 = N3346;
  assign N3351 = (N924)? 1'b0 : 
                 (N925)? N3350 : 1'b0;
  assign N924 = N3349;
  assign N925 = N3348;
  assign sent_n[308] = (N926)? 1'b1 : 
                       (N3353)? sent_r[308] : 1'b0;
  assign N926 = N3352;
  assign N3357 = (N927)? 1'b0 : 
                 (N928)? N3356 : 1'b0;
  assign N927 = N3355;
  assign N928 = N3354;
  assign sent_n[309] = (N929)? 1'b1 : 
                       (N3359)? sent_r[309] : 1'b0;
  assign N929 = N3358;
  assign N3363 = (N930)? 1'b0 : 
                 (N931)? N3362 : 1'b0;
  assign N930 = N3361;
  assign N931 = N3360;
  assign sent_n[310] = (N932)? 1'b1 : 
                       (N3365)? sent_r[310] : 1'b0;
  assign N932 = N3364;
  assign N3369 = (N933)? 1'b0 : 
                 (N934)? N3368 : 1'b0;
  assign N933 = N3367;
  assign N934 = N3366;
  assign sent_n[311] = (N935)? 1'b1 : 
                       (N3371)? sent_r[311] : 1'b0;
  assign N935 = N3370;
  assign N3375 = (N936)? 1'b0 : 
                 (N937)? N3374 : 1'b0;
  assign N936 = N3373;
  assign N937 = N3372;
  assign sent_n[312] = (N938)? 1'b1 : 
                       (N3377)? sent_r[312] : 1'b0;
  assign N938 = N3376;
  assign N3381 = (N939)? 1'b0 : 
                 (N940)? N3380 : 1'b0;
  assign N939 = N3379;
  assign N940 = N3378;
  assign sent_n[313] = (N941)? 1'b1 : 
                       (N3383)? sent_r[313] : 1'b0;
  assign N941 = N3382;
  assign N3387 = (N942)? 1'b0 : 
                 (N943)? N3386 : 1'b0;
  assign N942 = N3385;
  assign N943 = N3384;
  assign sent_n[314] = (N944)? 1'b1 : 
                       (N3389)? sent_r[314] : 1'b0;
  assign N944 = N3388;
  assign N3393 = (N945)? 1'b0 : 
                 (N946)? N3392 : 1'b0;
  assign N945 = N3391;
  assign N946 = N3390;
  assign sent_n[315] = (N947)? 1'b1 : 
                       (N3395)? sent_r[315] : 1'b0;
  assign N947 = N3394;
  assign N3399 = (N948)? 1'b0 : 
                 (N949)? N3398 : 1'b0;
  assign N948 = N3397;
  assign N949 = N3396;
  assign sent_n[316] = (N950)? 1'b1 : 
                       (N3401)? sent_r[316] : 1'b0;
  assign N950 = N3400;
  assign N3405 = (N951)? 1'b0 : 
                 (N952)? N3404 : 1'b0;
  assign N951 = N3403;
  assign N952 = N3402;
  assign sent_n[317] = (N953)? 1'b1 : 
                       (N3407)? sent_r[317] : 1'b0;
  assign N953 = N3406;
  assign N3411 = (N954)? 1'b0 : 
                 (N955)? N3410 : 1'b0;
  assign N954 = N3409;
  assign N955 = N3408;
  assign sent_n[318] = (N956)? 1'b1 : 
                       (N3413)? sent_r[318] : 1'b0;
  assign N956 = N3412;
  assign N3417 = (N957)? 1'b0 : 
                 (N958)? N3416 : 1'b0;
  assign N957 = N3415;
  assign N958 = N3414;
  assign sent_n[319] = (N959)? 1'b1 : 
                       (N3419)? sent_r[319] : 1'b0;
  assign N959 = N3418;
  assign N3423 = (N960)? 1'b0 : 
                 (N961)? N3422 : 1'b0;
  assign N960 = N3421;
  assign N961 = N3420;
  assign sent_n[320] = (N962)? 1'b1 : 
                       (N3425)? sent_r[320] : 1'b0;
  assign N962 = N3424;
  assign N3429 = (N963)? 1'b0 : 
                 (N964)? N3428 : 1'b0;
  assign N963 = N3427;
  assign N964 = N3426;
  assign sent_n[321] = (N965)? 1'b1 : 
                       (N3431)? sent_r[321] : 1'b0;
  assign N965 = N3430;
  assign N3435 = (N966)? 1'b0 : 
                 (N967)? N3434 : 1'b0;
  assign N966 = N3433;
  assign N967 = N3432;
  assign sent_n[322] = (N968)? 1'b1 : 
                       (N3437)? sent_r[322] : 1'b0;
  assign N968 = N3436;
  assign N3441 = (N969)? 1'b0 : 
                 (N970)? N3440 : 1'b0;
  assign N969 = N3439;
  assign N970 = N3438;
  assign sent_n[323] = (N971)? 1'b1 : 
                       (N3443)? sent_r[323] : 1'b0;
  assign N971 = N3442;
  assign N3447 = (N972)? 1'b0 : 
                 (N973)? N3446 : 1'b0;
  assign N972 = N3445;
  assign N973 = N3444;
  assign sent_n[324] = (N974)? 1'b1 : 
                       (N3449)? sent_r[324] : 1'b0;
  assign N974 = N3448;
  assign N3453 = (N975)? 1'b0 : 
                 (N976)? N3452 : 1'b0;
  assign N975 = N3451;
  assign N976 = N3450;
  assign sent_n[325] = (N977)? 1'b1 : 
                       (N3455)? sent_r[325] : 1'b0;
  assign N977 = N3454;
  assign N3459 = (N978)? 1'b0 : 
                 (N979)? N3458 : 1'b0;
  assign N978 = N3457;
  assign N979 = N3456;
  assign sent_n[326] = (N980)? 1'b1 : 
                       (N3461)? sent_r[326] : 1'b0;
  assign N980 = N3460;
  assign N3465 = (N981)? 1'b0 : 
                 (N982)? N3464 : 1'b0;
  assign N981 = N3463;
  assign N982 = N3462;
  assign sent_n[327] = (N983)? 1'b1 : 
                       (N3467)? sent_r[327] : 1'b0;
  assign N983 = N3466;
  assign N3471 = (N984)? 1'b0 : 
                 (N985)? N3470 : 1'b0;
  assign N984 = N3469;
  assign N985 = N3468;
  assign sent_n[328] = (N986)? 1'b1 : 
                       (N3473)? sent_r[328] : 1'b0;
  assign N986 = N3472;
  assign N3477 = (N987)? 1'b0 : 
                 (N988)? N3476 : 1'b0;
  assign N987 = N3475;
  assign N988 = N3474;
  assign sent_n[329] = (N989)? 1'b1 : 
                       (N3479)? sent_r[329] : 1'b0;
  assign N989 = N3478;
  assign N3483 = (N990)? 1'b0 : 
                 (N991)? N3482 : 1'b0;
  assign N990 = N3481;
  assign N991 = N3480;
  assign sent_n[330] = (N992)? 1'b1 : 
                       (N3485)? sent_r[330] : 1'b0;
  assign N992 = N3484;
  assign N3489 = (N993)? 1'b0 : 
                 (N994)? N3488 : 1'b0;
  assign N993 = N3487;
  assign N994 = N3486;
  assign sent_n[331] = (N995)? 1'b1 : 
                       (N3491)? sent_r[331] : 1'b0;
  assign N995 = N3490;
  assign N3495 = (N996)? 1'b0 : 
                 (N997)? N3494 : 1'b0;
  assign N996 = N3493;
  assign N997 = N3492;
  assign sent_n[332] = (N998)? 1'b1 : 
                       (N3497)? sent_r[332] : 1'b0;
  assign N998 = N3496;
  assign N3501 = (N999)? 1'b0 : 
                 (N1000)? N3500 : 1'b0;
  assign N999 = N3499;
  assign N1000 = N3498;
  assign sent_n[333] = (N1001)? 1'b1 : 
                       (N3503)? sent_r[333] : 1'b0;
  assign N1001 = N3502;
  assign N3507 = (N1002)? 1'b0 : 
                 (N1003)? N3506 : 1'b0;
  assign N1002 = N3505;
  assign N1003 = N3504;
  assign sent_n[334] = (N1004)? 1'b1 : 
                       (N3509)? sent_r[334] : 1'b0;
  assign N1004 = N3508;
  assign N3513 = (N1005)? 1'b0 : 
                 (N1006)? N3512 : 1'b0;
  assign N1005 = N3511;
  assign N1006 = N3510;
  assign sent_n[335] = (N1007)? 1'b1 : 
                       (N3515)? sent_r[335] : 1'b0;
  assign N1007 = N3514;
  assign N3519 = (N1008)? 1'b0 : 
                 (N1009)? N3518 : 1'b0;
  assign N1008 = N3517;
  assign N1009 = N3516;
  assign sent_n[336] = (N1010)? 1'b1 : 
                       (N3521)? sent_r[336] : 1'b0;
  assign N1010 = N3520;
  assign N3525 = (N1011)? 1'b0 : 
                 (N1012)? N3524 : 1'b0;
  assign N1011 = N3523;
  assign N1012 = N3522;
  assign sent_n[337] = (N1013)? 1'b1 : 
                       (N3527)? sent_r[337] : 1'b0;
  assign N1013 = N3526;
  assign N3531 = (N1014)? 1'b0 : 
                 (N1015)? N3530 : 1'b0;
  assign N1014 = N3529;
  assign N1015 = N3528;
  assign sent_n[338] = (N1016)? 1'b1 : 
                       (N3533)? sent_r[338] : 1'b0;
  assign N1016 = N3532;
  assign N3537 = (N1017)? 1'b0 : 
                 (N1018)? N3536 : 1'b0;
  assign N1017 = N3535;
  assign N1018 = N3534;
  assign sent_n[339] = (N1019)? 1'b1 : 
                       (N3539)? sent_r[339] : 1'b0;
  assign N1019 = N3538;
  assign N3543 = (N1020)? 1'b0 : 
                 (N1021)? N3542 : 1'b0;
  assign N1020 = N3541;
  assign N1021 = N3540;
  assign sent_n[340] = (N1022)? 1'b1 : 
                       (N3545)? sent_r[340] : 1'b0;
  assign N1022 = N3544;
  assign N3549 = (N1023)? 1'b0 : 
                 (N1024)? N3548 : 1'b0;
  assign N1023 = N3547;
  assign N1024 = N3546;
  assign sent_n[341] = (N1025)? 1'b1 : 
                       (N3551)? sent_r[341] : 1'b0;
  assign N1025 = N3550;
  assign N3555 = (N1026)? 1'b0 : 
                 (N1027)? N3554 : 1'b0;
  assign N1026 = N3553;
  assign N1027 = N3552;
  assign sent_n[342] = (N1028)? 1'b1 : 
                       (N3557)? sent_r[342] : 1'b0;
  assign N1028 = N3556;
  assign N3561 = (N1029)? 1'b0 : 
                 (N1030)? N3560 : 1'b0;
  assign N1029 = N3559;
  assign N1030 = N3558;
  assign sent_n[343] = (N1031)? 1'b1 : 
                       (N3563)? sent_r[343] : 1'b0;
  assign N1031 = N3562;
  assign N3567 = (N1032)? 1'b0 : 
                 (N1033)? N3566 : 1'b0;
  assign N1032 = N3565;
  assign N1033 = N3564;
  assign sent_n[344] = (N1034)? 1'b1 : 
                       (N3569)? sent_r[344] : 1'b0;
  assign N1034 = N3568;
  assign N3573 = (N1035)? 1'b0 : 
                 (N1036)? N3572 : 1'b0;
  assign N1035 = N3571;
  assign N1036 = N3570;
  assign sent_n[345] = (N1037)? 1'b1 : 
                       (N3575)? sent_r[345] : 1'b0;
  assign N1037 = N3574;
  assign N3579 = (N1038)? 1'b0 : 
                 (N1039)? N3578 : 1'b0;
  assign N1038 = N3577;
  assign N1039 = N3576;
  assign sent_n[346] = (N1040)? 1'b1 : 
                       (N3581)? sent_r[346] : 1'b0;
  assign N1040 = N3580;
  assign N3585 = (N1041)? 1'b0 : 
                 (N1042)? N3584 : 1'b0;
  assign N1041 = N3583;
  assign N1042 = N3582;
  assign sent_n[347] = (N1043)? 1'b1 : 
                       (N3587)? sent_r[347] : 1'b0;
  assign N1043 = N3586;
  assign N3591 = (N1044)? 1'b0 : 
                 (N1045)? N3590 : 1'b0;
  assign N1044 = N3589;
  assign N1045 = N3588;
  assign sent_n[348] = (N1046)? 1'b1 : 
                       (N3593)? sent_r[348] : 1'b0;
  assign N1046 = N3592;
  assign N3597 = (N1047)? 1'b0 : 
                 (N1048)? N3596 : 1'b0;
  assign N1047 = N3595;
  assign N1048 = N3594;
  assign sent_n[349] = (N1049)? 1'b1 : 
                       (N3599)? sent_r[349] : 1'b0;
  assign N1049 = N3598;
  assign N3603 = (N1050)? 1'b0 : 
                 (N1051)? N3602 : 1'b0;
  assign N1050 = N3601;
  assign N1051 = N3600;
  assign sent_n[350] = (N1052)? 1'b1 : 
                       (N3605)? sent_r[350] : 1'b0;
  assign N1052 = N3604;
  assign N3609 = (N1053)? 1'b0 : 
                 (N1054)? N3608 : 1'b0;
  assign N1053 = N3607;
  assign N1054 = N3606;
  assign sent_n[351] = (N1055)? 1'b1 : 
                       (N3611)? sent_r[351] : 1'b0;
  assign N1055 = N3610;
  assign N3615 = (N1056)? 1'b0 : 
                 (N1057)? N3614 : 1'b0;
  assign N1056 = N3613;
  assign N1057 = N3612;
  assign sent_n[352] = (N1058)? 1'b1 : 
                       (N3617)? sent_r[352] : 1'b0;
  assign N1058 = N3616;
  assign N3621 = (N1059)? 1'b0 : 
                 (N1060)? N3620 : 1'b0;
  assign N1059 = N3619;
  assign N1060 = N3618;
  assign sent_n[353] = (N1061)? 1'b1 : 
                       (N3623)? sent_r[353] : 1'b0;
  assign N1061 = N3622;
  assign N3627 = (N1062)? 1'b0 : 
                 (N1063)? N3626 : 1'b0;
  assign N1062 = N3625;
  assign N1063 = N3624;
  assign sent_n[354] = (N1064)? 1'b1 : 
                       (N3629)? sent_r[354] : 1'b0;
  assign N1064 = N3628;
  assign N3633 = (N1065)? 1'b0 : 
                 (N1066)? N3632 : 1'b0;
  assign N1065 = N3631;
  assign N1066 = N3630;
  assign sent_n[355] = (N1067)? 1'b1 : 
                       (N3635)? sent_r[355] : 1'b0;
  assign N1067 = N3634;
  assign N3639 = (N1068)? 1'b0 : 
                 (N1069)? N3638 : 1'b0;
  assign N1068 = N3637;
  assign N1069 = N3636;
  assign sent_n[356] = (N1070)? 1'b1 : 
                       (N3641)? sent_r[356] : 1'b0;
  assign N1070 = N3640;
  assign N3645 = (N1071)? 1'b0 : 
                 (N1072)? N3644 : 1'b0;
  assign N1071 = N3643;
  assign N1072 = N3642;
  assign sent_n[357] = (N1073)? 1'b1 : 
                       (N3647)? sent_r[357] : 1'b0;
  assign N1073 = N3646;
  assign N3651 = (N1074)? 1'b0 : 
                 (N1075)? N3650 : 1'b0;
  assign N1074 = N3649;
  assign N1075 = N3648;
  assign sent_n[358] = (N1076)? 1'b1 : 
                       (N3653)? sent_r[358] : 1'b0;
  assign N1076 = N3652;
  assign N3657 = (N1077)? 1'b0 : 
                 (N1078)? N3656 : 1'b0;
  assign N1077 = N3655;
  assign N1078 = N3654;
  assign sent_n[359] = (N1079)? 1'b1 : 
                       (N3659)? sent_r[359] : 1'b0;
  assign N1079 = N3658;
  assign N3663 = (N1080)? 1'b0 : 
                 (N1081)? N3662 : 1'b0;
  assign N1080 = N3661;
  assign N1081 = N3660;
  assign sent_n[360] = (N1082)? 1'b1 : 
                       (N3665)? sent_r[360] : 1'b0;
  assign N1082 = N3664;
  assign N3669 = (N1083)? 1'b0 : 
                 (N1084)? N3668 : 1'b0;
  assign N1083 = N3667;
  assign N1084 = N3666;
  assign sent_n[361] = (N1085)? 1'b1 : 
                       (N3671)? sent_r[361] : 1'b0;
  assign N1085 = N3670;
  assign N3675 = (N1086)? 1'b0 : 
                 (N1087)? N3674 : 1'b0;
  assign N1086 = N3673;
  assign N1087 = N3672;
  assign sent_n[362] = (N1088)? 1'b1 : 
                       (N3677)? sent_r[362] : 1'b0;
  assign N1088 = N3676;
  assign N3681 = (N1089)? 1'b0 : 
                 (N1090)? N3680 : 1'b0;
  assign N1089 = N3679;
  assign N1090 = N3678;
  assign sent_n[363] = (N1091)? 1'b1 : 
                       (N3683)? sent_r[363] : 1'b0;
  assign N1091 = N3682;
  assign N3687 = (N1092)? 1'b0 : 
                 (N1093)? N3686 : 1'b0;
  assign N1092 = N3685;
  assign N1093 = N3684;
  assign sent_n[364] = (N1094)? 1'b1 : 
                       (N3689)? sent_r[364] : 1'b0;
  assign N1094 = N3688;
  assign N3693 = (N1095)? 1'b0 : 
                 (N1096)? N3692 : 1'b0;
  assign N1095 = N3691;
  assign N1096 = N3690;
  assign sent_n[365] = (N1097)? 1'b1 : 
                       (N3695)? sent_r[365] : 1'b0;
  assign N1097 = N3694;
  assign N3699 = (N1098)? 1'b0 : 
                 (N1099)? N3698 : 1'b0;
  assign N1098 = N3697;
  assign N1099 = N3696;
  assign sent_n[366] = (N1100)? 1'b1 : 
                       (N3701)? sent_r[366] : 1'b0;
  assign N1100 = N3700;
  assign N3705 = (N1101)? 1'b0 : 
                 (N1102)? N3704 : 1'b0;
  assign N1101 = N3703;
  assign N1102 = N3702;
  assign sent_n[367] = (N1103)? 1'b1 : 
                       (N3707)? sent_r[367] : 1'b0;
  assign N1103 = N3706;
  assign N3711 = (N1104)? 1'b0 : 
                 (N1105)? N3710 : 1'b0;
  assign N1104 = N3709;
  assign N1105 = N3708;
  assign sent_n[368] = (N1106)? 1'b1 : 
                       (N3713)? sent_r[368] : 1'b0;
  assign N1106 = N3712;
  assign N3717 = (N1107)? 1'b0 : 
                 (N1108)? N3716 : 1'b0;
  assign N1107 = N3715;
  assign N1108 = N3714;
  assign sent_n[369] = (N1109)? 1'b1 : 
                       (N3719)? sent_r[369] : 1'b0;
  assign N1109 = N3718;
  assign N3723 = (N1110)? 1'b0 : 
                 (N1111)? N3722 : 1'b0;
  assign N1110 = N3721;
  assign N1111 = N3720;
  assign sent_n[370] = (N1112)? 1'b1 : 
                       (N3725)? sent_r[370] : 1'b0;
  assign N1112 = N3724;
  assign N3729 = (N1113)? 1'b0 : 
                 (N1114)? N3728 : 1'b0;
  assign N1113 = N3727;
  assign N1114 = N3726;
  assign sent_n[371] = (N1115)? 1'b1 : 
                       (N3731)? sent_r[371] : 1'b0;
  assign N1115 = N3730;
  assign N3735 = (N1116)? 1'b0 : 
                 (N1117)? N3734 : 1'b0;
  assign N1116 = N3733;
  assign N1117 = N3732;
  assign sent_n[372] = (N1118)? 1'b1 : 
                       (N3737)? sent_r[372] : 1'b0;
  assign N1118 = N3736;
  assign N3741 = (N1119)? 1'b0 : 
                 (N1120)? N3740 : 1'b0;
  assign N1119 = N3739;
  assign N1120 = N3738;
  assign sent_n[373] = (N1121)? 1'b1 : 
                       (N3743)? sent_r[373] : 1'b0;
  assign N1121 = N3742;
  assign N3747 = (N1122)? 1'b0 : 
                 (N1123)? N3746 : 1'b0;
  assign N1122 = N3745;
  assign N1123 = N3744;
  assign sent_n[374] = (N1124)? 1'b1 : 
                       (N3749)? sent_r[374] : 1'b0;
  assign N1124 = N3748;
  assign N3753 = (N1125)? 1'b0 : 
                 (N1126)? N3752 : 1'b0;
  assign N1125 = N3751;
  assign N1126 = N3750;
  assign sent_n[375] = (N1127)? 1'b1 : 
                       (N3755)? sent_r[375] : 1'b0;
  assign N1127 = N3754;
  assign N3759 = (N1128)? 1'b0 : 
                 (N1129)? N3758 : 1'b0;
  assign N1128 = N3757;
  assign N1129 = N3756;
  assign sent_n[376] = (N1130)? 1'b1 : 
                       (N3761)? sent_r[376] : 1'b0;
  assign N1130 = N3760;
  assign N3765 = (N1131)? 1'b0 : 
                 (N1132)? N3764 : 1'b0;
  assign N1131 = N3763;
  assign N1132 = N3762;
  assign sent_n[377] = (N1133)? 1'b1 : 
                       (N3767)? sent_r[377] : 1'b0;
  assign N1133 = N3766;
  assign N3771 = (N1134)? 1'b0 : 
                 (N1135)? N3770 : 1'b0;
  assign N1134 = N3769;
  assign N1135 = N3768;
  assign sent_n[378] = (N1136)? 1'b1 : 
                       (N3773)? sent_r[378] : 1'b0;
  assign N1136 = N3772;
  assign N3777 = (N1137)? 1'b0 : 
                 (N1138)? N3776 : 1'b0;
  assign N1137 = N3775;
  assign N1138 = N3774;
  assign sent_n[379] = (N1139)? 1'b1 : 
                       (N3779)? sent_r[379] : 1'b0;
  assign N1139 = N3778;
  assign N3783 = (N1140)? 1'b0 : 
                 (N1141)? N3782 : 1'b0;
  assign N1140 = N3781;
  assign N1141 = N3780;
  assign sent_n[380] = (N1142)? 1'b1 : 
                       (N3785)? sent_r[380] : 1'b0;
  assign N1142 = N3784;
  assign N3789 = (N1143)? 1'b0 : 
                 (N1144)? N3788 : 1'b0;
  assign N1143 = N3787;
  assign N1144 = N3786;
  assign sent_n[381] = (N1145)? 1'b1 : 
                       (N3791)? sent_r[381] : 1'b0;
  assign N1145 = N3790;
  assign N3795 = (N1146)? 1'b0 : 
                 (N1147)? N3794 : 1'b0;
  assign N1146 = N3793;
  assign N1147 = N3792;
  assign sent_n[382] = (N1148)? 1'b1 : 
                       (N3797)? sent_r[382] : 1'b0;
  assign N1148 = N3796;
  assign N3801 = (N1149)? 1'b0 : 
                 (N1150)? N3800 : 1'b0;
  assign N1149 = N3799;
  assign N1150 = N3798;
  assign sent_n[383] = (N1151)? 1'b1 : 
                       (N3803)? sent_r[383] : 1'b0;
  assign N1151 = N3802;
  assign N3807 = (N1152)? 1'b0 : 
                 (N1153)? N3806 : 1'b0;
  assign N1152 = N3805;
  assign N1153 = N3804;
  assign sent_n[384] = (N1154)? 1'b1 : 
                       (N3809)? sent_r[384] : 1'b0;
  assign N1154 = N3808;
  assign N3813 = (N1155)? 1'b0 : 
                 (N1156)? N3812 : 1'b0;
  assign N1155 = N3811;
  assign N1156 = N3810;
  assign sent_n[385] = (N1157)? 1'b1 : 
                       (N3815)? sent_r[385] : 1'b0;
  assign N1157 = N3814;
  assign N3819 = (N1158)? 1'b0 : 
                 (N1159)? N3818 : 1'b0;
  assign N1158 = N3817;
  assign N1159 = N3816;
  assign sent_n[386] = (N1160)? 1'b1 : 
                       (N3821)? sent_r[386] : 1'b0;
  assign N1160 = N3820;
  assign N3825 = (N1161)? 1'b0 : 
                 (N1162)? N3824 : 1'b0;
  assign N1161 = N3823;
  assign N1162 = N3822;
  assign sent_n[387] = (N1163)? 1'b1 : 
                       (N3827)? sent_r[387] : 1'b0;
  assign N1163 = N3826;
  assign N3831 = (N1164)? 1'b0 : 
                 (N1165)? N3830 : 1'b0;
  assign N1164 = N3829;
  assign N1165 = N3828;
  assign sent_n[388] = (N1166)? 1'b1 : 
                       (N3833)? sent_r[388] : 1'b0;
  assign N1166 = N3832;
  assign N3837 = (N1167)? 1'b0 : 
                 (N1168)? N3836 : 1'b0;
  assign N1167 = N3835;
  assign N1168 = N3834;
  assign sent_n[389] = (N1169)? 1'b1 : 
                       (N3839)? sent_r[389] : 1'b0;
  assign N1169 = N3838;
  assign N3843 = (N1170)? 1'b0 : 
                 (N1171)? N3842 : 1'b0;
  assign N1170 = N3841;
  assign N1171 = N3840;
  assign sent_n[390] = (N1172)? 1'b1 : 
                       (N3845)? sent_r[390] : 1'b0;
  assign N1172 = N3844;
  assign N3849 = (N1173)? 1'b0 : 
                 (N1174)? N3848 : 1'b0;
  assign N1173 = N3847;
  assign N1174 = N3846;
  assign sent_n[391] = (N1175)? 1'b1 : 
                       (N3851)? sent_r[391] : 1'b0;
  assign N1175 = N3850;
  assign N3855 = (N1176)? 1'b0 : 
                 (N1177)? N3854 : 1'b0;
  assign N1176 = N3853;
  assign N1177 = N3852;
  assign sent_n[392] = (N1178)? 1'b1 : 
                       (N3857)? sent_r[392] : 1'b0;
  assign N1178 = N3856;
  assign N3861 = (N1179)? 1'b0 : 
                 (N1180)? N3860 : 1'b0;
  assign N1179 = N3859;
  assign N1180 = N3858;
  assign sent_n[393] = (N1181)? 1'b1 : 
                       (N3863)? sent_r[393] : 1'b0;
  assign N1181 = N3862;
  assign N3867 = (N1182)? 1'b0 : 
                 (N1183)? N3866 : 1'b0;
  assign N1182 = N3865;
  assign N1183 = N3864;
  assign sent_n[394] = (N1184)? 1'b1 : 
                       (N3869)? sent_r[394] : 1'b0;
  assign N1184 = N3868;
  assign N3873 = (N1185)? 1'b0 : 
                 (N1186)? N3872 : 1'b0;
  assign N1185 = N3871;
  assign N1186 = N3870;
  assign sent_n[395] = (N1187)? 1'b1 : 
                       (N3875)? sent_r[395] : 1'b0;
  assign N1187 = N3874;
  assign N3879 = (N1188)? 1'b0 : 
                 (N1189)? N3878 : 1'b0;
  assign N1188 = N3877;
  assign N1189 = N3876;
  assign sent_n[396] = (N1190)? 1'b1 : 
                       (N3881)? sent_r[396] : 1'b0;
  assign N1190 = N3880;
  assign N3885 = (N1191)? 1'b0 : 
                 (N1192)? N3884 : 1'b0;
  assign N1191 = N3883;
  assign N1192 = N3882;
  assign sent_n[397] = (N1193)? 1'b1 : 
                       (N3887)? sent_r[397] : 1'b0;
  assign N1193 = N3886;
  assign N3891 = (N1194)? 1'b0 : 
                 (N1195)? N3890 : 1'b0;
  assign N1194 = N3889;
  assign N1195 = N3888;
  assign sent_n[398] = (N1196)? 1'b1 : 
                       (N3893)? sent_r[398] : 1'b0;
  assign N1196 = N3892;
  assign N3897 = (N1197)? 1'b0 : 
                 (N1198)? N3896 : 1'b0;
  assign N1197 = N3895;
  assign N1198 = N3894;
  assign sent_n[399] = (N1199)? 1'b1 : 
                       (N3899)? sent_r[399] : 1'b0;
  assign N1199 = N3898;
  assign N3903 = (N1200)? 1'b0 : 
                 (N1201)? N3902 : 1'b0;
  assign N1200 = N3901;
  assign N1201 = N3900;
  assign sent_n[400] = (N1202)? 1'b1 : 
                       (N3905)? sent_r[400] : 1'b0;
  assign N1202 = N3904;
  assign N3909 = (N1203)? 1'b0 : 
                 (N1204)? N3908 : 1'b0;
  assign N1203 = N3907;
  assign N1204 = N3906;
  assign sent_n[401] = (N1205)? 1'b1 : 
                       (N3911)? sent_r[401] : 1'b0;
  assign N1205 = N3910;
  assign N3915 = (N1206)? 1'b0 : 
                 (N1207)? N3914 : 1'b0;
  assign N1206 = N3913;
  assign N1207 = N3912;
  assign sent_n[402] = (N1208)? 1'b1 : 
                       (N3917)? sent_r[402] : 1'b0;
  assign N1208 = N3916;
  assign N3921 = (N1209)? 1'b0 : 
                 (N1210)? N3920 : 1'b0;
  assign N1209 = N3919;
  assign N1210 = N3918;
  assign sent_n[403] = (N1211)? 1'b1 : 
                       (N3923)? sent_r[403] : 1'b0;
  assign N1211 = N3922;
  assign N3927 = (N1212)? 1'b0 : 
                 (N1213)? N3926 : 1'b0;
  assign N1212 = N3925;
  assign N1213 = N3924;
  assign sent_n[404] = (N1214)? 1'b1 : 
                       (N3929)? sent_r[404] : 1'b0;
  assign N1214 = N3928;
  assign N3933 = (N1215)? 1'b0 : 
                 (N1216)? N3932 : 1'b0;
  assign N1215 = N3931;
  assign N1216 = N3930;
  assign sent_n[405] = (N1217)? 1'b1 : 
                       (N3935)? sent_r[405] : 1'b0;
  assign N1217 = N3934;
  assign N3939 = (N1218)? 1'b0 : 
                 (N1219)? N3938 : 1'b0;
  assign N1218 = N3937;
  assign N1219 = N3936;
  assign sent_n[406] = (N1220)? 1'b1 : 
                       (N3941)? sent_r[406] : 1'b0;
  assign N1220 = N3940;
  assign N3945 = (N1221)? 1'b0 : 
                 (N1222)? N3944 : 1'b0;
  assign N1221 = N3943;
  assign N1222 = N3942;
  assign sent_n[407] = (N1223)? 1'b1 : 
                       (N3947)? sent_r[407] : 1'b0;
  assign N1223 = N3946;
  assign N3951 = (N1224)? 1'b0 : 
                 (N1225)? N3950 : 1'b0;
  assign N1224 = N3949;
  assign N1225 = N3948;
  assign sent_n[408] = (N1226)? 1'b1 : 
                       (N3953)? sent_r[408] : 1'b0;
  assign N1226 = N3952;
  assign N3957 = (N1227)? 1'b0 : 
                 (N1228)? N3956 : 1'b0;
  assign N1227 = N3955;
  assign N1228 = N3954;
  assign sent_n[409] = (N1229)? 1'b1 : 
                       (N3959)? sent_r[409] : 1'b0;
  assign N1229 = N3958;
  assign N3963 = (N1230)? 1'b0 : 
                 (N1231)? N3962 : 1'b0;
  assign N1230 = N3961;
  assign N1231 = N3960;
  assign sent_n[410] = (N1232)? 1'b1 : 
                       (N3965)? sent_r[410] : 1'b0;
  assign N1232 = N3964;
  assign N3969 = (N1233)? 1'b0 : 
                 (N1234)? N3968 : 1'b0;
  assign N1233 = N3967;
  assign N1234 = N3966;
  assign sent_n[411] = (N1235)? 1'b1 : 
                       (N3971)? sent_r[411] : 1'b0;
  assign N1235 = N3970;
  assign N3975 = (N1236)? 1'b0 : 
                 (N1237)? N3974 : 1'b0;
  assign N1236 = N3973;
  assign N1237 = N3972;
  assign sent_n[412] = (N1238)? 1'b1 : 
                       (N3977)? sent_r[412] : 1'b0;
  assign N1238 = N3976;
  assign N3981 = (N1239)? 1'b0 : 
                 (N1240)? N3980 : 1'b0;
  assign N1239 = N3979;
  assign N1240 = N3978;
  assign sent_n[413] = (N1241)? 1'b1 : 
                       (N3983)? sent_r[413] : 1'b0;
  assign N1241 = N3982;
  assign N3987 = (N1242)? 1'b0 : 
                 (N1243)? N3986 : 1'b0;
  assign N1242 = N3985;
  assign N1243 = N3984;
  assign sent_n[414] = (N1244)? 1'b1 : 
                       (N3989)? sent_r[414] : 1'b0;
  assign N1244 = N3988;
  assign N3993 = (N1245)? 1'b0 : 
                 (N1246)? N3992 : 1'b0;
  assign N1245 = N3991;
  assign N1246 = N3990;
  assign sent_n[415] = (N1247)? 1'b1 : 
                       (N3995)? sent_r[415] : 1'b0;
  assign N1247 = N3994;
  assign N3999 = (N1248)? 1'b0 : 
                 (N1249)? N3998 : 1'b0;
  assign N1248 = N3997;
  assign N1249 = N3996;
  assign sent_n[416] = (N1250)? 1'b1 : 
                       (N4001)? sent_r[416] : 1'b0;
  assign N1250 = N4000;
  assign N4005 = (N1251)? 1'b0 : 
                 (N1252)? N4004 : 1'b0;
  assign N1251 = N4003;
  assign N1252 = N4002;
  assign sent_n[417] = (N1253)? 1'b1 : 
                       (N4007)? sent_r[417] : 1'b0;
  assign N1253 = N4006;
  assign N4011 = (N1254)? 1'b0 : 
                 (N1255)? N4010 : 1'b0;
  assign N1254 = N4009;
  assign N1255 = N4008;
  assign sent_n[418] = (N1256)? 1'b1 : 
                       (N4013)? sent_r[418] : 1'b0;
  assign N1256 = N4012;
  assign N4017 = (N1257)? 1'b0 : 
                 (N1258)? N4016 : 1'b0;
  assign N1257 = N4015;
  assign N1258 = N4014;
  assign sent_n[419] = (N1259)? 1'b1 : 
                       (N4019)? sent_r[419] : 1'b0;
  assign N1259 = N4018;
  assign N4023 = (N1260)? 1'b0 : 
                 (N1261)? N4022 : 1'b0;
  assign N1260 = N4021;
  assign N1261 = N4020;
  assign sent_n[420] = (N1262)? 1'b1 : 
                       (N4025)? sent_r[420] : 1'b0;
  assign N1262 = N4024;
  assign N4029 = (N1263)? 1'b0 : 
                 (N1264)? N4028 : 1'b0;
  assign N1263 = N4027;
  assign N1264 = N4026;
  assign sent_n[421] = (N1265)? 1'b1 : 
                       (N4031)? sent_r[421] : 1'b0;
  assign N1265 = N4030;
  assign N4035 = (N1266)? 1'b0 : 
                 (N1267)? N4034 : 1'b0;
  assign N1266 = N4033;
  assign N1267 = N4032;
  assign sent_n[422] = (N1268)? 1'b1 : 
                       (N4037)? sent_r[422] : 1'b0;
  assign N1268 = N4036;
  assign N4041 = (N1269)? 1'b0 : 
                 (N1270)? N4040 : 1'b0;
  assign N1269 = N4039;
  assign N1270 = N4038;
  assign sent_n[423] = (N1271)? 1'b1 : 
                       (N4043)? sent_r[423] : 1'b0;
  assign N1271 = N4042;
  assign N4047 = (N1272)? 1'b0 : 
                 (N1273)? N4046 : 1'b0;
  assign N1272 = N4045;
  assign N1273 = N4044;
  assign sent_n[424] = (N1274)? 1'b1 : 
                       (N4049)? sent_r[424] : 1'b0;
  assign N1274 = N4048;
  assign N4053 = (N1275)? 1'b0 : 
                 (N1276)? N4052 : 1'b0;
  assign N1275 = N4051;
  assign N1276 = N4050;
  assign sent_n[425] = (N1277)? 1'b1 : 
                       (N4055)? sent_r[425] : 1'b0;
  assign N1277 = N4054;
  assign N4059 = (N1278)? 1'b0 : 
                 (N1279)? N4058 : 1'b0;
  assign N1278 = N4057;
  assign N1279 = N4056;
  assign sent_n[426] = (N1280)? 1'b1 : 
                       (N4061)? sent_r[426] : 1'b0;
  assign N1280 = N4060;
  assign N4065 = (N1281)? 1'b0 : 
                 (N1282)? N4064 : 1'b0;
  assign N1281 = N4063;
  assign N1282 = N4062;
  assign sent_n[427] = (N1283)? 1'b1 : 
                       (N4067)? sent_r[427] : 1'b0;
  assign N1283 = N4066;
  assign N4071 = (N1284)? 1'b0 : 
                 (N1285)? N4070 : 1'b0;
  assign N1284 = N4069;
  assign N1285 = N4068;
  assign sent_n[428] = (N1286)? 1'b1 : 
                       (N4073)? sent_r[428] : 1'b0;
  assign N1286 = N4072;
  assign N4077 = (N1287)? 1'b0 : 
                 (N1288)? N4076 : 1'b0;
  assign N1287 = N4075;
  assign N1288 = N4074;
  assign sent_n[429] = (N1289)? 1'b1 : 
                       (N4079)? sent_r[429] : 1'b0;
  assign N1289 = N4078;
  assign N4083 = (N1290)? 1'b0 : 
                 (N1291)? N4082 : 1'b0;
  assign N1290 = N4081;
  assign N1291 = N4080;
  assign sent_n[430] = (N1292)? 1'b1 : 
                       (N4085)? sent_r[430] : 1'b0;
  assign N1292 = N4084;
  assign N4089 = (N1293)? 1'b0 : 
                 (N1294)? N4088 : 1'b0;
  assign N1293 = N4087;
  assign N1294 = N4086;
  assign sent_n[431] = (N1295)? 1'b1 : 
                       (N4091)? sent_r[431] : 1'b0;
  assign N1295 = N4090;
  assign N4095 = (N1296)? 1'b0 : 
                 (N1297)? N4094 : 1'b0;
  assign N1296 = N4093;
  assign N1297 = N4092;
  assign sent_n[432] = (N1298)? 1'b1 : 
                       (N4097)? sent_r[432] : 1'b0;
  assign N1298 = N4096;
  assign N4101 = (N1299)? 1'b0 : 
                 (N1300)? N4100 : 1'b0;
  assign N1299 = N4099;
  assign N1300 = N4098;
  assign sent_n[433] = (N1301)? 1'b1 : 
                       (N4103)? sent_r[433] : 1'b0;
  assign N1301 = N4102;
  assign N4107 = (N1302)? 1'b0 : 
                 (N1303)? N4106 : 1'b0;
  assign N1302 = N4105;
  assign N1303 = N4104;
  assign sent_n[434] = (N1304)? 1'b1 : 
                       (N4109)? sent_r[434] : 1'b0;
  assign N1304 = N4108;
  assign N4113 = (N1305)? 1'b0 : 
                 (N1306)? N4112 : 1'b0;
  assign N1305 = N4111;
  assign N1306 = N4110;
  assign sent_n[435] = (N1307)? 1'b1 : 
                       (N4115)? sent_r[435] : 1'b0;
  assign N1307 = N4114;
  assign N4119 = (N1308)? 1'b0 : 
                 (N1309)? N4118 : 1'b0;
  assign N1308 = N4117;
  assign N1309 = N4116;
  assign sent_n[436] = (N1310)? 1'b1 : 
                       (N4121)? sent_r[436] : 1'b0;
  assign N1310 = N4120;
  assign N4125 = (N1311)? 1'b0 : 
                 (N1312)? N4124 : 1'b0;
  assign N1311 = N4123;
  assign N1312 = N4122;
  assign sent_n[437] = (N1313)? 1'b1 : 
                       (N4127)? sent_r[437] : 1'b0;
  assign N1313 = N4126;
  assign N4131 = (N1314)? 1'b0 : 
                 (N1315)? N4130 : 1'b0;
  assign N1314 = N4129;
  assign N1315 = N4128;
  assign sent_n[438] = (N1316)? 1'b1 : 
                       (N4133)? sent_r[438] : 1'b0;
  assign N1316 = N4132;
  assign N4137 = (N1317)? 1'b0 : 
                 (N1318)? N4136 : 1'b0;
  assign N1317 = N4135;
  assign N1318 = N4134;
  assign sent_n[439] = (N1319)? 1'b1 : 
                       (N4139)? sent_r[439] : 1'b0;
  assign N1319 = N4138;
  assign N4143 = (N1320)? 1'b0 : 
                 (N1321)? N4142 : 1'b0;
  assign N1320 = N4141;
  assign N1321 = N4140;
  assign sent_n[440] = (N1322)? 1'b1 : 
                       (N4145)? sent_r[440] : 1'b0;
  assign N1322 = N4144;
  assign N4149 = (N1323)? 1'b0 : 
                 (N1324)? N4148 : 1'b0;
  assign N1323 = N4147;
  assign N1324 = N4146;
  assign sent_n[441] = (N1325)? 1'b1 : 
                       (N4151)? sent_r[441] : 1'b0;
  assign N1325 = N4150;
  assign N4155 = (N1326)? 1'b0 : 
                 (N1327)? N4154 : 1'b0;
  assign N1326 = N4153;
  assign N1327 = N4152;
  assign sent_n[442] = (N1328)? 1'b1 : 
                       (N4157)? sent_r[442] : 1'b0;
  assign N1328 = N4156;
  assign N4161 = (N1329)? 1'b0 : 
                 (N1330)? N4160 : 1'b0;
  assign N1329 = N4159;
  assign N1330 = N4158;
  assign sent_n[443] = (N1331)? 1'b1 : 
                       (N4163)? sent_r[443] : 1'b0;
  assign N1331 = N4162;
  assign N4167 = (N1332)? 1'b0 : 
                 (N1333)? N4166 : 1'b0;
  assign N1332 = N4165;
  assign N1333 = N4164;
  assign sent_n[444] = (N1334)? 1'b1 : 
                       (N4169)? sent_r[444] : 1'b0;
  assign N1334 = N4168;
  assign N4173 = (N1335)? 1'b0 : 
                 (N1336)? N4172 : 1'b0;
  assign N1335 = N4171;
  assign N1336 = N4170;
  assign sent_n[445] = (N1337)? 1'b1 : 
                       (N4175)? sent_r[445] : 1'b0;
  assign N1337 = N4174;
  assign N4179 = (N1338)? 1'b0 : 
                 (N1339)? N4178 : 1'b0;
  assign N1338 = N4177;
  assign N1339 = N4176;
  assign sent_n[446] = (N1340)? 1'b1 : 
                       (N4181)? sent_r[446] : 1'b0;
  assign N1340 = N4180;
  assign N4185 = (N1341)? 1'b0 : 
                 (N1342)? N4184 : 1'b0;
  assign N1341 = N4183;
  assign N1342 = N4182;
  assign sent_n[447] = (N1343)? 1'b1 : 
                       (N4187)? sent_r[447] : 1'b0;
  assign N1343 = N4186;
  assign N4191 = (N1344)? 1'b0 : 
                 (N1345)? N4190 : 1'b0;
  assign N1344 = N4189;
  assign N1345 = N4188;
  assign sent_n[448] = (N1346)? 1'b1 : 
                       (N4193)? sent_r[448] : 1'b0;
  assign N1346 = N4192;
  assign N4197 = (N1347)? 1'b0 : 
                 (N1348)? N4196 : 1'b0;
  assign N1347 = N4195;
  assign N1348 = N4194;
  assign sent_n[449] = (N1349)? 1'b1 : 
                       (N4199)? sent_r[449] : 1'b0;
  assign N1349 = N4198;
  assign N4203 = (N1350)? 1'b0 : 
                 (N1351)? N4202 : 1'b0;
  assign N1350 = N4201;
  assign N1351 = N4200;
  assign sent_n[450] = (N1352)? 1'b1 : 
                       (N4205)? sent_r[450] : 1'b0;
  assign N1352 = N4204;
  assign N4209 = (N1353)? 1'b0 : 
                 (N1354)? N4208 : 1'b0;
  assign N1353 = N4207;
  assign N1354 = N4206;
  assign sent_n[451] = (N1355)? 1'b1 : 
                       (N4211)? sent_r[451] : 1'b0;
  assign N1355 = N4210;
  assign N4215 = (N1356)? 1'b0 : 
                 (N1357)? N4214 : 1'b0;
  assign N1356 = N4213;
  assign N1357 = N4212;
  assign sent_n[452] = (N1358)? 1'b1 : 
                       (N4217)? sent_r[452] : 1'b0;
  assign N1358 = N4216;
  assign N4221 = (N1359)? 1'b0 : 
                 (N1360)? N4220 : 1'b0;
  assign N1359 = N4219;
  assign N1360 = N4218;
  assign sent_n[453] = (N1361)? 1'b1 : 
                       (N4223)? sent_r[453] : 1'b0;
  assign N1361 = N4222;
  assign N4227 = (N1362)? 1'b0 : 
                 (N1363)? N4226 : 1'b0;
  assign N1362 = N4225;
  assign N1363 = N4224;
  assign sent_n[454] = (N1364)? 1'b1 : 
                       (N4229)? sent_r[454] : 1'b0;
  assign N1364 = N4228;
  assign N4233 = (N1365)? 1'b0 : 
                 (N1366)? N4232 : 1'b0;
  assign N1365 = N4231;
  assign N1366 = N4230;
  assign sent_n[455] = (N1367)? 1'b1 : 
                       (N4235)? sent_r[455] : 1'b0;
  assign N1367 = N4234;
  assign N4239 = (N1368)? 1'b0 : 
                 (N1369)? N4238 : 1'b0;
  assign N1368 = N4237;
  assign N1369 = N4236;
  assign sent_n[456] = (N1370)? 1'b1 : 
                       (N4241)? sent_r[456] : 1'b0;
  assign N1370 = N4240;
  assign N4245 = (N1371)? 1'b0 : 
                 (N1372)? N4244 : 1'b0;
  assign N1371 = N4243;
  assign N1372 = N4242;
  assign sent_n[457] = (N1373)? 1'b1 : 
                       (N4247)? sent_r[457] : 1'b0;
  assign N1373 = N4246;
  assign N4251 = (N1374)? 1'b0 : 
                 (N1375)? N4250 : 1'b0;
  assign N1374 = N4249;
  assign N1375 = N4248;
  assign sent_n[458] = (N1376)? 1'b1 : 
                       (N4253)? sent_r[458] : 1'b0;
  assign N1376 = N4252;
  assign N4257 = (N1377)? 1'b0 : 
                 (N1378)? N4256 : 1'b0;
  assign N1377 = N4255;
  assign N1378 = N4254;
  assign sent_n[459] = (N1379)? 1'b1 : 
                       (N4259)? sent_r[459] : 1'b0;
  assign N1379 = N4258;
  assign N4263 = (N1380)? 1'b0 : 
                 (N1381)? N4262 : 1'b0;
  assign N1380 = N4261;
  assign N1381 = N4260;
  assign sent_n[460] = (N1382)? 1'b1 : 
                       (N4265)? sent_r[460] : 1'b0;
  assign N1382 = N4264;
  assign N4269 = (N1383)? 1'b0 : 
                 (N1384)? N4268 : 1'b0;
  assign N1383 = N4267;
  assign N1384 = N4266;
  assign sent_n[461] = (N1385)? 1'b1 : 
                       (N4271)? sent_r[461] : 1'b0;
  assign N1385 = N4270;
  assign N4275 = (N1386)? 1'b0 : 
                 (N1387)? N4274 : 1'b0;
  assign N1386 = N4273;
  assign N1387 = N4272;
  assign sent_n[462] = (N1388)? 1'b1 : 
                       (N4277)? sent_r[462] : 1'b0;
  assign N1388 = N4276;
  assign N4281 = (N1389)? 1'b0 : 
                 (N1390)? N4280 : 1'b0;
  assign N1389 = N4279;
  assign N1390 = N4278;
  assign sent_n[463] = (N1391)? 1'b1 : 
                       (N4283)? sent_r[463] : 1'b0;
  assign N1391 = N4282;
  assign N4287 = (N1392)? 1'b0 : 
                 (N1393)? N4286 : 1'b0;
  assign N1392 = N4285;
  assign N1393 = N4284;
  assign sent_n[464] = (N1394)? 1'b1 : 
                       (N4289)? sent_r[464] : 1'b0;
  assign N1394 = N4288;
  assign N4293 = (N1395)? 1'b0 : 
                 (N1396)? N4292 : 1'b0;
  assign N1395 = N4291;
  assign N1396 = N4290;
  assign sent_n[465] = (N1397)? 1'b1 : 
                       (N4295)? sent_r[465] : 1'b0;
  assign N1397 = N4294;
  assign N4299 = (N1398)? 1'b0 : 
                 (N1399)? N4298 : 1'b0;
  assign N1398 = N4297;
  assign N1399 = N4296;
  assign sent_n[466] = (N1400)? 1'b1 : 
                       (N4301)? sent_r[466] : 1'b0;
  assign N1400 = N4300;
  assign N4305 = (N1401)? 1'b0 : 
                 (N1402)? N4304 : 1'b0;
  assign N1401 = N4303;
  assign N1402 = N4302;
  assign sent_n[467] = (N1403)? 1'b1 : 
                       (N4307)? sent_r[467] : 1'b0;
  assign N1403 = N4306;
  assign N4311 = (N1404)? 1'b0 : 
                 (N1405)? N4310 : 1'b0;
  assign N1404 = N4309;
  assign N1405 = N4308;
  assign sent_n[468] = (N1406)? 1'b1 : 
                       (N4313)? sent_r[468] : 1'b0;
  assign N1406 = N4312;
  assign N4317 = (N1407)? 1'b0 : 
                 (N1408)? N4316 : 1'b0;
  assign N1407 = N4315;
  assign N1408 = N4314;
  assign sent_n[469] = (N1409)? 1'b1 : 
                       (N4319)? sent_r[469] : 1'b0;
  assign N1409 = N4318;
  assign N4323 = (N1410)? 1'b0 : 
                 (N1411)? N4322 : 1'b0;
  assign N1410 = N4321;
  assign N1411 = N4320;
  assign sent_n[470] = (N1412)? 1'b1 : 
                       (N4325)? sent_r[470] : 1'b0;
  assign N1412 = N4324;
  assign N4329 = (N1413)? 1'b0 : 
                 (N1414)? N4328 : 1'b0;
  assign N1413 = N4327;
  assign N1414 = N4326;
  assign sent_n[471] = (N1415)? 1'b1 : 
                       (N4331)? sent_r[471] : 1'b0;
  assign N1415 = N4330;
  assign N4335 = (N1416)? 1'b0 : 
                 (N1417)? N4334 : 1'b0;
  assign N1416 = N4333;
  assign N1417 = N4332;
  assign sent_n[472] = (N1418)? 1'b1 : 
                       (N4337)? sent_r[472] : 1'b0;
  assign N1418 = N4336;
  assign N4341 = (N1419)? 1'b0 : 
                 (N1420)? N4340 : 1'b0;
  assign N1419 = N4339;
  assign N1420 = N4338;
  assign sent_n[473] = (N1421)? 1'b1 : 
                       (N4343)? sent_r[473] : 1'b0;
  assign N1421 = N4342;
  assign N4347 = (N1422)? 1'b0 : 
                 (N1423)? N4346 : 1'b0;
  assign N1422 = N4345;
  assign N1423 = N4344;
  assign sent_n[474] = (N1424)? 1'b1 : 
                       (N4349)? sent_r[474] : 1'b0;
  assign N1424 = N4348;
  assign N4353 = (N1425)? 1'b0 : 
                 (N1426)? N4352 : 1'b0;
  assign N1425 = N4351;
  assign N1426 = N4350;
  assign sent_n[475] = (N1427)? 1'b1 : 
                       (N4355)? sent_r[475] : 1'b0;
  assign N1427 = N4354;
  assign N4359 = (N1428)? 1'b0 : 
                 (N1429)? N4358 : 1'b0;
  assign N1428 = N4357;
  assign N1429 = N4356;
  assign sent_n[476] = (N1430)? 1'b1 : 
                       (N4361)? sent_r[476] : 1'b0;
  assign N1430 = N4360;
  assign N4365 = (N1431)? 1'b0 : 
                 (N1432)? N4364 : 1'b0;
  assign N1431 = N4363;
  assign N1432 = N4362;
  assign sent_n[477] = (N1433)? 1'b1 : 
                       (N4367)? sent_r[477] : 1'b0;
  assign N1433 = N4366;
  assign N4371 = (N1434)? 1'b0 : 
                 (N1435)? N4370 : 1'b0;
  assign N1434 = N4369;
  assign N1435 = N4368;
  assign sent_n[478] = (N1436)? 1'b1 : 
                       (N4373)? sent_r[478] : 1'b0;
  assign N1436 = N4372;
  assign N4377 = (N1437)? 1'b0 : 
                 (N1438)? N4376 : 1'b0;
  assign N1437 = N4375;
  assign N1438 = N4374;
  assign sent_n[479] = (N1439)? 1'b1 : 
                       (N4379)? sent_r[479] : 1'b0;
  assign N1439 = N4378;
  assign N4383 = (N1440)? 1'b0 : 
                 (N1441)? N4382 : 1'b0;
  assign N1440 = N4381;
  assign N1441 = N4380;
  assign sent_n[480] = (N1442)? 1'b1 : 
                       (N4385)? sent_r[480] : 1'b0;
  assign N1442 = N4384;
  assign N4389 = (N1443)? 1'b0 : 
                 (N1444)? N4388 : 1'b0;
  assign N1443 = N4387;
  assign N1444 = N4386;
  assign sent_n[481] = (N1445)? 1'b1 : 
                       (N4391)? sent_r[481] : 1'b0;
  assign N1445 = N4390;
  assign N4395 = (N1446)? 1'b0 : 
                 (N1447)? N4394 : 1'b0;
  assign N1446 = N4393;
  assign N1447 = N4392;
  assign sent_n[482] = (N1448)? 1'b1 : 
                       (N4397)? sent_r[482] : 1'b0;
  assign N1448 = N4396;
  assign N4401 = (N1449)? 1'b0 : 
                 (N1450)? N4400 : 1'b0;
  assign N1449 = N4399;
  assign N1450 = N4398;
  assign sent_n[483] = (N1451)? 1'b1 : 
                       (N4403)? sent_r[483] : 1'b0;
  assign N1451 = N4402;
  assign N4407 = (N1452)? 1'b0 : 
                 (N1453)? N4406 : 1'b0;
  assign N1452 = N4405;
  assign N1453 = N4404;
  assign sent_n[484] = (N1454)? 1'b1 : 
                       (N4409)? sent_r[484] : 1'b0;
  assign N1454 = N4408;
  assign N4413 = (N1455)? 1'b0 : 
                 (N1456)? N4412 : 1'b0;
  assign N1455 = N4411;
  assign N1456 = N4410;
  assign sent_n[485] = (N1457)? 1'b1 : 
                       (N4415)? sent_r[485] : 1'b0;
  assign N1457 = N4414;
  assign N4419 = (N1458)? 1'b0 : 
                 (N1459)? N4418 : 1'b0;
  assign N1458 = N4417;
  assign N1459 = N4416;
  assign sent_n[486] = (N1460)? 1'b1 : 
                       (N4421)? sent_r[486] : 1'b0;
  assign N1460 = N4420;
  assign N4425 = (N1461)? 1'b0 : 
                 (N1462)? N4424 : 1'b0;
  assign N1461 = N4423;
  assign N1462 = N4422;
  assign sent_n[487] = (N1463)? 1'b1 : 
                       (N4427)? sent_r[487] : 1'b0;
  assign N1463 = N4426;
  assign N4431 = (N1464)? 1'b0 : 
                 (N1465)? N4430 : 1'b0;
  assign N1464 = N4429;
  assign N1465 = N4428;
  assign sent_n[488] = (N1466)? 1'b1 : 
                       (N4433)? sent_r[488] : 1'b0;
  assign N1466 = N4432;
  assign N4437 = (N1467)? 1'b0 : 
                 (N1468)? N4436 : 1'b0;
  assign N1467 = N4435;
  assign N1468 = N4434;
  assign sent_n[489] = (N1469)? 1'b1 : 
                       (N4439)? sent_r[489] : 1'b0;
  assign N1469 = N4438;
  assign N4443 = (N1470)? 1'b0 : 
                 (N1471)? N4442 : 1'b0;
  assign N1470 = N4441;
  assign N1471 = N4440;
  assign sent_n[490] = (N1472)? 1'b1 : 
                       (N4445)? sent_r[490] : 1'b0;
  assign N1472 = N4444;
  assign N4449 = (N1473)? 1'b0 : 
                 (N1474)? N4448 : 1'b0;
  assign N1473 = N4447;
  assign N1474 = N4446;
  assign sent_n[491] = (N1475)? 1'b1 : 
                       (N4451)? sent_r[491] : 1'b0;
  assign N1475 = N4450;
  assign N4455 = (N1476)? 1'b0 : 
                 (N1477)? N4454 : 1'b0;
  assign N1476 = N4453;
  assign N1477 = N4452;
  assign sent_n[492] = (N1478)? 1'b1 : 
                       (N4457)? sent_r[492] : 1'b0;
  assign N1478 = N4456;
  assign N4461 = (N1479)? 1'b0 : 
                 (N1480)? N4460 : 1'b0;
  assign N1479 = N4459;
  assign N1480 = N4458;
  assign sent_n[493] = (N1481)? 1'b1 : 
                       (N4463)? sent_r[493] : 1'b0;
  assign N1481 = N4462;
  assign N4467 = (N1482)? 1'b0 : 
                 (N1483)? N4466 : 1'b0;
  assign N1482 = N4465;
  assign N1483 = N4464;
  assign sent_n[494] = (N1484)? 1'b1 : 
                       (N4469)? sent_r[494] : 1'b0;
  assign N1484 = N4468;
  assign N4473 = (N1485)? 1'b0 : 
                 (N1486)? N4472 : 1'b0;
  assign N1485 = N4471;
  assign N1486 = N4470;
  assign sent_n[495] = (N1487)? 1'b1 : 
                       (N4475)? sent_r[495] : 1'b0;
  assign N1487 = N4474;
  assign N4479 = (N1488)? 1'b0 : 
                 (N1489)? N4478 : 1'b0;
  assign N1488 = N4477;
  assign N1489 = N4476;
  assign sent_n[496] = (N1490)? 1'b1 : 
                       (N4481)? sent_r[496] : 1'b0;
  assign N1490 = N4480;
  assign N4485 = (N1491)? 1'b0 : 
                 (N1492)? N4484 : 1'b0;
  assign N1491 = N4483;
  assign N1492 = N4482;
  assign sent_n[497] = (N1493)? 1'b1 : 
                       (N4487)? sent_r[497] : 1'b0;
  assign N1493 = N4486;
  assign N4491 = (N1494)? 1'b0 : 
                 (N1495)? N4490 : 1'b0;
  assign N1494 = N4489;
  assign N1495 = N4488;
  assign sent_n[498] = (N1496)? 1'b1 : 
                       (N4493)? sent_r[498] : 1'b0;
  assign N1496 = N4492;
  assign N4497 = (N1497)? 1'b0 : 
                 (N1498)? N4496 : 1'b0;
  assign N1497 = N4495;
  assign N1498 = N4494;
  assign sent_n[499] = (N1499)? 1'b1 : 
                       (N4499)? sent_r[499] : 1'b0;
  assign N1499 = N4498;
  assign v_o[0] = fifo_v & N4500;
  assign N4500 = ~sent_r[0];
  assign N1500 = ~reset_i;
  assign N1501 = reset_i;
  assign N1502 = sent_n[0] & N4501;
  assign N4501 = ~fifo_yumi;
  assign N1504 = v_o[0] & ready_i[0];
  assign N1505 = ~N1504;
  assign v_o[1] = fifo_v & N4502;
  assign N4502 = ~sent_r[1];
  assign N1506 = ~reset_i;
  assign N1507 = reset_i;
  assign N1508 = sent_n[1] & N4503;
  assign N4503 = ~fifo_yumi;
  assign N1510 = v_o[1] & ready_i[1];
  assign N1511 = ~N1510;
  assign v_o[2] = fifo_v & N4504;
  assign N4504 = ~sent_r[2];
  assign N1512 = ~reset_i;
  assign N1513 = reset_i;
  assign N1514 = sent_n[2] & N4505;
  assign N4505 = ~fifo_yumi;
  assign N1516 = v_o[2] & ready_i[2];
  assign N1517 = ~N1516;
  assign v_o[3] = fifo_v & N4506;
  assign N4506 = ~sent_r[3];
  assign N1518 = ~reset_i;
  assign N1519 = reset_i;
  assign N1520 = sent_n[3] & N4507;
  assign N4507 = ~fifo_yumi;
  assign N1522 = v_o[3] & ready_i[3];
  assign N1523 = ~N1522;
  assign v_o[4] = fifo_v & N4508;
  assign N4508 = ~sent_r[4];
  assign N1524 = ~reset_i;
  assign N1525 = reset_i;
  assign N1526 = sent_n[4] & N4509;
  assign N4509 = ~fifo_yumi;
  assign N1528 = v_o[4] & ready_i[4];
  assign N1529 = ~N1528;
  assign v_o[5] = fifo_v & N4510;
  assign N4510 = ~sent_r[5];
  assign N1530 = ~reset_i;
  assign N1531 = reset_i;
  assign N1532 = sent_n[5] & N4511;
  assign N4511 = ~fifo_yumi;
  assign N1534 = v_o[5] & ready_i[5];
  assign N1535 = ~N1534;
  assign v_o[6] = fifo_v & N4512;
  assign N4512 = ~sent_r[6];
  assign N1536 = ~reset_i;
  assign N1537 = reset_i;
  assign N1538 = sent_n[6] & N4513;
  assign N4513 = ~fifo_yumi;
  assign N1540 = v_o[6] & ready_i[6];
  assign N1541 = ~N1540;
  assign v_o[7] = fifo_v & N4514;
  assign N4514 = ~sent_r[7];
  assign N1542 = ~reset_i;
  assign N1543 = reset_i;
  assign N1544 = sent_n[7] & N4515;
  assign N4515 = ~fifo_yumi;
  assign N1546 = v_o[7] & ready_i[7];
  assign N1547 = ~N1546;
  assign v_o[8] = fifo_v & N4516;
  assign N4516 = ~sent_r[8];
  assign N1548 = ~reset_i;
  assign N1549 = reset_i;
  assign N1550 = sent_n[8] & N4517;
  assign N4517 = ~fifo_yumi;
  assign N1552 = v_o[8] & ready_i[8];
  assign N1553 = ~N1552;
  assign v_o[9] = fifo_v & N4518;
  assign N4518 = ~sent_r[9];
  assign N1554 = ~reset_i;
  assign N1555 = reset_i;
  assign N1556 = sent_n[9] & N4519;
  assign N4519 = ~fifo_yumi;
  assign N1558 = v_o[9] & ready_i[9];
  assign N1559 = ~N1558;
  assign v_o[10] = fifo_v & N4520;
  assign N4520 = ~sent_r[10];
  assign N1560 = ~reset_i;
  assign N1561 = reset_i;
  assign N1562 = sent_n[10] & N4521;
  assign N4521 = ~fifo_yumi;
  assign N1564 = v_o[10] & ready_i[10];
  assign N1565 = ~N1564;
  assign v_o[11] = fifo_v & N4522;
  assign N4522 = ~sent_r[11];
  assign N1566 = ~reset_i;
  assign N1567 = reset_i;
  assign N1568 = sent_n[11] & N4523;
  assign N4523 = ~fifo_yumi;
  assign N1570 = v_o[11] & ready_i[11];
  assign N1571 = ~N1570;
  assign v_o[12] = fifo_v & N4524;
  assign N4524 = ~sent_r[12];
  assign N1572 = ~reset_i;
  assign N1573 = reset_i;
  assign N1574 = sent_n[12] & N4525;
  assign N4525 = ~fifo_yumi;
  assign N1576 = v_o[12] & ready_i[12];
  assign N1577 = ~N1576;
  assign v_o[13] = fifo_v & N4526;
  assign N4526 = ~sent_r[13];
  assign N1578 = ~reset_i;
  assign N1579 = reset_i;
  assign N1580 = sent_n[13] & N4527;
  assign N4527 = ~fifo_yumi;
  assign N1582 = v_o[13] & ready_i[13];
  assign N1583 = ~N1582;
  assign v_o[14] = fifo_v & N4528;
  assign N4528 = ~sent_r[14];
  assign N1584 = ~reset_i;
  assign N1585 = reset_i;
  assign N1586 = sent_n[14] & N4529;
  assign N4529 = ~fifo_yumi;
  assign N1588 = v_o[14] & ready_i[14];
  assign N1589 = ~N1588;
  assign v_o[15] = fifo_v & N4530;
  assign N4530 = ~sent_r[15];
  assign N1590 = ~reset_i;
  assign N1591 = reset_i;
  assign N1592 = sent_n[15] & N4531;
  assign N4531 = ~fifo_yumi;
  assign N1594 = v_o[15] & ready_i[15];
  assign N1595 = ~N1594;
  assign v_o[16] = fifo_v & N4532;
  assign N4532 = ~sent_r[16];
  assign N1596 = ~reset_i;
  assign N1597 = reset_i;
  assign N1598 = sent_n[16] & N4533;
  assign N4533 = ~fifo_yumi;
  assign N1600 = v_o[16] & ready_i[16];
  assign N1601 = ~N1600;
  assign v_o[17] = fifo_v & N4534;
  assign N4534 = ~sent_r[17];
  assign N1602 = ~reset_i;
  assign N1603 = reset_i;
  assign N1604 = sent_n[17] & N4535;
  assign N4535 = ~fifo_yumi;
  assign N1606 = v_o[17] & ready_i[17];
  assign N1607 = ~N1606;
  assign v_o[18] = fifo_v & N4536;
  assign N4536 = ~sent_r[18];
  assign N1608 = ~reset_i;
  assign N1609 = reset_i;
  assign N1610 = sent_n[18] & N4537;
  assign N4537 = ~fifo_yumi;
  assign N1612 = v_o[18] & ready_i[18];
  assign N1613 = ~N1612;
  assign v_o[19] = fifo_v & N4538;
  assign N4538 = ~sent_r[19];
  assign N1614 = ~reset_i;
  assign N1615 = reset_i;
  assign N1616 = sent_n[19] & N4539;
  assign N4539 = ~fifo_yumi;
  assign N1618 = v_o[19] & ready_i[19];
  assign N1619 = ~N1618;
  assign v_o[20] = fifo_v & N4540;
  assign N4540 = ~sent_r[20];
  assign N1620 = ~reset_i;
  assign N1621 = reset_i;
  assign N1622 = sent_n[20] & N4541;
  assign N4541 = ~fifo_yumi;
  assign N1624 = v_o[20] & ready_i[20];
  assign N1625 = ~N1624;
  assign v_o[21] = fifo_v & N4542;
  assign N4542 = ~sent_r[21];
  assign N1626 = ~reset_i;
  assign N1627 = reset_i;
  assign N1628 = sent_n[21] & N4543;
  assign N4543 = ~fifo_yumi;
  assign N1630 = v_o[21] & ready_i[21];
  assign N1631 = ~N1630;
  assign v_o[22] = fifo_v & N4544;
  assign N4544 = ~sent_r[22];
  assign N1632 = ~reset_i;
  assign N1633 = reset_i;
  assign N1634 = sent_n[22] & N4545;
  assign N4545 = ~fifo_yumi;
  assign N1636 = v_o[22] & ready_i[22];
  assign N1637 = ~N1636;
  assign v_o[23] = fifo_v & N4546;
  assign N4546 = ~sent_r[23];
  assign N1638 = ~reset_i;
  assign N1639 = reset_i;
  assign N1640 = sent_n[23] & N4547;
  assign N4547 = ~fifo_yumi;
  assign N1642 = v_o[23] & ready_i[23];
  assign N1643 = ~N1642;
  assign v_o[24] = fifo_v & N4548;
  assign N4548 = ~sent_r[24];
  assign N1644 = ~reset_i;
  assign N1645 = reset_i;
  assign N1646 = sent_n[24] & N4549;
  assign N4549 = ~fifo_yumi;
  assign N1648 = v_o[24] & ready_i[24];
  assign N1649 = ~N1648;
  assign v_o[25] = fifo_v & N4550;
  assign N4550 = ~sent_r[25];
  assign N1650 = ~reset_i;
  assign N1651 = reset_i;
  assign N1652 = sent_n[25] & N4551;
  assign N4551 = ~fifo_yumi;
  assign N1654 = v_o[25] & ready_i[25];
  assign N1655 = ~N1654;
  assign v_o[26] = fifo_v & N4552;
  assign N4552 = ~sent_r[26];
  assign N1656 = ~reset_i;
  assign N1657 = reset_i;
  assign N1658 = sent_n[26] & N4553;
  assign N4553 = ~fifo_yumi;
  assign N1660 = v_o[26] & ready_i[26];
  assign N1661 = ~N1660;
  assign v_o[27] = fifo_v & N4554;
  assign N4554 = ~sent_r[27];
  assign N1662 = ~reset_i;
  assign N1663 = reset_i;
  assign N1664 = sent_n[27] & N4555;
  assign N4555 = ~fifo_yumi;
  assign N1666 = v_o[27] & ready_i[27];
  assign N1667 = ~N1666;
  assign v_o[28] = fifo_v & N4556;
  assign N4556 = ~sent_r[28];
  assign N1668 = ~reset_i;
  assign N1669 = reset_i;
  assign N1670 = sent_n[28] & N4557;
  assign N4557 = ~fifo_yumi;
  assign N1672 = v_o[28] & ready_i[28];
  assign N1673 = ~N1672;
  assign v_o[29] = fifo_v & N4558;
  assign N4558 = ~sent_r[29];
  assign N1674 = ~reset_i;
  assign N1675 = reset_i;
  assign N1676 = sent_n[29] & N4559;
  assign N4559 = ~fifo_yumi;
  assign N1678 = v_o[29] & ready_i[29];
  assign N1679 = ~N1678;
  assign v_o[30] = fifo_v & N4560;
  assign N4560 = ~sent_r[30];
  assign N1680 = ~reset_i;
  assign N1681 = reset_i;
  assign N1682 = sent_n[30] & N4561;
  assign N4561 = ~fifo_yumi;
  assign N1684 = v_o[30] & ready_i[30];
  assign N1685 = ~N1684;
  assign v_o[31] = fifo_v & N4562;
  assign N4562 = ~sent_r[31];
  assign N1686 = ~reset_i;
  assign N1687 = reset_i;
  assign N1688 = sent_n[31] & N4563;
  assign N4563 = ~fifo_yumi;
  assign N1690 = v_o[31] & ready_i[31];
  assign N1691 = ~N1690;
  assign v_o[32] = fifo_v & N4564;
  assign N4564 = ~sent_r[32];
  assign N1692 = ~reset_i;
  assign N1693 = reset_i;
  assign N1694 = sent_n[32] & N4565;
  assign N4565 = ~fifo_yumi;
  assign N1696 = v_o[32] & ready_i[32];
  assign N1697 = ~N1696;
  assign v_o[33] = fifo_v & N4566;
  assign N4566 = ~sent_r[33];
  assign N1698 = ~reset_i;
  assign N1699 = reset_i;
  assign N1700 = sent_n[33] & N4567;
  assign N4567 = ~fifo_yumi;
  assign N1702 = v_o[33] & ready_i[33];
  assign N1703 = ~N1702;
  assign v_o[34] = fifo_v & N4568;
  assign N4568 = ~sent_r[34];
  assign N1704 = ~reset_i;
  assign N1705 = reset_i;
  assign N1706 = sent_n[34] & N4569;
  assign N4569 = ~fifo_yumi;
  assign N1708 = v_o[34] & ready_i[34];
  assign N1709 = ~N1708;
  assign v_o[35] = fifo_v & N4570;
  assign N4570 = ~sent_r[35];
  assign N1710 = ~reset_i;
  assign N1711 = reset_i;
  assign N1712 = sent_n[35] & N4571;
  assign N4571 = ~fifo_yumi;
  assign N1714 = v_o[35] & ready_i[35];
  assign N1715 = ~N1714;
  assign v_o[36] = fifo_v & N4572;
  assign N4572 = ~sent_r[36];
  assign N1716 = ~reset_i;
  assign N1717 = reset_i;
  assign N1718 = sent_n[36] & N4573;
  assign N4573 = ~fifo_yumi;
  assign N1720 = v_o[36] & ready_i[36];
  assign N1721 = ~N1720;
  assign v_o[37] = fifo_v & N4574;
  assign N4574 = ~sent_r[37];
  assign N1722 = ~reset_i;
  assign N1723 = reset_i;
  assign N1724 = sent_n[37] & N4575;
  assign N4575 = ~fifo_yumi;
  assign N1726 = v_o[37] & ready_i[37];
  assign N1727 = ~N1726;
  assign v_o[38] = fifo_v & N4576;
  assign N4576 = ~sent_r[38];
  assign N1728 = ~reset_i;
  assign N1729 = reset_i;
  assign N1730 = sent_n[38] & N4577;
  assign N4577 = ~fifo_yumi;
  assign N1732 = v_o[38] & ready_i[38];
  assign N1733 = ~N1732;
  assign v_o[39] = fifo_v & N4578;
  assign N4578 = ~sent_r[39];
  assign N1734 = ~reset_i;
  assign N1735 = reset_i;
  assign N1736 = sent_n[39] & N4579;
  assign N4579 = ~fifo_yumi;
  assign N1738 = v_o[39] & ready_i[39];
  assign N1739 = ~N1738;
  assign v_o[40] = fifo_v & N4580;
  assign N4580 = ~sent_r[40];
  assign N1740 = ~reset_i;
  assign N1741 = reset_i;
  assign N1742 = sent_n[40] & N4581;
  assign N4581 = ~fifo_yumi;
  assign N1744 = v_o[40] & ready_i[40];
  assign N1745 = ~N1744;
  assign v_o[41] = fifo_v & N4582;
  assign N4582 = ~sent_r[41];
  assign N1746 = ~reset_i;
  assign N1747 = reset_i;
  assign N1748 = sent_n[41] & N4583;
  assign N4583 = ~fifo_yumi;
  assign N1750 = v_o[41] & ready_i[41];
  assign N1751 = ~N1750;
  assign v_o[42] = fifo_v & N4584;
  assign N4584 = ~sent_r[42];
  assign N1752 = ~reset_i;
  assign N1753 = reset_i;
  assign N1754 = sent_n[42] & N4585;
  assign N4585 = ~fifo_yumi;
  assign N1756 = v_o[42] & ready_i[42];
  assign N1757 = ~N1756;
  assign v_o[43] = fifo_v & N4586;
  assign N4586 = ~sent_r[43];
  assign N1758 = ~reset_i;
  assign N1759 = reset_i;
  assign N1760 = sent_n[43] & N4587;
  assign N4587 = ~fifo_yumi;
  assign N1762 = v_o[43] & ready_i[43];
  assign N1763 = ~N1762;
  assign v_o[44] = fifo_v & N4588;
  assign N4588 = ~sent_r[44];
  assign N1764 = ~reset_i;
  assign N1765 = reset_i;
  assign N1766 = sent_n[44] & N4589;
  assign N4589 = ~fifo_yumi;
  assign N1768 = v_o[44] & ready_i[44];
  assign N1769 = ~N1768;
  assign v_o[45] = fifo_v & N4590;
  assign N4590 = ~sent_r[45];
  assign N1770 = ~reset_i;
  assign N1771 = reset_i;
  assign N1772 = sent_n[45] & N4591;
  assign N4591 = ~fifo_yumi;
  assign N1774 = v_o[45] & ready_i[45];
  assign N1775 = ~N1774;
  assign v_o[46] = fifo_v & N4592;
  assign N4592 = ~sent_r[46];
  assign N1776 = ~reset_i;
  assign N1777 = reset_i;
  assign N1778 = sent_n[46] & N4593;
  assign N4593 = ~fifo_yumi;
  assign N1780 = v_o[46] & ready_i[46];
  assign N1781 = ~N1780;
  assign v_o[47] = fifo_v & N4594;
  assign N4594 = ~sent_r[47];
  assign N1782 = ~reset_i;
  assign N1783 = reset_i;
  assign N1784 = sent_n[47] & N4595;
  assign N4595 = ~fifo_yumi;
  assign N1786 = v_o[47] & ready_i[47];
  assign N1787 = ~N1786;
  assign v_o[48] = fifo_v & N4596;
  assign N4596 = ~sent_r[48];
  assign N1788 = ~reset_i;
  assign N1789 = reset_i;
  assign N1790 = sent_n[48] & N4597;
  assign N4597 = ~fifo_yumi;
  assign N1792 = v_o[48] & ready_i[48];
  assign N1793 = ~N1792;
  assign v_o[49] = fifo_v & N4598;
  assign N4598 = ~sent_r[49];
  assign N1794 = ~reset_i;
  assign N1795 = reset_i;
  assign N1796 = sent_n[49] & N4599;
  assign N4599 = ~fifo_yumi;
  assign N1798 = v_o[49] & ready_i[49];
  assign N1799 = ~N1798;
  assign v_o[50] = fifo_v & N4600;
  assign N4600 = ~sent_r[50];
  assign N1800 = ~reset_i;
  assign N1801 = reset_i;
  assign N1802 = sent_n[50] & N4601;
  assign N4601 = ~fifo_yumi;
  assign N1804 = v_o[50] & ready_i[50];
  assign N1805 = ~N1804;
  assign v_o[51] = fifo_v & N4602;
  assign N4602 = ~sent_r[51];
  assign N1806 = ~reset_i;
  assign N1807 = reset_i;
  assign N1808 = sent_n[51] & N4603;
  assign N4603 = ~fifo_yumi;
  assign N1810 = v_o[51] & ready_i[51];
  assign N1811 = ~N1810;
  assign v_o[52] = fifo_v & N4604;
  assign N4604 = ~sent_r[52];
  assign N1812 = ~reset_i;
  assign N1813 = reset_i;
  assign N1814 = sent_n[52] & N4605;
  assign N4605 = ~fifo_yumi;
  assign N1816 = v_o[52] & ready_i[52];
  assign N1817 = ~N1816;
  assign v_o[53] = fifo_v & N4606;
  assign N4606 = ~sent_r[53];
  assign N1818 = ~reset_i;
  assign N1819 = reset_i;
  assign N1820 = sent_n[53] & N4607;
  assign N4607 = ~fifo_yumi;
  assign N1822 = v_o[53] & ready_i[53];
  assign N1823 = ~N1822;
  assign v_o[54] = fifo_v & N4608;
  assign N4608 = ~sent_r[54];
  assign N1824 = ~reset_i;
  assign N1825 = reset_i;
  assign N1826 = sent_n[54] & N4609;
  assign N4609 = ~fifo_yumi;
  assign N1828 = v_o[54] & ready_i[54];
  assign N1829 = ~N1828;
  assign v_o[55] = fifo_v & N4610;
  assign N4610 = ~sent_r[55];
  assign N1830 = ~reset_i;
  assign N1831 = reset_i;
  assign N1832 = sent_n[55] & N4611;
  assign N4611 = ~fifo_yumi;
  assign N1834 = v_o[55] & ready_i[55];
  assign N1835 = ~N1834;
  assign v_o[56] = fifo_v & N4612;
  assign N4612 = ~sent_r[56];
  assign N1836 = ~reset_i;
  assign N1837 = reset_i;
  assign N1838 = sent_n[56] & N4613;
  assign N4613 = ~fifo_yumi;
  assign N1840 = v_o[56] & ready_i[56];
  assign N1841 = ~N1840;
  assign v_o[57] = fifo_v & N4614;
  assign N4614 = ~sent_r[57];
  assign N1842 = ~reset_i;
  assign N1843 = reset_i;
  assign N1844 = sent_n[57] & N4615;
  assign N4615 = ~fifo_yumi;
  assign N1846 = v_o[57] & ready_i[57];
  assign N1847 = ~N1846;
  assign v_o[58] = fifo_v & N4616;
  assign N4616 = ~sent_r[58];
  assign N1848 = ~reset_i;
  assign N1849 = reset_i;
  assign N1850 = sent_n[58] & N4617;
  assign N4617 = ~fifo_yumi;
  assign N1852 = v_o[58] & ready_i[58];
  assign N1853 = ~N1852;
  assign v_o[59] = fifo_v & N4618;
  assign N4618 = ~sent_r[59];
  assign N1854 = ~reset_i;
  assign N1855 = reset_i;
  assign N1856 = sent_n[59] & N4619;
  assign N4619 = ~fifo_yumi;
  assign N1858 = v_o[59] & ready_i[59];
  assign N1859 = ~N1858;
  assign v_o[60] = fifo_v & N4620;
  assign N4620 = ~sent_r[60];
  assign N1860 = ~reset_i;
  assign N1861 = reset_i;
  assign N1862 = sent_n[60] & N4621;
  assign N4621 = ~fifo_yumi;
  assign N1864 = v_o[60] & ready_i[60];
  assign N1865 = ~N1864;
  assign v_o[61] = fifo_v & N4622;
  assign N4622 = ~sent_r[61];
  assign N1866 = ~reset_i;
  assign N1867 = reset_i;
  assign N1868 = sent_n[61] & N4623;
  assign N4623 = ~fifo_yumi;
  assign N1870 = v_o[61] & ready_i[61];
  assign N1871 = ~N1870;
  assign v_o[62] = fifo_v & N4624;
  assign N4624 = ~sent_r[62];
  assign N1872 = ~reset_i;
  assign N1873 = reset_i;
  assign N1874 = sent_n[62] & N4625;
  assign N4625 = ~fifo_yumi;
  assign N1876 = v_o[62] & ready_i[62];
  assign N1877 = ~N1876;
  assign v_o[63] = fifo_v & N4626;
  assign N4626 = ~sent_r[63];
  assign N1878 = ~reset_i;
  assign N1879 = reset_i;
  assign N1880 = sent_n[63] & N4627;
  assign N4627 = ~fifo_yumi;
  assign N1882 = v_o[63] & ready_i[63];
  assign N1883 = ~N1882;
  assign v_o[64] = fifo_v & N4628;
  assign N4628 = ~sent_r[64];
  assign N1884 = ~reset_i;
  assign N1885 = reset_i;
  assign N1886 = sent_n[64] & N4629;
  assign N4629 = ~fifo_yumi;
  assign N1888 = v_o[64] & ready_i[64];
  assign N1889 = ~N1888;
  assign v_o[65] = fifo_v & N4630;
  assign N4630 = ~sent_r[65];
  assign N1890 = ~reset_i;
  assign N1891 = reset_i;
  assign N1892 = sent_n[65] & N4631;
  assign N4631 = ~fifo_yumi;
  assign N1894 = v_o[65] & ready_i[65];
  assign N1895 = ~N1894;
  assign v_o[66] = fifo_v & N4632;
  assign N4632 = ~sent_r[66];
  assign N1896 = ~reset_i;
  assign N1897 = reset_i;
  assign N1898 = sent_n[66] & N4633;
  assign N4633 = ~fifo_yumi;
  assign N1900 = v_o[66] & ready_i[66];
  assign N1901 = ~N1900;
  assign v_o[67] = fifo_v & N4634;
  assign N4634 = ~sent_r[67];
  assign N1902 = ~reset_i;
  assign N1903 = reset_i;
  assign N1904 = sent_n[67] & N4635;
  assign N4635 = ~fifo_yumi;
  assign N1906 = v_o[67] & ready_i[67];
  assign N1907 = ~N1906;
  assign v_o[68] = fifo_v & N4636;
  assign N4636 = ~sent_r[68];
  assign N1908 = ~reset_i;
  assign N1909 = reset_i;
  assign N1910 = sent_n[68] & N4637;
  assign N4637 = ~fifo_yumi;
  assign N1912 = v_o[68] & ready_i[68];
  assign N1913 = ~N1912;
  assign v_o[69] = fifo_v & N4638;
  assign N4638 = ~sent_r[69];
  assign N1914 = ~reset_i;
  assign N1915 = reset_i;
  assign N1916 = sent_n[69] & N4639;
  assign N4639 = ~fifo_yumi;
  assign N1918 = v_o[69] & ready_i[69];
  assign N1919 = ~N1918;
  assign v_o[70] = fifo_v & N4640;
  assign N4640 = ~sent_r[70];
  assign N1920 = ~reset_i;
  assign N1921 = reset_i;
  assign N1922 = sent_n[70] & N4641;
  assign N4641 = ~fifo_yumi;
  assign N1924 = v_o[70] & ready_i[70];
  assign N1925 = ~N1924;
  assign v_o[71] = fifo_v & N4642;
  assign N4642 = ~sent_r[71];
  assign N1926 = ~reset_i;
  assign N1927 = reset_i;
  assign N1928 = sent_n[71] & N4643;
  assign N4643 = ~fifo_yumi;
  assign N1930 = v_o[71] & ready_i[71];
  assign N1931 = ~N1930;
  assign v_o[72] = fifo_v & N4644;
  assign N4644 = ~sent_r[72];
  assign N1932 = ~reset_i;
  assign N1933 = reset_i;
  assign N1934 = sent_n[72] & N4645;
  assign N4645 = ~fifo_yumi;
  assign N1936 = v_o[72] & ready_i[72];
  assign N1937 = ~N1936;
  assign v_o[73] = fifo_v & N4646;
  assign N4646 = ~sent_r[73];
  assign N1938 = ~reset_i;
  assign N1939 = reset_i;
  assign N1940 = sent_n[73] & N4647;
  assign N4647 = ~fifo_yumi;
  assign N1942 = v_o[73] & ready_i[73];
  assign N1943 = ~N1942;
  assign v_o[74] = fifo_v & N4648;
  assign N4648 = ~sent_r[74];
  assign N1944 = ~reset_i;
  assign N1945 = reset_i;
  assign N1946 = sent_n[74] & N4649;
  assign N4649 = ~fifo_yumi;
  assign N1948 = v_o[74] & ready_i[74];
  assign N1949 = ~N1948;
  assign v_o[75] = fifo_v & N4650;
  assign N4650 = ~sent_r[75];
  assign N1950 = ~reset_i;
  assign N1951 = reset_i;
  assign N1952 = sent_n[75] & N4651;
  assign N4651 = ~fifo_yumi;
  assign N1954 = v_o[75] & ready_i[75];
  assign N1955 = ~N1954;
  assign v_o[76] = fifo_v & N4652;
  assign N4652 = ~sent_r[76];
  assign N1956 = ~reset_i;
  assign N1957 = reset_i;
  assign N1958 = sent_n[76] & N4653;
  assign N4653 = ~fifo_yumi;
  assign N1960 = v_o[76] & ready_i[76];
  assign N1961 = ~N1960;
  assign v_o[77] = fifo_v & N4654;
  assign N4654 = ~sent_r[77];
  assign N1962 = ~reset_i;
  assign N1963 = reset_i;
  assign N1964 = sent_n[77] & N4655;
  assign N4655 = ~fifo_yumi;
  assign N1966 = v_o[77] & ready_i[77];
  assign N1967 = ~N1966;
  assign v_o[78] = fifo_v & N4656;
  assign N4656 = ~sent_r[78];
  assign N1968 = ~reset_i;
  assign N1969 = reset_i;
  assign N1970 = sent_n[78] & N4657;
  assign N4657 = ~fifo_yumi;
  assign N1972 = v_o[78] & ready_i[78];
  assign N1973 = ~N1972;
  assign v_o[79] = fifo_v & N4658;
  assign N4658 = ~sent_r[79];
  assign N1974 = ~reset_i;
  assign N1975 = reset_i;
  assign N1976 = sent_n[79] & N4659;
  assign N4659 = ~fifo_yumi;
  assign N1978 = v_o[79] & ready_i[79];
  assign N1979 = ~N1978;
  assign v_o[80] = fifo_v & N4660;
  assign N4660 = ~sent_r[80];
  assign N1980 = ~reset_i;
  assign N1981 = reset_i;
  assign N1982 = sent_n[80] & N4661;
  assign N4661 = ~fifo_yumi;
  assign N1984 = v_o[80] & ready_i[80];
  assign N1985 = ~N1984;
  assign v_o[81] = fifo_v & N4662;
  assign N4662 = ~sent_r[81];
  assign N1986 = ~reset_i;
  assign N1987 = reset_i;
  assign N1988 = sent_n[81] & N4663;
  assign N4663 = ~fifo_yumi;
  assign N1990 = v_o[81] & ready_i[81];
  assign N1991 = ~N1990;
  assign v_o[82] = fifo_v & N4664;
  assign N4664 = ~sent_r[82];
  assign N1992 = ~reset_i;
  assign N1993 = reset_i;
  assign N1994 = sent_n[82] & N4665;
  assign N4665 = ~fifo_yumi;
  assign N1996 = v_o[82] & ready_i[82];
  assign N1997 = ~N1996;
  assign v_o[83] = fifo_v & N4666;
  assign N4666 = ~sent_r[83];
  assign N1998 = ~reset_i;
  assign N1999 = reset_i;
  assign N2000 = sent_n[83] & N4667;
  assign N4667 = ~fifo_yumi;
  assign N2002 = v_o[83] & ready_i[83];
  assign N2003 = ~N2002;
  assign v_o[84] = fifo_v & N4668;
  assign N4668 = ~sent_r[84];
  assign N2004 = ~reset_i;
  assign N2005 = reset_i;
  assign N2006 = sent_n[84] & N4669;
  assign N4669 = ~fifo_yumi;
  assign N2008 = v_o[84] & ready_i[84];
  assign N2009 = ~N2008;
  assign v_o[85] = fifo_v & N4670;
  assign N4670 = ~sent_r[85];
  assign N2010 = ~reset_i;
  assign N2011 = reset_i;
  assign N2012 = sent_n[85] & N4671;
  assign N4671 = ~fifo_yumi;
  assign N2014 = v_o[85] & ready_i[85];
  assign N2015 = ~N2014;
  assign v_o[86] = fifo_v & N4672;
  assign N4672 = ~sent_r[86];
  assign N2016 = ~reset_i;
  assign N2017 = reset_i;
  assign N2018 = sent_n[86] & N4673;
  assign N4673 = ~fifo_yumi;
  assign N2020 = v_o[86] & ready_i[86];
  assign N2021 = ~N2020;
  assign v_o[87] = fifo_v & N4674;
  assign N4674 = ~sent_r[87];
  assign N2022 = ~reset_i;
  assign N2023 = reset_i;
  assign N2024 = sent_n[87] & N4675;
  assign N4675 = ~fifo_yumi;
  assign N2026 = v_o[87] & ready_i[87];
  assign N2027 = ~N2026;
  assign v_o[88] = fifo_v & N4676;
  assign N4676 = ~sent_r[88];
  assign N2028 = ~reset_i;
  assign N2029 = reset_i;
  assign N2030 = sent_n[88] & N4677;
  assign N4677 = ~fifo_yumi;
  assign N2032 = v_o[88] & ready_i[88];
  assign N2033 = ~N2032;
  assign v_o[89] = fifo_v & N4678;
  assign N4678 = ~sent_r[89];
  assign N2034 = ~reset_i;
  assign N2035 = reset_i;
  assign N2036 = sent_n[89] & N4679;
  assign N4679 = ~fifo_yumi;
  assign N2038 = v_o[89] & ready_i[89];
  assign N2039 = ~N2038;
  assign v_o[90] = fifo_v & N4680;
  assign N4680 = ~sent_r[90];
  assign N2040 = ~reset_i;
  assign N2041 = reset_i;
  assign N2042 = sent_n[90] & N4681;
  assign N4681 = ~fifo_yumi;
  assign N2044 = v_o[90] & ready_i[90];
  assign N2045 = ~N2044;
  assign v_o[91] = fifo_v & N4682;
  assign N4682 = ~sent_r[91];
  assign N2046 = ~reset_i;
  assign N2047 = reset_i;
  assign N2048 = sent_n[91] & N4683;
  assign N4683 = ~fifo_yumi;
  assign N2050 = v_o[91] & ready_i[91];
  assign N2051 = ~N2050;
  assign v_o[92] = fifo_v & N4684;
  assign N4684 = ~sent_r[92];
  assign N2052 = ~reset_i;
  assign N2053 = reset_i;
  assign N2054 = sent_n[92] & N4685;
  assign N4685 = ~fifo_yumi;
  assign N2056 = v_o[92] & ready_i[92];
  assign N2057 = ~N2056;
  assign v_o[93] = fifo_v & N4686;
  assign N4686 = ~sent_r[93];
  assign N2058 = ~reset_i;
  assign N2059 = reset_i;
  assign N2060 = sent_n[93] & N4687;
  assign N4687 = ~fifo_yumi;
  assign N2062 = v_o[93] & ready_i[93];
  assign N2063 = ~N2062;
  assign v_o[94] = fifo_v & N4688;
  assign N4688 = ~sent_r[94];
  assign N2064 = ~reset_i;
  assign N2065 = reset_i;
  assign N2066 = sent_n[94] & N4689;
  assign N4689 = ~fifo_yumi;
  assign N2068 = v_o[94] & ready_i[94];
  assign N2069 = ~N2068;
  assign v_o[95] = fifo_v & N4690;
  assign N4690 = ~sent_r[95];
  assign N2070 = ~reset_i;
  assign N2071 = reset_i;
  assign N2072 = sent_n[95] & N4691;
  assign N4691 = ~fifo_yumi;
  assign N2074 = v_o[95] & ready_i[95];
  assign N2075 = ~N2074;
  assign v_o[96] = fifo_v & N4692;
  assign N4692 = ~sent_r[96];
  assign N2076 = ~reset_i;
  assign N2077 = reset_i;
  assign N2078 = sent_n[96] & N4693;
  assign N4693 = ~fifo_yumi;
  assign N2080 = v_o[96] & ready_i[96];
  assign N2081 = ~N2080;
  assign v_o[97] = fifo_v & N4694;
  assign N4694 = ~sent_r[97];
  assign N2082 = ~reset_i;
  assign N2083 = reset_i;
  assign N2084 = sent_n[97] & N4695;
  assign N4695 = ~fifo_yumi;
  assign N2086 = v_o[97] & ready_i[97];
  assign N2087 = ~N2086;
  assign v_o[98] = fifo_v & N4696;
  assign N4696 = ~sent_r[98];
  assign N2088 = ~reset_i;
  assign N2089 = reset_i;
  assign N2090 = sent_n[98] & N4697;
  assign N4697 = ~fifo_yumi;
  assign N2092 = v_o[98] & ready_i[98];
  assign N2093 = ~N2092;
  assign v_o[99] = fifo_v & N4698;
  assign N4698 = ~sent_r[99];
  assign N2094 = ~reset_i;
  assign N2095 = reset_i;
  assign N2096 = sent_n[99] & N4699;
  assign N4699 = ~fifo_yumi;
  assign N2098 = v_o[99] & ready_i[99];
  assign N2099 = ~N2098;
  assign v_o[100] = fifo_v & N4700;
  assign N4700 = ~sent_r[100];
  assign N2100 = ~reset_i;
  assign N2101 = reset_i;
  assign N2102 = sent_n[100] & N4701;
  assign N4701 = ~fifo_yumi;
  assign N2104 = v_o[100] & ready_i[100];
  assign N2105 = ~N2104;
  assign v_o[101] = fifo_v & N4702;
  assign N4702 = ~sent_r[101];
  assign N2106 = ~reset_i;
  assign N2107 = reset_i;
  assign N2108 = sent_n[101] & N4703;
  assign N4703 = ~fifo_yumi;
  assign N2110 = v_o[101] & ready_i[101];
  assign N2111 = ~N2110;
  assign v_o[102] = fifo_v & N4704;
  assign N4704 = ~sent_r[102];
  assign N2112 = ~reset_i;
  assign N2113 = reset_i;
  assign N2114 = sent_n[102] & N4705;
  assign N4705 = ~fifo_yumi;
  assign N2116 = v_o[102] & ready_i[102];
  assign N2117 = ~N2116;
  assign v_o[103] = fifo_v & N4706;
  assign N4706 = ~sent_r[103];
  assign N2118 = ~reset_i;
  assign N2119 = reset_i;
  assign N2120 = sent_n[103] & N4707;
  assign N4707 = ~fifo_yumi;
  assign N2122 = v_o[103] & ready_i[103];
  assign N2123 = ~N2122;
  assign v_o[104] = fifo_v & N4708;
  assign N4708 = ~sent_r[104];
  assign N2124 = ~reset_i;
  assign N2125 = reset_i;
  assign N2126 = sent_n[104] & N4709;
  assign N4709 = ~fifo_yumi;
  assign N2128 = v_o[104] & ready_i[104];
  assign N2129 = ~N2128;
  assign v_o[105] = fifo_v & N4710;
  assign N4710 = ~sent_r[105];
  assign N2130 = ~reset_i;
  assign N2131 = reset_i;
  assign N2132 = sent_n[105] & N4711;
  assign N4711 = ~fifo_yumi;
  assign N2134 = v_o[105] & ready_i[105];
  assign N2135 = ~N2134;
  assign v_o[106] = fifo_v & N4712;
  assign N4712 = ~sent_r[106];
  assign N2136 = ~reset_i;
  assign N2137 = reset_i;
  assign N2138 = sent_n[106] & N4713;
  assign N4713 = ~fifo_yumi;
  assign N2140 = v_o[106] & ready_i[106];
  assign N2141 = ~N2140;
  assign v_o[107] = fifo_v & N4714;
  assign N4714 = ~sent_r[107];
  assign N2142 = ~reset_i;
  assign N2143 = reset_i;
  assign N2144 = sent_n[107] & N4715;
  assign N4715 = ~fifo_yumi;
  assign N2146 = v_o[107] & ready_i[107];
  assign N2147 = ~N2146;
  assign v_o[108] = fifo_v & N4716;
  assign N4716 = ~sent_r[108];
  assign N2148 = ~reset_i;
  assign N2149 = reset_i;
  assign N2150 = sent_n[108] & N4717;
  assign N4717 = ~fifo_yumi;
  assign N2152 = v_o[108] & ready_i[108];
  assign N2153 = ~N2152;
  assign v_o[109] = fifo_v & N4718;
  assign N4718 = ~sent_r[109];
  assign N2154 = ~reset_i;
  assign N2155 = reset_i;
  assign N2156 = sent_n[109] & N4719;
  assign N4719 = ~fifo_yumi;
  assign N2158 = v_o[109] & ready_i[109];
  assign N2159 = ~N2158;
  assign v_o[110] = fifo_v & N4720;
  assign N4720 = ~sent_r[110];
  assign N2160 = ~reset_i;
  assign N2161 = reset_i;
  assign N2162 = sent_n[110] & N4721;
  assign N4721 = ~fifo_yumi;
  assign N2164 = v_o[110] & ready_i[110];
  assign N2165 = ~N2164;
  assign v_o[111] = fifo_v & N4722;
  assign N4722 = ~sent_r[111];
  assign N2166 = ~reset_i;
  assign N2167 = reset_i;
  assign N2168 = sent_n[111] & N4723;
  assign N4723 = ~fifo_yumi;
  assign N2170 = v_o[111] & ready_i[111];
  assign N2171 = ~N2170;
  assign v_o[112] = fifo_v & N4724;
  assign N4724 = ~sent_r[112];
  assign N2172 = ~reset_i;
  assign N2173 = reset_i;
  assign N2174 = sent_n[112] & N4725;
  assign N4725 = ~fifo_yumi;
  assign N2176 = v_o[112] & ready_i[112];
  assign N2177 = ~N2176;
  assign v_o[113] = fifo_v & N4726;
  assign N4726 = ~sent_r[113];
  assign N2178 = ~reset_i;
  assign N2179 = reset_i;
  assign N2180 = sent_n[113] & N4727;
  assign N4727 = ~fifo_yumi;
  assign N2182 = v_o[113] & ready_i[113];
  assign N2183 = ~N2182;
  assign v_o[114] = fifo_v & N4728;
  assign N4728 = ~sent_r[114];
  assign N2184 = ~reset_i;
  assign N2185 = reset_i;
  assign N2186 = sent_n[114] & N4729;
  assign N4729 = ~fifo_yumi;
  assign N2188 = v_o[114] & ready_i[114];
  assign N2189 = ~N2188;
  assign v_o[115] = fifo_v & N4730;
  assign N4730 = ~sent_r[115];
  assign N2190 = ~reset_i;
  assign N2191 = reset_i;
  assign N2192 = sent_n[115] & N4731;
  assign N4731 = ~fifo_yumi;
  assign N2194 = v_o[115] & ready_i[115];
  assign N2195 = ~N2194;
  assign v_o[116] = fifo_v & N4732;
  assign N4732 = ~sent_r[116];
  assign N2196 = ~reset_i;
  assign N2197 = reset_i;
  assign N2198 = sent_n[116] & N4733;
  assign N4733 = ~fifo_yumi;
  assign N2200 = v_o[116] & ready_i[116];
  assign N2201 = ~N2200;
  assign v_o[117] = fifo_v & N4734;
  assign N4734 = ~sent_r[117];
  assign N2202 = ~reset_i;
  assign N2203 = reset_i;
  assign N2204 = sent_n[117] & N4735;
  assign N4735 = ~fifo_yumi;
  assign N2206 = v_o[117] & ready_i[117];
  assign N2207 = ~N2206;
  assign v_o[118] = fifo_v & N4736;
  assign N4736 = ~sent_r[118];
  assign N2208 = ~reset_i;
  assign N2209 = reset_i;
  assign N2210 = sent_n[118] & N4737;
  assign N4737 = ~fifo_yumi;
  assign N2212 = v_o[118] & ready_i[118];
  assign N2213 = ~N2212;
  assign v_o[119] = fifo_v & N4738;
  assign N4738 = ~sent_r[119];
  assign N2214 = ~reset_i;
  assign N2215 = reset_i;
  assign N2216 = sent_n[119] & N4739;
  assign N4739 = ~fifo_yumi;
  assign N2218 = v_o[119] & ready_i[119];
  assign N2219 = ~N2218;
  assign v_o[120] = fifo_v & N4740;
  assign N4740 = ~sent_r[120];
  assign N2220 = ~reset_i;
  assign N2221 = reset_i;
  assign N2222 = sent_n[120] & N4741;
  assign N4741 = ~fifo_yumi;
  assign N2224 = v_o[120] & ready_i[120];
  assign N2225 = ~N2224;
  assign v_o[121] = fifo_v & N4742;
  assign N4742 = ~sent_r[121];
  assign N2226 = ~reset_i;
  assign N2227 = reset_i;
  assign N2228 = sent_n[121] & N4743;
  assign N4743 = ~fifo_yumi;
  assign N2230 = v_o[121] & ready_i[121];
  assign N2231 = ~N2230;
  assign v_o[122] = fifo_v & N4744;
  assign N4744 = ~sent_r[122];
  assign N2232 = ~reset_i;
  assign N2233 = reset_i;
  assign N2234 = sent_n[122] & N4745;
  assign N4745 = ~fifo_yumi;
  assign N2236 = v_o[122] & ready_i[122];
  assign N2237 = ~N2236;
  assign v_o[123] = fifo_v & N4746;
  assign N4746 = ~sent_r[123];
  assign N2238 = ~reset_i;
  assign N2239 = reset_i;
  assign N2240 = sent_n[123] & N4747;
  assign N4747 = ~fifo_yumi;
  assign N2242 = v_o[123] & ready_i[123];
  assign N2243 = ~N2242;
  assign v_o[124] = fifo_v & N4748;
  assign N4748 = ~sent_r[124];
  assign N2244 = ~reset_i;
  assign N2245 = reset_i;
  assign N2246 = sent_n[124] & N4749;
  assign N4749 = ~fifo_yumi;
  assign N2248 = v_o[124] & ready_i[124];
  assign N2249 = ~N2248;
  assign v_o[125] = fifo_v & N4750;
  assign N4750 = ~sent_r[125];
  assign N2250 = ~reset_i;
  assign N2251 = reset_i;
  assign N2252 = sent_n[125] & N4751;
  assign N4751 = ~fifo_yumi;
  assign N2254 = v_o[125] & ready_i[125];
  assign N2255 = ~N2254;
  assign v_o[126] = fifo_v & N4752;
  assign N4752 = ~sent_r[126];
  assign N2256 = ~reset_i;
  assign N2257 = reset_i;
  assign N2258 = sent_n[126] & N4753;
  assign N4753 = ~fifo_yumi;
  assign N2260 = v_o[126] & ready_i[126];
  assign N2261 = ~N2260;
  assign v_o[127] = fifo_v & N4754;
  assign N4754 = ~sent_r[127];
  assign N2262 = ~reset_i;
  assign N2263 = reset_i;
  assign N2264 = sent_n[127] & N4755;
  assign N4755 = ~fifo_yumi;
  assign N2266 = v_o[127] & ready_i[127];
  assign N2267 = ~N2266;
  assign v_o[128] = fifo_v & N4756;
  assign N4756 = ~sent_r[128];
  assign N2268 = ~reset_i;
  assign N2269 = reset_i;
  assign N2270 = sent_n[128] & N4757;
  assign N4757 = ~fifo_yumi;
  assign N2272 = v_o[128] & ready_i[128];
  assign N2273 = ~N2272;
  assign v_o[129] = fifo_v & N4758;
  assign N4758 = ~sent_r[129];
  assign N2274 = ~reset_i;
  assign N2275 = reset_i;
  assign N2276 = sent_n[129] & N4759;
  assign N4759 = ~fifo_yumi;
  assign N2278 = v_o[129] & ready_i[129];
  assign N2279 = ~N2278;
  assign v_o[130] = fifo_v & N4760;
  assign N4760 = ~sent_r[130];
  assign N2280 = ~reset_i;
  assign N2281 = reset_i;
  assign N2282 = sent_n[130] & N4761;
  assign N4761 = ~fifo_yumi;
  assign N2284 = v_o[130] & ready_i[130];
  assign N2285 = ~N2284;
  assign v_o[131] = fifo_v & N4762;
  assign N4762 = ~sent_r[131];
  assign N2286 = ~reset_i;
  assign N2287 = reset_i;
  assign N2288 = sent_n[131] & N4763;
  assign N4763 = ~fifo_yumi;
  assign N2290 = v_o[131] & ready_i[131];
  assign N2291 = ~N2290;
  assign v_o[132] = fifo_v & N4764;
  assign N4764 = ~sent_r[132];
  assign N2292 = ~reset_i;
  assign N2293 = reset_i;
  assign N2294 = sent_n[132] & N4765;
  assign N4765 = ~fifo_yumi;
  assign N2296 = v_o[132] & ready_i[132];
  assign N2297 = ~N2296;
  assign v_o[133] = fifo_v & N4766;
  assign N4766 = ~sent_r[133];
  assign N2298 = ~reset_i;
  assign N2299 = reset_i;
  assign N2300 = sent_n[133] & N4767;
  assign N4767 = ~fifo_yumi;
  assign N2302 = v_o[133] & ready_i[133];
  assign N2303 = ~N2302;
  assign v_o[134] = fifo_v & N4768;
  assign N4768 = ~sent_r[134];
  assign N2304 = ~reset_i;
  assign N2305 = reset_i;
  assign N2306 = sent_n[134] & N4769;
  assign N4769 = ~fifo_yumi;
  assign N2308 = v_o[134] & ready_i[134];
  assign N2309 = ~N2308;
  assign v_o[135] = fifo_v & N4770;
  assign N4770 = ~sent_r[135];
  assign N2310 = ~reset_i;
  assign N2311 = reset_i;
  assign N2312 = sent_n[135] & N4771;
  assign N4771 = ~fifo_yumi;
  assign N2314 = v_o[135] & ready_i[135];
  assign N2315 = ~N2314;
  assign v_o[136] = fifo_v & N4772;
  assign N4772 = ~sent_r[136];
  assign N2316 = ~reset_i;
  assign N2317 = reset_i;
  assign N2318 = sent_n[136] & N4773;
  assign N4773 = ~fifo_yumi;
  assign N2320 = v_o[136] & ready_i[136];
  assign N2321 = ~N2320;
  assign v_o[137] = fifo_v & N4774;
  assign N4774 = ~sent_r[137];
  assign N2322 = ~reset_i;
  assign N2323 = reset_i;
  assign N2324 = sent_n[137] & N4775;
  assign N4775 = ~fifo_yumi;
  assign N2326 = v_o[137] & ready_i[137];
  assign N2327 = ~N2326;
  assign v_o[138] = fifo_v & N4776;
  assign N4776 = ~sent_r[138];
  assign N2328 = ~reset_i;
  assign N2329 = reset_i;
  assign N2330 = sent_n[138] & N4777;
  assign N4777 = ~fifo_yumi;
  assign N2332 = v_o[138] & ready_i[138];
  assign N2333 = ~N2332;
  assign v_o[139] = fifo_v & N4778;
  assign N4778 = ~sent_r[139];
  assign N2334 = ~reset_i;
  assign N2335 = reset_i;
  assign N2336 = sent_n[139] & N4779;
  assign N4779 = ~fifo_yumi;
  assign N2338 = v_o[139] & ready_i[139];
  assign N2339 = ~N2338;
  assign v_o[140] = fifo_v & N4780;
  assign N4780 = ~sent_r[140];
  assign N2340 = ~reset_i;
  assign N2341 = reset_i;
  assign N2342 = sent_n[140] & N4781;
  assign N4781 = ~fifo_yumi;
  assign N2344 = v_o[140] & ready_i[140];
  assign N2345 = ~N2344;
  assign v_o[141] = fifo_v & N4782;
  assign N4782 = ~sent_r[141];
  assign N2346 = ~reset_i;
  assign N2347 = reset_i;
  assign N2348 = sent_n[141] & N4783;
  assign N4783 = ~fifo_yumi;
  assign N2350 = v_o[141] & ready_i[141];
  assign N2351 = ~N2350;
  assign v_o[142] = fifo_v & N4784;
  assign N4784 = ~sent_r[142];
  assign N2352 = ~reset_i;
  assign N2353 = reset_i;
  assign N2354 = sent_n[142] & N4785;
  assign N4785 = ~fifo_yumi;
  assign N2356 = v_o[142] & ready_i[142];
  assign N2357 = ~N2356;
  assign v_o[143] = fifo_v & N4786;
  assign N4786 = ~sent_r[143];
  assign N2358 = ~reset_i;
  assign N2359 = reset_i;
  assign N2360 = sent_n[143] & N4787;
  assign N4787 = ~fifo_yumi;
  assign N2362 = v_o[143] & ready_i[143];
  assign N2363 = ~N2362;
  assign v_o[144] = fifo_v & N4788;
  assign N4788 = ~sent_r[144];
  assign N2364 = ~reset_i;
  assign N2365 = reset_i;
  assign N2366 = sent_n[144] & N4789;
  assign N4789 = ~fifo_yumi;
  assign N2368 = v_o[144] & ready_i[144];
  assign N2369 = ~N2368;
  assign v_o[145] = fifo_v & N4790;
  assign N4790 = ~sent_r[145];
  assign N2370 = ~reset_i;
  assign N2371 = reset_i;
  assign N2372 = sent_n[145] & N4791;
  assign N4791 = ~fifo_yumi;
  assign N2374 = v_o[145] & ready_i[145];
  assign N2375 = ~N2374;
  assign v_o[146] = fifo_v & N4792;
  assign N4792 = ~sent_r[146];
  assign N2376 = ~reset_i;
  assign N2377 = reset_i;
  assign N2378 = sent_n[146] & N4793;
  assign N4793 = ~fifo_yumi;
  assign N2380 = v_o[146] & ready_i[146];
  assign N2381 = ~N2380;
  assign v_o[147] = fifo_v & N4794;
  assign N4794 = ~sent_r[147];
  assign N2382 = ~reset_i;
  assign N2383 = reset_i;
  assign N2384 = sent_n[147] & N4795;
  assign N4795 = ~fifo_yumi;
  assign N2386 = v_o[147] & ready_i[147];
  assign N2387 = ~N2386;
  assign v_o[148] = fifo_v & N4796;
  assign N4796 = ~sent_r[148];
  assign N2388 = ~reset_i;
  assign N2389 = reset_i;
  assign N2390 = sent_n[148] & N4797;
  assign N4797 = ~fifo_yumi;
  assign N2392 = v_o[148] & ready_i[148];
  assign N2393 = ~N2392;
  assign v_o[149] = fifo_v & N4798;
  assign N4798 = ~sent_r[149];
  assign N2394 = ~reset_i;
  assign N2395 = reset_i;
  assign N2396 = sent_n[149] & N4799;
  assign N4799 = ~fifo_yumi;
  assign N2398 = v_o[149] & ready_i[149];
  assign N2399 = ~N2398;
  assign v_o[150] = fifo_v & N4800;
  assign N4800 = ~sent_r[150];
  assign N2400 = ~reset_i;
  assign N2401 = reset_i;
  assign N2402 = sent_n[150] & N4801;
  assign N4801 = ~fifo_yumi;
  assign N2404 = v_o[150] & ready_i[150];
  assign N2405 = ~N2404;
  assign v_o[151] = fifo_v & N4802;
  assign N4802 = ~sent_r[151];
  assign N2406 = ~reset_i;
  assign N2407 = reset_i;
  assign N2408 = sent_n[151] & N4803;
  assign N4803 = ~fifo_yumi;
  assign N2410 = v_o[151] & ready_i[151];
  assign N2411 = ~N2410;
  assign v_o[152] = fifo_v & N4804;
  assign N4804 = ~sent_r[152];
  assign N2412 = ~reset_i;
  assign N2413 = reset_i;
  assign N2414 = sent_n[152] & N4805;
  assign N4805 = ~fifo_yumi;
  assign N2416 = v_o[152] & ready_i[152];
  assign N2417 = ~N2416;
  assign v_o[153] = fifo_v & N4806;
  assign N4806 = ~sent_r[153];
  assign N2418 = ~reset_i;
  assign N2419 = reset_i;
  assign N2420 = sent_n[153] & N4807;
  assign N4807 = ~fifo_yumi;
  assign N2422 = v_o[153] & ready_i[153];
  assign N2423 = ~N2422;
  assign v_o[154] = fifo_v & N4808;
  assign N4808 = ~sent_r[154];
  assign N2424 = ~reset_i;
  assign N2425 = reset_i;
  assign N2426 = sent_n[154] & N4809;
  assign N4809 = ~fifo_yumi;
  assign N2428 = v_o[154] & ready_i[154];
  assign N2429 = ~N2428;
  assign v_o[155] = fifo_v & N4810;
  assign N4810 = ~sent_r[155];
  assign N2430 = ~reset_i;
  assign N2431 = reset_i;
  assign N2432 = sent_n[155] & N4811;
  assign N4811 = ~fifo_yumi;
  assign N2434 = v_o[155] & ready_i[155];
  assign N2435 = ~N2434;
  assign v_o[156] = fifo_v & N4812;
  assign N4812 = ~sent_r[156];
  assign N2436 = ~reset_i;
  assign N2437 = reset_i;
  assign N2438 = sent_n[156] & N4813;
  assign N4813 = ~fifo_yumi;
  assign N2440 = v_o[156] & ready_i[156];
  assign N2441 = ~N2440;
  assign v_o[157] = fifo_v & N4814;
  assign N4814 = ~sent_r[157];
  assign N2442 = ~reset_i;
  assign N2443 = reset_i;
  assign N2444 = sent_n[157] & N4815;
  assign N4815 = ~fifo_yumi;
  assign N2446 = v_o[157] & ready_i[157];
  assign N2447 = ~N2446;
  assign v_o[158] = fifo_v & N4816;
  assign N4816 = ~sent_r[158];
  assign N2448 = ~reset_i;
  assign N2449 = reset_i;
  assign N2450 = sent_n[158] & N4817;
  assign N4817 = ~fifo_yumi;
  assign N2452 = v_o[158] & ready_i[158];
  assign N2453 = ~N2452;
  assign v_o[159] = fifo_v & N4818;
  assign N4818 = ~sent_r[159];
  assign N2454 = ~reset_i;
  assign N2455 = reset_i;
  assign N2456 = sent_n[159] & N4819;
  assign N4819 = ~fifo_yumi;
  assign N2458 = v_o[159] & ready_i[159];
  assign N2459 = ~N2458;
  assign v_o[160] = fifo_v & N4820;
  assign N4820 = ~sent_r[160];
  assign N2460 = ~reset_i;
  assign N2461 = reset_i;
  assign N2462 = sent_n[160] & N4821;
  assign N4821 = ~fifo_yumi;
  assign N2464 = v_o[160] & ready_i[160];
  assign N2465 = ~N2464;
  assign v_o[161] = fifo_v & N4822;
  assign N4822 = ~sent_r[161];
  assign N2466 = ~reset_i;
  assign N2467 = reset_i;
  assign N2468 = sent_n[161] & N4823;
  assign N4823 = ~fifo_yumi;
  assign N2470 = v_o[161] & ready_i[161];
  assign N2471 = ~N2470;
  assign v_o[162] = fifo_v & N4824;
  assign N4824 = ~sent_r[162];
  assign N2472 = ~reset_i;
  assign N2473 = reset_i;
  assign N2474 = sent_n[162] & N4825;
  assign N4825 = ~fifo_yumi;
  assign N2476 = v_o[162] & ready_i[162];
  assign N2477 = ~N2476;
  assign v_o[163] = fifo_v & N4826;
  assign N4826 = ~sent_r[163];
  assign N2478 = ~reset_i;
  assign N2479 = reset_i;
  assign N2480 = sent_n[163] & N4827;
  assign N4827 = ~fifo_yumi;
  assign N2482 = v_o[163] & ready_i[163];
  assign N2483 = ~N2482;
  assign v_o[164] = fifo_v & N4828;
  assign N4828 = ~sent_r[164];
  assign N2484 = ~reset_i;
  assign N2485 = reset_i;
  assign N2486 = sent_n[164] & N4829;
  assign N4829 = ~fifo_yumi;
  assign N2488 = v_o[164] & ready_i[164];
  assign N2489 = ~N2488;
  assign v_o[165] = fifo_v & N4830;
  assign N4830 = ~sent_r[165];
  assign N2490 = ~reset_i;
  assign N2491 = reset_i;
  assign N2492 = sent_n[165] & N4831;
  assign N4831 = ~fifo_yumi;
  assign N2494 = v_o[165] & ready_i[165];
  assign N2495 = ~N2494;
  assign v_o[166] = fifo_v & N4832;
  assign N4832 = ~sent_r[166];
  assign N2496 = ~reset_i;
  assign N2497 = reset_i;
  assign N2498 = sent_n[166] & N4833;
  assign N4833 = ~fifo_yumi;
  assign N2500 = v_o[166] & ready_i[166];
  assign N2501 = ~N2500;
  assign v_o[167] = fifo_v & N4834;
  assign N4834 = ~sent_r[167];
  assign N2502 = ~reset_i;
  assign N2503 = reset_i;
  assign N2504 = sent_n[167] & N4835;
  assign N4835 = ~fifo_yumi;
  assign N2506 = v_o[167] & ready_i[167];
  assign N2507 = ~N2506;
  assign v_o[168] = fifo_v & N4836;
  assign N4836 = ~sent_r[168];
  assign N2508 = ~reset_i;
  assign N2509 = reset_i;
  assign N2510 = sent_n[168] & N4837;
  assign N4837 = ~fifo_yumi;
  assign N2512 = v_o[168] & ready_i[168];
  assign N2513 = ~N2512;
  assign v_o[169] = fifo_v & N4838;
  assign N4838 = ~sent_r[169];
  assign N2514 = ~reset_i;
  assign N2515 = reset_i;
  assign N2516 = sent_n[169] & N4839;
  assign N4839 = ~fifo_yumi;
  assign N2518 = v_o[169] & ready_i[169];
  assign N2519 = ~N2518;
  assign v_o[170] = fifo_v & N4840;
  assign N4840 = ~sent_r[170];
  assign N2520 = ~reset_i;
  assign N2521 = reset_i;
  assign N2522 = sent_n[170] & N4841;
  assign N4841 = ~fifo_yumi;
  assign N2524 = v_o[170] & ready_i[170];
  assign N2525 = ~N2524;
  assign v_o[171] = fifo_v & N4842;
  assign N4842 = ~sent_r[171];
  assign N2526 = ~reset_i;
  assign N2527 = reset_i;
  assign N2528 = sent_n[171] & N4843;
  assign N4843 = ~fifo_yumi;
  assign N2530 = v_o[171] & ready_i[171];
  assign N2531 = ~N2530;
  assign v_o[172] = fifo_v & N4844;
  assign N4844 = ~sent_r[172];
  assign N2532 = ~reset_i;
  assign N2533 = reset_i;
  assign N2534 = sent_n[172] & N4845;
  assign N4845 = ~fifo_yumi;
  assign N2536 = v_o[172] & ready_i[172];
  assign N2537 = ~N2536;
  assign v_o[173] = fifo_v & N4846;
  assign N4846 = ~sent_r[173];
  assign N2538 = ~reset_i;
  assign N2539 = reset_i;
  assign N2540 = sent_n[173] & N4847;
  assign N4847 = ~fifo_yumi;
  assign N2542 = v_o[173] & ready_i[173];
  assign N2543 = ~N2542;
  assign v_o[174] = fifo_v & N4848;
  assign N4848 = ~sent_r[174];
  assign N2544 = ~reset_i;
  assign N2545 = reset_i;
  assign N2546 = sent_n[174] & N4849;
  assign N4849 = ~fifo_yumi;
  assign N2548 = v_o[174] & ready_i[174];
  assign N2549 = ~N2548;
  assign v_o[175] = fifo_v & N4850;
  assign N4850 = ~sent_r[175];
  assign N2550 = ~reset_i;
  assign N2551 = reset_i;
  assign N2552 = sent_n[175] & N4851;
  assign N4851 = ~fifo_yumi;
  assign N2554 = v_o[175] & ready_i[175];
  assign N2555 = ~N2554;
  assign v_o[176] = fifo_v & N4852;
  assign N4852 = ~sent_r[176];
  assign N2556 = ~reset_i;
  assign N2557 = reset_i;
  assign N2558 = sent_n[176] & N4853;
  assign N4853 = ~fifo_yumi;
  assign N2560 = v_o[176] & ready_i[176];
  assign N2561 = ~N2560;
  assign v_o[177] = fifo_v & N4854;
  assign N4854 = ~sent_r[177];
  assign N2562 = ~reset_i;
  assign N2563 = reset_i;
  assign N2564 = sent_n[177] & N4855;
  assign N4855 = ~fifo_yumi;
  assign N2566 = v_o[177] & ready_i[177];
  assign N2567 = ~N2566;
  assign v_o[178] = fifo_v & N4856;
  assign N4856 = ~sent_r[178];
  assign N2568 = ~reset_i;
  assign N2569 = reset_i;
  assign N2570 = sent_n[178] & N4857;
  assign N4857 = ~fifo_yumi;
  assign N2572 = v_o[178] & ready_i[178];
  assign N2573 = ~N2572;
  assign v_o[179] = fifo_v & N4858;
  assign N4858 = ~sent_r[179];
  assign N2574 = ~reset_i;
  assign N2575 = reset_i;
  assign N2576 = sent_n[179] & N4859;
  assign N4859 = ~fifo_yumi;
  assign N2578 = v_o[179] & ready_i[179];
  assign N2579 = ~N2578;
  assign v_o[180] = fifo_v & N4860;
  assign N4860 = ~sent_r[180];
  assign N2580 = ~reset_i;
  assign N2581 = reset_i;
  assign N2582 = sent_n[180] & N4861;
  assign N4861 = ~fifo_yumi;
  assign N2584 = v_o[180] & ready_i[180];
  assign N2585 = ~N2584;
  assign v_o[181] = fifo_v & N4862;
  assign N4862 = ~sent_r[181];
  assign N2586 = ~reset_i;
  assign N2587 = reset_i;
  assign N2588 = sent_n[181] & N4863;
  assign N4863 = ~fifo_yumi;
  assign N2590 = v_o[181] & ready_i[181];
  assign N2591 = ~N2590;
  assign v_o[182] = fifo_v & N4864;
  assign N4864 = ~sent_r[182];
  assign N2592 = ~reset_i;
  assign N2593 = reset_i;
  assign N2594 = sent_n[182] & N4865;
  assign N4865 = ~fifo_yumi;
  assign N2596 = v_o[182] & ready_i[182];
  assign N2597 = ~N2596;
  assign v_o[183] = fifo_v & N4866;
  assign N4866 = ~sent_r[183];
  assign N2598 = ~reset_i;
  assign N2599 = reset_i;
  assign N2600 = sent_n[183] & N4867;
  assign N4867 = ~fifo_yumi;
  assign N2602 = v_o[183] & ready_i[183];
  assign N2603 = ~N2602;
  assign v_o[184] = fifo_v & N4868;
  assign N4868 = ~sent_r[184];
  assign N2604 = ~reset_i;
  assign N2605 = reset_i;
  assign N2606 = sent_n[184] & N4869;
  assign N4869 = ~fifo_yumi;
  assign N2608 = v_o[184] & ready_i[184];
  assign N2609 = ~N2608;
  assign v_o[185] = fifo_v & N4870;
  assign N4870 = ~sent_r[185];
  assign N2610 = ~reset_i;
  assign N2611 = reset_i;
  assign N2612 = sent_n[185] & N4871;
  assign N4871 = ~fifo_yumi;
  assign N2614 = v_o[185] & ready_i[185];
  assign N2615 = ~N2614;
  assign v_o[186] = fifo_v & N4872;
  assign N4872 = ~sent_r[186];
  assign N2616 = ~reset_i;
  assign N2617 = reset_i;
  assign N2618 = sent_n[186] & N4873;
  assign N4873 = ~fifo_yumi;
  assign N2620 = v_o[186] & ready_i[186];
  assign N2621 = ~N2620;
  assign v_o[187] = fifo_v & N4874;
  assign N4874 = ~sent_r[187];
  assign N2622 = ~reset_i;
  assign N2623 = reset_i;
  assign N2624 = sent_n[187] & N4875;
  assign N4875 = ~fifo_yumi;
  assign N2626 = v_o[187] & ready_i[187];
  assign N2627 = ~N2626;
  assign v_o[188] = fifo_v & N4876;
  assign N4876 = ~sent_r[188];
  assign N2628 = ~reset_i;
  assign N2629 = reset_i;
  assign N2630 = sent_n[188] & N4877;
  assign N4877 = ~fifo_yumi;
  assign N2632 = v_o[188] & ready_i[188];
  assign N2633 = ~N2632;
  assign v_o[189] = fifo_v & N4878;
  assign N4878 = ~sent_r[189];
  assign N2634 = ~reset_i;
  assign N2635 = reset_i;
  assign N2636 = sent_n[189] & N4879;
  assign N4879 = ~fifo_yumi;
  assign N2638 = v_o[189] & ready_i[189];
  assign N2639 = ~N2638;
  assign v_o[190] = fifo_v & N4880;
  assign N4880 = ~sent_r[190];
  assign N2640 = ~reset_i;
  assign N2641 = reset_i;
  assign N2642 = sent_n[190] & N4881;
  assign N4881 = ~fifo_yumi;
  assign N2644 = v_o[190] & ready_i[190];
  assign N2645 = ~N2644;
  assign v_o[191] = fifo_v & N4882;
  assign N4882 = ~sent_r[191];
  assign N2646 = ~reset_i;
  assign N2647 = reset_i;
  assign N2648 = sent_n[191] & N4883;
  assign N4883 = ~fifo_yumi;
  assign N2650 = v_o[191] & ready_i[191];
  assign N2651 = ~N2650;
  assign v_o[192] = fifo_v & N4884;
  assign N4884 = ~sent_r[192];
  assign N2652 = ~reset_i;
  assign N2653 = reset_i;
  assign N2654 = sent_n[192] & N4885;
  assign N4885 = ~fifo_yumi;
  assign N2656 = v_o[192] & ready_i[192];
  assign N2657 = ~N2656;
  assign v_o[193] = fifo_v & N4886;
  assign N4886 = ~sent_r[193];
  assign N2658 = ~reset_i;
  assign N2659 = reset_i;
  assign N2660 = sent_n[193] & N4887;
  assign N4887 = ~fifo_yumi;
  assign N2662 = v_o[193] & ready_i[193];
  assign N2663 = ~N2662;
  assign v_o[194] = fifo_v & N4888;
  assign N4888 = ~sent_r[194];
  assign N2664 = ~reset_i;
  assign N2665 = reset_i;
  assign N2666 = sent_n[194] & N4889;
  assign N4889 = ~fifo_yumi;
  assign N2668 = v_o[194] & ready_i[194];
  assign N2669 = ~N2668;
  assign v_o[195] = fifo_v & N4890;
  assign N4890 = ~sent_r[195];
  assign N2670 = ~reset_i;
  assign N2671 = reset_i;
  assign N2672 = sent_n[195] & N4891;
  assign N4891 = ~fifo_yumi;
  assign N2674 = v_o[195] & ready_i[195];
  assign N2675 = ~N2674;
  assign v_o[196] = fifo_v & N4892;
  assign N4892 = ~sent_r[196];
  assign N2676 = ~reset_i;
  assign N2677 = reset_i;
  assign N2678 = sent_n[196] & N4893;
  assign N4893 = ~fifo_yumi;
  assign N2680 = v_o[196] & ready_i[196];
  assign N2681 = ~N2680;
  assign v_o[197] = fifo_v & N4894;
  assign N4894 = ~sent_r[197];
  assign N2682 = ~reset_i;
  assign N2683 = reset_i;
  assign N2684 = sent_n[197] & N4895;
  assign N4895 = ~fifo_yumi;
  assign N2686 = v_o[197] & ready_i[197];
  assign N2687 = ~N2686;
  assign v_o[198] = fifo_v & N4896;
  assign N4896 = ~sent_r[198];
  assign N2688 = ~reset_i;
  assign N2689 = reset_i;
  assign N2690 = sent_n[198] & N4897;
  assign N4897 = ~fifo_yumi;
  assign N2692 = v_o[198] & ready_i[198];
  assign N2693 = ~N2692;
  assign v_o[199] = fifo_v & N4898;
  assign N4898 = ~sent_r[199];
  assign N2694 = ~reset_i;
  assign N2695 = reset_i;
  assign N2696 = sent_n[199] & N4899;
  assign N4899 = ~fifo_yumi;
  assign N2698 = v_o[199] & ready_i[199];
  assign N2699 = ~N2698;
  assign v_o[200] = fifo_v & N4900;
  assign N4900 = ~sent_r[200];
  assign N2700 = ~reset_i;
  assign N2701 = reset_i;
  assign N2702 = sent_n[200] & N4901;
  assign N4901 = ~fifo_yumi;
  assign N2704 = v_o[200] & ready_i[200];
  assign N2705 = ~N2704;
  assign v_o[201] = fifo_v & N4902;
  assign N4902 = ~sent_r[201];
  assign N2706 = ~reset_i;
  assign N2707 = reset_i;
  assign N2708 = sent_n[201] & N4903;
  assign N4903 = ~fifo_yumi;
  assign N2710 = v_o[201] & ready_i[201];
  assign N2711 = ~N2710;
  assign v_o[202] = fifo_v & N4904;
  assign N4904 = ~sent_r[202];
  assign N2712 = ~reset_i;
  assign N2713 = reset_i;
  assign N2714 = sent_n[202] & N4905;
  assign N4905 = ~fifo_yumi;
  assign N2716 = v_o[202] & ready_i[202];
  assign N2717 = ~N2716;
  assign v_o[203] = fifo_v & N4906;
  assign N4906 = ~sent_r[203];
  assign N2718 = ~reset_i;
  assign N2719 = reset_i;
  assign N2720 = sent_n[203] & N4907;
  assign N4907 = ~fifo_yumi;
  assign N2722 = v_o[203] & ready_i[203];
  assign N2723 = ~N2722;
  assign v_o[204] = fifo_v & N4908;
  assign N4908 = ~sent_r[204];
  assign N2724 = ~reset_i;
  assign N2725 = reset_i;
  assign N2726 = sent_n[204] & N4909;
  assign N4909 = ~fifo_yumi;
  assign N2728 = v_o[204] & ready_i[204];
  assign N2729 = ~N2728;
  assign v_o[205] = fifo_v & N4910;
  assign N4910 = ~sent_r[205];
  assign N2730 = ~reset_i;
  assign N2731 = reset_i;
  assign N2732 = sent_n[205] & N4911;
  assign N4911 = ~fifo_yumi;
  assign N2734 = v_o[205] & ready_i[205];
  assign N2735 = ~N2734;
  assign v_o[206] = fifo_v & N4912;
  assign N4912 = ~sent_r[206];
  assign N2736 = ~reset_i;
  assign N2737 = reset_i;
  assign N2738 = sent_n[206] & N4913;
  assign N4913 = ~fifo_yumi;
  assign N2740 = v_o[206] & ready_i[206];
  assign N2741 = ~N2740;
  assign v_o[207] = fifo_v & N4914;
  assign N4914 = ~sent_r[207];
  assign N2742 = ~reset_i;
  assign N2743 = reset_i;
  assign N2744 = sent_n[207] & N4915;
  assign N4915 = ~fifo_yumi;
  assign N2746 = v_o[207] & ready_i[207];
  assign N2747 = ~N2746;
  assign v_o[208] = fifo_v & N4916;
  assign N4916 = ~sent_r[208];
  assign N2748 = ~reset_i;
  assign N2749 = reset_i;
  assign N2750 = sent_n[208] & N4917;
  assign N4917 = ~fifo_yumi;
  assign N2752 = v_o[208] & ready_i[208];
  assign N2753 = ~N2752;
  assign v_o[209] = fifo_v & N4918;
  assign N4918 = ~sent_r[209];
  assign N2754 = ~reset_i;
  assign N2755 = reset_i;
  assign N2756 = sent_n[209] & N4919;
  assign N4919 = ~fifo_yumi;
  assign N2758 = v_o[209] & ready_i[209];
  assign N2759 = ~N2758;
  assign v_o[210] = fifo_v & N4920;
  assign N4920 = ~sent_r[210];
  assign N2760 = ~reset_i;
  assign N2761 = reset_i;
  assign N2762 = sent_n[210] & N4921;
  assign N4921 = ~fifo_yumi;
  assign N2764 = v_o[210] & ready_i[210];
  assign N2765 = ~N2764;
  assign v_o[211] = fifo_v & N4922;
  assign N4922 = ~sent_r[211];
  assign N2766 = ~reset_i;
  assign N2767 = reset_i;
  assign N2768 = sent_n[211] & N4923;
  assign N4923 = ~fifo_yumi;
  assign N2770 = v_o[211] & ready_i[211];
  assign N2771 = ~N2770;
  assign v_o[212] = fifo_v & N4924;
  assign N4924 = ~sent_r[212];
  assign N2772 = ~reset_i;
  assign N2773 = reset_i;
  assign N2774 = sent_n[212] & N4925;
  assign N4925 = ~fifo_yumi;
  assign N2776 = v_o[212] & ready_i[212];
  assign N2777 = ~N2776;
  assign v_o[213] = fifo_v & N4926;
  assign N4926 = ~sent_r[213];
  assign N2778 = ~reset_i;
  assign N2779 = reset_i;
  assign N2780 = sent_n[213] & N4927;
  assign N4927 = ~fifo_yumi;
  assign N2782 = v_o[213] & ready_i[213];
  assign N2783 = ~N2782;
  assign v_o[214] = fifo_v & N4928;
  assign N4928 = ~sent_r[214];
  assign N2784 = ~reset_i;
  assign N2785 = reset_i;
  assign N2786 = sent_n[214] & N4929;
  assign N4929 = ~fifo_yumi;
  assign N2788 = v_o[214] & ready_i[214];
  assign N2789 = ~N2788;
  assign v_o[215] = fifo_v & N4930;
  assign N4930 = ~sent_r[215];
  assign N2790 = ~reset_i;
  assign N2791 = reset_i;
  assign N2792 = sent_n[215] & N4931;
  assign N4931 = ~fifo_yumi;
  assign N2794 = v_o[215] & ready_i[215];
  assign N2795 = ~N2794;
  assign v_o[216] = fifo_v & N4932;
  assign N4932 = ~sent_r[216];
  assign N2796 = ~reset_i;
  assign N2797 = reset_i;
  assign N2798 = sent_n[216] & N4933;
  assign N4933 = ~fifo_yumi;
  assign N2800 = v_o[216] & ready_i[216];
  assign N2801 = ~N2800;
  assign v_o[217] = fifo_v & N4934;
  assign N4934 = ~sent_r[217];
  assign N2802 = ~reset_i;
  assign N2803 = reset_i;
  assign N2804 = sent_n[217] & N4935;
  assign N4935 = ~fifo_yumi;
  assign N2806 = v_o[217] & ready_i[217];
  assign N2807 = ~N2806;
  assign v_o[218] = fifo_v & N4936;
  assign N4936 = ~sent_r[218];
  assign N2808 = ~reset_i;
  assign N2809 = reset_i;
  assign N2810 = sent_n[218] & N4937;
  assign N4937 = ~fifo_yumi;
  assign N2812 = v_o[218] & ready_i[218];
  assign N2813 = ~N2812;
  assign v_o[219] = fifo_v & N4938;
  assign N4938 = ~sent_r[219];
  assign N2814 = ~reset_i;
  assign N2815 = reset_i;
  assign N2816 = sent_n[219] & N4939;
  assign N4939 = ~fifo_yumi;
  assign N2818 = v_o[219] & ready_i[219];
  assign N2819 = ~N2818;
  assign v_o[220] = fifo_v & N4940;
  assign N4940 = ~sent_r[220];
  assign N2820 = ~reset_i;
  assign N2821 = reset_i;
  assign N2822 = sent_n[220] & N4941;
  assign N4941 = ~fifo_yumi;
  assign N2824 = v_o[220] & ready_i[220];
  assign N2825 = ~N2824;
  assign v_o[221] = fifo_v & N4942;
  assign N4942 = ~sent_r[221];
  assign N2826 = ~reset_i;
  assign N2827 = reset_i;
  assign N2828 = sent_n[221] & N4943;
  assign N4943 = ~fifo_yumi;
  assign N2830 = v_o[221] & ready_i[221];
  assign N2831 = ~N2830;
  assign v_o[222] = fifo_v & N4944;
  assign N4944 = ~sent_r[222];
  assign N2832 = ~reset_i;
  assign N2833 = reset_i;
  assign N2834 = sent_n[222] & N4945;
  assign N4945 = ~fifo_yumi;
  assign N2836 = v_o[222] & ready_i[222];
  assign N2837 = ~N2836;
  assign v_o[223] = fifo_v & N4946;
  assign N4946 = ~sent_r[223];
  assign N2838 = ~reset_i;
  assign N2839 = reset_i;
  assign N2840 = sent_n[223] & N4947;
  assign N4947 = ~fifo_yumi;
  assign N2842 = v_o[223] & ready_i[223];
  assign N2843 = ~N2842;
  assign v_o[224] = fifo_v & N4948;
  assign N4948 = ~sent_r[224];
  assign N2844 = ~reset_i;
  assign N2845 = reset_i;
  assign N2846 = sent_n[224] & N4949;
  assign N4949 = ~fifo_yumi;
  assign N2848 = v_o[224] & ready_i[224];
  assign N2849 = ~N2848;
  assign v_o[225] = fifo_v & N4950;
  assign N4950 = ~sent_r[225];
  assign N2850 = ~reset_i;
  assign N2851 = reset_i;
  assign N2852 = sent_n[225] & N4951;
  assign N4951 = ~fifo_yumi;
  assign N2854 = v_o[225] & ready_i[225];
  assign N2855 = ~N2854;
  assign v_o[226] = fifo_v & N4952;
  assign N4952 = ~sent_r[226];
  assign N2856 = ~reset_i;
  assign N2857 = reset_i;
  assign N2858 = sent_n[226] & N4953;
  assign N4953 = ~fifo_yumi;
  assign N2860 = v_o[226] & ready_i[226];
  assign N2861 = ~N2860;
  assign v_o[227] = fifo_v & N4954;
  assign N4954 = ~sent_r[227];
  assign N2862 = ~reset_i;
  assign N2863 = reset_i;
  assign N2864 = sent_n[227] & N4955;
  assign N4955 = ~fifo_yumi;
  assign N2866 = v_o[227] & ready_i[227];
  assign N2867 = ~N2866;
  assign v_o[228] = fifo_v & N4956;
  assign N4956 = ~sent_r[228];
  assign N2868 = ~reset_i;
  assign N2869 = reset_i;
  assign N2870 = sent_n[228] & N4957;
  assign N4957 = ~fifo_yumi;
  assign N2872 = v_o[228] & ready_i[228];
  assign N2873 = ~N2872;
  assign v_o[229] = fifo_v & N4958;
  assign N4958 = ~sent_r[229];
  assign N2874 = ~reset_i;
  assign N2875 = reset_i;
  assign N2876 = sent_n[229] & N4959;
  assign N4959 = ~fifo_yumi;
  assign N2878 = v_o[229] & ready_i[229];
  assign N2879 = ~N2878;
  assign v_o[230] = fifo_v & N4960;
  assign N4960 = ~sent_r[230];
  assign N2880 = ~reset_i;
  assign N2881 = reset_i;
  assign N2882 = sent_n[230] & N4961;
  assign N4961 = ~fifo_yumi;
  assign N2884 = v_o[230] & ready_i[230];
  assign N2885 = ~N2884;
  assign v_o[231] = fifo_v & N4962;
  assign N4962 = ~sent_r[231];
  assign N2886 = ~reset_i;
  assign N2887 = reset_i;
  assign N2888 = sent_n[231] & N4963;
  assign N4963 = ~fifo_yumi;
  assign N2890 = v_o[231] & ready_i[231];
  assign N2891 = ~N2890;
  assign v_o[232] = fifo_v & N4964;
  assign N4964 = ~sent_r[232];
  assign N2892 = ~reset_i;
  assign N2893 = reset_i;
  assign N2894 = sent_n[232] & N4965;
  assign N4965 = ~fifo_yumi;
  assign N2896 = v_o[232] & ready_i[232];
  assign N2897 = ~N2896;
  assign v_o[233] = fifo_v & N4966;
  assign N4966 = ~sent_r[233];
  assign N2898 = ~reset_i;
  assign N2899 = reset_i;
  assign N2900 = sent_n[233] & N4967;
  assign N4967 = ~fifo_yumi;
  assign N2902 = v_o[233] & ready_i[233];
  assign N2903 = ~N2902;
  assign v_o[234] = fifo_v & N4968;
  assign N4968 = ~sent_r[234];
  assign N2904 = ~reset_i;
  assign N2905 = reset_i;
  assign N2906 = sent_n[234] & N4969;
  assign N4969 = ~fifo_yumi;
  assign N2908 = v_o[234] & ready_i[234];
  assign N2909 = ~N2908;
  assign v_o[235] = fifo_v & N4970;
  assign N4970 = ~sent_r[235];
  assign N2910 = ~reset_i;
  assign N2911 = reset_i;
  assign N2912 = sent_n[235] & N4971;
  assign N4971 = ~fifo_yumi;
  assign N2914 = v_o[235] & ready_i[235];
  assign N2915 = ~N2914;
  assign v_o[236] = fifo_v & N4972;
  assign N4972 = ~sent_r[236];
  assign N2916 = ~reset_i;
  assign N2917 = reset_i;
  assign N2918 = sent_n[236] & N4973;
  assign N4973 = ~fifo_yumi;
  assign N2920 = v_o[236] & ready_i[236];
  assign N2921 = ~N2920;
  assign v_o[237] = fifo_v & N4974;
  assign N4974 = ~sent_r[237];
  assign N2922 = ~reset_i;
  assign N2923 = reset_i;
  assign N2924 = sent_n[237] & N4975;
  assign N4975 = ~fifo_yumi;
  assign N2926 = v_o[237] & ready_i[237];
  assign N2927 = ~N2926;
  assign v_o[238] = fifo_v & N4976;
  assign N4976 = ~sent_r[238];
  assign N2928 = ~reset_i;
  assign N2929 = reset_i;
  assign N2930 = sent_n[238] & N4977;
  assign N4977 = ~fifo_yumi;
  assign N2932 = v_o[238] & ready_i[238];
  assign N2933 = ~N2932;
  assign v_o[239] = fifo_v & N4978;
  assign N4978 = ~sent_r[239];
  assign N2934 = ~reset_i;
  assign N2935 = reset_i;
  assign N2936 = sent_n[239] & N4979;
  assign N4979 = ~fifo_yumi;
  assign N2938 = v_o[239] & ready_i[239];
  assign N2939 = ~N2938;
  assign v_o[240] = fifo_v & N4980;
  assign N4980 = ~sent_r[240];
  assign N2940 = ~reset_i;
  assign N2941 = reset_i;
  assign N2942 = sent_n[240] & N4981;
  assign N4981 = ~fifo_yumi;
  assign N2944 = v_o[240] & ready_i[240];
  assign N2945 = ~N2944;
  assign v_o[241] = fifo_v & N4982;
  assign N4982 = ~sent_r[241];
  assign N2946 = ~reset_i;
  assign N2947 = reset_i;
  assign N2948 = sent_n[241] & N4983;
  assign N4983 = ~fifo_yumi;
  assign N2950 = v_o[241] & ready_i[241];
  assign N2951 = ~N2950;
  assign v_o[242] = fifo_v & N4984;
  assign N4984 = ~sent_r[242];
  assign N2952 = ~reset_i;
  assign N2953 = reset_i;
  assign N2954 = sent_n[242] & N4985;
  assign N4985 = ~fifo_yumi;
  assign N2956 = v_o[242] & ready_i[242];
  assign N2957 = ~N2956;
  assign v_o[243] = fifo_v & N4986;
  assign N4986 = ~sent_r[243];
  assign N2958 = ~reset_i;
  assign N2959 = reset_i;
  assign N2960 = sent_n[243] & N4987;
  assign N4987 = ~fifo_yumi;
  assign N2962 = v_o[243] & ready_i[243];
  assign N2963 = ~N2962;
  assign v_o[244] = fifo_v & N4988;
  assign N4988 = ~sent_r[244];
  assign N2964 = ~reset_i;
  assign N2965 = reset_i;
  assign N2966 = sent_n[244] & N4989;
  assign N4989 = ~fifo_yumi;
  assign N2968 = v_o[244] & ready_i[244];
  assign N2969 = ~N2968;
  assign v_o[245] = fifo_v & N4990;
  assign N4990 = ~sent_r[245];
  assign N2970 = ~reset_i;
  assign N2971 = reset_i;
  assign N2972 = sent_n[245] & N4991;
  assign N4991 = ~fifo_yumi;
  assign N2974 = v_o[245] & ready_i[245];
  assign N2975 = ~N2974;
  assign v_o[246] = fifo_v & N4992;
  assign N4992 = ~sent_r[246];
  assign N2976 = ~reset_i;
  assign N2977 = reset_i;
  assign N2978 = sent_n[246] & N4993;
  assign N4993 = ~fifo_yumi;
  assign N2980 = v_o[246] & ready_i[246];
  assign N2981 = ~N2980;
  assign v_o[247] = fifo_v & N4994;
  assign N4994 = ~sent_r[247];
  assign N2982 = ~reset_i;
  assign N2983 = reset_i;
  assign N2984 = sent_n[247] & N4995;
  assign N4995 = ~fifo_yumi;
  assign N2986 = v_o[247] & ready_i[247];
  assign N2987 = ~N2986;
  assign v_o[248] = fifo_v & N4996;
  assign N4996 = ~sent_r[248];
  assign N2988 = ~reset_i;
  assign N2989 = reset_i;
  assign N2990 = sent_n[248] & N4997;
  assign N4997 = ~fifo_yumi;
  assign N2992 = v_o[248] & ready_i[248];
  assign N2993 = ~N2992;
  assign v_o[249] = fifo_v & N4998;
  assign N4998 = ~sent_r[249];
  assign N2994 = ~reset_i;
  assign N2995 = reset_i;
  assign N2996 = sent_n[249] & N4999;
  assign N4999 = ~fifo_yumi;
  assign N2998 = v_o[249] & ready_i[249];
  assign N2999 = ~N2998;
  assign v_o[250] = fifo_v & N5000;
  assign N5000 = ~sent_r[250];
  assign N3000 = ~reset_i;
  assign N3001 = reset_i;
  assign N3002 = sent_n[250] & N5001;
  assign N5001 = ~fifo_yumi;
  assign N3004 = v_o[250] & ready_i[250];
  assign N3005 = ~N3004;
  assign v_o[251] = fifo_v & N5002;
  assign N5002 = ~sent_r[251];
  assign N3006 = ~reset_i;
  assign N3007 = reset_i;
  assign N3008 = sent_n[251] & N5003;
  assign N5003 = ~fifo_yumi;
  assign N3010 = v_o[251] & ready_i[251];
  assign N3011 = ~N3010;
  assign v_o[252] = fifo_v & N5004;
  assign N5004 = ~sent_r[252];
  assign N3012 = ~reset_i;
  assign N3013 = reset_i;
  assign N3014 = sent_n[252] & N5005;
  assign N5005 = ~fifo_yumi;
  assign N3016 = v_o[252] & ready_i[252];
  assign N3017 = ~N3016;
  assign v_o[253] = fifo_v & N5006;
  assign N5006 = ~sent_r[253];
  assign N3018 = ~reset_i;
  assign N3019 = reset_i;
  assign N3020 = sent_n[253] & N5007;
  assign N5007 = ~fifo_yumi;
  assign N3022 = v_o[253] & ready_i[253];
  assign N3023 = ~N3022;
  assign v_o[254] = fifo_v & N5008;
  assign N5008 = ~sent_r[254];
  assign N3024 = ~reset_i;
  assign N3025 = reset_i;
  assign N3026 = sent_n[254] & N5009;
  assign N5009 = ~fifo_yumi;
  assign N3028 = v_o[254] & ready_i[254];
  assign N3029 = ~N3028;
  assign v_o[255] = fifo_v & N5010;
  assign N5010 = ~sent_r[255];
  assign N3030 = ~reset_i;
  assign N3031 = reset_i;
  assign N3032 = sent_n[255] & N5011;
  assign N5011 = ~fifo_yumi;
  assign N3034 = v_o[255] & ready_i[255];
  assign N3035 = ~N3034;
  assign v_o[256] = fifo_v & N5012;
  assign N5012 = ~sent_r[256];
  assign N3036 = ~reset_i;
  assign N3037 = reset_i;
  assign N3038 = sent_n[256] & N5013;
  assign N5013 = ~fifo_yumi;
  assign N3040 = v_o[256] & ready_i[256];
  assign N3041 = ~N3040;
  assign v_o[257] = fifo_v & N5014;
  assign N5014 = ~sent_r[257];
  assign N3042 = ~reset_i;
  assign N3043 = reset_i;
  assign N3044 = sent_n[257] & N5015;
  assign N5015 = ~fifo_yumi;
  assign N3046 = v_o[257] & ready_i[257];
  assign N3047 = ~N3046;
  assign v_o[258] = fifo_v & N5016;
  assign N5016 = ~sent_r[258];
  assign N3048 = ~reset_i;
  assign N3049 = reset_i;
  assign N3050 = sent_n[258] & N5017;
  assign N5017 = ~fifo_yumi;
  assign N3052 = v_o[258] & ready_i[258];
  assign N3053 = ~N3052;
  assign v_o[259] = fifo_v & N5018;
  assign N5018 = ~sent_r[259];
  assign N3054 = ~reset_i;
  assign N3055 = reset_i;
  assign N3056 = sent_n[259] & N5019;
  assign N5019 = ~fifo_yumi;
  assign N3058 = v_o[259] & ready_i[259];
  assign N3059 = ~N3058;
  assign v_o[260] = fifo_v & N5020;
  assign N5020 = ~sent_r[260];
  assign N3060 = ~reset_i;
  assign N3061 = reset_i;
  assign N3062 = sent_n[260] & N5021;
  assign N5021 = ~fifo_yumi;
  assign N3064 = v_o[260] & ready_i[260];
  assign N3065 = ~N3064;
  assign v_o[261] = fifo_v & N5022;
  assign N5022 = ~sent_r[261];
  assign N3066 = ~reset_i;
  assign N3067 = reset_i;
  assign N3068 = sent_n[261] & N5023;
  assign N5023 = ~fifo_yumi;
  assign N3070 = v_o[261] & ready_i[261];
  assign N3071 = ~N3070;
  assign v_o[262] = fifo_v & N5024;
  assign N5024 = ~sent_r[262];
  assign N3072 = ~reset_i;
  assign N3073 = reset_i;
  assign N3074 = sent_n[262] & N5025;
  assign N5025 = ~fifo_yumi;
  assign N3076 = v_o[262] & ready_i[262];
  assign N3077 = ~N3076;
  assign v_o[263] = fifo_v & N5026;
  assign N5026 = ~sent_r[263];
  assign N3078 = ~reset_i;
  assign N3079 = reset_i;
  assign N3080 = sent_n[263] & N5027;
  assign N5027 = ~fifo_yumi;
  assign N3082 = v_o[263] & ready_i[263];
  assign N3083 = ~N3082;
  assign v_o[264] = fifo_v & N5028;
  assign N5028 = ~sent_r[264];
  assign N3084 = ~reset_i;
  assign N3085 = reset_i;
  assign N3086 = sent_n[264] & N5029;
  assign N5029 = ~fifo_yumi;
  assign N3088 = v_o[264] & ready_i[264];
  assign N3089 = ~N3088;
  assign v_o[265] = fifo_v & N5030;
  assign N5030 = ~sent_r[265];
  assign N3090 = ~reset_i;
  assign N3091 = reset_i;
  assign N3092 = sent_n[265] & N5031;
  assign N5031 = ~fifo_yumi;
  assign N3094 = v_o[265] & ready_i[265];
  assign N3095 = ~N3094;
  assign v_o[266] = fifo_v & N5032;
  assign N5032 = ~sent_r[266];
  assign N3096 = ~reset_i;
  assign N3097 = reset_i;
  assign N3098 = sent_n[266] & N5033;
  assign N5033 = ~fifo_yumi;
  assign N3100 = v_o[266] & ready_i[266];
  assign N3101 = ~N3100;
  assign v_o[267] = fifo_v & N5034;
  assign N5034 = ~sent_r[267];
  assign N3102 = ~reset_i;
  assign N3103 = reset_i;
  assign N3104 = sent_n[267] & N5035;
  assign N5035 = ~fifo_yumi;
  assign N3106 = v_o[267] & ready_i[267];
  assign N3107 = ~N3106;
  assign v_o[268] = fifo_v & N5036;
  assign N5036 = ~sent_r[268];
  assign N3108 = ~reset_i;
  assign N3109 = reset_i;
  assign N3110 = sent_n[268] & N5037;
  assign N5037 = ~fifo_yumi;
  assign N3112 = v_o[268] & ready_i[268];
  assign N3113 = ~N3112;
  assign v_o[269] = fifo_v & N5038;
  assign N5038 = ~sent_r[269];
  assign N3114 = ~reset_i;
  assign N3115 = reset_i;
  assign N3116 = sent_n[269] & N5039;
  assign N5039 = ~fifo_yumi;
  assign N3118 = v_o[269] & ready_i[269];
  assign N3119 = ~N3118;
  assign v_o[270] = fifo_v & N5040;
  assign N5040 = ~sent_r[270];
  assign N3120 = ~reset_i;
  assign N3121 = reset_i;
  assign N3122 = sent_n[270] & N5041;
  assign N5041 = ~fifo_yumi;
  assign N3124 = v_o[270] & ready_i[270];
  assign N3125 = ~N3124;
  assign v_o[271] = fifo_v & N5042;
  assign N5042 = ~sent_r[271];
  assign N3126 = ~reset_i;
  assign N3127 = reset_i;
  assign N3128 = sent_n[271] & N5043;
  assign N5043 = ~fifo_yumi;
  assign N3130 = v_o[271] & ready_i[271];
  assign N3131 = ~N3130;
  assign v_o[272] = fifo_v & N5044;
  assign N5044 = ~sent_r[272];
  assign N3132 = ~reset_i;
  assign N3133 = reset_i;
  assign N3134 = sent_n[272] & N5045;
  assign N5045 = ~fifo_yumi;
  assign N3136 = v_o[272] & ready_i[272];
  assign N3137 = ~N3136;
  assign v_o[273] = fifo_v & N5046;
  assign N5046 = ~sent_r[273];
  assign N3138 = ~reset_i;
  assign N3139 = reset_i;
  assign N3140 = sent_n[273] & N5047;
  assign N5047 = ~fifo_yumi;
  assign N3142 = v_o[273] & ready_i[273];
  assign N3143 = ~N3142;
  assign v_o[274] = fifo_v & N5048;
  assign N5048 = ~sent_r[274];
  assign N3144 = ~reset_i;
  assign N3145 = reset_i;
  assign N3146 = sent_n[274] & N5049;
  assign N5049 = ~fifo_yumi;
  assign N3148 = v_o[274] & ready_i[274];
  assign N3149 = ~N3148;
  assign v_o[275] = fifo_v & N5050;
  assign N5050 = ~sent_r[275];
  assign N3150 = ~reset_i;
  assign N3151 = reset_i;
  assign N3152 = sent_n[275] & N5051;
  assign N5051 = ~fifo_yumi;
  assign N3154 = v_o[275] & ready_i[275];
  assign N3155 = ~N3154;
  assign v_o[276] = fifo_v & N5052;
  assign N5052 = ~sent_r[276];
  assign N3156 = ~reset_i;
  assign N3157 = reset_i;
  assign N3158 = sent_n[276] & N5053;
  assign N5053 = ~fifo_yumi;
  assign N3160 = v_o[276] & ready_i[276];
  assign N3161 = ~N3160;
  assign v_o[277] = fifo_v & N5054;
  assign N5054 = ~sent_r[277];
  assign N3162 = ~reset_i;
  assign N3163 = reset_i;
  assign N3164 = sent_n[277] & N5055;
  assign N5055 = ~fifo_yumi;
  assign N3166 = v_o[277] & ready_i[277];
  assign N3167 = ~N3166;
  assign v_o[278] = fifo_v & N5056;
  assign N5056 = ~sent_r[278];
  assign N3168 = ~reset_i;
  assign N3169 = reset_i;
  assign N3170 = sent_n[278] & N5057;
  assign N5057 = ~fifo_yumi;
  assign N3172 = v_o[278] & ready_i[278];
  assign N3173 = ~N3172;
  assign v_o[279] = fifo_v & N5058;
  assign N5058 = ~sent_r[279];
  assign N3174 = ~reset_i;
  assign N3175 = reset_i;
  assign N3176 = sent_n[279] & N5059;
  assign N5059 = ~fifo_yumi;
  assign N3178 = v_o[279] & ready_i[279];
  assign N3179 = ~N3178;
  assign v_o[280] = fifo_v & N5060;
  assign N5060 = ~sent_r[280];
  assign N3180 = ~reset_i;
  assign N3181 = reset_i;
  assign N3182 = sent_n[280] & N5061;
  assign N5061 = ~fifo_yumi;
  assign N3184 = v_o[280] & ready_i[280];
  assign N3185 = ~N3184;
  assign v_o[281] = fifo_v & N5062;
  assign N5062 = ~sent_r[281];
  assign N3186 = ~reset_i;
  assign N3187 = reset_i;
  assign N3188 = sent_n[281] & N5063;
  assign N5063 = ~fifo_yumi;
  assign N3190 = v_o[281] & ready_i[281];
  assign N3191 = ~N3190;
  assign v_o[282] = fifo_v & N5064;
  assign N5064 = ~sent_r[282];
  assign N3192 = ~reset_i;
  assign N3193 = reset_i;
  assign N3194 = sent_n[282] & N5065;
  assign N5065 = ~fifo_yumi;
  assign N3196 = v_o[282] & ready_i[282];
  assign N3197 = ~N3196;
  assign v_o[283] = fifo_v & N5066;
  assign N5066 = ~sent_r[283];
  assign N3198 = ~reset_i;
  assign N3199 = reset_i;
  assign N3200 = sent_n[283] & N5067;
  assign N5067 = ~fifo_yumi;
  assign N3202 = v_o[283] & ready_i[283];
  assign N3203 = ~N3202;
  assign v_o[284] = fifo_v & N5068;
  assign N5068 = ~sent_r[284];
  assign N3204 = ~reset_i;
  assign N3205 = reset_i;
  assign N3206 = sent_n[284] & N5069;
  assign N5069 = ~fifo_yumi;
  assign N3208 = v_o[284] & ready_i[284];
  assign N3209 = ~N3208;
  assign v_o[285] = fifo_v & N5070;
  assign N5070 = ~sent_r[285];
  assign N3210 = ~reset_i;
  assign N3211 = reset_i;
  assign N3212 = sent_n[285] & N5071;
  assign N5071 = ~fifo_yumi;
  assign N3214 = v_o[285] & ready_i[285];
  assign N3215 = ~N3214;
  assign v_o[286] = fifo_v & N5072;
  assign N5072 = ~sent_r[286];
  assign N3216 = ~reset_i;
  assign N3217 = reset_i;
  assign N3218 = sent_n[286] & N5073;
  assign N5073 = ~fifo_yumi;
  assign N3220 = v_o[286] & ready_i[286];
  assign N3221 = ~N3220;
  assign v_o[287] = fifo_v & N5074;
  assign N5074 = ~sent_r[287];
  assign N3222 = ~reset_i;
  assign N3223 = reset_i;
  assign N3224 = sent_n[287] & N5075;
  assign N5075 = ~fifo_yumi;
  assign N3226 = v_o[287] & ready_i[287];
  assign N3227 = ~N3226;
  assign v_o[288] = fifo_v & N5076;
  assign N5076 = ~sent_r[288];
  assign N3228 = ~reset_i;
  assign N3229 = reset_i;
  assign N3230 = sent_n[288] & N5077;
  assign N5077 = ~fifo_yumi;
  assign N3232 = v_o[288] & ready_i[288];
  assign N3233 = ~N3232;
  assign v_o[289] = fifo_v & N5078;
  assign N5078 = ~sent_r[289];
  assign N3234 = ~reset_i;
  assign N3235 = reset_i;
  assign N3236 = sent_n[289] & N5079;
  assign N5079 = ~fifo_yumi;
  assign N3238 = v_o[289] & ready_i[289];
  assign N3239 = ~N3238;
  assign v_o[290] = fifo_v & N5080;
  assign N5080 = ~sent_r[290];
  assign N3240 = ~reset_i;
  assign N3241 = reset_i;
  assign N3242 = sent_n[290] & N5081;
  assign N5081 = ~fifo_yumi;
  assign N3244 = v_o[290] & ready_i[290];
  assign N3245 = ~N3244;
  assign v_o[291] = fifo_v & N5082;
  assign N5082 = ~sent_r[291];
  assign N3246 = ~reset_i;
  assign N3247 = reset_i;
  assign N3248 = sent_n[291] & N5083;
  assign N5083 = ~fifo_yumi;
  assign N3250 = v_o[291] & ready_i[291];
  assign N3251 = ~N3250;
  assign v_o[292] = fifo_v & N5084;
  assign N5084 = ~sent_r[292];
  assign N3252 = ~reset_i;
  assign N3253 = reset_i;
  assign N3254 = sent_n[292] & N5085;
  assign N5085 = ~fifo_yumi;
  assign N3256 = v_o[292] & ready_i[292];
  assign N3257 = ~N3256;
  assign v_o[293] = fifo_v & N5086;
  assign N5086 = ~sent_r[293];
  assign N3258 = ~reset_i;
  assign N3259 = reset_i;
  assign N3260 = sent_n[293] & N5087;
  assign N5087 = ~fifo_yumi;
  assign N3262 = v_o[293] & ready_i[293];
  assign N3263 = ~N3262;
  assign v_o[294] = fifo_v & N5088;
  assign N5088 = ~sent_r[294];
  assign N3264 = ~reset_i;
  assign N3265 = reset_i;
  assign N3266 = sent_n[294] & N5089;
  assign N5089 = ~fifo_yumi;
  assign N3268 = v_o[294] & ready_i[294];
  assign N3269 = ~N3268;
  assign v_o[295] = fifo_v & N5090;
  assign N5090 = ~sent_r[295];
  assign N3270 = ~reset_i;
  assign N3271 = reset_i;
  assign N3272 = sent_n[295] & N5091;
  assign N5091 = ~fifo_yumi;
  assign N3274 = v_o[295] & ready_i[295];
  assign N3275 = ~N3274;
  assign v_o[296] = fifo_v & N5092;
  assign N5092 = ~sent_r[296];
  assign N3276 = ~reset_i;
  assign N3277 = reset_i;
  assign N3278 = sent_n[296] & N5093;
  assign N5093 = ~fifo_yumi;
  assign N3280 = v_o[296] & ready_i[296];
  assign N3281 = ~N3280;
  assign v_o[297] = fifo_v & N5094;
  assign N5094 = ~sent_r[297];
  assign N3282 = ~reset_i;
  assign N3283 = reset_i;
  assign N3284 = sent_n[297] & N5095;
  assign N5095 = ~fifo_yumi;
  assign N3286 = v_o[297] & ready_i[297];
  assign N3287 = ~N3286;
  assign v_o[298] = fifo_v & N5096;
  assign N5096 = ~sent_r[298];
  assign N3288 = ~reset_i;
  assign N3289 = reset_i;
  assign N3290 = sent_n[298] & N5097;
  assign N5097 = ~fifo_yumi;
  assign N3292 = v_o[298] & ready_i[298];
  assign N3293 = ~N3292;
  assign v_o[299] = fifo_v & N5098;
  assign N5098 = ~sent_r[299];
  assign N3294 = ~reset_i;
  assign N3295 = reset_i;
  assign N3296 = sent_n[299] & N5099;
  assign N5099 = ~fifo_yumi;
  assign N3298 = v_o[299] & ready_i[299];
  assign N3299 = ~N3298;
  assign v_o[300] = fifo_v & N5100;
  assign N5100 = ~sent_r[300];
  assign N3300 = ~reset_i;
  assign N3301 = reset_i;
  assign N3302 = sent_n[300] & N5101;
  assign N5101 = ~fifo_yumi;
  assign N3304 = v_o[300] & ready_i[300];
  assign N3305 = ~N3304;
  assign v_o[301] = fifo_v & N5102;
  assign N5102 = ~sent_r[301];
  assign N3306 = ~reset_i;
  assign N3307 = reset_i;
  assign N3308 = sent_n[301] & N5103;
  assign N5103 = ~fifo_yumi;
  assign N3310 = v_o[301] & ready_i[301];
  assign N3311 = ~N3310;
  assign v_o[302] = fifo_v & N5104;
  assign N5104 = ~sent_r[302];
  assign N3312 = ~reset_i;
  assign N3313 = reset_i;
  assign N3314 = sent_n[302] & N5105;
  assign N5105 = ~fifo_yumi;
  assign N3316 = v_o[302] & ready_i[302];
  assign N3317 = ~N3316;
  assign v_o[303] = fifo_v & N5106;
  assign N5106 = ~sent_r[303];
  assign N3318 = ~reset_i;
  assign N3319 = reset_i;
  assign N3320 = sent_n[303] & N5107;
  assign N5107 = ~fifo_yumi;
  assign N3322 = v_o[303] & ready_i[303];
  assign N3323 = ~N3322;
  assign v_o[304] = fifo_v & N5108;
  assign N5108 = ~sent_r[304];
  assign N3324 = ~reset_i;
  assign N3325 = reset_i;
  assign N3326 = sent_n[304] & N5109;
  assign N5109 = ~fifo_yumi;
  assign N3328 = v_o[304] & ready_i[304];
  assign N3329 = ~N3328;
  assign v_o[305] = fifo_v & N5110;
  assign N5110 = ~sent_r[305];
  assign N3330 = ~reset_i;
  assign N3331 = reset_i;
  assign N3332 = sent_n[305] & N5111;
  assign N5111 = ~fifo_yumi;
  assign N3334 = v_o[305] & ready_i[305];
  assign N3335 = ~N3334;
  assign v_o[306] = fifo_v & N5112;
  assign N5112 = ~sent_r[306];
  assign N3336 = ~reset_i;
  assign N3337 = reset_i;
  assign N3338 = sent_n[306] & N5113;
  assign N5113 = ~fifo_yumi;
  assign N3340 = v_o[306] & ready_i[306];
  assign N3341 = ~N3340;
  assign v_o[307] = fifo_v & N5114;
  assign N5114 = ~sent_r[307];
  assign N3342 = ~reset_i;
  assign N3343 = reset_i;
  assign N3344 = sent_n[307] & N5115;
  assign N5115 = ~fifo_yumi;
  assign N3346 = v_o[307] & ready_i[307];
  assign N3347 = ~N3346;
  assign v_o[308] = fifo_v & N5116;
  assign N5116 = ~sent_r[308];
  assign N3348 = ~reset_i;
  assign N3349 = reset_i;
  assign N3350 = sent_n[308] & N5117;
  assign N5117 = ~fifo_yumi;
  assign N3352 = v_o[308] & ready_i[308];
  assign N3353 = ~N3352;
  assign v_o[309] = fifo_v & N5118;
  assign N5118 = ~sent_r[309];
  assign N3354 = ~reset_i;
  assign N3355 = reset_i;
  assign N3356 = sent_n[309] & N5119;
  assign N5119 = ~fifo_yumi;
  assign N3358 = v_o[309] & ready_i[309];
  assign N3359 = ~N3358;
  assign v_o[310] = fifo_v & N5120;
  assign N5120 = ~sent_r[310];
  assign N3360 = ~reset_i;
  assign N3361 = reset_i;
  assign N3362 = sent_n[310] & N5121;
  assign N5121 = ~fifo_yumi;
  assign N3364 = v_o[310] & ready_i[310];
  assign N3365 = ~N3364;
  assign v_o[311] = fifo_v & N5122;
  assign N5122 = ~sent_r[311];
  assign N3366 = ~reset_i;
  assign N3367 = reset_i;
  assign N3368 = sent_n[311] & N5123;
  assign N5123 = ~fifo_yumi;
  assign N3370 = v_o[311] & ready_i[311];
  assign N3371 = ~N3370;
  assign v_o[312] = fifo_v & N5124;
  assign N5124 = ~sent_r[312];
  assign N3372 = ~reset_i;
  assign N3373 = reset_i;
  assign N3374 = sent_n[312] & N5125;
  assign N5125 = ~fifo_yumi;
  assign N3376 = v_o[312] & ready_i[312];
  assign N3377 = ~N3376;
  assign v_o[313] = fifo_v & N5126;
  assign N5126 = ~sent_r[313];
  assign N3378 = ~reset_i;
  assign N3379 = reset_i;
  assign N3380 = sent_n[313] & N5127;
  assign N5127 = ~fifo_yumi;
  assign N3382 = v_o[313] & ready_i[313];
  assign N3383 = ~N3382;
  assign v_o[314] = fifo_v & N5128;
  assign N5128 = ~sent_r[314];
  assign N3384 = ~reset_i;
  assign N3385 = reset_i;
  assign N3386 = sent_n[314] & N5129;
  assign N5129 = ~fifo_yumi;
  assign N3388 = v_o[314] & ready_i[314];
  assign N3389 = ~N3388;
  assign v_o[315] = fifo_v & N5130;
  assign N5130 = ~sent_r[315];
  assign N3390 = ~reset_i;
  assign N3391 = reset_i;
  assign N3392 = sent_n[315] & N5131;
  assign N5131 = ~fifo_yumi;
  assign N3394 = v_o[315] & ready_i[315];
  assign N3395 = ~N3394;
  assign v_o[316] = fifo_v & N5132;
  assign N5132 = ~sent_r[316];
  assign N3396 = ~reset_i;
  assign N3397 = reset_i;
  assign N3398 = sent_n[316] & N5133;
  assign N5133 = ~fifo_yumi;
  assign N3400 = v_o[316] & ready_i[316];
  assign N3401 = ~N3400;
  assign v_o[317] = fifo_v & N5134;
  assign N5134 = ~sent_r[317];
  assign N3402 = ~reset_i;
  assign N3403 = reset_i;
  assign N3404 = sent_n[317] & N5135;
  assign N5135 = ~fifo_yumi;
  assign N3406 = v_o[317] & ready_i[317];
  assign N3407 = ~N3406;
  assign v_o[318] = fifo_v & N5136;
  assign N5136 = ~sent_r[318];
  assign N3408 = ~reset_i;
  assign N3409 = reset_i;
  assign N3410 = sent_n[318] & N5137;
  assign N5137 = ~fifo_yumi;
  assign N3412 = v_o[318] & ready_i[318];
  assign N3413 = ~N3412;
  assign v_o[319] = fifo_v & N5138;
  assign N5138 = ~sent_r[319];
  assign N3414 = ~reset_i;
  assign N3415 = reset_i;
  assign N3416 = sent_n[319] & N5139;
  assign N5139 = ~fifo_yumi;
  assign N3418 = v_o[319] & ready_i[319];
  assign N3419 = ~N3418;
  assign v_o[320] = fifo_v & N5140;
  assign N5140 = ~sent_r[320];
  assign N3420 = ~reset_i;
  assign N3421 = reset_i;
  assign N3422 = sent_n[320] & N5141;
  assign N5141 = ~fifo_yumi;
  assign N3424 = v_o[320] & ready_i[320];
  assign N3425 = ~N3424;
  assign v_o[321] = fifo_v & N5142;
  assign N5142 = ~sent_r[321];
  assign N3426 = ~reset_i;
  assign N3427 = reset_i;
  assign N3428 = sent_n[321] & N5143;
  assign N5143 = ~fifo_yumi;
  assign N3430 = v_o[321] & ready_i[321];
  assign N3431 = ~N3430;
  assign v_o[322] = fifo_v & N5144;
  assign N5144 = ~sent_r[322];
  assign N3432 = ~reset_i;
  assign N3433 = reset_i;
  assign N3434 = sent_n[322] & N5145;
  assign N5145 = ~fifo_yumi;
  assign N3436 = v_o[322] & ready_i[322];
  assign N3437 = ~N3436;
  assign v_o[323] = fifo_v & N5146;
  assign N5146 = ~sent_r[323];
  assign N3438 = ~reset_i;
  assign N3439 = reset_i;
  assign N3440 = sent_n[323] & N5147;
  assign N5147 = ~fifo_yumi;
  assign N3442 = v_o[323] & ready_i[323];
  assign N3443 = ~N3442;
  assign v_o[324] = fifo_v & N5148;
  assign N5148 = ~sent_r[324];
  assign N3444 = ~reset_i;
  assign N3445 = reset_i;
  assign N3446 = sent_n[324] & N5149;
  assign N5149 = ~fifo_yumi;
  assign N3448 = v_o[324] & ready_i[324];
  assign N3449 = ~N3448;
  assign v_o[325] = fifo_v & N5150;
  assign N5150 = ~sent_r[325];
  assign N3450 = ~reset_i;
  assign N3451 = reset_i;
  assign N3452 = sent_n[325] & N5151;
  assign N5151 = ~fifo_yumi;
  assign N3454 = v_o[325] & ready_i[325];
  assign N3455 = ~N3454;
  assign v_o[326] = fifo_v & N5152;
  assign N5152 = ~sent_r[326];
  assign N3456 = ~reset_i;
  assign N3457 = reset_i;
  assign N3458 = sent_n[326] & N5153;
  assign N5153 = ~fifo_yumi;
  assign N3460 = v_o[326] & ready_i[326];
  assign N3461 = ~N3460;
  assign v_o[327] = fifo_v & N5154;
  assign N5154 = ~sent_r[327];
  assign N3462 = ~reset_i;
  assign N3463 = reset_i;
  assign N3464 = sent_n[327] & N5155;
  assign N5155 = ~fifo_yumi;
  assign N3466 = v_o[327] & ready_i[327];
  assign N3467 = ~N3466;
  assign v_o[328] = fifo_v & N5156;
  assign N5156 = ~sent_r[328];
  assign N3468 = ~reset_i;
  assign N3469 = reset_i;
  assign N3470 = sent_n[328] & N5157;
  assign N5157 = ~fifo_yumi;
  assign N3472 = v_o[328] & ready_i[328];
  assign N3473 = ~N3472;
  assign v_o[329] = fifo_v & N5158;
  assign N5158 = ~sent_r[329];
  assign N3474 = ~reset_i;
  assign N3475 = reset_i;
  assign N3476 = sent_n[329] & N5159;
  assign N5159 = ~fifo_yumi;
  assign N3478 = v_o[329] & ready_i[329];
  assign N3479 = ~N3478;
  assign v_o[330] = fifo_v & N5160;
  assign N5160 = ~sent_r[330];
  assign N3480 = ~reset_i;
  assign N3481 = reset_i;
  assign N3482 = sent_n[330] & N5161;
  assign N5161 = ~fifo_yumi;
  assign N3484 = v_o[330] & ready_i[330];
  assign N3485 = ~N3484;
  assign v_o[331] = fifo_v & N5162;
  assign N5162 = ~sent_r[331];
  assign N3486 = ~reset_i;
  assign N3487 = reset_i;
  assign N3488 = sent_n[331] & N5163;
  assign N5163 = ~fifo_yumi;
  assign N3490 = v_o[331] & ready_i[331];
  assign N3491 = ~N3490;
  assign v_o[332] = fifo_v & N5164;
  assign N5164 = ~sent_r[332];
  assign N3492 = ~reset_i;
  assign N3493 = reset_i;
  assign N3494 = sent_n[332] & N5165;
  assign N5165 = ~fifo_yumi;
  assign N3496 = v_o[332] & ready_i[332];
  assign N3497 = ~N3496;
  assign v_o[333] = fifo_v & N5166;
  assign N5166 = ~sent_r[333];
  assign N3498 = ~reset_i;
  assign N3499 = reset_i;
  assign N3500 = sent_n[333] & N5167;
  assign N5167 = ~fifo_yumi;
  assign N3502 = v_o[333] & ready_i[333];
  assign N3503 = ~N3502;
  assign v_o[334] = fifo_v & N5168;
  assign N5168 = ~sent_r[334];
  assign N3504 = ~reset_i;
  assign N3505 = reset_i;
  assign N3506 = sent_n[334] & N5169;
  assign N5169 = ~fifo_yumi;
  assign N3508 = v_o[334] & ready_i[334];
  assign N3509 = ~N3508;
  assign v_o[335] = fifo_v & N5170;
  assign N5170 = ~sent_r[335];
  assign N3510 = ~reset_i;
  assign N3511 = reset_i;
  assign N3512 = sent_n[335] & N5171;
  assign N5171 = ~fifo_yumi;
  assign N3514 = v_o[335] & ready_i[335];
  assign N3515 = ~N3514;
  assign v_o[336] = fifo_v & N5172;
  assign N5172 = ~sent_r[336];
  assign N3516 = ~reset_i;
  assign N3517 = reset_i;
  assign N3518 = sent_n[336] & N5173;
  assign N5173 = ~fifo_yumi;
  assign N3520 = v_o[336] & ready_i[336];
  assign N3521 = ~N3520;
  assign v_o[337] = fifo_v & N5174;
  assign N5174 = ~sent_r[337];
  assign N3522 = ~reset_i;
  assign N3523 = reset_i;
  assign N3524 = sent_n[337] & N5175;
  assign N5175 = ~fifo_yumi;
  assign N3526 = v_o[337] & ready_i[337];
  assign N3527 = ~N3526;
  assign v_o[338] = fifo_v & N5176;
  assign N5176 = ~sent_r[338];
  assign N3528 = ~reset_i;
  assign N3529 = reset_i;
  assign N3530 = sent_n[338] & N5177;
  assign N5177 = ~fifo_yumi;
  assign N3532 = v_o[338] & ready_i[338];
  assign N3533 = ~N3532;
  assign v_o[339] = fifo_v & N5178;
  assign N5178 = ~sent_r[339];
  assign N3534 = ~reset_i;
  assign N3535 = reset_i;
  assign N3536 = sent_n[339] & N5179;
  assign N5179 = ~fifo_yumi;
  assign N3538 = v_o[339] & ready_i[339];
  assign N3539 = ~N3538;
  assign v_o[340] = fifo_v & N5180;
  assign N5180 = ~sent_r[340];
  assign N3540 = ~reset_i;
  assign N3541 = reset_i;
  assign N3542 = sent_n[340] & N5181;
  assign N5181 = ~fifo_yumi;
  assign N3544 = v_o[340] & ready_i[340];
  assign N3545 = ~N3544;
  assign v_o[341] = fifo_v & N5182;
  assign N5182 = ~sent_r[341];
  assign N3546 = ~reset_i;
  assign N3547 = reset_i;
  assign N3548 = sent_n[341] & N5183;
  assign N5183 = ~fifo_yumi;
  assign N3550 = v_o[341] & ready_i[341];
  assign N3551 = ~N3550;
  assign v_o[342] = fifo_v & N5184;
  assign N5184 = ~sent_r[342];
  assign N3552 = ~reset_i;
  assign N3553 = reset_i;
  assign N3554 = sent_n[342] & N5185;
  assign N5185 = ~fifo_yumi;
  assign N3556 = v_o[342] & ready_i[342];
  assign N3557 = ~N3556;
  assign v_o[343] = fifo_v & N5186;
  assign N5186 = ~sent_r[343];
  assign N3558 = ~reset_i;
  assign N3559 = reset_i;
  assign N3560 = sent_n[343] & N5187;
  assign N5187 = ~fifo_yumi;
  assign N3562 = v_o[343] & ready_i[343];
  assign N3563 = ~N3562;
  assign v_o[344] = fifo_v & N5188;
  assign N5188 = ~sent_r[344];
  assign N3564 = ~reset_i;
  assign N3565 = reset_i;
  assign N3566 = sent_n[344] & N5189;
  assign N5189 = ~fifo_yumi;
  assign N3568 = v_o[344] & ready_i[344];
  assign N3569 = ~N3568;
  assign v_o[345] = fifo_v & N5190;
  assign N5190 = ~sent_r[345];
  assign N3570 = ~reset_i;
  assign N3571 = reset_i;
  assign N3572 = sent_n[345] & N5191;
  assign N5191 = ~fifo_yumi;
  assign N3574 = v_o[345] & ready_i[345];
  assign N3575 = ~N3574;
  assign v_o[346] = fifo_v & N5192;
  assign N5192 = ~sent_r[346];
  assign N3576 = ~reset_i;
  assign N3577 = reset_i;
  assign N3578 = sent_n[346] & N5193;
  assign N5193 = ~fifo_yumi;
  assign N3580 = v_o[346] & ready_i[346];
  assign N3581 = ~N3580;
  assign v_o[347] = fifo_v & N5194;
  assign N5194 = ~sent_r[347];
  assign N3582 = ~reset_i;
  assign N3583 = reset_i;
  assign N3584 = sent_n[347] & N5195;
  assign N5195 = ~fifo_yumi;
  assign N3586 = v_o[347] & ready_i[347];
  assign N3587 = ~N3586;
  assign v_o[348] = fifo_v & N5196;
  assign N5196 = ~sent_r[348];
  assign N3588 = ~reset_i;
  assign N3589 = reset_i;
  assign N3590 = sent_n[348] & N5197;
  assign N5197 = ~fifo_yumi;
  assign N3592 = v_o[348] & ready_i[348];
  assign N3593 = ~N3592;
  assign v_o[349] = fifo_v & N5198;
  assign N5198 = ~sent_r[349];
  assign N3594 = ~reset_i;
  assign N3595 = reset_i;
  assign N3596 = sent_n[349] & N5199;
  assign N5199 = ~fifo_yumi;
  assign N3598 = v_o[349] & ready_i[349];
  assign N3599 = ~N3598;
  assign v_o[350] = fifo_v & N5200;
  assign N5200 = ~sent_r[350];
  assign N3600 = ~reset_i;
  assign N3601 = reset_i;
  assign N3602 = sent_n[350] & N5201;
  assign N5201 = ~fifo_yumi;
  assign N3604 = v_o[350] & ready_i[350];
  assign N3605 = ~N3604;
  assign v_o[351] = fifo_v & N5202;
  assign N5202 = ~sent_r[351];
  assign N3606 = ~reset_i;
  assign N3607 = reset_i;
  assign N3608 = sent_n[351] & N5203;
  assign N5203 = ~fifo_yumi;
  assign N3610 = v_o[351] & ready_i[351];
  assign N3611 = ~N3610;
  assign v_o[352] = fifo_v & N5204;
  assign N5204 = ~sent_r[352];
  assign N3612 = ~reset_i;
  assign N3613 = reset_i;
  assign N3614 = sent_n[352] & N5205;
  assign N5205 = ~fifo_yumi;
  assign N3616 = v_o[352] & ready_i[352];
  assign N3617 = ~N3616;
  assign v_o[353] = fifo_v & N5206;
  assign N5206 = ~sent_r[353];
  assign N3618 = ~reset_i;
  assign N3619 = reset_i;
  assign N3620 = sent_n[353] & N5207;
  assign N5207 = ~fifo_yumi;
  assign N3622 = v_o[353] & ready_i[353];
  assign N3623 = ~N3622;
  assign v_o[354] = fifo_v & N5208;
  assign N5208 = ~sent_r[354];
  assign N3624 = ~reset_i;
  assign N3625 = reset_i;
  assign N3626 = sent_n[354] & N5209;
  assign N5209 = ~fifo_yumi;
  assign N3628 = v_o[354] & ready_i[354];
  assign N3629 = ~N3628;
  assign v_o[355] = fifo_v & N5210;
  assign N5210 = ~sent_r[355];
  assign N3630 = ~reset_i;
  assign N3631 = reset_i;
  assign N3632 = sent_n[355] & N5211;
  assign N5211 = ~fifo_yumi;
  assign N3634 = v_o[355] & ready_i[355];
  assign N3635 = ~N3634;
  assign v_o[356] = fifo_v & N5212;
  assign N5212 = ~sent_r[356];
  assign N3636 = ~reset_i;
  assign N3637 = reset_i;
  assign N3638 = sent_n[356] & N5213;
  assign N5213 = ~fifo_yumi;
  assign N3640 = v_o[356] & ready_i[356];
  assign N3641 = ~N3640;
  assign v_o[357] = fifo_v & N5214;
  assign N5214 = ~sent_r[357];
  assign N3642 = ~reset_i;
  assign N3643 = reset_i;
  assign N3644 = sent_n[357] & N5215;
  assign N5215 = ~fifo_yumi;
  assign N3646 = v_o[357] & ready_i[357];
  assign N3647 = ~N3646;
  assign v_o[358] = fifo_v & N5216;
  assign N5216 = ~sent_r[358];
  assign N3648 = ~reset_i;
  assign N3649 = reset_i;
  assign N3650 = sent_n[358] & N5217;
  assign N5217 = ~fifo_yumi;
  assign N3652 = v_o[358] & ready_i[358];
  assign N3653 = ~N3652;
  assign v_o[359] = fifo_v & N5218;
  assign N5218 = ~sent_r[359];
  assign N3654 = ~reset_i;
  assign N3655 = reset_i;
  assign N3656 = sent_n[359] & N5219;
  assign N5219 = ~fifo_yumi;
  assign N3658 = v_o[359] & ready_i[359];
  assign N3659 = ~N3658;
  assign v_o[360] = fifo_v & N5220;
  assign N5220 = ~sent_r[360];
  assign N3660 = ~reset_i;
  assign N3661 = reset_i;
  assign N3662 = sent_n[360] & N5221;
  assign N5221 = ~fifo_yumi;
  assign N3664 = v_o[360] & ready_i[360];
  assign N3665 = ~N3664;
  assign v_o[361] = fifo_v & N5222;
  assign N5222 = ~sent_r[361];
  assign N3666 = ~reset_i;
  assign N3667 = reset_i;
  assign N3668 = sent_n[361] & N5223;
  assign N5223 = ~fifo_yumi;
  assign N3670 = v_o[361] & ready_i[361];
  assign N3671 = ~N3670;
  assign v_o[362] = fifo_v & N5224;
  assign N5224 = ~sent_r[362];
  assign N3672 = ~reset_i;
  assign N3673 = reset_i;
  assign N3674 = sent_n[362] & N5225;
  assign N5225 = ~fifo_yumi;
  assign N3676 = v_o[362] & ready_i[362];
  assign N3677 = ~N3676;
  assign v_o[363] = fifo_v & N5226;
  assign N5226 = ~sent_r[363];
  assign N3678 = ~reset_i;
  assign N3679 = reset_i;
  assign N3680 = sent_n[363] & N5227;
  assign N5227 = ~fifo_yumi;
  assign N3682 = v_o[363] & ready_i[363];
  assign N3683 = ~N3682;
  assign v_o[364] = fifo_v & N5228;
  assign N5228 = ~sent_r[364];
  assign N3684 = ~reset_i;
  assign N3685 = reset_i;
  assign N3686 = sent_n[364] & N5229;
  assign N5229 = ~fifo_yumi;
  assign N3688 = v_o[364] & ready_i[364];
  assign N3689 = ~N3688;
  assign v_o[365] = fifo_v & N5230;
  assign N5230 = ~sent_r[365];
  assign N3690 = ~reset_i;
  assign N3691 = reset_i;
  assign N3692 = sent_n[365] & N5231;
  assign N5231 = ~fifo_yumi;
  assign N3694 = v_o[365] & ready_i[365];
  assign N3695 = ~N3694;
  assign v_o[366] = fifo_v & N5232;
  assign N5232 = ~sent_r[366];
  assign N3696 = ~reset_i;
  assign N3697 = reset_i;
  assign N3698 = sent_n[366] & N5233;
  assign N5233 = ~fifo_yumi;
  assign N3700 = v_o[366] & ready_i[366];
  assign N3701 = ~N3700;
  assign v_o[367] = fifo_v & N5234;
  assign N5234 = ~sent_r[367];
  assign N3702 = ~reset_i;
  assign N3703 = reset_i;
  assign N3704 = sent_n[367] & N5235;
  assign N5235 = ~fifo_yumi;
  assign N3706 = v_o[367] & ready_i[367];
  assign N3707 = ~N3706;
  assign v_o[368] = fifo_v & N5236;
  assign N5236 = ~sent_r[368];
  assign N3708 = ~reset_i;
  assign N3709 = reset_i;
  assign N3710 = sent_n[368] & N5237;
  assign N5237 = ~fifo_yumi;
  assign N3712 = v_o[368] & ready_i[368];
  assign N3713 = ~N3712;
  assign v_o[369] = fifo_v & N5238;
  assign N5238 = ~sent_r[369];
  assign N3714 = ~reset_i;
  assign N3715 = reset_i;
  assign N3716 = sent_n[369] & N5239;
  assign N5239 = ~fifo_yumi;
  assign N3718 = v_o[369] & ready_i[369];
  assign N3719 = ~N3718;
  assign v_o[370] = fifo_v & N5240;
  assign N5240 = ~sent_r[370];
  assign N3720 = ~reset_i;
  assign N3721 = reset_i;
  assign N3722 = sent_n[370] & N5241;
  assign N5241 = ~fifo_yumi;
  assign N3724 = v_o[370] & ready_i[370];
  assign N3725 = ~N3724;
  assign v_o[371] = fifo_v & N5242;
  assign N5242 = ~sent_r[371];
  assign N3726 = ~reset_i;
  assign N3727 = reset_i;
  assign N3728 = sent_n[371] & N5243;
  assign N5243 = ~fifo_yumi;
  assign N3730 = v_o[371] & ready_i[371];
  assign N3731 = ~N3730;
  assign v_o[372] = fifo_v & N5244;
  assign N5244 = ~sent_r[372];
  assign N3732 = ~reset_i;
  assign N3733 = reset_i;
  assign N3734 = sent_n[372] & N5245;
  assign N5245 = ~fifo_yumi;
  assign N3736 = v_o[372] & ready_i[372];
  assign N3737 = ~N3736;
  assign v_o[373] = fifo_v & N5246;
  assign N5246 = ~sent_r[373];
  assign N3738 = ~reset_i;
  assign N3739 = reset_i;
  assign N3740 = sent_n[373] & N5247;
  assign N5247 = ~fifo_yumi;
  assign N3742 = v_o[373] & ready_i[373];
  assign N3743 = ~N3742;
  assign v_o[374] = fifo_v & N5248;
  assign N5248 = ~sent_r[374];
  assign N3744 = ~reset_i;
  assign N3745 = reset_i;
  assign N3746 = sent_n[374] & N5249;
  assign N5249 = ~fifo_yumi;
  assign N3748 = v_o[374] & ready_i[374];
  assign N3749 = ~N3748;
  assign v_o[375] = fifo_v & N5250;
  assign N5250 = ~sent_r[375];
  assign N3750 = ~reset_i;
  assign N3751 = reset_i;
  assign N3752 = sent_n[375] & N5251;
  assign N5251 = ~fifo_yumi;
  assign N3754 = v_o[375] & ready_i[375];
  assign N3755 = ~N3754;
  assign v_o[376] = fifo_v & N5252;
  assign N5252 = ~sent_r[376];
  assign N3756 = ~reset_i;
  assign N3757 = reset_i;
  assign N3758 = sent_n[376] & N5253;
  assign N5253 = ~fifo_yumi;
  assign N3760 = v_o[376] & ready_i[376];
  assign N3761 = ~N3760;
  assign v_o[377] = fifo_v & N5254;
  assign N5254 = ~sent_r[377];
  assign N3762 = ~reset_i;
  assign N3763 = reset_i;
  assign N3764 = sent_n[377] & N5255;
  assign N5255 = ~fifo_yumi;
  assign N3766 = v_o[377] & ready_i[377];
  assign N3767 = ~N3766;
  assign v_o[378] = fifo_v & N5256;
  assign N5256 = ~sent_r[378];
  assign N3768 = ~reset_i;
  assign N3769 = reset_i;
  assign N3770 = sent_n[378] & N5257;
  assign N5257 = ~fifo_yumi;
  assign N3772 = v_o[378] & ready_i[378];
  assign N3773 = ~N3772;
  assign v_o[379] = fifo_v & N5258;
  assign N5258 = ~sent_r[379];
  assign N3774 = ~reset_i;
  assign N3775 = reset_i;
  assign N3776 = sent_n[379] & N5259;
  assign N5259 = ~fifo_yumi;
  assign N3778 = v_o[379] & ready_i[379];
  assign N3779 = ~N3778;
  assign v_o[380] = fifo_v & N5260;
  assign N5260 = ~sent_r[380];
  assign N3780 = ~reset_i;
  assign N3781 = reset_i;
  assign N3782 = sent_n[380] & N5261;
  assign N5261 = ~fifo_yumi;
  assign N3784 = v_o[380] & ready_i[380];
  assign N3785 = ~N3784;
  assign v_o[381] = fifo_v & N5262;
  assign N5262 = ~sent_r[381];
  assign N3786 = ~reset_i;
  assign N3787 = reset_i;
  assign N3788 = sent_n[381] & N5263;
  assign N5263 = ~fifo_yumi;
  assign N3790 = v_o[381] & ready_i[381];
  assign N3791 = ~N3790;
  assign v_o[382] = fifo_v & N5264;
  assign N5264 = ~sent_r[382];
  assign N3792 = ~reset_i;
  assign N3793 = reset_i;
  assign N3794 = sent_n[382] & N5265;
  assign N5265 = ~fifo_yumi;
  assign N3796 = v_o[382] & ready_i[382];
  assign N3797 = ~N3796;
  assign v_o[383] = fifo_v & N5266;
  assign N5266 = ~sent_r[383];
  assign N3798 = ~reset_i;
  assign N3799 = reset_i;
  assign N3800 = sent_n[383] & N5267;
  assign N5267 = ~fifo_yumi;
  assign N3802 = v_o[383] & ready_i[383];
  assign N3803 = ~N3802;
  assign v_o[384] = fifo_v & N5268;
  assign N5268 = ~sent_r[384];
  assign N3804 = ~reset_i;
  assign N3805 = reset_i;
  assign N3806 = sent_n[384] & N5269;
  assign N5269 = ~fifo_yumi;
  assign N3808 = v_o[384] & ready_i[384];
  assign N3809 = ~N3808;
  assign v_o[385] = fifo_v & N5270;
  assign N5270 = ~sent_r[385];
  assign N3810 = ~reset_i;
  assign N3811 = reset_i;
  assign N3812 = sent_n[385] & N5271;
  assign N5271 = ~fifo_yumi;
  assign N3814 = v_o[385] & ready_i[385];
  assign N3815 = ~N3814;
  assign v_o[386] = fifo_v & N5272;
  assign N5272 = ~sent_r[386];
  assign N3816 = ~reset_i;
  assign N3817 = reset_i;
  assign N3818 = sent_n[386] & N5273;
  assign N5273 = ~fifo_yumi;
  assign N3820 = v_o[386] & ready_i[386];
  assign N3821 = ~N3820;
  assign v_o[387] = fifo_v & N5274;
  assign N5274 = ~sent_r[387];
  assign N3822 = ~reset_i;
  assign N3823 = reset_i;
  assign N3824 = sent_n[387] & N5275;
  assign N5275 = ~fifo_yumi;
  assign N3826 = v_o[387] & ready_i[387];
  assign N3827 = ~N3826;
  assign v_o[388] = fifo_v & N5276;
  assign N5276 = ~sent_r[388];
  assign N3828 = ~reset_i;
  assign N3829 = reset_i;
  assign N3830 = sent_n[388] & N5277;
  assign N5277 = ~fifo_yumi;
  assign N3832 = v_o[388] & ready_i[388];
  assign N3833 = ~N3832;
  assign v_o[389] = fifo_v & N5278;
  assign N5278 = ~sent_r[389];
  assign N3834 = ~reset_i;
  assign N3835 = reset_i;
  assign N3836 = sent_n[389] & N5279;
  assign N5279 = ~fifo_yumi;
  assign N3838 = v_o[389] & ready_i[389];
  assign N3839 = ~N3838;
  assign v_o[390] = fifo_v & N5280;
  assign N5280 = ~sent_r[390];
  assign N3840 = ~reset_i;
  assign N3841 = reset_i;
  assign N3842 = sent_n[390] & N5281;
  assign N5281 = ~fifo_yumi;
  assign N3844 = v_o[390] & ready_i[390];
  assign N3845 = ~N3844;
  assign v_o[391] = fifo_v & N5282;
  assign N5282 = ~sent_r[391];
  assign N3846 = ~reset_i;
  assign N3847 = reset_i;
  assign N3848 = sent_n[391] & N5283;
  assign N5283 = ~fifo_yumi;
  assign N3850 = v_o[391] & ready_i[391];
  assign N3851 = ~N3850;
  assign v_o[392] = fifo_v & N5284;
  assign N5284 = ~sent_r[392];
  assign N3852 = ~reset_i;
  assign N3853 = reset_i;
  assign N3854 = sent_n[392] & N5285;
  assign N5285 = ~fifo_yumi;
  assign N3856 = v_o[392] & ready_i[392];
  assign N3857 = ~N3856;
  assign v_o[393] = fifo_v & N5286;
  assign N5286 = ~sent_r[393];
  assign N3858 = ~reset_i;
  assign N3859 = reset_i;
  assign N3860 = sent_n[393] & N5287;
  assign N5287 = ~fifo_yumi;
  assign N3862 = v_o[393] & ready_i[393];
  assign N3863 = ~N3862;
  assign v_o[394] = fifo_v & N5288;
  assign N5288 = ~sent_r[394];
  assign N3864 = ~reset_i;
  assign N3865 = reset_i;
  assign N3866 = sent_n[394] & N5289;
  assign N5289 = ~fifo_yumi;
  assign N3868 = v_o[394] & ready_i[394];
  assign N3869 = ~N3868;
  assign v_o[395] = fifo_v & N5290;
  assign N5290 = ~sent_r[395];
  assign N3870 = ~reset_i;
  assign N3871 = reset_i;
  assign N3872 = sent_n[395] & N5291;
  assign N5291 = ~fifo_yumi;
  assign N3874 = v_o[395] & ready_i[395];
  assign N3875 = ~N3874;
  assign v_o[396] = fifo_v & N5292;
  assign N5292 = ~sent_r[396];
  assign N3876 = ~reset_i;
  assign N3877 = reset_i;
  assign N3878 = sent_n[396] & N5293;
  assign N5293 = ~fifo_yumi;
  assign N3880 = v_o[396] & ready_i[396];
  assign N3881 = ~N3880;
  assign v_o[397] = fifo_v & N5294;
  assign N5294 = ~sent_r[397];
  assign N3882 = ~reset_i;
  assign N3883 = reset_i;
  assign N3884 = sent_n[397] & N5295;
  assign N5295 = ~fifo_yumi;
  assign N3886 = v_o[397] & ready_i[397];
  assign N3887 = ~N3886;
  assign v_o[398] = fifo_v & N5296;
  assign N5296 = ~sent_r[398];
  assign N3888 = ~reset_i;
  assign N3889 = reset_i;
  assign N3890 = sent_n[398] & N5297;
  assign N5297 = ~fifo_yumi;
  assign N3892 = v_o[398] & ready_i[398];
  assign N3893 = ~N3892;
  assign v_o[399] = fifo_v & N5298;
  assign N5298 = ~sent_r[399];
  assign N3894 = ~reset_i;
  assign N3895 = reset_i;
  assign N3896 = sent_n[399] & N5299;
  assign N5299 = ~fifo_yumi;
  assign N3898 = v_o[399] & ready_i[399];
  assign N3899 = ~N3898;
  assign v_o[400] = fifo_v & N5300;
  assign N5300 = ~sent_r[400];
  assign N3900 = ~reset_i;
  assign N3901 = reset_i;
  assign N3902 = sent_n[400] & N5301;
  assign N5301 = ~fifo_yumi;
  assign N3904 = v_o[400] & ready_i[400];
  assign N3905 = ~N3904;
  assign v_o[401] = fifo_v & N5302;
  assign N5302 = ~sent_r[401];
  assign N3906 = ~reset_i;
  assign N3907 = reset_i;
  assign N3908 = sent_n[401] & N5303;
  assign N5303 = ~fifo_yumi;
  assign N3910 = v_o[401] & ready_i[401];
  assign N3911 = ~N3910;
  assign v_o[402] = fifo_v & N5304;
  assign N5304 = ~sent_r[402];
  assign N3912 = ~reset_i;
  assign N3913 = reset_i;
  assign N3914 = sent_n[402] & N5305;
  assign N5305 = ~fifo_yumi;
  assign N3916 = v_o[402] & ready_i[402];
  assign N3917 = ~N3916;
  assign v_o[403] = fifo_v & N5306;
  assign N5306 = ~sent_r[403];
  assign N3918 = ~reset_i;
  assign N3919 = reset_i;
  assign N3920 = sent_n[403] & N5307;
  assign N5307 = ~fifo_yumi;
  assign N3922 = v_o[403] & ready_i[403];
  assign N3923 = ~N3922;
  assign v_o[404] = fifo_v & N5308;
  assign N5308 = ~sent_r[404];
  assign N3924 = ~reset_i;
  assign N3925 = reset_i;
  assign N3926 = sent_n[404] & N5309;
  assign N5309 = ~fifo_yumi;
  assign N3928 = v_o[404] & ready_i[404];
  assign N3929 = ~N3928;
  assign v_o[405] = fifo_v & N5310;
  assign N5310 = ~sent_r[405];
  assign N3930 = ~reset_i;
  assign N3931 = reset_i;
  assign N3932 = sent_n[405] & N5311;
  assign N5311 = ~fifo_yumi;
  assign N3934 = v_o[405] & ready_i[405];
  assign N3935 = ~N3934;
  assign v_o[406] = fifo_v & N5312;
  assign N5312 = ~sent_r[406];
  assign N3936 = ~reset_i;
  assign N3937 = reset_i;
  assign N3938 = sent_n[406] & N5313;
  assign N5313 = ~fifo_yumi;
  assign N3940 = v_o[406] & ready_i[406];
  assign N3941 = ~N3940;
  assign v_o[407] = fifo_v & N5314;
  assign N5314 = ~sent_r[407];
  assign N3942 = ~reset_i;
  assign N3943 = reset_i;
  assign N3944 = sent_n[407] & N5315;
  assign N5315 = ~fifo_yumi;
  assign N3946 = v_o[407] & ready_i[407];
  assign N3947 = ~N3946;
  assign v_o[408] = fifo_v & N5316;
  assign N5316 = ~sent_r[408];
  assign N3948 = ~reset_i;
  assign N3949 = reset_i;
  assign N3950 = sent_n[408] & N5317;
  assign N5317 = ~fifo_yumi;
  assign N3952 = v_o[408] & ready_i[408];
  assign N3953 = ~N3952;
  assign v_o[409] = fifo_v & N5318;
  assign N5318 = ~sent_r[409];
  assign N3954 = ~reset_i;
  assign N3955 = reset_i;
  assign N3956 = sent_n[409] & N5319;
  assign N5319 = ~fifo_yumi;
  assign N3958 = v_o[409] & ready_i[409];
  assign N3959 = ~N3958;
  assign v_o[410] = fifo_v & N5320;
  assign N5320 = ~sent_r[410];
  assign N3960 = ~reset_i;
  assign N3961 = reset_i;
  assign N3962 = sent_n[410] & N5321;
  assign N5321 = ~fifo_yumi;
  assign N3964 = v_o[410] & ready_i[410];
  assign N3965 = ~N3964;
  assign v_o[411] = fifo_v & N5322;
  assign N5322 = ~sent_r[411];
  assign N3966 = ~reset_i;
  assign N3967 = reset_i;
  assign N3968 = sent_n[411] & N5323;
  assign N5323 = ~fifo_yumi;
  assign N3970 = v_o[411] & ready_i[411];
  assign N3971 = ~N3970;
  assign v_o[412] = fifo_v & N5324;
  assign N5324 = ~sent_r[412];
  assign N3972 = ~reset_i;
  assign N3973 = reset_i;
  assign N3974 = sent_n[412] & N5325;
  assign N5325 = ~fifo_yumi;
  assign N3976 = v_o[412] & ready_i[412];
  assign N3977 = ~N3976;
  assign v_o[413] = fifo_v & N5326;
  assign N5326 = ~sent_r[413];
  assign N3978 = ~reset_i;
  assign N3979 = reset_i;
  assign N3980 = sent_n[413] & N5327;
  assign N5327 = ~fifo_yumi;
  assign N3982 = v_o[413] & ready_i[413];
  assign N3983 = ~N3982;
  assign v_o[414] = fifo_v & N5328;
  assign N5328 = ~sent_r[414];
  assign N3984 = ~reset_i;
  assign N3985 = reset_i;
  assign N3986 = sent_n[414] & N5329;
  assign N5329 = ~fifo_yumi;
  assign N3988 = v_o[414] & ready_i[414];
  assign N3989 = ~N3988;
  assign v_o[415] = fifo_v & N5330;
  assign N5330 = ~sent_r[415];
  assign N3990 = ~reset_i;
  assign N3991 = reset_i;
  assign N3992 = sent_n[415] & N5331;
  assign N5331 = ~fifo_yumi;
  assign N3994 = v_o[415] & ready_i[415];
  assign N3995 = ~N3994;
  assign v_o[416] = fifo_v & N5332;
  assign N5332 = ~sent_r[416];
  assign N3996 = ~reset_i;
  assign N3997 = reset_i;
  assign N3998 = sent_n[416] & N5333;
  assign N5333 = ~fifo_yumi;
  assign N4000 = v_o[416] & ready_i[416];
  assign N4001 = ~N4000;
  assign v_o[417] = fifo_v & N5334;
  assign N5334 = ~sent_r[417];
  assign N4002 = ~reset_i;
  assign N4003 = reset_i;
  assign N4004 = sent_n[417] & N5335;
  assign N5335 = ~fifo_yumi;
  assign N4006 = v_o[417] & ready_i[417];
  assign N4007 = ~N4006;
  assign v_o[418] = fifo_v & N5336;
  assign N5336 = ~sent_r[418];
  assign N4008 = ~reset_i;
  assign N4009 = reset_i;
  assign N4010 = sent_n[418] & N5337;
  assign N5337 = ~fifo_yumi;
  assign N4012 = v_o[418] & ready_i[418];
  assign N4013 = ~N4012;
  assign v_o[419] = fifo_v & N5338;
  assign N5338 = ~sent_r[419];
  assign N4014 = ~reset_i;
  assign N4015 = reset_i;
  assign N4016 = sent_n[419] & N5339;
  assign N5339 = ~fifo_yumi;
  assign N4018 = v_o[419] & ready_i[419];
  assign N4019 = ~N4018;
  assign v_o[420] = fifo_v & N5340;
  assign N5340 = ~sent_r[420];
  assign N4020 = ~reset_i;
  assign N4021 = reset_i;
  assign N4022 = sent_n[420] & N5341;
  assign N5341 = ~fifo_yumi;
  assign N4024 = v_o[420] & ready_i[420];
  assign N4025 = ~N4024;
  assign v_o[421] = fifo_v & N5342;
  assign N5342 = ~sent_r[421];
  assign N4026 = ~reset_i;
  assign N4027 = reset_i;
  assign N4028 = sent_n[421] & N5343;
  assign N5343 = ~fifo_yumi;
  assign N4030 = v_o[421] & ready_i[421];
  assign N4031 = ~N4030;
  assign v_o[422] = fifo_v & N5344;
  assign N5344 = ~sent_r[422];
  assign N4032 = ~reset_i;
  assign N4033 = reset_i;
  assign N4034 = sent_n[422] & N5345;
  assign N5345 = ~fifo_yumi;
  assign N4036 = v_o[422] & ready_i[422];
  assign N4037 = ~N4036;
  assign v_o[423] = fifo_v & N5346;
  assign N5346 = ~sent_r[423];
  assign N4038 = ~reset_i;
  assign N4039 = reset_i;
  assign N4040 = sent_n[423] & N5347;
  assign N5347 = ~fifo_yumi;
  assign N4042 = v_o[423] & ready_i[423];
  assign N4043 = ~N4042;
  assign v_o[424] = fifo_v & N5348;
  assign N5348 = ~sent_r[424];
  assign N4044 = ~reset_i;
  assign N4045 = reset_i;
  assign N4046 = sent_n[424] & N5349;
  assign N5349 = ~fifo_yumi;
  assign N4048 = v_o[424] & ready_i[424];
  assign N4049 = ~N4048;
  assign v_o[425] = fifo_v & N5350;
  assign N5350 = ~sent_r[425];
  assign N4050 = ~reset_i;
  assign N4051 = reset_i;
  assign N4052 = sent_n[425] & N5351;
  assign N5351 = ~fifo_yumi;
  assign N4054 = v_o[425] & ready_i[425];
  assign N4055 = ~N4054;
  assign v_o[426] = fifo_v & N5352;
  assign N5352 = ~sent_r[426];
  assign N4056 = ~reset_i;
  assign N4057 = reset_i;
  assign N4058 = sent_n[426] & N5353;
  assign N5353 = ~fifo_yumi;
  assign N4060 = v_o[426] & ready_i[426];
  assign N4061 = ~N4060;
  assign v_o[427] = fifo_v & N5354;
  assign N5354 = ~sent_r[427];
  assign N4062 = ~reset_i;
  assign N4063 = reset_i;
  assign N4064 = sent_n[427] & N5355;
  assign N5355 = ~fifo_yumi;
  assign N4066 = v_o[427] & ready_i[427];
  assign N4067 = ~N4066;
  assign v_o[428] = fifo_v & N5356;
  assign N5356 = ~sent_r[428];
  assign N4068 = ~reset_i;
  assign N4069 = reset_i;
  assign N4070 = sent_n[428] & N5357;
  assign N5357 = ~fifo_yumi;
  assign N4072 = v_o[428] & ready_i[428];
  assign N4073 = ~N4072;
  assign v_o[429] = fifo_v & N5358;
  assign N5358 = ~sent_r[429];
  assign N4074 = ~reset_i;
  assign N4075 = reset_i;
  assign N4076 = sent_n[429] & N5359;
  assign N5359 = ~fifo_yumi;
  assign N4078 = v_o[429] & ready_i[429];
  assign N4079 = ~N4078;
  assign v_o[430] = fifo_v & N5360;
  assign N5360 = ~sent_r[430];
  assign N4080 = ~reset_i;
  assign N4081 = reset_i;
  assign N4082 = sent_n[430] & N5361;
  assign N5361 = ~fifo_yumi;
  assign N4084 = v_o[430] & ready_i[430];
  assign N4085 = ~N4084;
  assign v_o[431] = fifo_v & N5362;
  assign N5362 = ~sent_r[431];
  assign N4086 = ~reset_i;
  assign N4087 = reset_i;
  assign N4088 = sent_n[431] & N5363;
  assign N5363 = ~fifo_yumi;
  assign N4090 = v_o[431] & ready_i[431];
  assign N4091 = ~N4090;
  assign v_o[432] = fifo_v & N5364;
  assign N5364 = ~sent_r[432];
  assign N4092 = ~reset_i;
  assign N4093 = reset_i;
  assign N4094 = sent_n[432] & N5365;
  assign N5365 = ~fifo_yumi;
  assign N4096 = v_o[432] & ready_i[432];
  assign N4097 = ~N4096;
  assign v_o[433] = fifo_v & N5366;
  assign N5366 = ~sent_r[433];
  assign N4098 = ~reset_i;
  assign N4099 = reset_i;
  assign N4100 = sent_n[433] & N5367;
  assign N5367 = ~fifo_yumi;
  assign N4102 = v_o[433] & ready_i[433];
  assign N4103 = ~N4102;
  assign v_o[434] = fifo_v & N5368;
  assign N5368 = ~sent_r[434];
  assign N4104 = ~reset_i;
  assign N4105 = reset_i;
  assign N4106 = sent_n[434] & N5369;
  assign N5369 = ~fifo_yumi;
  assign N4108 = v_o[434] & ready_i[434];
  assign N4109 = ~N4108;
  assign v_o[435] = fifo_v & N5370;
  assign N5370 = ~sent_r[435];
  assign N4110 = ~reset_i;
  assign N4111 = reset_i;
  assign N4112 = sent_n[435] & N5371;
  assign N5371 = ~fifo_yumi;
  assign N4114 = v_o[435] & ready_i[435];
  assign N4115 = ~N4114;
  assign v_o[436] = fifo_v & N5372;
  assign N5372 = ~sent_r[436];
  assign N4116 = ~reset_i;
  assign N4117 = reset_i;
  assign N4118 = sent_n[436] & N5373;
  assign N5373 = ~fifo_yumi;
  assign N4120 = v_o[436] & ready_i[436];
  assign N4121 = ~N4120;
  assign v_o[437] = fifo_v & N5374;
  assign N5374 = ~sent_r[437];
  assign N4122 = ~reset_i;
  assign N4123 = reset_i;
  assign N4124 = sent_n[437] & N5375;
  assign N5375 = ~fifo_yumi;
  assign N4126 = v_o[437] & ready_i[437];
  assign N4127 = ~N4126;
  assign v_o[438] = fifo_v & N5376;
  assign N5376 = ~sent_r[438];
  assign N4128 = ~reset_i;
  assign N4129 = reset_i;
  assign N4130 = sent_n[438] & N5377;
  assign N5377 = ~fifo_yumi;
  assign N4132 = v_o[438] & ready_i[438];
  assign N4133 = ~N4132;
  assign v_o[439] = fifo_v & N5378;
  assign N5378 = ~sent_r[439];
  assign N4134 = ~reset_i;
  assign N4135 = reset_i;
  assign N4136 = sent_n[439] & N5379;
  assign N5379 = ~fifo_yumi;
  assign N4138 = v_o[439] & ready_i[439];
  assign N4139 = ~N4138;
  assign v_o[440] = fifo_v & N5380;
  assign N5380 = ~sent_r[440];
  assign N4140 = ~reset_i;
  assign N4141 = reset_i;
  assign N4142 = sent_n[440] & N5381;
  assign N5381 = ~fifo_yumi;
  assign N4144 = v_o[440] & ready_i[440];
  assign N4145 = ~N4144;
  assign v_o[441] = fifo_v & N5382;
  assign N5382 = ~sent_r[441];
  assign N4146 = ~reset_i;
  assign N4147 = reset_i;
  assign N4148 = sent_n[441] & N5383;
  assign N5383 = ~fifo_yumi;
  assign N4150 = v_o[441] & ready_i[441];
  assign N4151 = ~N4150;
  assign v_o[442] = fifo_v & N5384;
  assign N5384 = ~sent_r[442];
  assign N4152 = ~reset_i;
  assign N4153 = reset_i;
  assign N4154 = sent_n[442] & N5385;
  assign N5385 = ~fifo_yumi;
  assign N4156 = v_o[442] & ready_i[442];
  assign N4157 = ~N4156;
  assign v_o[443] = fifo_v & N5386;
  assign N5386 = ~sent_r[443];
  assign N4158 = ~reset_i;
  assign N4159 = reset_i;
  assign N4160 = sent_n[443] & N5387;
  assign N5387 = ~fifo_yumi;
  assign N4162 = v_o[443] & ready_i[443];
  assign N4163 = ~N4162;
  assign v_o[444] = fifo_v & N5388;
  assign N5388 = ~sent_r[444];
  assign N4164 = ~reset_i;
  assign N4165 = reset_i;
  assign N4166 = sent_n[444] & N5389;
  assign N5389 = ~fifo_yumi;
  assign N4168 = v_o[444] & ready_i[444];
  assign N4169 = ~N4168;
  assign v_o[445] = fifo_v & N5390;
  assign N5390 = ~sent_r[445];
  assign N4170 = ~reset_i;
  assign N4171 = reset_i;
  assign N4172 = sent_n[445] & N5391;
  assign N5391 = ~fifo_yumi;
  assign N4174 = v_o[445] & ready_i[445];
  assign N4175 = ~N4174;
  assign v_o[446] = fifo_v & N5392;
  assign N5392 = ~sent_r[446];
  assign N4176 = ~reset_i;
  assign N4177 = reset_i;
  assign N4178 = sent_n[446] & N5393;
  assign N5393 = ~fifo_yumi;
  assign N4180 = v_o[446] & ready_i[446];
  assign N4181 = ~N4180;
  assign v_o[447] = fifo_v & N5394;
  assign N5394 = ~sent_r[447];
  assign N4182 = ~reset_i;
  assign N4183 = reset_i;
  assign N4184 = sent_n[447] & N5395;
  assign N5395 = ~fifo_yumi;
  assign N4186 = v_o[447] & ready_i[447];
  assign N4187 = ~N4186;
  assign v_o[448] = fifo_v & N5396;
  assign N5396 = ~sent_r[448];
  assign N4188 = ~reset_i;
  assign N4189 = reset_i;
  assign N4190 = sent_n[448] & N5397;
  assign N5397 = ~fifo_yumi;
  assign N4192 = v_o[448] & ready_i[448];
  assign N4193 = ~N4192;
  assign v_o[449] = fifo_v & N5398;
  assign N5398 = ~sent_r[449];
  assign N4194 = ~reset_i;
  assign N4195 = reset_i;
  assign N4196 = sent_n[449] & N5399;
  assign N5399 = ~fifo_yumi;
  assign N4198 = v_o[449] & ready_i[449];
  assign N4199 = ~N4198;
  assign v_o[450] = fifo_v & N5400;
  assign N5400 = ~sent_r[450];
  assign N4200 = ~reset_i;
  assign N4201 = reset_i;
  assign N4202 = sent_n[450] & N5401;
  assign N5401 = ~fifo_yumi;
  assign N4204 = v_o[450] & ready_i[450];
  assign N4205 = ~N4204;
  assign v_o[451] = fifo_v & N5402;
  assign N5402 = ~sent_r[451];
  assign N4206 = ~reset_i;
  assign N4207 = reset_i;
  assign N4208 = sent_n[451] & N5403;
  assign N5403 = ~fifo_yumi;
  assign N4210 = v_o[451] & ready_i[451];
  assign N4211 = ~N4210;
  assign v_o[452] = fifo_v & N5404;
  assign N5404 = ~sent_r[452];
  assign N4212 = ~reset_i;
  assign N4213 = reset_i;
  assign N4214 = sent_n[452] & N5405;
  assign N5405 = ~fifo_yumi;
  assign N4216 = v_o[452] & ready_i[452];
  assign N4217 = ~N4216;
  assign v_o[453] = fifo_v & N5406;
  assign N5406 = ~sent_r[453];
  assign N4218 = ~reset_i;
  assign N4219 = reset_i;
  assign N4220 = sent_n[453] & N5407;
  assign N5407 = ~fifo_yumi;
  assign N4222 = v_o[453] & ready_i[453];
  assign N4223 = ~N4222;
  assign v_o[454] = fifo_v & N5408;
  assign N5408 = ~sent_r[454];
  assign N4224 = ~reset_i;
  assign N4225 = reset_i;
  assign N4226 = sent_n[454] & N5409;
  assign N5409 = ~fifo_yumi;
  assign N4228 = v_o[454] & ready_i[454];
  assign N4229 = ~N4228;
  assign v_o[455] = fifo_v & N5410;
  assign N5410 = ~sent_r[455];
  assign N4230 = ~reset_i;
  assign N4231 = reset_i;
  assign N4232 = sent_n[455] & N5411;
  assign N5411 = ~fifo_yumi;
  assign N4234 = v_o[455] & ready_i[455];
  assign N4235 = ~N4234;
  assign v_o[456] = fifo_v & N5412;
  assign N5412 = ~sent_r[456];
  assign N4236 = ~reset_i;
  assign N4237 = reset_i;
  assign N4238 = sent_n[456] & N5413;
  assign N5413 = ~fifo_yumi;
  assign N4240 = v_o[456] & ready_i[456];
  assign N4241 = ~N4240;
  assign v_o[457] = fifo_v & N5414;
  assign N5414 = ~sent_r[457];
  assign N4242 = ~reset_i;
  assign N4243 = reset_i;
  assign N4244 = sent_n[457] & N5415;
  assign N5415 = ~fifo_yumi;
  assign N4246 = v_o[457] & ready_i[457];
  assign N4247 = ~N4246;
  assign v_o[458] = fifo_v & N5416;
  assign N5416 = ~sent_r[458];
  assign N4248 = ~reset_i;
  assign N4249 = reset_i;
  assign N4250 = sent_n[458] & N5417;
  assign N5417 = ~fifo_yumi;
  assign N4252 = v_o[458] & ready_i[458];
  assign N4253 = ~N4252;
  assign v_o[459] = fifo_v & N5418;
  assign N5418 = ~sent_r[459];
  assign N4254 = ~reset_i;
  assign N4255 = reset_i;
  assign N4256 = sent_n[459] & N5419;
  assign N5419 = ~fifo_yumi;
  assign N4258 = v_o[459] & ready_i[459];
  assign N4259 = ~N4258;
  assign v_o[460] = fifo_v & N5420;
  assign N5420 = ~sent_r[460];
  assign N4260 = ~reset_i;
  assign N4261 = reset_i;
  assign N4262 = sent_n[460] & N5421;
  assign N5421 = ~fifo_yumi;
  assign N4264 = v_o[460] & ready_i[460];
  assign N4265 = ~N4264;
  assign v_o[461] = fifo_v & N5422;
  assign N5422 = ~sent_r[461];
  assign N4266 = ~reset_i;
  assign N4267 = reset_i;
  assign N4268 = sent_n[461] & N5423;
  assign N5423 = ~fifo_yumi;
  assign N4270 = v_o[461] & ready_i[461];
  assign N4271 = ~N4270;
  assign v_o[462] = fifo_v & N5424;
  assign N5424 = ~sent_r[462];
  assign N4272 = ~reset_i;
  assign N4273 = reset_i;
  assign N4274 = sent_n[462] & N5425;
  assign N5425 = ~fifo_yumi;
  assign N4276 = v_o[462] & ready_i[462];
  assign N4277 = ~N4276;
  assign v_o[463] = fifo_v & N5426;
  assign N5426 = ~sent_r[463];
  assign N4278 = ~reset_i;
  assign N4279 = reset_i;
  assign N4280 = sent_n[463] & N5427;
  assign N5427 = ~fifo_yumi;
  assign N4282 = v_o[463] & ready_i[463];
  assign N4283 = ~N4282;
  assign v_o[464] = fifo_v & N5428;
  assign N5428 = ~sent_r[464];
  assign N4284 = ~reset_i;
  assign N4285 = reset_i;
  assign N4286 = sent_n[464] & N5429;
  assign N5429 = ~fifo_yumi;
  assign N4288 = v_o[464] & ready_i[464];
  assign N4289 = ~N4288;
  assign v_o[465] = fifo_v & N5430;
  assign N5430 = ~sent_r[465];
  assign N4290 = ~reset_i;
  assign N4291 = reset_i;
  assign N4292 = sent_n[465] & N5431;
  assign N5431 = ~fifo_yumi;
  assign N4294 = v_o[465] & ready_i[465];
  assign N4295 = ~N4294;
  assign v_o[466] = fifo_v & N5432;
  assign N5432 = ~sent_r[466];
  assign N4296 = ~reset_i;
  assign N4297 = reset_i;
  assign N4298 = sent_n[466] & N5433;
  assign N5433 = ~fifo_yumi;
  assign N4300 = v_o[466] & ready_i[466];
  assign N4301 = ~N4300;
  assign v_o[467] = fifo_v & N5434;
  assign N5434 = ~sent_r[467];
  assign N4302 = ~reset_i;
  assign N4303 = reset_i;
  assign N4304 = sent_n[467] & N5435;
  assign N5435 = ~fifo_yumi;
  assign N4306 = v_o[467] & ready_i[467];
  assign N4307 = ~N4306;
  assign v_o[468] = fifo_v & N5436;
  assign N5436 = ~sent_r[468];
  assign N4308 = ~reset_i;
  assign N4309 = reset_i;
  assign N4310 = sent_n[468] & N5437;
  assign N5437 = ~fifo_yumi;
  assign N4312 = v_o[468] & ready_i[468];
  assign N4313 = ~N4312;
  assign v_o[469] = fifo_v & N5438;
  assign N5438 = ~sent_r[469];
  assign N4314 = ~reset_i;
  assign N4315 = reset_i;
  assign N4316 = sent_n[469] & N5439;
  assign N5439 = ~fifo_yumi;
  assign N4318 = v_o[469] & ready_i[469];
  assign N4319 = ~N4318;
  assign v_o[470] = fifo_v & N5440;
  assign N5440 = ~sent_r[470];
  assign N4320 = ~reset_i;
  assign N4321 = reset_i;
  assign N4322 = sent_n[470] & N5441;
  assign N5441 = ~fifo_yumi;
  assign N4324 = v_o[470] & ready_i[470];
  assign N4325 = ~N4324;
  assign v_o[471] = fifo_v & N5442;
  assign N5442 = ~sent_r[471];
  assign N4326 = ~reset_i;
  assign N4327 = reset_i;
  assign N4328 = sent_n[471] & N5443;
  assign N5443 = ~fifo_yumi;
  assign N4330 = v_o[471] & ready_i[471];
  assign N4331 = ~N4330;
  assign v_o[472] = fifo_v & N5444;
  assign N5444 = ~sent_r[472];
  assign N4332 = ~reset_i;
  assign N4333 = reset_i;
  assign N4334 = sent_n[472] & N5445;
  assign N5445 = ~fifo_yumi;
  assign N4336 = v_o[472] & ready_i[472];
  assign N4337 = ~N4336;
  assign v_o[473] = fifo_v & N5446;
  assign N5446 = ~sent_r[473];
  assign N4338 = ~reset_i;
  assign N4339 = reset_i;
  assign N4340 = sent_n[473] & N5447;
  assign N5447 = ~fifo_yumi;
  assign N4342 = v_o[473] & ready_i[473];
  assign N4343 = ~N4342;
  assign v_o[474] = fifo_v & N5448;
  assign N5448 = ~sent_r[474];
  assign N4344 = ~reset_i;
  assign N4345 = reset_i;
  assign N4346 = sent_n[474] & N5449;
  assign N5449 = ~fifo_yumi;
  assign N4348 = v_o[474] & ready_i[474];
  assign N4349 = ~N4348;
  assign v_o[475] = fifo_v & N5450;
  assign N5450 = ~sent_r[475];
  assign N4350 = ~reset_i;
  assign N4351 = reset_i;
  assign N4352 = sent_n[475] & N5451;
  assign N5451 = ~fifo_yumi;
  assign N4354 = v_o[475] & ready_i[475];
  assign N4355 = ~N4354;
  assign v_o[476] = fifo_v & N5452;
  assign N5452 = ~sent_r[476];
  assign N4356 = ~reset_i;
  assign N4357 = reset_i;
  assign N4358 = sent_n[476] & N5453;
  assign N5453 = ~fifo_yumi;
  assign N4360 = v_o[476] & ready_i[476];
  assign N4361 = ~N4360;
  assign v_o[477] = fifo_v & N5454;
  assign N5454 = ~sent_r[477];
  assign N4362 = ~reset_i;
  assign N4363 = reset_i;
  assign N4364 = sent_n[477] & N5455;
  assign N5455 = ~fifo_yumi;
  assign N4366 = v_o[477] & ready_i[477];
  assign N4367 = ~N4366;
  assign v_o[478] = fifo_v & N5456;
  assign N5456 = ~sent_r[478];
  assign N4368 = ~reset_i;
  assign N4369 = reset_i;
  assign N4370 = sent_n[478] & N5457;
  assign N5457 = ~fifo_yumi;
  assign N4372 = v_o[478] & ready_i[478];
  assign N4373 = ~N4372;
  assign v_o[479] = fifo_v & N5458;
  assign N5458 = ~sent_r[479];
  assign N4374 = ~reset_i;
  assign N4375 = reset_i;
  assign N4376 = sent_n[479] & N5459;
  assign N5459 = ~fifo_yumi;
  assign N4378 = v_o[479] & ready_i[479];
  assign N4379 = ~N4378;
  assign v_o[480] = fifo_v & N5460;
  assign N5460 = ~sent_r[480];
  assign N4380 = ~reset_i;
  assign N4381 = reset_i;
  assign N4382 = sent_n[480] & N5461;
  assign N5461 = ~fifo_yumi;
  assign N4384 = v_o[480] & ready_i[480];
  assign N4385 = ~N4384;
  assign v_o[481] = fifo_v & N5462;
  assign N5462 = ~sent_r[481];
  assign N4386 = ~reset_i;
  assign N4387 = reset_i;
  assign N4388 = sent_n[481] & N5463;
  assign N5463 = ~fifo_yumi;
  assign N4390 = v_o[481] & ready_i[481];
  assign N4391 = ~N4390;
  assign v_o[482] = fifo_v & N5464;
  assign N5464 = ~sent_r[482];
  assign N4392 = ~reset_i;
  assign N4393 = reset_i;
  assign N4394 = sent_n[482] & N5465;
  assign N5465 = ~fifo_yumi;
  assign N4396 = v_o[482] & ready_i[482];
  assign N4397 = ~N4396;
  assign v_o[483] = fifo_v & N5466;
  assign N5466 = ~sent_r[483];
  assign N4398 = ~reset_i;
  assign N4399 = reset_i;
  assign N4400 = sent_n[483] & N5467;
  assign N5467 = ~fifo_yumi;
  assign N4402 = v_o[483] & ready_i[483];
  assign N4403 = ~N4402;
  assign v_o[484] = fifo_v & N5468;
  assign N5468 = ~sent_r[484];
  assign N4404 = ~reset_i;
  assign N4405 = reset_i;
  assign N4406 = sent_n[484] & N5469;
  assign N5469 = ~fifo_yumi;
  assign N4408 = v_o[484] & ready_i[484];
  assign N4409 = ~N4408;
  assign v_o[485] = fifo_v & N5470;
  assign N5470 = ~sent_r[485];
  assign N4410 = ~reset_i;
  assign N4411 = reset_i;
  assign N4412 = sent_n[485] & N5471;
  assign N5471 = ~fifo_yumi;
  assign N4414 = v_o[485] & ready_i[485];
  assign N4415 = ~N4414;
  assign v_o[486] = fifo_v & N5472;
  assign N5472 = ~sent_r[486];
  assign N4416 = ~reset_i;
  assign N4417 = reset_i;
  assign N4418 = sent_n[486] & N5473;
  assign N5473 = ~fifo_yumi;
  assign N4420 = v_o[486] & ready_i[486];
  assign N4421 = ~N4420;
  assign v_o[487] = fifo_v & N5474;
  assign N5474 = ~sent_r[487];
  assign N4422 = ~reset_i;
  assign N4423 = reset_i;
  assign N4424 = sent_n[487] & N5475;
  assign N5475 = ~fifo_yumi;
  assign N4426 = v_o[487] & ready_i[487];
  assign N4427 = ~N4426;
  assign v_o[488] = fifo_v & N5476;
  assign N5476 = ~sent_r[488];
  assign N4428 = ~reset_i;
  assign N4429 = reset_i;
  assign N4430 = sent_n[488] & N5477;
  assign N5477 = ~fifo_yumi;
  assign N4432 = v_o[488] & ready_i[488];
  assign N4433 = ~N4432;
  assign v_o[489] = fifo_v & N5478;
  assign N5478 = ~sent_r[489];
  assign N4434 = ~reset_i;
  assign N4435 = reset_i;
  assign N4436 = sent_n[489] & N5479;
  assign N5479 = ~fifo_yumi;
  assign N4438 = v_o[489] & ready_i[489];
  assign N4439 = ~N4438;
  assign v_o[490] = fifo_v & N5480;
  assign N5480 = ~sent_r[490];
  assign N4440 = ~reset_i;
  assign N4441 = reset_i;
  assign N4442 = sent_n[490] & N5481;
  assign N5481 = ~fifo_yumi;
  assign N4444 = v_o[490] & ready_i[490];
  assign N4445 = ~N4444;
  assign v_o[491] = fifo_v & N5482;
  assign N5482 = ~sent_r[491];
  assign N4446 = ~reset_i;
  assign N4447 = reset_i;
  assign N4448 = sent_n[491] & N5483;
  assign N5483 = ~fifo_yumi;
  assign N4450 = v_o[491] & ready_i[491];
  assign N4451 = ~N4450;
  assign v_o[492] = fifo_v & N5484;
  assign N5484 = ~sent_r[492];
  assign N4452 = ~reset_i;
  assign N4453 = reset_i;
  assign N4454 = sent_n[492] & N5485;
  assign N5485 = ~fifo_yumi;
  assign N4456 = v_o[492] & ready_i[492];
  assign N4457 = ~N4456;
  assign v_o[493] = fifo_v & N5486;
  assign N5486 = ~sent_r[493];
  assign N4458 = ~reset_i;
  assign N4459 = reset_i;
  assign N4460 = sent_n[493] & N5487;
  assign N5487 = ~fifo_yumi;
  assign N4462 = v_o[493] & ready_i[493];
  assign N4463 = ~N4462;
  assign v_o[494] = fifo_v & N5488;
  assign N5488 = ~sent_r[494];
  assign N4464 = ~reset_i;
  assign N4465 = reset_i;
  assign N4466 = sent_n[494] & N5489;
  assign N5489 = ~fifo_yumi;
  assign N4468 = v_o[494] & ready_i[494];
  assign N4469 = ~N4468;
  assign v_o[495] = fifo_v & N5490;
  assign N5490 = ~sent_r[495];
  assign N4470 = ~reset_i;
  assign N4471 = reset_i;
  assign N4472 = sent_n[495] & N5491;
  assign N5491 = ~fifo_yumi;
  assign N4474 = v_o[495] & ready_i[495];
  assign N4475 = ~N4474;
  assign v_o[496] = fifo_v & N5492;
  assign N5492 = ~sent_r[496];
  assign N4476 = ~reset_i;
  assign N4477 = reset_i;
  assign N4478 = sent_n[496] & N5493;
  assign N5493 = ~fifo_yumi;
  assign N4480 = v_o[496] & ready_i[496];
  assign N4481 = ~N4480;
  assign v_o[497] = fifo_v & N5494;
  assign N5494 = ~sent_r[497];
  assign N4482 = ~reset_i;
  assign N4483 = reset_i;
  assign N4484 = sent_n[497] & N5495;
  assign N5495 = ~fifo_yumi;
  assign N4486 = v_o[497] & ready_i[497];
  assign N4487 = ~N4486;
  assign v_o[498] = fifo_v & N5496;
  assign N5496 = ~sent_r[498];
  assign N4488 = ~reset_i;
  assign N4489 = reset_i;
  assign N4490 = sent_n[498] & N5497;
  assign N5497 = ~fifo_yumi;
  assign N4492 = v_o[498] & ready_i[498];
  assign N4493 = ~N4492;
  assign v_o[499] = fifo_v & N5498;
  assign N5498 = ~sent_r[499];
  assign N4494 = ~reset_i;
  assign N4495 = reset_i;
  assign N4496 = sent_n[499] & N5499;
  assign N5499 = ~fifo_yumi;
  assign N4498 = v_o[499] & ready_i[499];
  assign N4499 = ~N4498;
  assign fifo_yumi = N5997 & sent_n[0];
  assign N5997 = N5996 & sent_n[1];
  assign N5996 = N5995 & sent_n[2];
  assign N5995 = N5994 & sent_n[3];
  assign N5994 = N5993 & sent_n[4];
  assign N5993 = N5992 & sent_n[5];
  assign N5992 = N5991 & sent_n[6];
  assign N5991 = N5990 & sent_n[7];
  assign N5990 = N5989 & sent_n[8];
  assign N5989 = N5988 & sent_n[9];
  assign N5988 = N5987 & sent_n[10];
  assign N5987 = N5986 & sent_n[11];
  assign N5986 = N5985 & sent_n[12];
  assign N5985 = N5984 & sent_n[13];
  assign N5984 = N5983 & sent_n[14];
  assign N5983 = N5982 & sent_n[15];
  assign N5982 = N5981 & sent_n[16];
  assign N5981 = N5980 & sent_n[17];
  assign N5980 = N5979 & sent_n[18];
  assign N5979 = N5978 & sent_n[19];
  assign N5978 = N5977 & sent_n[20];
  assign N5977 = N5976 & sent_n[21];
  assign N5976 = N5975 & sent_n[22];
  assign N5975 = N5974 & sent_n[23];
  assign N5974 = N5973 & sent_n[24];
  assign N5973 = N5972 & sent_n[25];
  assign N5972 = N5971 & sent_n[26];
  assign N5971 = N5970 & sent_n[27];
  assign N5970 = N5969 & sent_n[28];
  assign N5969 = N5968 & sent_n[29];
  assign N5968 = N5967 & sent_n[30];
  assign N5967 = N5966 & sent_n[31];
  assign N5966 = N5965 & sent_n[32];
  assign N5965 = N5964 & sent_n[33];
  assign N5964 = N5963 & sent_n[34];
  assign N5963 = N5962 & sent_n[35];
  assign N5962 = N5961 & sent_n[36];
  assign N5961 = N5960 & sent_n[37];
  assign N5960 = N5959 & sent_n[38];
  assign N5959 = N5958 & sent_n[39];
  assign N5958 = N5957 & sent_n[40];
  assign N5957 = N5956 & sent_n[41];
  assign N5956 = N5955 & sent_n[42];
  assign N5955 = N5954 & sent_n[43];
  assign N5954 = N5953 & sent_n[44];
  assign N5953 = N5952 & sent_n[45];
  assign N5952 = N5951 & sent_n[46];
  assign N5951 = N5950 & sent_n[47];
  assign N5950 = N5949 & sent_n[48];
  assign N5949 = N5948 & sent_n[49];
  assign N5948 = N5947 & sent_n[50];
  assign N5947 = N5946 & sent_n[51];
  assign N5946 = N5945 & sent_n[52];
  assign N5945 = N5944 & sent_n[53];
  assign N5944 = N5943 & sent_n[54];
  assign N5943 = N5942 & sent_n[55];
  assign N5942 = N5941 & sent_n[56];
  assign N5941 = N5940 & sent_n[57];
  assign N5940 = N5939 & sent_n[58];
  assign N5939 = N5938 & sent_n[59];
  assign N5938 = N5937 & sent_n[60];
  assign N5937 = N5936 & sent_n[61];
  assign N5936 = N5935 & sent_n[62];
  assign N5935 = N5934 & sent_n[63];
  assign N5934 = N5933 & sent_n[64];
  assign N5933 = N5932 & sent_n[65];
  assign N5932 = N5931 & sent_n[66];
  assign N5931 = N5930 & sent_n[67];
  assign N5930 = N5929 & sent_n[68];
  assign N5929 = N5928 & sent_n[69];
  assign N5928 = N5927 & sent_n[70];
  assign N5927 = N5926 & sent_n[71];
  assign N5926 = N5925 & sent_n[72];
  assign N5925 = N5924 & sent_n[73];
  assign N5924 = N5923 & sent_n[74];
  assign N5923 = N5922 & sent_n[75];
  assign N5922 = N5921 & sent_n[76];
  assign N5921 = N5920 & sent_n[77];
  assign N5920 = N5919 & sent_n[78];
  assign N5919 = N5918 & sent_n[79];
  assign N5918 = N5917 & sent_n[80];
  assign N5917 = N5916 & sent_n[81];
  assign N5916 = N5915 & sent_n[82];
  assign N5915 = N5914 & sent_n[83];
  assign N5914 = N5913 & sent_n[84];
  assign N5913 = N5912 & sent_n[85];
  assign N5912 = N5911 & sent_n[86];
  assign N5911 = N5910 & sent_n[87];
  assign N5910 = N5909 & sent_n[88];
  assign N5909 = N5908 & sent_n[89];
  assign N5908 = N5907 & sent_n[90];
  assign N5907 = N5906 & sent_n[91];
  assign N5906 = N5905 & sent_n[92];
  assign N5905 = N5904 & sent_n[93];
  assign N5904 = N5903 & sent_n[94];
  assign N5903 = N5902 & sent_n[95];
  assign N5902 = N5901 & sent_n[96];
  assign N5901 = N5900 & sent_n[97];
  assign N5900 = N5899 & sent_n[98];
  assign N5899 = N5898 & sent_n[99];
  assign N5898 = N5897 & sent_n[100];
  assign N5897 = N5896 & sent_n[101];
  assign N5896 = N5895 & sent_n[102];
  assign N5895 = N5894 & sent_n[103];
  assign N5894 = N5893 & sent_n[104];
  assign N5893 = N5892 & sent_n[105];
  assign N5892 = N5891 & sent_n[106];
  assign N5891 = N5890 & sent_n[107];
  assign N5890 = N5889 & sent_n[108];
  assign N5889 = N5888 & sent_n[109];
  assign N5888 = N5887 & sent_n[110];
  assign N5887 = N5886 & sent_n[111];
  assign N5886 = N5885 & sent_n[112];
  assign N5885 = N5884 & sent_n[113];
  assign N5884 = N5883 & sent_n[114];
  assign N5883 = N5882 & sent_n[115];
  assign N5882 = N5881 & sent_n[116];
  assign N5881 = N5880 & sent_n[117];
  assign N5880 = N5879 & sent_n[118];
  assign N5879 = N5878 & sent_n[119];
  assign N5878 = N5877 & sent_n[120];
  assign N5877 = N5876 & sent_n[121];
  assign N5876 = N5875 & sent_n[122];
  assign N5875 = N5874 & sent_n[123];
  assign N5874 = N5873 & sent_n[124];
  assign N5873 = N5872 & sent_n[125];
  assign N5872 = N5871 & sent_n[126];
  assign N5871 = N5870 & sent_n[127];
  assign N5870 = N5869 & sent_n[128];
  assign N5869 = N5868 & sent_n[129];
  assign N5868 = N5867 & sent_n[130];
  assign N5867 = N5866 & sent_n[131];
  assign N5866 = N5865 & sent_n[132];
  assign N5865 = N5864 & sent_n[133];
  assign N5864 = N5863 & sent_n[134];
  assign N5863 = N5862 & sent_n[135];
  assign N5862 = N5861 & sent_n[136];
  assign N5861 = N5860 & sent_n[137];
  assign N5860 = N5859 & sent_n[138];
  assign N5859 = N5858 & sent_n[139];
  assign N5858 = N5857 & sent_n[140];
  assign N5857 = N5856 & sent_n[141];
  assign N5856 = N5855 & sent_n[142];
  assign N5855 = N5854 & sent_n[143];
  assign N5854 = N5853 & sent_n[144];
  assign N5853 = N5852 & sent_n[145];
  assign N5852 = N5851 & sent_n[146];
  assign N5851 = N5850 & sent_n[147];
  assign N5850 = N5849 & sent_n[148];
  assign N5849 = N5848 & sent_n[149];
  assign N5848 = N5847 & sent_n[150];
  assign N5847 = N5846 & sent_n[151];
  assign N5846 = N5845 & sent_n[152];
  assign N5845 = N5844 & sent_n[153];
  assign N5844 = N5843 & sent_n[154];
  assign N5843 = N5842 & sent_n[155];
  assign N5842 = N5841 & sent_n[156];
  assign N5841 = N5840 & sent_n[157];
  assign N5840 = N5839 & sent_n[158];
  assign N5839 = N5838 & sent_n[159];
  assign N5838 = N5837 & sent_n[160];
  assign N5837 = N5836 & sent_n[161];
  assign N5836 = N5835 & sent_n[162];
  assign N5835 = N5834 & sent_n[163];
  assign N5834 = N5833 & sent_n[164];
  assign N5833 = N5832 & sent_n[165];
  assign N5832 = N5831 & sent_n[166];
  assign N5831 = N5830 & sent_n[167];
  assign N5830 = N5829 & sent_n[168];
  assign N5829 = N5828 & sent_n[169];
  assign N5828 = N5827 & sent_n[170];
  assign N5827 = N5826 & sent_n[171];
  assign N5826 = N5825 & sent_n[172];
  assign N5825 = N5824 & sent_n[173];
  assign N5824 = N5823 & sent_n[174];
  assign N5823 = N5822 & sent_n[175];
  assign N5822 = N5821 & sent_n[176];
  assign N5821 = N5820 & sent_n[177];
  assign N5820 = N5819 & sent_n[178];
  assign N5819 = N5818 & sent_n[179];
  assign N5818 = N5817 & sent_n[180];
  assign N5817 = N5816 & sent_n[181];
  assign N5816 = N5815 & sent_n[182];
  assign N5815 = N5814 & sent_n[183];
  assign N5814 = N5813 & sent_n[184];
  assign N5813 = N5812 & sent_n[185];
  assign N5812 = N5811 & sent_n[186];
  assign N5811 = N5810 & sent_n[187];
  assign N5810 = N5809 & sent_n[188];
  assign N5809 = N5808 & sent_n[189];
  assign N5808 = N5807 & sent_n[190];
  assign N5807 = N5806 & sent_n[191];
  assign N5806 = N5805 & sent_n[192];
  assign N5805 = N5804 & sent_n[193];
  assign N5804 = N5803 & sent_n[194];
  assign N5803 = N5802 & sent_n[195];
  assign N5802 = N5801 & sent_n[196];
  assign N5801 = N5800 & sent_n[197];
  assign N5800 = N5799 & sent_n[198];
  assign N5799 = N5798 & sent_n[199];
  assign N5798 = N5797 & sent_n[200];
  assign N5797 = N5796 & sent_n[201];
  assign N5796 = N5795 & sent_n[202];
  assign N5795 = N5794 & sent_n[203];
  assign N5794 = N5793 & sent_n[204];
  assign N5793 = N5792 & sent_n[205];
  assign N5792 = N5791 & sent_n[206];
  assign N5791 = N5790 & sent_n[207];
  assign N5790 = N5789 & sent_n[208];
  assign N5789 = N5788 & sent_n[209];
  assign N5788 = N5787 & sent_n[210];
  assign N5787 = N5786 & sent_n[211];
  assign N5786 = N5785 & sent_n[212];
  assign N5785 = N5784 & sent_n[213];
  assign N5784 = N5783 & sent_n[214];
  assign N5783 = N5782 & sent_n[215];
  assign N5782 = N5781 & sent_n[216];
  assign N5781 = N5780 & sent_n[217];
  assign N5780 = N5779 & sent_n[218];
  assign N5779 = N5778 & sent_n[219];
  assign N5778 = N5777 & sent_n[220];
  assign N5777 = N5776 & sent_n[221];
  assign N5776 = N5775 & sent_n[222];
  assign N5775 = N5774 & sent_n[223];
  assign N5774 = N5773 & sent_n[224];
  assign N5773 = N5772 & sent_n[225];
  assign N5772 = N5771 & sent_n[226];
  assign N5771 = N5770 & sent_n[227];
  assign N5770 = N5769 & sent_n[228];
  assign N5769 = N5768 & sent_n[229];
  assign N5768 = N5767 & sent_n[230];
  assign N5767 = N5766 & sent_n[231];
  assign N5766 = N5765 & sent_n[232];
  assign N5765 = N5764 & sent_n[233];
  assign N5764 = N5763 & sent_n[234];
  assign N5763 = N5762 & sent_n[235];
  assign N5762 = N5761 & sent_n[236];
  assign N5761 = N5760 & sent_n[237];
  assign N5760 = N5759 & sent_n[238];
  assign N5759 = N5758 & sent_n[239];
  assign N5758 = N5757 & sent_n[240];
  assign N5757 = N5756 & sent_n[241];
  assign N5756 = N5755 & sent_n[242];
  assign N5755 = N5754 & sent_n[243];
  assign N5754 = N5753 & sent_n[244];
  assign N5753 = N5752 & sent_n[245];
  assign N5752 = N5751 & sent_n[246];
  assign N5751 = N5750 & sent_n[247];
  assign N5750 = N5749 & sent_n[248];
  assign N5749 = N5748 & sent_n[249];
  assign N5748 = N5747 & sent_n[250];
  assign N5747 = N5746 & sent_n[251];
  assign N5746 = N5745 & sent_n[252];
  assign N5745 = N5744 & sent_n[253];
  assign N5744 = N5743 & sent_n[254];
  assign N5743 = N5742 & sent_n[255];
  assign N5742 = N5741 & sent_n[256];
  assign N5741 = N5740 & sent_n[257];
  assign N5740 = N5739 & sent_n[258];
  assign N5739 = N5738 & sent_n[259];
  assign N5738 = N5737 & sent_n[260];
  assign N5737 = N5736 & sent_n[261];
  assign N5736 = N5735 & sent_n[262];
  assign N5735 = N5734 & sent_n[263];
  assign N5734 = N5733 & sent_n[264];
  assign N5733 = N5732 & sent_n[265];
  assign N5732 = N5731 & sent_n[266];
  assign N5731 = N5730 & sent_n[267];
  assign N5730 = N5729 & sent_n[268];
  assign N5729 = N5728 & sent_n[269];
  assign N5728 = N5727 & sent_n[270];
  assign N5727 = N5726 & sent_n[271];
  assign N5726 = N5725 & sent_n[272];
  assign N5725 = N5724 & sent_n[273];
  assign N5724 = N5723 & sent_n[274];
  assign N5723 = N5722 & sent_n[275];
  assign N5722 = N5721 & sent_n[276];
  assign N5721 = N5720 & sent_n[277];
  assign N5720 = N5719 & sent_n[278];
  assign N5719 = N5718 & sent_n[279];
  assign N5718 = N5717 & sent_n[280];
  assign N5717 = N5716 & sent_n[281];
  assign N5716 = N5715 & sent_n[282];
  assign N5715 = N5714 & sent_n[283];
  assign N5714 = N5713 & sent_n[284];
  assign N5713 = N5712 & sent_n[285];
  assign N5712 = N5711 & sent_n[286];
  assign N5711 = N5710 & sent_n[287];
  assign N5710 = N5709 & sent_n[288];
  assign N5709 = N5708 & sent_n[289];
  assign N5708 = N5707 & sent_n[290];
  assign N5707 = N5706 & sent_n[291];
  assign N5706 = N5705 & sent_n[292];
  assign N5705 = N5704 & sent_n[293];
  assign N5704 = N5703 & sent_n[294];
  assign N5703 = N5702 & sent_n[295];
  assign N5702 = N5701 & sent_n[296];
  assign N5701 = N5700 & sent_n[297];
  assign N5700 = N5699 & sent_n[298];
  assign N5699 = N5698 & sent_n[299];
  assign N5698 = N5697 & sent_n[300];
  assign N5697 = N5696 & sent_n[301];
  assign N5696 = N5695 & sent_n[302];
  assign N5695 = N5694 & sent_n[303];
  assign N5694 = N5693 & sent_n[304];
  assign N5693 = N5692 & sent_n[305];
  assign N5692 = N5691 & sent_n[306];
  assign N5691 = N5690 & sent_n[307];
  assign N5690 = N5689 & sent_n[308];
  assign N5689 = N5688 & sent_n[309];
  assign N5688 = N5687 & sent_n[310];
  assign N5687 = N5686 & sent_n[311];
  assign N5686 = N5685 & sent_n[312];
  assign N5685 = N5684 & sent_n[313];
  assign N5684 = N5683 & sent_n[314];
  assign N5683 = N5682 & sent_n[315];
  assign N5682 = N5681 & sent_n[316];
  assign N5681 = N5680 & sent_n[317];
  assign N5680 = N5679 & sent_n[318];
  assign N5679 = N5678 & sent_n[319];
  assign N5678 = N5677 & sent_n[320];
  assign N5677 = N5676 & sent_n[321];
  assign N5676 = N5675 & sent_n[322];
  assign N5675 = N5674 & sent_n[323];
  assign N5674 = N5673 & sent_n[324];
  assign N5673 = N5672 & sent_n[325];
  assign N5672 = N5671 & sent_n[326];
  assign N5671 = N5670 & sent_n[327];
  assign N5670 = N5669 & sent_n[328];
  assign N5669 = N5668 & sent_n[329];
  assign N5668 = N5667 & sent_n[330];
  assign N5667 = N5666 & sent_n[331];
  assign N5666 = N5665 & sent_n[332];
  assign N5665 = N5664 & sent_n[333];
  assign N5664 = N5663 & sent_n[334];
  assign N5663 = N5662 & sent_n[335];
  assign N5662 = N5661 & sent_n[336];
  assign N5661 = N5660 & sent_n[337];
  assign N5660 = N5659 & sent_n[338];
  assign N5659 = N5658 & sent_n[339];
  assign N5658 = N5657 & sent_n[340];
  assign N5657 = N5656 & sent_n[341];
  assign N5656 = N5655 & sent_n[342];
  assign N5655 = N5654 & sent_n[343];
  assign N5654 = N5653 & sent_n[344];
  assign N5653 = N5652 & sent_n[345];
  assign N5652 = N5651 & sent_n[346];
  assign N5651 = N5650 & sent_n[347];
  assign N5650 = N5649 & sent_n[348];
  assign N5649 = N5648 & sent_n[349];
  assign N5648 = N5647 & sent_n[350];
  assign N5647 = N5646 & sent_n[351];
  assign N5646 = N5645 & sent_n[352];
  assign N5645 = N5644 & sent_n[353];
  assign N5644 = N5643 & sent_n[354];
  assign N5643 = N5642 & sent_n[355];
  assign N5642 = N5641 & sent_n[356];
  assign N5641 = N5640 & sent_n[357];
  assign N5640 = N5639 & sent_n[358];
  assign N5639 = N5638 & sent_n[359];
  assign N5638 = N5637 & sent_n[360];
  assign N5637 = N5636 & sent_n[361];
  assign N5636 = N5635 & sent_n[362];
  assign N5635 = N5634 & sent_n[363];
  assign N5634 = N5633 & sent_n[364];
  assign N5633 = N5632 & sent_n[365];
  assign N5632 = N5631 & sent_n[366];
  assign N5631 = N5630 & sent_n[367];
  assign N5630 = N5629 & sent_n[368];
  assign N5629 = N5628 & sent_n[369];
  assign N5628 = N5627 & sent_n[370];
  assign N5627 = N5626 & sent_n[371];
  assign N5626 = N5625 & sent_n[372];
  assign N5625 = N5624 & sent_n[373];
  assign N5624 = N5623 & sent_n[374];
  assign N5623 = N5622 & sent_n[375];
  assign N5622 = N5621 & sent_n[376];
  assign N5621 = N5620 & sent_n[377];
  assign N5620 = N5619 & sent_n[378];
  assign N5619 = N5618 & sent_n[379];
  assign N5618 = N5617 & sent_n[380];
  assign N5617 = N5616 & sent_n[381];
  assign N5616 = N5615 & sent_n[382];
  assign N5615 = N5614 & sent_n[383];
  assign N5614 = N5613 & sent_n[384];
  assign N5613 = N5612 & sent_n[385];
  assign N5612 = N5611 & sent_n[386];
  assign N5611 = N5610 & sent_n[387];
  assign N5610 = N5609 & sent_n[388];
  assign N5609 = N5608 & sent_n[389];
  assign N5608 = N5607 & sent_n[390];
  assign N5607 = N5606 & sent_n[391];
  assign N5606 = N5605 & sent_n[392];
  assign N5605 = N5604 & sent_n[393];
  assign N5604 = N5603 & sent_n[394];
  assign N5603 = N5602 & sent_n[395];
  assign N5602 = N5601 & sent_n[396];
  assign N5601 = N5600 & sent_n[397];
  assign N5600 = N5599 & sent_n[398];
  assign N5599 = N5598 & sent_n[399];
  assign N5598 = N5597 & sent_n[400];
  assign N5597 = N5596 & sent_n[401];
  assign N5596 = N5595 & sent_n[402];
  assign N5595 = N5594 & sent_n[403];
  assign N5594 = N5593 & sent_n[404];
  assign N5593 = N5592 & sent_n[405];
  assign N5592 = N5591 & sent_n[406];
  assign N5591 = N5590 & sent_n[407];
  assign N5590 = N5589 & sent_n[408];
  assign N5589 = N5588 & sent_n[409];
  assign N5588 = N5587 & sent_n[410];
  assign N5587 = N5586 & sent_n[411];
  assign N5586 = N5585 & sent_n[412];
  assign N5585 = N5584 & sent_n[413];
  assign N5584 = N5583 & sent_n[414];
  assign N5583 = N5582 & sent_n[415];
  assign N5582 = N5581 & sent_n[416];
  assign N5581 = N5580 & sent_n[417];
  assign N5580 = N5579 & sent_n[418];
  assign N5579 = N5578 & sent_n[419];
  assign N5578 = N5577 & sent_n[420];
  assign N5577 = N5576 & sent_n[421];
  assign N5576 = N5575 & sent_n[422];
  assign N5575 = N5574 & sent_n[423];
  assign N5574 = N5573 & sent_n[424];
  assign N5573 = N5572 & sent_n[425];
  assign N5572 = N5571 & sent_n[426];
  assign N5571 = N5570 & sent_n[427];
  assign N5570 = N5569 & sent_n[428];
  assign N5569 = N5568 & sent_n[429];
  assign N5568 = N5567 & sent_n[430];
  assign N5567 = N5566 & sent_n[431];
  assign N5566 = N5565 & sent_n[432];
  assign N5565 = N5564 & sent_n[433];
  assign N5564 = N5563 & sent_n[434];
  assign N5563 = N5562 & sent_n[435];
  assign N5562 = N5561 & sent_n[436];
  assign N5561 = N5560 & sent_n[437];
  assign N5560 = N5559 & sent_n[438];
  assign N5559 = N5558 & sent_n[439];
  assign N5558 = N5557 & sent_n[440];
  assign N5557 = N5556 & sent_n[441];
  assign N5556 = N5555 & sent_n[442];
  assign N5555 = N5554 & sent_n[443];
  assign N5554 = N5553 & sent_n[444];
  assign N5553 = N5552 & sent_n[445];
  assign N5552 = N5551 & sent_n[446];
  assign N5551 = N5550 & sent_n[447];
  assign N5550 = N5549 & sent_n[448];
  assign N5549 = N5548 & sent_n[449];
  assign N5548 = N5547 & sent_n[450];
  assign N5547 = N5546 & sent_n[451];
  assign N5546 = N5545 & sent_n[452];
  assign N5545 = N5544 & sent_n[453];
  assign N5544 = N5543 & sent_n[454];
  assign N5543 = N5542 & sent_n[455];
  assign N5542 = N5541 & sent_n[456];
  assign N5541 = N5540 & sent_n[457];
  assign N5540 = N5539 & sent_n[458];
  assign N5539 = N5538 & sent_n[459];
  assign N5538 = N5537 & sent_n[460];
  assign N5537 = N5536 & sent_n[461];
  assign N5536 = N5535 & sent_n[462];
  assign N5535 = N5534 & sent_n[463];
  assign N5534 = N5533 & sent_n[464];
  assign N5533 = N5532 & sent_n[465];
  assign N5532 = N5531 & sent_n[466];
  assign N5531 = N5530 & sent_n[467];
  assign N5530 = N5529 & sent_n[468];
  assign N5529 = N5528 & sent_n[469];
  assign N5528 = N5527 & sent_n[470];
  assign N5527 = N5526 & sent_n[471];
  assign N5526 = N5525 & sent_n[472];
  assign N5525 = N5524 & sent_n[473];
  assign N5524 = N5523 & sent_n[474];
  assign N5523 = N5522 & sent_n[475];
  assign N5522 = N5521 & sent_n[476];
  assign N5521 = N5520 & sent_n[477];
  assign N5520 = N5519 & sent_n[478];
  assign N5519 = N5518 & sent_n[479];
  assign N5518 = N5517 & sent_n[480];
  assign N5517 = N5516 & sent_n[481];
  assign N5516 = N5515 & sent_n[482];
  assign N5515 = N5514 & sent_n[483];
  assign N5514 = N5513 & sent_n[484];
  assign N5513 = N5512 & sent_n[485];
  assign N5512 = N5511 & sent_n[486];
  assign N5511 = N5510 & sent_n[487];
  assign N5510 = N5509 & sent_n[488];
  assign N5509 = N5508 & sent_n[489];
  assign N5508 = N5507 & sent_n[490];
  assign N5507 = N5506 & sent_n[491];
  assign N5506 = N5505 & sent_n[492];
  assign N5505 = N5504 & sent_n[493];
  assign N5504 = N5503 & sent_n[494];
  assign N5503 = N5502 & sent_n[495];
  assign N5502 = N5501 & sent_n[496];
  assign N5501 = N5500 & sent_n[497];
  assign N5500 = sent_n[499] & sent_n[498];

  always @(posedge clk_i) begin
    if(1'b1) begin
      { sent_r[499:0] } <= { N4497, N4491, N4485, N4479, N4473, N4467, N4461, N4455, N4449, N4443, N4437, N4431, N4425, N4419, N4413, N4407, N4401, N4395, N4389, N4383, N4377, N4371, N4365, N4359, N4353, N4347, N4341, N4335, N4329, N4323, N4317, N4311, N4305, N4299, N4293, N4287, N4281, N4275, N4269, N4263, N4257, N4251, N4245, N4239, N4233, N4227, N4221, N4215, N4209, N4203, N4197, N4191, N4185, N4179, N4173, N4167, N4161, N4155, N4149, N4143, N4137, N4131, N4125, N4119, N4113, N4107, N4101, N4095, N4089, N4083, N4077, N4071, N4065, N4059, N4053, N4047, N4041, N4035, N4029, N4023, N4017, N4011, N4005, N3999, N3993, N3987, N3981, N3975, N3969, N3963, N3957, N3951, N3945, N3939, N3933, N3927, N3921, N3915, N3909, N3903, N3897, N3891, N3885, N3879, N3873, N3867, N3861, N3855, N3849, N3843, N3837, N3831, N3825, N3819, N3813, N3807, N3801, N3795, N3789, N3783, N3777, N3771, N3765, N3759, N3753, N3747, N3741, N3735, N3729, N3723, N3717, N3711, N3705, N3699, N3693, N3687, N3681, N3675, N3669, N3663, N3657, N3651, N3645, N3639, N3633, N3627, N3621, N3615, N3609, N3603, N3597, N3591, N3585, N3579, N3573, N3567, N3561, N3555, N3549, N3543, N3537, N3531, N3525, N3519, N3513, N3507, N3501, N3495, N3489, N3483, N3477, N3471, N3465, N3459, N3453, N3447, N3441, N3435, N3429, N3423, N3417, N3411, N3405, N3399, N3393, N3387, N3381, N3375, N3369, N3363, N3357, N3351, N3345, N3339, N3333, N3327, N3321, N3315, N3309, N3303, N3297, N3291, N3285, N3279, N3273, N3267, N3261, N3255, N3249, N3243, N3237, N3231, N3225, N3219, N3213, N3207, N3201, N3195, N3189, N3183, N3177, N3171, N3165, N3159, N3153, N3147, N3141, N3135, N3129, N3123, N3117, N3111, N3105, N3099, N3093, N3087, N3081, N3075, N3069, N3063, N3057, N3051, N3045, N3039, N3033, N3027, N3021, N3015, N3009, N3003, N2997, N2991, N2985, N2979, N2973, N2967, N2961, N2955, N2949, N2943, N2937, N2931, N2925, N2919, N2913, N2907, N2901, N2895, N2889, N2883, N2877, N2871, N2865, N2859, N2853, N2847, N2841, N2835, N2829, N2823, N2817, N2811, N2805, N2799, N2793, N2787, N2781, N2775, N2769, N2763, N2757, N2751, N2745, N2739, N2733, N2727, N2721, N2715, N2709, N2703, N2697, N2691, N2685, N2679, N2673, N2667, N2661, N2655, N2649, N2643, N2637, N2631, N2625, N2619, N2613, N2607, N2601, N2595, N2589, N2583, N2577, N2571, N2565, N2559, N2553, N2547, N2541, N2535, N2529, N2523, N2517, N2511, N2505, N2499, N2493, N2487, N2481, N2475, N2469, N2463, N2457, N2451, N2445, N2439, N2433, N2427, N2421, N2415, N2409, N2403, N2397, N2391, N2385, N2379, N2373, N2367, N2361, N2355, N2349, N2343, N2337, N2331, N2325, N2319, N2313, N2307, N2301, N2295, N2289, N2283, N2277, N2271, N2265, N2259, N2253, N2247, N2241, N2235, N2229, N2223, N2217, N2211, N2205, N2199, N2193, N2187, N2181, N2175, N2169, N2163, N2157, N2151, N2145, N2139, N2133, N2127, N2121, N2115, N2109, N2103, N2097, N2091, N2085, N2079, N2073, N2067, N2061, N2055, N2049, N2043, N2037, N2031, N2025, N2019, N2013, N2007, N2001, N1995, N1989, N1983, N1977, N1971, N1965, N1959, N1953, N1947, N1941, N1935, N1929, N1923, N1917, N1911, N1905, N1899, N1893, N1887, N1881, N1875, N1869, N1863, N1857, N1851, N1845, N1839, N1833, N1827, N1821, N1815, N1809, N1803, N1797, N1791, N1785, N1779, N1773, N1767, N1761, N1755, N1749, N1743, N1737, N1731, N1725, N1719, N1713, N1707, N1701, N1695, N1689, N1683, N1677, N1671, N1665, N1659, N1653, N1647, N1641, N1635, N1629, N1623, N1617, N1611, N1605, N1599, N1593, N1587, N1581, N1575, N1569, N1563, N1557, N1551, N1545, N1539, N1533, N1527, N1521, N1515, N1509, N1503 };
    end 
  end


endmodule

