

module top
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [127:0] sel_i;
  output [15:0] data_o;
  input clk_i;

  bsg_fifo_shift_datapath
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_fifo_shift_datapath
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [127:0] sel_i;
  output [15:0] data_o;
  input clk_i;
  wire [15:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,r_63__15_,r_63__14_,r_63__13_,r_63__12_,
  r_63__11_,r_63__10_,r_63__9_,r_63__8_,r_63__7_,r_63__6_,r_63__5_,r_63__4_,
  r_63__3_,r_63__2_,r_63__1_,r_63__0_,r_62__15_,r_62__14_,r_62__13_,r_62__12_,r_62__11_,
  r_62__10_,r_62__9_,r_62__8_,r_62__7_,r_62__6_,r_62__5_,r_62__4_,r_62__3_,
  r_62__2_,r_62__1_,r_62__0_,r_61__15_,r_61__14_,r_61__13_,r_61__12_,r_61__11_,r_61__10_,
  r_61__9_,r_61__8_,r_61__7_,r_61__6_,r_61__5_,r_61__4_,r_61__3_,r_61__2_,
  r_61__1_,r_61__0_,r_60__15_,r_60__14_,r_60__13_,r_60__12_,r_60__11_,r_60__10_,r_60__9_,
  r_60__8_,r_60__7_,r_60__6_,r_60__5_,r_60__4_,r_60__3_,r_60__2_,r_60__1_,r_60__0_,
  r_59__15_,r_59__14_,r_59__13_,r_59__12_,r_59__11_,r_59__10_,r_59__9_,r_59__8_,
  r_59__7_,r_59__6_,r_59__5_,r_59__4_,r_59__3_,r_59__2_,r_59__1_,r_59__0_,r_58__15_,
  r_58__14_,r_58__13_,r_58__12_,r_58__11_,r_58__10_,r_58__9_,r_58__8_,r_58__7_,
  r_58__6_,r_58__5_,r_58__4_,r_58__3_,r_58__2_,r_58__1_,r_58__0_,r_57__15_,r_57__14_,
  r_57__13_,r_57__12_,r_57__11_,r_57__10_,r_57__9_,r_57__8_,r_57__7_,r_57__6_,
  r_57__5_,r_57__4_,r_57__3_,r_57__2_,r_57__1_,r_57__0_,r_56__15_,r_56__14_,r_56__13_,
  r_56__12_,r_56__11_,r_56__10_,r_56__9_,r_56__8_,r_56__7_,r_56__6_,r_56__5_,
  r_56__4_,r_56__3_,r_56__2_,r_56__1_,r_56__0_,r_55__15_,r_55__14_,r_55__13_,r_55__12_,
  r_55__11_,r_55__10_,r_55__9_,r_55__8_,r_55__7_,r_55__6_,r_55__5_,r_55__4_,
  r_55__3_,r_55__2_,r_55__1_,r_55__0_,r_54__15_,r_54__14_,r_54__13_,r_54__12_,r_54__11_,
  r_54__10_,r_54__9_,r_54__8_,r_54__7_,r_54__6_,r_54__5_,r_54__4_,r_54__3_,
  r_54__2_,r_54__1_,r_54__0_,r_53__15_,r_53__14_,r_53__13_,r_53__12_,r_53__11_,r_53__10_,
  r_53__9_,r_53__8_,r_53__7_,r_53__6_,r_53__5_,r_53__4_,r_53__3_,r_53__2_,
  r_53__1_,r_53__0_,r_52__15_,r_52__14_,r_52__13_,r_52__12_,r_52__11_,r_52__10_,r_52__9_,
  r_52__8_,r_52__7_,r_52__6_,r_52__5_,r_52__4_,r_52__3_,r_52__2_,r_52__1_,r_52__0_,
  r_51__15_,r_51__14_,r_51__13_,r_51__12_,r_51__11_,r_51__10_,r_51__9_,r_51__8_,
  r_51__7_,r_51__6_,r_51__5_,r_51__4_,r_51__3_,r_51__2_,r_51__1_,r_51__0_,r_50__15_,
  r_50__14_,r_50__13_,r_50__12_,r_50__11_,r_50__10_,r_50__9_,r_50__8_,r_50__7_,
  r_50__6_,r_50__5_,r_50__4_,r_50__3_,r_50__2_,r_50__1_,r_50__0_,r_49__15_,r_49__14_,
  r_49__13_,r_49__12_,r_49__11_,r_49__10_,r_49__9_,r_49__8_,r_49__7_,r_49__6_,
  r_49__5_,r_49__4_,r_49__3_,r_49__2_,r_49__1_,r_49__0_,r_48__15_,r_48__14_,r_48__13_,
  r_48__12_,r_48__11_,r_48__10_,r_48__9_,r_48__8_,r_48__7_,r_48__6_,r_48__5_,
  r_48__4_,r_48__3_,r_48__2_,r_48__1_,r_48__0_,r_47__15_,r_47__14_,r_47__13_,r_47__12_,
  r_47__11_,r_47__10_,r_47__9_,r_47__8_,r_47__7_,r_47__6_,r_47__5_,r_47__4_,
  r_47__3_,r_47__2_,r_47__1_,r_47__0_,r_46__15_,r_46__14_,r_46__13_,r_46__12_,r_46__11_,
  r_46__10_,r_46__9_,r_46__8_,r_46__7_,r_46__6_,r_46__5_,r_46__4_,r_46__3_,
  r_46__2_,r_46__1_,r_46__0_,r_45__15_,r_45__14_,r_45__13_,r_45__12_,r_45__11_,r_45__10_,
  r_45__9_,r_45__8_,r_45__7_,r_45__6_,r_45__5_,r_45__4_,r_45__3_,r_45__2_,
  r_45__1_,r_45__0_,r_44__15_,r_44__14_,r_44__13_,r_44__12_,r_44__11_,r_44__10_,r_44__9_,
  r_44__8_,r_44__7_,r_44__6_,r_44__5_,r_44__4_,r_44__3_,r_44__2_,r_44__1_,r_44__0_,
  r_43__15_,r_43__14_,r_43__13_,r_43__12_,r_43__11_,r_43__10_,r_43__9_,r_43__8_,
  r_43__7_,r_43__6_,r_43__5_,r_43__4_,r_43__3_,r_43__2_,r_43__1_,r_43__0_,r_42__15_,
  r_42__14_,r_42__13_,r_42__12_,r_42__11_,r_42__10_,r_42__9_,r_42__8_,r_42__7_,
  r_42__6_,r_42__5_,r_42__4_,r_42__3_,r_42__2_,r_42__1_,r_42__0_,r_41__15_,r_41__14_,
  r_41__13_,r_41__12_,r_41__11_,r_41__10_,r_41__9_,r_41__8_,r_41__7_,r_41__6_,
  r_41__5_,r_41__4_,r_41__3_,r_41__2_,r_41__1_,r_41__0_,r_40__15_,r_40__14_,r_40__13_,
  r_40__12_,r_40__11_,r_40__10_,r_40__9_,r_40__8_,r_40__7_,r_40__6_,r_40__5_,
  r_40__4_,r_40__3_,r_40__2_,r_40__1_,r_40__0_,r_39__15_,r_39__14_,r_39__13_,r_39__12_,
  r_39__11_,r_39__10_,r_39__9_,r_39__8_,r_39__7_,r_39__6_,r_39__5_,r_39__4_,
  r_39__3_,r_39__2_,r_39__1_,r_39__0_,r_38__15_,r_38__14_,r_38__13_,r_38__12_,r_38__11_,
  r_38__10_,r_38__9_,r_38__8_,r_38__7_,r_38__6_,r_38__5_,r_38__4_,r_38__3_,
  r_38__2_,r_38__1_,r_38__0_,r_37__15_,r_37__14_,r_37__13_,r_37__12_,r_37__11_,r_37__10_,
  r_37__9_,r_37__8_,r_37__7_,r_37__6_,r_37__5_,r_37__4_,r_37__3_,r_37__2_,
  r_37__1_,r_37__0_,r_36__15_,r_36__14_,r_36__13_,r_36__12_,r_36__11_,r_36__10_,r_36__9_,
  r_36__8_,r_36__7_,r_36__6_,r_36__5_,r_36__4_,r_36__3_,r_36__2_,r_36__1_,r_36__0_,
  r_35__15_,r_35__14_,r_35__13_,r_35__12_,r_35__11_,r_35__10_,r_35__9_,r_35__8_,
  r_35__7_,r_35__6_,r_35__5_,r_35__4_,r_35__3_,r_35__2_,r_35__1_,r_35__0_,r_34__15_,
  r_34__14_,r_34__13_,r_34__12_,r_34__11_,r_34__10_,r_34__9_,r_34__8_,r_34__7_,
  r_34__6_,r_34__5_,r_34__4_,r_34__3_,r_34__2_,r_34__1_,r_34__0_,r_33__15_,r_33__14_,
  r_33__13_,r_33__12_,r_33__11_,r_33__10_,r_33__9_,r_33__8_,r_33__7_,r_33__6_,
  r_33__5_,r_33__4_,r_33__3_,r_33__2_,r_33__1_,r_33__0_,N126,N127,N128,N129,N130,
  r_32__15_,r_32__14_,r_32__13_,r_32__12_,r_32__11_,r_32__10_,r_32__9_,r_32__8_,
  r_32__7_,r_32__6_,r_32__5_,r_32__4_,r_32__3_,r_32__2_,r_32__1_,r_32__0_,r_31__15_,
  r_31__14_,r_31__13_,r_31__12_,r_31__11_,r_31__10_,r_31__9_,r_31__8_,r_31__7_,
  r_31__6_,r_31__5_,r_31__4_,r_31__3_,r_31__2_,r_31__1_,r_31__0_,r_30__15_,r_30__14_,
  r_30__13_,r_30__12_,r_30__11_,r_30__10_,r_30__9_,r_30__8_,r_30__7_,r_30__6_,r_30__5_,
  r_30__4_,r_30__3_,r_30__2_,r_30__1_,r_30__0_,r_29__15_,r_29__14_,r_29__13_,
  r_29__12_,r_29__11_,r_29__10_,r_29__9_,r_29__8_,r_29__7_,r_29__6_,r_29__5_,r_29__4_,
  r_29__3_,r_29__2_,r_29__1_,r_29__0_,r_28__15_,r_28__14_,r_28__13_,r_28__12_,
  r_28__11_,r_28__10_,r_28__9_,r_28__8_,r_28__7_,r_28__6_,r_28__5_,r_28__4_,r_28__3_,
  r_28__2_,r_28__1_,r_28__0_,r_27__15_,r_27__14_,r_27__13_,r_27__12_,r_27__11_,
  r_27__10_,r_27__9_,r_27__8_,r_27__7_,r_27__6_,r_27__5_,r_27__4_,r_27__3_,r_27__2_,
  r_27__1_,r_27__0_,r_26__15_,r_26__14_,r_26__13_,r_26__12_,r_26__11_,r_26__10_,
  r_26__9_,r_26__8_,r_26__7_,r_26__6_,r_26__5_,r_26__4_,r_26__3_,r_26__2_,r_26__1_,
  r_26__0_,r_25__15_,r_25__14_,r_25__13_,r_25__12_,r_25__11_,r_25__10_,r_25__9_,
  r_25__8_,r_25__7_,r_25__6_,r_25__5_,r_25__4_,r_25__3_,r_25__2_,r_25__1_,r_25__0_,
  r_24__15_,r_24__14_,r_24__13_,r_24__12_,r_24__11_,r_24__10_,r_24__9_,r_24__8_,
  r_24__7_,r_24__6_,r_24__5_,r_24__4_,r_24__3_,r_24__2_,r_24__1_,r_24__0_,r_23__15_,
  r_23__14_,r_23__13_,r_23__12_,r_23__11_,r_23__10_,r_23__9_,r_23__8_,r_23__7_,
  r_23__6_,r_23__5_,r_23__4_,r_23__3_,r_23__2_,r_23__1_,r_23__0_,r_22__15_,r_22__14_,
  r_22__13_,r_22__12_,r_22__11_,r_22__10_,r_22__9_,r_22__8_,r_22__7_,r_22__6_,r_22__5_,
  r_22__4_,r_22__3_,r_22__2_,r_22__1_,r_22__0_,r_21__15_,r_21__14_,r_21__13_,
  r_21__12_,r_21__11_,r_21__10_,r_21__9_,r_21__8_,r_21__7_,r_21__6_,r_21__5_,r_21__4_,
  r_21__3_,r_21__2_,r_21__1_,r_21__0_,r_20__15_,r_20__14_,r_20__13_,r_20__12_,
  r_20__11_,r_20__10_,r_20__9_,r_20__8_,r_20__7_,r_20__6_,r_20__5_,r_20__4_,r_20__3_,
  r_20__2_,r_20__1_,r_20__0_,r_19__15_,r_19__14_,r_19__13_,r_19__12_,r_19__11_,
  r_19__10_,r_19__9_,r_19__8_,r_19__7_,r_19__6_,r_19__5_,r_19__4_,r_19__3_,r_19__2_,
  r_19__1_,r_19__0_,r_18__15_,r_18__14_,r_18__13_,r_18__12_,r_18__11_,r_18__10_,
  r_18__9_,r_18__8_,r_18__7_,r_18__6_,r_18__5_,r_18__4_,r_18__3_,r_18__2_,r_18__1_,
  r_18__0_,r_17__15_,r_17__14_,r_17__13_,r_17__12_,r_17__11_,r_17__10_,r_17__9_,
  r_17__8_,r_17__7_,r_17__6_,r_17__5_,r_17__4_,r_17__3_,r_17__2_,r_17__1_,r_17__0_,
  r_16__15_,r_16__14_,r_16__13_,r_16__12_,r_16__11_,r_16__10_,r_16__9_,r_16__8_,
  r_16__7_,r_16__6_,r_16__5_,r_16__4_,r_16__3_,r_16__2_,r_16__1_,r_16__0_,r_15__15_,
  r_15__14_,r_15__13_,r_15__12_,r_15__11_,r_15__10_,r_15__9_,r_15__8_,r_15__7_,
  r_15__6_,r_15__5_,r_15__4_,r_15__3_,r_15__2_,r_15__1_,r_15__0_,r_14__15_,r_14__14_,
  r_14__13_,r_14__12_,r_14__11_,r_14__10_,r_14__9_,r_14__8_,r_14__7_,r_14__6_,r_14__5_,
  r_14__4_,r_14__3_,r_14__2_,r_14__1_,r_14__0_,r_13__15_,r_13__14_,r_13__13_,
  r_13__12_,r_13__11_,r_13__10_,r_13__9_,r_13__8_,r_13__7_,r_13__6_,r_13__5_,r_13__4_,
  r_13__3_,r_13__2_,r_13__1_,r_13__0_,r_12__15_,r_12__14_,r_12__13_,r_12__12_,
  r_12__11_,r_12__10_,r_12__9_,r_12__8_,r_12__7_,r_12__6_,r_12__5_,r_12__4_,r_12__3_,
  r_12__2_,r_12__1_,r_12__0_,r_11__15_,r_11__14_,r_11__13_,r_11__12_,r_11__11_,
  r_11__10_,r_11__9_,r_11__8_,r_11__7_,r_11__6_,r_11__5_,r_11__4_,r_11__3_,r_11__2_,
  r_11__1_,r_11__0_,r_10__15_,r_10__14_,r_10__13_,r_10__12_,r_10__11_,r_10__10_,
  r_10__9_,r_10__8_,r_10__7_,r_10__6_,r_10__5_,r_10__4_,r_10__3_,r_10__2_,r_10__1_,
  r_10__0_,r_9__15_,r_9__14_,r_9__13_,r_9__12_,r_9__11_,r_9__10_,r_9__9_,r_9__8_,
  r_9__7_,r_9__6_,r_9__5_,r_9__4_,r_9__3_,r_9__2_,r_9__1_,r_9__0_,r_8__15_,r_8__14_,
  r_8__13_,r_8__12_,r_8__11_,r_8__10_,r_8__9_,r_8__8_,r_8__7_,r_8__6_,r_8__5_,
  r_8__4_,r_8__3_,r_8__2_,r_8__1_,r_8__0_,r_7__15_,r_7__14_,r_7__13_,r_7__12_,r_7__11_,
  r_7__10_,r_7__9_,r_7__8_,r_7__7_,r_7__6_,r_7__5_,r_7__4_,r_7__3_,r_7__2_,r_7__1_,
  r_7__0_,r_6__15_,r_6__14_,r_6__13_,r_6__12_,r_6__11_,r_6__10_,r_6__9_,r_6__8_,
  r_6__7_,r_6__6_,r_6__5_,r_6__4_,r_6__3_,r_6__2_,r_6__1_,r_6__0_,r_5__15_,r_5__14_,
  r_5__13_,r_5__12_,r_5__11_,r_5__10_,r_5__9_,r_5__8_,r_5__7_,r_5__6_,r_5__5_,
  r_5__4_,r_5__3_,r_5__2_,r_5__1_,r_5__0_,r_4__15_,r_4__14_,r_4__13_,r_4__12_,r_4__11_,
  r_4__10_,r_4__9_,r_4__8_,r_4__7_,r_4__6_,r_4__5_,r_4__4_,r_4__3_,r_4__2_,
  r_4__1_,r_4__0_,r_3__15_,r_3__14_,r_3__13_,r_3__12_,r_3__11_,r_3__10_,r_3__9_,r_3__8_,
  r_3__7_,r_3__6_,r_3__5_,r_3__4_,r_3__3_,r_3__2_,r_3__1_,r_3__0_,r_2__15_,
  r_2__14_,r_2__13_,r_2__12_,r_2__11_,r_2__10_,r_2__9_,r_2__8_,r_2__7_,r_2__6_,r_2__5_,
  r_2__4_,r_2__3_,r_2__2_,r_2__1_,r_2__0_,r_1__15_,r_1__14_,r_1__13_,r_1__12_,
  r_1__11_,r_1__10_,r_1__9_,r_1__8_,r_1__7_,r_1__6_,r_1__5_,r_1__4_,r_1__3_,r_1__2_,
  r_1__1_,r_1__0_,r_n_0__15_,r_n_0__14_,r_n_0__13_,r_n_0__12_,r_n_0__11_,r_n_0__10_,
  r_n_0__9_,r_n_0__8_,r_n_0__7_,r_n_0__6_,r_n_0__5_,r_n_0__4_,r_n_0__3_,r_n_0__2_,
  r_n_0__1_,r_n_0__0_,r_n_32__15_,r_n_32__14_,r_n_32__13_,r_n_32__12_,r_n_32__11_,
  r_n_32__10_,r_n_32__9_,r_n_32__8_,r_n_32__7_,r_n_32__6_,r_n_32__5_,r_n_32__4_,
  r_n_32__3_,r_n_32__2_,r_n_32__1_,r_n_32__0_,r_n_31__15_,r_n_31__14_,r_n_31__13_,
  r_n_31__12_,r_n_31__11_,r_n_31__10_,r_n_31__9_,r_n_31__8_,r_n_31__7_,r_n_31__6_,
  r_n_31__5_,r_n_31__4_,r_n_31__3_,r_n_31__2_,r_n_31__1_,r_n_31__0_,r_n_30__15_,
  r_n_30__14_,r_n_30__13_,r_n_30__12_,r_n_30__11_,r_n_30__10_,r_n_30__9_,r_n_30__8_,
  r_n_30__7_,r_n_30__6_,r_n_30__5_,r_n_30__4_,r_n_30__3_,r_n_30__2_,r_n_30__1_,
  r_n_30__0_,r_n_29__15_,r_n_29__14_,r_n_29__13_,r_n_29__12_,r_n_29__11_,r_n_29__10_,
  r_n_29__9_,r_n_29__8_,r_n_29__7_,r_n_29__6_,r_n_29__5_,r_n_29__4_,r_n_29__3_,
  r_n_29__2_,r_n_29__1_,r_n_29__0_,r_n_28__15_,r_n_28__14_,r_n_28__13_,r_n_28__12_,
  r_n_28__11_,r_n_28__10_,r_n_28__9_,r_n_28__8_,r_n_28__7_,r_n_28__6_,r_n_28__5_,
  r_n_28__4_,r_n_28__3_,r_n_28__2_,r_n_28__1_,r_n_28__0_,r_n_27__15_,r_n_27__14_,
  r_n_27__13_,r_n_27__12_,r_n_27__11_,r_n_27__10_,r_n_27__9_,r_n_27__8_,r_n_27__7_,
  r_n_27__6_,r_n_27__5_,r_n_27__4_,r_n_27__3_,r_n_27__2_,r_n_27__1_,r_n_27__0_,
  r_n_26__15_,r_n_26__14_,r_n_26__13_,r_n_26__12_,r_n_26__11_,r_n_26__10_,r_n_26__9_,
  r_n_26__8_,r_n_26__7_,r_n_26__6_,r_n_26__5_,r_n_26__4_,r_n_26__3_,r_n_26__2_,r_n_26__1_,
  r_n_26__0_,r_n_25__15_,r_n_25__14_,r_n_25__13_,r_n_25__12_,r_n_25__11_,
  r_n_25__10_,r_n_25__9_,r_n_25__8_,r_n_25__7_,r_n_25__6_,r_n_25__5_,r_n_25__4_,r_n_25__3_,
  r_n_25__2_,r_n_25__1_,r_n_25__0_,r_n_24__15_,r_n_24__14_,r_n_24__13_,
  r_n_24__12_,r_n_24__11_,r_n_24__10_,r_n_24__9_,r_n_24__8_,r_n_24__7_,r_n_24__6_,r_n_24__5_,
  r_n_24__4_,r_n_24__3_,r_n_24__2_,r_n_24__1_,r_n_24__0_,r_n_23__15_,r_n_23__14_,
  r_n_23__13_,r_n_23__12_,r_n_23__11_,r_n_23__10_,r_n_23__9_,r_n_23__8_,r_n_23__7_,
  r_n_23__6_,r_n_23__5_,r_n_23__4_,r_n_23__3_,r_n_23__2_,r_n_23__1_,r_n_23__0_,
  r_n_22__15_,r_n_22__14_,r_n_22__13_,r_n_22__12_,r_n_22__11_,r_n_22__10_,r_n_22__9_,
  r_n_22__8_,r_n_22__7_,r_n_22__6_,r_n_22__5_,r_n_22__4_,r_n_22__3_,r_n_22__2_,
  r_n_22__1_,r_n_22__0_,r_n_21__15_,r_n_21__14_,r_n_21__13_,r_n_21__12_,r_n_21__11_,
  r_n_21__10_,r_n_21__9_,r_n_21__8_,r_n_21__7_,r_n_21__6_,r_n_21__5_,r_n_21__4_,
  r_n_21__3_,r_n_21__2_,r_n_21__1_,r_n_21__0_,r_n_20__15_,r_n_20__14_,r_n_20__13_,
  r_n_20__12_,r_n_20__11_,r_n_20__10_,r_n_20__9_,r_n_20__8_,r_n_20__7_,r_n_20__6_,
  r_n_20__5_,r_n_20__4_,r_n_20__3_,r_n_20__2_,r_n_20__1_,r_n_20__0_,r_n_19__15_,
  r_n_19__14_,r_n_19__13_,r_n_19__12_,r_n_19__11_,r_n_19__10_,r_n_19__9_,r_n_19__8_,
  r_n_19__7_,r_n_19__6_,r_n_19__5_,r_n_19__4_,r_n_19__3_,r_n_19__2_,r_n_19__1_,
  r_n_19__0_,r_n_18__15_,r_n_18__14_,r_n_18__13_,r_n_18__12_,r_n_18__11_,r_n_18__10_,
  r_n_18__9_,r_n_18__8_,r_n_18__7_,r_n_18__6_,r_n_18__5_,r_n_18__4_,r_n_18__3_,
  r_n_18__2_,r_n_18__1_,r_n_18__0_,r_n_17__15_,r_n_17__14_,r_n_17__13_,r_n_17__12_,
  r_n_17__11_,r_n_17__10_,r_n_17__9_,r_n_17__8_,r_n_17__7_,r_n_17__6_,r_n_17__5_,
  r_n_17__4_,r_n_17__3_,r_n_17__2_,r_n_17__1_,r_n_17__0_,r_n_16__15_,r_n_16__14_,
  r_n_16__13_,r_n_16__12_,r_n_16__11_,r_n_16__10_,r_n_16__9_,r_n_16__8_,r_n_16__7_,
  r_n_16__6_,r_n_16__5_,r_n_16__4_,r_n_16__3_,r_n_16__2_,r_n_16__1_,r_n_16__0_,
  r_n_15__15_,r_n_15__14_,r_n_15__13_,r_n_15__12_,r_n_15__11_,r_n_15__10_,r_n_15__9_,
  r_n_15__8_,r_n_15__7_,r_n_15__6_,r_n_15__5_,r_n_15__4_,r_n_15__3_,r_n_15__2_,
  r_n_15__1_,r_n_15__0_,r_n_14__15_,r_n_14__14_,r_n_14__13_,r_n_14__12_,r_n_14__11_,
  r_n_14__10_,r_n_14__9_,r_n_14__8_,r_n_14__7_,r_n_14__6_,r_n_14__5_,r_n_14__4_,
  r_n_14__3_,r_n_14__2_,r_n_14__1_,r_n_14__0_,r_n_13__15_,r_n_13__14_,r_n_13__13_,
  r_n_13__12_,r_n_13__11_,r_n_13__10_,r_n_13__9_,r_n_13__8_,r_n_13__7_,r_n_13__6_,
  r_n_13__5_,r_n_13__4_,r_n_13__3_,r_n_13__2_,r_n_13__1_,r_n_13__0_,r_n_12__15_,
  r_n_12__14_,r_n_12__13_,r_n_12__12_,r_n_12__11_,r_n_12__10_,r_n_12__9_,r_n_12__8_,
  r_n_12__7_,r_n_12__6_,r_n_12__5_,r_n_12__4_,r_n_12__3_,r_n_12__2_,r_n_12__1_,r_n_12__0_,
  r_n_11__15_,r_n_11__14_,r_n_11__13_,r_n_11__12_,r_n_11__11_,r_n_11__10_,
  r_n_11__9_,r_n_11__8_,r_n_11__7_,r_n_11__6_,r_n_11__5_,r_n_11__4_,r_n_11__3_,r_n_11__2_,
  r_n_11__1_,r_n_11__0_,r_n_10__15_,r_n_10__14_,r_n_10__13_,r_n_10__12_,
  r_n_10__11_,r_n_10__10_,r_n_10__9_,r_n_10__8_,r_n_10__7_,r_n_10__6_,r_n_10__5_,r_n_10__4_,
  r_n_10__3_,r_n_10__2_,r_n_10__1_,r_n_10__0_,r_n_9__15_,r_n_9__14_,r_n_9__13_,
  r_n_9__12_,r_n_9__11_,r_n_9__10_,r_n_9__9_,r_n_9__8_,r_n_9__7_,r_n_9__6_,r_n_9__5_,
  r_n_9__4_,r_n_9__3_,r_n_9__2_,r_n_9__1_,r_n_9__0_,r_n_8__15_,r_n_8__14_,
  r_n_8__13_,r_n_8__12_,r_n_8__11_,r_n_8__10_,r_n_8__9_,r_n_8__8_,r_n_8__7_,r_n_8__6_,
  r_n_8__5_,r_n_8__4_,r_n_8__3_,r_n_8__2_,r_n_8__1_,r_n_8__0_,r_n_7__15_,r_n_7__14_,
  r_n_7__13_,r_n_7__12_,r_n_7__11_,r_n_7__10_,r_n_7__9_,r_n_7__8_,r_n_7__7_,
  r_n_7__6_,r_n_7__5_,r_n_7__4_,r_n_7__3_,r_n_7__2_,r_n_7__1_,r_n_7__0_,r_n_6__15_,
  r_n_6__14_,r_n_6__13_,r_n_6__12_,r_n_6__11_,r_n_6__10_,r_n_6__9_,r_n_6__8_,r_n_6__7_,
  r_n_6__6_,r_n_6__5_,r_n_6__4_,r_n_6__3_,r_n_6__2_,r_n_6__1_,r_n_6__0_,r_n_5__15_,
  r_n_5__14_,r_n_5__13_,r_n_5__12_,r_n_5__11_,r_n_5__10_,r_n_5__9_,r_n_5__8_,
  r_n_5__7_,r_n_5__6_,r_n_5__5_,r_n_5__4_,r_n_5__3_,r_n_5__2_,r_n_5__1_,r_n_5__0_,
  r_n_4__15_,r_n_4__14_,r_n_4__13_,r_n_4__12_,r_n_4__11_,r_n_4__10_,r_n_4__9_,r_n_4__8_,
  r_n_4__7_,r_n_4__6_,r_n_4__5_,r_n_4__4_,r_n_4__3_,r_n_4__2_,r_n_4__1_,r_n_4__0_,
  r_n_3__15_,r_n_3__14_,r_n_3__13_,r_n_3__12_,r_n_3__11_,r_n_3__10_,r_n_3__9_,
  r_n_3__8_,r_n_3__7_,r_n_3__6_,r_n_3__5_,r_n_3__4_,r_n_3__3_,r_n_3__2_,r_n_3__1_,
  r_n_3__0_,r_n_2__15_,r_n_2__14_,r_n_2__13_,r_n_2__12_,r_n_2__11_,r_n_2__10_,
  r_n_2__9_,r_n_2__8_,r_n_2__7_,r_n_2__6_,r_n_2__5_,r_n_2__4_,r_n_2__3_,r_n_2__2_,
  r_n_2__1_,r_n_2__0_,r_n_1__15_,r_n_1__14_,r_n_1__13_,r_n_1__12_,r_n_1__11_,r_n_1__10_,
  r_n_1__9_,r_n_1__8_,r_n_1__7_,r_n_1__6_,r_n_1__5_,r_n_1__4_,r_n_1__3_,r_n_1__2_,
  r_n_1__1_,r_n_1__0_,r_n_62__15_,r_n_62__14_,r_n_62__13_,r_n_62__12_,r_n_62__11_,
  r_n_62__10_,r_n_62__9_,r_n_62__8_,r_n_62__7_,r_n_62__6_,r_n_62__5_,r_n_62__4_,
  r_n_62__3_,r_n_62__2_,r_n_62__1_,r_n_62__0_,r_n_61__15_,r_n_61__14_,r_n_61__13_,
  r_n_61__12_,r_n_61__11_,r_n_61__10_,r_n_61__9_,r_n_61__8_,r_n_61__7_,r_n_61__6_,
  r_n_61__5_,r_n_61__4_,r_n_61__3_,r_n_61__2_,r_n_61__1_,r_n_61__0_,r_n_60__15_,
  r_n_60__14_,r_n_60__13_,r_n_60__12_,r_n_60__11_,r_n_60__10_,r_n_60__9_,r_n_60__8_,
  r_n_60__7_,r_n_60__6_,r_n_60__5_,r_n_60__4_,r_n_60__3_,r_n_60__2_,r_n_60__1_,
  r_n_60__0_,r_n_59__15_,r_n_59__14_,r_n_59__13_,r_n_59__12_,r_n_59__11_,r_n_59__10_,
  r_n_59__9_,r_n_59__8_,r_n_59__7_,r_n_59__6_,r_n_59__5_,r_n_59__4_,r_n_59__3_,
  r_n_59__2_,r_n_59__1_,r_n_59__0_,r_n_58__15_,r_n_58__14_,r_n_58__13_,r_n_58__12_,
  r_n_58__11_,r_n_58__10_,r_n_58__9_,r_n_58__8_,r_n_58__7_,r_n_58__6_,r_n_58__5_,
  r_n_58__4_,r_n_58__3_,r_n_58__2_,r_n_58__1_,r_n_58__0_,r_n_57__15_,r_n_57__14_,
  r_n_57__13_,r_n_57__12_,r_n_57__11_,r_n_57__10_,r_n_57__9_,r_n_57__8_,r_n_57__7_,
  r_n_57__6_,r_n_57__5_,r_n_57__4_,r_n_57__3_,r_n_57__2_,r_n_57__1_,r_n_57__0_,
  r_n_56__15_,r_n_56__14_,r_n_56__13_,r_n_56__12_,r_n_56__11_,r_n_56__10_,r_n_56__9_,
  r_n_56__8_,r_n_56__7_,r_n_56__6_,r_n_56__5_,r_n_56__4_,r_n_56__3_,r_n_56__2_,r_n_56__1_,
  r_n_56__0_,r_n_55__15_,r_n_55__14_,r_n_55__13_,r_n_55__12_,r_n_55__11_,
  r_n_55__10_,r_n_55__9_,r_n_55__8_,r_n_55__7_,r_n_55__6_,r_n_55__5_,r_n_55__4_,r_n_55__3_,
  r_n_55__2_,r_n_55__1_,r_n_55__0_,r_n_54__15_,r_n_54__14_,r_n_54__13_,
  r_n_54__12_,r_n_54__11_,r_n_54__10_,r_n_54__9_,r_n_54__8_,r_n_54__7_,r_n_54__6_,r_n_54__5_,
  r_n_54__4_,r_n_54__3_,r_n_54__2_,r_n_54__1_,r_n_54__0_,r_n_53__15_,r_n_53__14_,
  r_n_53__13_,r_n_53__12_,r_n_53__11_,r_n_53__10_,r_n_53__9_,r_n_53__8_,r_n_53__7_,
  r_n_53__6_,r_n_53__5_,r_n_53__4_,r_n_53__3_,r_n_53__2_,r_n_53__1_,r_n_53__0_,
  r_n_52__15_,r_n_52__14_,r_n_52__13_,r_n_52__12_,r_n_52__11_,r_n_52__10_,r_n_52__9_,
  r_n_52__8_,r_n_52__7_,r_n_52__6_,r_n_52__5_,r_n_52__4_,r_n_52__3_,r_n_52__2_,
  r_n_52__1_,r_n_52__0_,r_n_51__15_,r_n_51__14_,r_n_51__13_,r_n_51__12_,r_n_51__11_,
  r_n_51__10_,r_n_51__9_,r_n_51__8_,r_n_51__7_,r_n_51__6_,r_n_51__5_,r_n_51__4_,
  r_n_51__3_,r_n_51__2_,r_n_51__1_,r_n_51__0_,r_n_50__15_,r_n_50__14_,r_n_50__13_,
  r_n_50__12_,r_n_50__11_,r_n_50__10_,r_n_50__9_,r_n_50__8_,r_n_50__7_,r_n_50__6_,
  r_n_50__5_,r_n_50__4_,r_n_50__3_,r_n_50__2_,r_n_50__1_,r_n_50__0_,r_n_49__15_,
  r_n_49__14_,r_n_49__13_,r_n_49__12_,r_n_49__11_,r_n_49__10_,r_n_49__9_,r_n_49__8_,
  r_n_49__7_,r_n_49__6_,r_n_49__5_,r_n_49__4_,r_n_49__3_,r_n_49__2_,r_n_49__1_,
  r_n_49__0_,r_n_48__15_,r_n_48__14_,r_n_48__13_,r_n_48__12_,r_n_48__11_,r_n_48__10_,
  r_n_48__9_,r_n_48__8_,r_n_48__7_,r_n_48__6_,r_n_48__5_,r_n_48__4_,r_n_48__3_,
  r_n_48__2_,r_n_48__1_,r_n_48__0_,r_n_47__15_,r_n_47__14_,r_n_47__13_,r_n_47__12_,
  r_n_47__11_,r_n_47__10_,r_n_47__9_,r_n_47__8_,r_n_47__7_,r_n_47__6_,r_n_47__5_,
  r_n_47__4_,r_n_47__3_,r_n_47__2_,r_n_47__1_,r_n_47__0_,r_n_46__15_,r_n_46__14_,
  r_n_46__13_,r_n_46__12_,r_n_46__11_,r_n_46__10_,r_n_46__9_,r_n_46__8_,r_n_46__7_,
  r_n_46__6_,r_n_46__5_,r_n_46__4_,r_n_46__3_,r_n_46__2_,r_n_46__1_,r_n_46__0_,
  r_n_45__15_,r_n_45__14_,r_n_45__13_,r_n_45__12_,r_n_45__11_,r_n_45__10_,r_n_45__9_,
  r_n_45__8_,r_n_45__7_,r_n_45__6_,r_n_45__5_,r_n_45__4_,r_n_45__3_,r_n_45__2_,
  r_n_45__1_,r_n_45__0_,r_n_44__15_,r_n_44__14_,r_n_44__13_,r_n_44__12_,r_n_44__11_,
  r_n_44__10_,r_n_44__9_,r_n_44__8_,r_n_44__7_,r_n_44__6_,r_n_44__5_,r_n_44__4_,
  r_n_44__3_,r_n_44__2_,r_n_44__1_,r_n_44__0_,r_n_43__15_,r_n_43__14_,r_n_43__13_,
  r_n_43__12_,r_n_43__11_,r_n_43__10_,r_n_43__9_,r_n_43__8_,r_n_43__7_,r_n_43__6_,
  r_n_43__5_,r_n_43__4_,r_n_43__3_,r_n_43__2_,r_n_43__1_,r_n_43__0_,r_n_42__15_,
  r_n_42__14_,r_n_42__13_,r_n_42__12_,r_n_42__11_,r_n_42__10_,r_n_42__9_,r_n_42__8_,
  r_n_42__7_,r_n_42__6_,r_n_42__5_,r_n_42__4_,r_n_42__3_,r_n_42__2_,r_n_42__1_,r_n_42__0_,
  r_n_41__15_,r_n_41__14_,r_n_41__13_,r_n_41__12_,r_n_41__11_,r_n_41__10_,
  r_n_41__9_,r_n_41__8_,r_n_41__7_,r_n_41__6_,r_n_41__5_,r_n_41__4_,r_n_41__3_,r_n_41__2_,
  r_n_41__1_,r_n_41__0_,r_n_40__15_,r_n_40__14_,r_n_40__13_,r_n_40__12_,
  r_n_40__11_,r_n_40__10_,r_n_40__9_,r_n_40__8_,r_n_40__7_,r_n_40__6_,r_n_40__5_,r_n_40__4_,
  r_n_40__3_,r_n_40__2_,r_n_40__1_,r_n_40__0_,r_n_39__15_,r_n_39__14_,r_n_39__13_,
  r_n_39__12_,r_n_39__11_,r_n_39__10_,r_n_39__9_,r_n_39__8_,r_n_39__7_,r_n_39__6_,
  r_n_39__5_,r_n_39__4_,r_n_39__3_,r_n_39__2_,r_n_39__1_,r_n_39__0_,r_n_38__15_,
  r_n_38__14_,r_n_38__13_,r_n_38__12_,r_n_38__11_,r_n_38__10_,r_n_38__9_,r_n_38__8_,
  r_n_38__7_,r_n_38__6_,r_n_38__5_,r_n_38__4_,r_n_38__3_,r_n_38__2_,r_n_38__1_,
  r_n_38__0_,r_n_37__15_,r_n_37__14_,r_n_37__13_,r_n_37__12_,r_n_37__11_,r_n_37__10_,
  r_n_37__9_,r_n_37__8_,r_n_37__7_,r_n_37__6_,r_n_37__5_,r_n_37__4_,r_n_37__3_,
  r_n_37__2_,r_n_37__1_,r_n_37__0_,r_n_36__15_,r_n_36__14_,r_n_36__13_,r_n_36__12_,
  r_n_36__11_,r_n_36__10_,r_n_36__9_,r_n_36__8_,r_n_36__7_,r_n_36__6_,r_n_36__5_,
  r_n_36__4_,r_n_36__3_,r_n_36__2_,r_n_36__1_,r_n_36__0_,r_n_35__15_,r_n_35__14_,
  r_n_35__13_,r_n_35__12_,r_n_35__11_,r_n_35__10_,r_n_35__9_,r_n_35__8_,r_n_35__7_,
  r_n_35__6_,r_n_35__5_,r_n_35__4_,r_n_35__3_,r_n_35__2_,r_n_35__1_,r_n_35__0_,
  r_n_34__15_,r_n_34__14_,r_n_34__13_,r_n_34__12_,r_n_34__11_,r_n_34__10_,r_n_34__9_,
  r_n_34__8_,r_n_34__7_,r_n_34__6_,r_n_34__5_,r_n_34__4_,r_n_34__3_,r_n_34__2_,
  r_n_34__1_,r_n_34__0_,r_n_33__15_,r_n_33__14_,r_n_33__13_,r_n_33__12_,r_n_33__11_,
  r_n_33__10_,r_n_33__9_,r_n_33__8_,r_n_33__7_,r_n_33__6_,r_n_33__5_,r_n_33__4_,
  r_n_33__3_,r_n_33__2_,r_n_33__1_,r_n_33__0_,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,
  N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,
  N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,
  N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
  N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,
  N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,
  N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,
  N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,
  N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
  N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,
  N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,
  N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,
  N507,N508,N509,N510,N511;
  reg data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg,r_1__15__sv2v_reg,
  r_1__14__sv2v_reg,r_1__13__sv2v_reg,r_1__12__sv2v_reg,r_1__11__sv2v_reg,
  r_1__10__sv2v_reg,r_1__9__sv2v_reg,r_1__8__sv2v_reg,r_1__7__sv2v_reg,r_1__6__sv2v_reg,
  r_1__5__sv2v_reg,r_1__4__sv2v_reg,r_1__3__sv2v_reg,r_1__2__sv2v_reg,r_1__1__sv2v_reg,
  r_1__0__sv2v_reg,r_2__15__sv2v_reg,r_2__14__sv2v_reg,r_2__13__sv2v_reg,
  r_2__12__sv2v_reg,r_2__11__sv2v_reg,r_2__10__sv2v_reg,r_2__9__sv2v_reg,r_2__8__sv2v_reg,
  r_2__7__sv2v_reg,r_2__6__sv2v_reg,r_2__5__sv2v_reg,r_2__4__sv2v_reg,r_2__3__sv2v_reg,
  r_2__2__sv2v_reg,r_2__1__sv2v_reg,r_2__0__sv2v_reg,r_3__15__sv2v_reg,
  r_3__14__sv2v_reg,r_3__13__sv2v_reg,r_3__12__sv2v_reg,r_3__11__sv2v_reg,r_3__10__sv2v_reg,
  r_3__9__sv2v_reg,r_3__8__sv2v_reg,r_3__7__sv2v_reg,r_3__6__sv2v_reg,
  r_3__5__sv2v_reg,r_3__4__sv2v_reg,r_3__3__sv2v_reg,r_3__2__sv2v_reg,r_3__1__sv2v_reg,
  r_3__0__sv2v_reg,r_4__15__sv2v_reg,r_4__14__sv2v_reg,r_4__13__sv2v_reg,r_4__12__sv2v_reg,
  r_4__11__sv2v_reg,r_4__10__sv2v_reg,r_4__9__sv2v_reg,r_4__8__sv2v_reg,
  r_4__7__sv2v_reg,r_4__6__sv2v_reg,r_4__5__sv2v_reg,r_4__4__sv2v_reg,r_4__3__sv2v_reg,
  r_4__2__sv2v_reg,r_4__1__sv2v_reg,r_4__0__sv2v_reg,r_5__15__sv2v_reg,
  r_5__14__sv2v_reg,r_5__13__sv2v_reg,r_5__12__sv2v_reg,r_5__11__sv2v_reg,r_5__10__sv2v_reg,
  r_5__9__sv2v_reg,r_5__8__sv2v_reg,r_5__7__sv2v_reg,r_5__6__sv2v_reg,r_5__5__sv2v_reg,
  r_5__4__sv2v_reg,r_5__3__sv2v_reg,r_5__2__sv2v_reg,r_5__1__sv2v_reg,
  r_5__0__sv2v_reg,r_6__15__sv2v_reg,r_6__14__sv2v_reg,r_6__13__sv2v_reg,r_6__12__sv2v_reg,
  r_6__11__sv2v_reg,r_6__10__sv2v_reg,r_6__9__sv2v_reg,r_6__8__sv2v_reg,
  r_6__7__sv2v_reg,r_6__6__sv2v_reg,r_6__5__sv2v_reg,r_6__4__sv2v_reg,r_6__3__sv2v_reg,
  r_6__2__sv2v_reg,r_6__1__sv2v_reg,r_6__0__sv2v_reg,r_7__15__sv2v_reg,r_7__14__sv2v_reg,
  r_7__13__sv2v_reg,r_7__12__sv2v_reg,r_7__11__sv2v_reg,r_7__10__sv2v_reg,
  r_7__9__sv2v_reg,r_7__8__sv2v_reg,r_7__7__sv2v_reg,r_7__6__sv2v_reg,r_7__5__sv2v_reg,
  r_7__4__sv2v_reg,r_7__3__sv2v_reg,r_7__2__sv2v_reg,r_7__1__sv2v_reg,r_7__0__sv2v_reg,
  r_8__15__sv2v_reg,r_8__14__sv2v_reg,r_8__13__sv2v_reg,r_8__12__sv2v_reg,
  r_8__11__sv2v_reg,r_8__10__sv2v_reg,r_8__9__sv2v_reg,r_8__8__sv2v_reg,r_8__7__sv2v_reg,
  r_8__6__sv2v_reg,r_8__5__sv2v_reg,r_8__4__sv2v_reg,r_8__3__sv2v_reg,
  r_8__2__sv2v_reg,r_8__1__sv2v_reg,r_8__0__sv2v_reg,r_9__15__sv2v_reg,r_9__14__sv2v_reg,
  r_9__13__sv2v_reg,r_9__12__sv2v_reg,r_9__11__sv2v_reg,r_9__10__sv2v_reg,
  r_9__9__sv2v_reg,r_9__8__sv2v_reg,r_9__7__sv2v_reg,r_9__6__sv2v_reg,r_9__5__sv2v_reg,
  r_9__4__sv2v_reg,r_9__3__sv2v_reg,r_9__2__sv2v_reg,r_9__1__sv2v_reg,r_9__0__sv2v_reg,
  r_10__15__sv2v_reg,r_10__14__sv2v_reg,r_10__13__sv2v_reg,r_10__12__sv2v_reg,
  r_10__11__sv2v_reg,r_10__10__sv2v_reg,r_10__9__sv2v_reg,r_10__8__sv2v_reg,
  r_10__7__sv2v_reg,r_10__6__sv2v_reg,r_10__5__sv2v_reg,r_10__4__sv2v_reg,r_10__3__sv2v_reg,
  r_10__2__sv2v_reg,r_10__1__sv2v_reg,r_10__0__sv2v_reg,r_11__15__sv2v_reg,
  r_11__14__sv2v_reg,r_11__13__sv2v_reg,r_11__12__sv2v_reg,r_11__11__sv2v_reg,
  r_11__10__sv2v_reg,r_11__9__sv2v_reg,r_11__8__sv2v_reg,r_11__7__sv2v_reg,r_11__6__sv2v_reg,
  r_11__5__sv2v_reg,r_11__4__sv2v_reg,r_11__3__sv2v_reg,r_11__2__sv2v_reg,
  r_11__1__sv2v_reg,r_11__0__sv2v_reg,r_12__15__sv2v_reg,r_12__14__sv2v_reg,
  r_12__13__sv2v_reg,r_12__12__sv2v_reg,r_12__11__sv2v_reg,r_12__10__sv2v_reg,r_12__9__sv2v_reg,
  r_12__8__sv2v_reg,r_12__7__sv2v_reg,r_12__6__sv2v_reg,r_12__5__sv2v_reg,
  r_12__4__sv2v_reg,r_12__3__sv2v_reg,r_12__2__sv2v_reg,r_12__1__sv2v_reg,r_12__0__sv2v_reg,
  r_13__15__sv2v_reg,r_13__14__sv2v_reg,r_13__13__sv2v_reg,r_13__12__sv2v_reg,
  r_13__11__sv2v_reg,r_13__10__sv2v_reg,r_13__9__sv2v_reg,r_13__8__sv2v_reg,
  r_13__7__sv2v_reg,r_13__6__sv2v_reg,r_13__5__sv2v_reg,r_13__4__sv2v_reg,r_13__3__sv2v_reg,
  r_13__2__sv2v_reg,r_13__1__sv2v_reg,r_13__0__sv2v_reg,r_14__15__sv2v_reg,
  r_14__14__sv2v_reg,r_14__13__sv2v_reg,r_14__12__sv2v_reg,r_14__11__sv2v_reg,
  r_14__10__sv2v_reg,r_14__9__sv2v_reg,r_14__8__sv2v_reg,r_14__7__sv2v_reg,r_14__6__sv2v_reg,
  r_14__5__sv2v_reg,r_14__4__sv2v_reg,r_14__3__sv2v_reg,r_14__2__sv2v_reg,
  r_14__1__sv2v_reg,r_14__0__sv2v_reg,r_15__15__sv2v_reg,r_15__14__sv2v_reg,
  r_15__13__sv2v_reg,r_15__12__sv2v_reg,r_15__11__sv2v_reg,r_15__10__sv2v_reg,r_15__9__sv2v_reg,
  r_15__8__sv2v_reg,r_15__7__sv2v_reg,r_15__6__sv2v_reg,r_15__5__sv2v_reg,
  r_15__4__sv2v_reg,r_15__3__sv2v_reg,r_15__2__sv2v_reg,r_15__1__sv2v_reg,r_15__0__sv2v_reg,
  r_16__15__sv2v_reg,r_16__14__sv2v_reg,r_16__13__sv2v_reg,r_16__12__sv2v_reg,
  r_16__11__sv2v_reg,r_16__10__sv2v_reg,r_16__9__sv2v_reg,r_16__8__sv2v_reg,
  r_16__7__sv2v_reg,r_16__6__sv2v_reg,r_16__5__sv2v_reg,r_16__4__sv2v_reg,r_16__3__sv2v_reg,
  r_16__2__sv2v_reg,r_16__1__sv2v_reg,r_16__0__sv2v_reg,r_17__15__sv2v_reg,
  r_17__14__sv2v_reg,r_17__13__sv2v_reg,r_17__12__sv2v_reg,r_17__11__sv2v_reg,
  r_17__10__sv2v_reg,r_17__9__sv2v_reg,r_17__8__sv2v_reg,r_17__7__sv2v_reg,r_17__6__sv2v_reg,
  r_17__5__sv2v_reg,r_17__4__sv2v_reg,r_17__3__sv2v_reg,r_17__2__sv2v_reg,
  r_17__1__sv2v_reg,r_17__0__sv2v_reg,r_18__15__sv2v_reg,r_18__14__sv2v_reg,
  r_18__13__sv2v_reg,r_18__12__sv2v_reg,r_18__11__sv2v_reg,r_18__10__sv2v_reg,r_18__9__sv2v_reg,
  r_18__8__sv2v_reg,r_18__7__sv2v_reg,r_18__6__sv2v_reg,r_18__5__sv2v_reg,
  r_18__4__sv2v_reg,r_18__3__sv2v_reg,r_18__2__sv2v_reg,r_18__1__sv2v_reg,
  r_18__0__sv2v_reg,r_19__15__sv2v_reg,r_19__14__sv2v_reg,r_19__13__sv2v_reg,r_19__12__sv2v_reg,
  r_19__11__sv2v_reg,r_19__10__sv2v_reg,r_19__9__sv2v_reg,r_19__8__sv2v_reg,
  r_19__7__sv2v_reg,r_19__6__sv2v_reg,r_19__5__sv2v_reg,r_19__4__sv2v_reg,
  r_19__3__sv2v_reg,r_19__2__sv2v_reg,r_19__1__sv2v_reg,r_19__0__sv2v_reg,r_20__15__sv2v_reg,
  r_20__14__sv2v_reg,r_20__13__sv2v_reg,r_20__12__sv2v_reg,r_20__11__sv2v_reg,
  r_20__10__sv2v_reg,r_20__9__sv2v_reg,r_20__8__sv2v_reg,r_20__7__sv2v_reg,
  r_20__6__sv2v_reg,r_20__5__sv2v_reg,r_20__4__sv2v_reg,r_20__3__sv2v_reg,r_20__2__sv2v_reg,
  r_20__1__sv2v_reg,r_20__0__sv2v_reg,r_21__15__sv2v_reg,r_21__14__sv2v_reg,
  r_21__13__sv2v_reg,r_21__12__sv2v_reg,r_21__11__sv2v_reg,r_21__10__sv2v_reg,
  r_21__9__sv2v_reg,r_21__8__sv2v_reg,r_21__7__sv2v_reg,r_21__6__sv2v_reg,r_21__5__sv2v_reg,
  r_21__4__sv2v_reg,r_21__3__sv2v_reg,r_21__2__sv2v_reg,r_21__1__sv2v_reg,
  r_21__0__sv2v_reg,r_22__15__sv2v_reg,r_22__14__sv2v_reg,r_22__13__sv2v_reg,r_22__12__sv2v_reg,
  r_22__11__sv2v_reg,r_22__10__sv2v_reg,r_22__9__sv2v_reg,r_22__8__sv2v_reg,
  r_22__7__sv2v_reg,r_22__6__sv2v_reg,r_22__5__sv2v_reg,r_22__4__sv2v_reg,
  r_22__3__sv2v_reg,r_22__2__sv2v_reg,r_22__1__sv2v_reg,r_22__0__sv2v_reg,r_23__15__sv2v_reg,
  r_23__14__sv2v_reg,r_23__13__sv2v_reg,r_23__12__sv2v_reg,r_23__11__sv2v_reg,
  r_23__10__sv2v_reg,r_23__9__sv2v_reg,r_23__8__sv2v_reg,r_23__7__sv2v_reg,
  r_23__6__sv2v_reg,r_23__5__sv2v_reg,r_23__4__sv2v_reg,r_23__3__sv2v_reg,r_23__2__sv2v_reg,
  r_23__1__sv2v_reg,r_23__0__sv2v_reg,r_24__15__sv2v_reg,r_24__14__sv2v_reg,
  r_24__13__sv2v_reg,r_24__12__sv2v_reg,r_24__11__sv2v_reg,r_24__10__sv2v_reg,
  r_24__9__sv2v_reg,r_24__8__sv2v_reg,r_24__7__sv2v_reg,r_24__6__sv2v_reg,r_24__5__sv2v_reg,
  r_24__4__sv2v_reg,r_24__3__sv2v_reg,r_24__2__sv2v_reg,r_24__1__sv2v_reg,
  r_24__0__sv2v_reg,r_25__15__sv2v_reg,r_25__14__sv2v_reg,r_25__13__sv2v_reg,
  r_25__12__sv2v_reg,r_25__11__sv2v_reg,r_25__10__sv2v_reg,r_25__9__sv2v_reg,r_25__8__sv2v_reg,
  r_25__7__sv2v_reg,r_25__6__sv2v_reg,r_25__5__sv2v_reg,r_25__4__sv2v_reg,
  r_25__3__sv2v_reg,r_25__2__sv2v_reg,r_25__1__sv2v_reg,r_25__0__sv2v_reg,r_26__15__sv2v_reg,
  r_26__14__sv2v_reg,r_26__13__sv2v_reg,r_26__12__sv2v_reg,r_26__11__sv2v_reg,
  r_26__10__sv2v_reg,r_26__9__sv2v_reg,r_26__8__sv2v_reg,r_26__7__sv2v_reg,
  r_26__6__sv2v_reg,r_26__5__sv2v_reg,r_26__4__sv2v_reg,r_26__3__sv2v_reg,r_26__2__sv2v_reg,
  r_26__1__sv2v_reg,r_26__0__sv2v_reg,r_27__15__sv2v_reg,r_27__14__sv2v_reg,
  r_27__13__sv2v_reg,r_27__12__sv2v_reg,r_27__11__sv2v_reg,r_27__10__sv2v_reg,
  r_27__9__sv2v_reg,r_27__8__sv2v_reg,r_27__7__sv2v_reg,r_27__6__sv2v_reg,r_27__5__sv2v_reg,
  r_27__4__sv2v_reg,r_27__3__sv2v_reg,r_27__2__sv2v_reg,r_27__1__sv2v_reg,
  r_27__0__sv2v_reg,r_28__15__sv2v_reg,r_28__14__sv2v_reg,r_28__13__sv2v_reg,
  r_28__12__sv2v_reg,r_28__11__sv2v_reg,r_28__10__sv2v_reg,r_28__9__sv2v_reg,r_28__8__sv2v_reg,
  r_28__7__sv2v_reg,r_28__6__sv2v_reg,r_28__5__sv2v_reg,r_28__4__sv2v_reg,
  r_28__3__sv2v_reg,r_28__2__sv2v_reg,r_28__1__sv2v_reg,r_28__0__sv2v_reg,
  r_29__15__sv2v_reg,r_29__14__sv2v_reg,r_29__13__sv2v_reg,r_29__12__sv2v_reg,r_29__11__sv2v_reg,
  r_29__10__sv2v_reg,r_29__9__sv2v_reg,r_29__8__sv2v_reg,r_29__7__sv2v_reg,
  r_29__6__sv2v_reg,r_29__5__sv2v_reg,r_29__4__sv2v_reg,r_29__3__sv2v_reg,r_29__2__sv2v_reg,
  r_29__1__sv2v_reg,r_29__0__sv2v_reg,r_30__15__sv2v_reg,r_30__14__sv2v_reg,
  r_30__13__sv2v_reg,r_30__12__sv2v_reg,r_30__11__sv2v_reg,r_30__10__sv2v_reg,
  r_30__9__sv2v_reg,r_30__8__sv2v_reg,r_30__7__sv2v_reg,r_30__6__sv2v_reg,r_30__5__sv2v_reg,
  r_30__4__sv2v_reg,r_30__3__sv2v_reg,r_30__2__sv2v_reg,r_30__1__sv2v_reg,
  r_30__0__sv2v_reg,r_31__15__sv2v_reg,r_31__14__sv2v_reg,r_31__13__sv2v_reg,
  r_31__12__sv2v_reg,r_31__11__sv2v_reg,r_31__10__sv2v_reg,r_31__9__sv2v_reg,r_31__8__sv2v_reg,
  r_31__7__sv2v_reg,r_31__6__sv2v_reg,r_31__5__sv2v_reg,r_31__4__sv2v_reg,
  r_31__3__sv2v_reg,r_31__2__sv2v_reg,r_31__1__sv2v_reg,r_31__0__sv2v_reg,
  r_32__15__sv2v_reg,r_32__14__sv2v_reg,r_32__13__sv2v_reg,r_32__12__sv2v_reg,r_32__11__sv2v_reg,
  r_32__10__sv2v_reg,r_32__9__sv2v_reg,r_32__8__sv2v_reg,r_32__7__sv2v_reg,
  r_32__6__sv2v_reg,r_32__5__sv2v_reg,r_32__4__sv2v_reg,r_32__3__sv2v_reg,
  r_32__2__sv2v_reg,r_32__1__sv2v_reg,r_32__0__sv2v_reg,r_33__15__sv2v_reg,r_33__14__sv2v_reg,
  r_33__13__sv2v_reg,r_33__12__sv2v_reg,r_33__11__sv2v_reg,r_33__10__sv2v_reg,
  r_33__9__sv2v_reg,r_33__8__sv2v_reg,r_33__7__sv2v_reg,r_33__6__sv2v_reg,
  r_33__5__sv2v_reg,r_33__4__sv2v_reg,r_33__3__sv2v_reg,r_33__2__sv2v_reg,r_33__1__sv2v_reg,
  r_33__0__sv2v_reg,r_34__15__sv2v_reg,r_34__14__sv2v_reg,r_34__13__sv2v_reg,
  r_34__12__sv2v_reg,r_34__11__sv2v_reg,r_34__10__sv2v_reg,r_34__9__sv2v_reg,
  r_34__8__sv2v_reg,r_34__7__sv2v_reg,r_34__6__sv2v_reg,r_34__5__sv2v_reg,r_34__4__sv2v_reg,
  r_34__3__sv2v_reg,r_34__2__sv2v_reg,r_34__1__sv2v_reg,r_34__0__sv2v_reg,
  r_35__15__sv2v_reg,r_35__14__sv2v_reg,r_35__13__sv2v_reg,r_35__12__sv2v_reg,
  r_35__11__sv2v_reg,r_35__10__sv2v_reg,r_35__9__sv2v_reg,r_35__8__sv2v_reg,r_35__7__sv2v_reg,
  r_35__6__sv2v_reg,r_35__5__sv2v_reg,r_35__4__sv2v_reg,r_35__3__sv2v_reg,
  r_35__2__sv2v_reg,r_35__1__sv2v_reg,r_35__0__sv2v_reg,r_36__15__sv2v_reg,r_36__14__sv2v_reg,
  r_36__13__sv2v_reg,r_36__12__sv2v_reg,r_36__11__sv2v_reg,r_36__10__sv2v_reg,
  r_36__9__sv2v_reg,r_36__8__sv2v_reg,r_36__7__sv2v_reg,r_36__6__sv2v_reg,
  r_36__5__sv2v_reg,r_36__4__sv2v_reg,r_36__3__sv2v_reg,r_36__2__sv2v_reg,r_36__1__sv2v_reg,
  r_36__0__sv2v_reg,r_37__15__sv2v_reg,r_37__14__sv2v_reg,r_37__13__sv2v_reg,
  r_37__12__sv2v_reg,r_37__11__sv2v_reg,r_37__10__sv2v_reg,r_37__9__sv2v_reg,
  r_37__8__sv2v_reg,r_37__7__sv2v_reg,r_37__6__sv2v_reg,r_37__5__sv2v_reg,r_37__4__sv2v_reg,
  r_37__3__sv2v_reg,r_37__2__sv2v_reg,r_37__1__sv2v_reg,r_37__0__sv2v_reg,
  r_38__15__sv2v_reg,r_38__14__sv2v_reg,r_38__13__sv2v_reg,r_38__12__sv2v_reg,
  r_38__11__sv2v_reg,r_38__10__sv2v_reg,r_38__9__sv2v_reg,r_38__8__sv2v_reg,r_38__7__sv2v_reg,
  r_38__6__sv2v_reg,r_38__5__sv2v_reg,r_38__4__sv2v_reg,r_38__3__sv2v_reg,
  r_38__2__sv2v_reg,r_38__1__sv2v_reg,r_38__0__sv2v_reg,r_39__15__sv2v_reg,r_39__14__sv2v_reg,
  r_39__13__sv2v_reg,r_39__12__sv2v_reg,r_39__11__sv2v_reg,r_39__10__sv2v_reg,
  r_39__9__sv2v_reg,r_39__8__sv2v_reg,r_39__7__sv2v_reg,r_39__6__sv2v_reg,
  r_39__5__sv2v_reg,r_39__4__sv2v_reg,r_39__3__sv2v_reg,r_39__2__sv2v_reg,r_39__1__sv2v_reg,
  r_39__0__sv2v_reg,r_40__15__sv2v_reg,r_40__14__sv2v_reg,r_40__13__sv2v_reg,
  r_40__12__sv2v_reg,r_40__11__sv2v_reg,r_40__10__sv2v_reg,r_40__9__sv2v_reg,
  r_40__8__sv2v_reg,r_40__7__sv2v_reg,r_40__6__sv2v_reg,r_40__5__sv2v_reg,r_40__4__sv2v_reg,
  r_40__3__sv2v_reg,r_40__2__sv2v_reg,r_40__1__sv2v_reg,r_40__0__sv2v_reg,
  r_41__15__sv2v_reg,r_41__14__sv2v_reg,r_41__13__sv2v_reg,r_41__12__sv2v_reg,
  r_41__11__sv2v_reg,r_41__10__sv2v_reg,r_41__9__sv2v_reg,r_41__8__sv2v_reg,r_41__7__sv2v_reg,
  r_41__6__sv2v_reg,r_41__5__sv2v_reg,r_41__4__sv2v_reg,r_41__3__sv2v_reg,
  r_41__2__sv2v_reg,r_41__1__sv2v_reg,r_41__0__sv2v_reg,r_42__15__sv2v_reg,
  r_42__14__sv2v_reg,r_42__13__sv2v_reg,r_42__12__sv2v_reg,r_42__11__sv2v_reg,r_42__10__sv2v_reg,
  r_42__9__sv2v_reg,r_42__8__sv2v_reg,r_42__7__sv2v_reg,r_42__6__sv2v_reg,
  r_42__5__sv2v_reg,r_42__4__sv2v_reg,r_42__3__sv2v_reg,r_42__2__sv2v_reg,r_42__1__sv2v_reg,
  r_42__0__sv2v_reg,r_43__15__sv2v_reg,r_43__14__sv2v_reg,r_43__13__sv2v_reg,
  r_43__12__sv2v_reg,r_43__11__sv2v_reg,r_43__10__sv2v_reg,r_43__9__sv2v_reg,
  r_43__8__sv2v_reg,r_43__7__sv2v_reg,r_43__6__sv2v_reg,r_43__5__sv2v_reg,r_43__4__sv2v_reg,
  r_43__3__sv2v_reg,r_43__2__sv2v_reg,r_43__1__sv2v_reg,r_43__0__sv2v_reg,
  r_44__15__sv2v_reg,r_44__14__sv2v_reg,r_44__13__sv2v_reg,r_44__12__sv2v_reg,
  r_44__11__sv2v_reg,r_44__10__sv2v_reg,r_44__9__sv2v_reg,r_44__8__sv2v_reg,r_44__7__sv2v_reg,
  r_44__6__sv2v_reg,r_44__5__sv2v_reg,r_44__4__sv2v_reg,r_44__3__sv2v_reg,
  r_44__2__sv2v_reg,r_44__1__sv2v_reg,r_44__0__sv2v_reg,r_45__15__sv2v_reg,
  r_45__14__sv2v_reg,r_45__13__sv2v_reg,r_45__12__sv2v_reg,r_45__11__sv2v_reg,r_45__10__sv2v_reg,
  r_45__9__sv2v_reg,r_45__8__sv2v_reg,r_45__7__sv2v_reg,r_45__6__sv2v_reg,
  r_45__5__sv2v_reg,r_45__4__sv2v_reg,r_45__3__sv2v_reg,r_45__2__sv2v_reg,
  r_45__1__sv2v_reg,r_45__0__sv2v_reg,r_46__15__sv2v_reg,r_46__14__sv2v_reg,r_46__13__sv2v_reg,
  r_46__12__sv2v_reg,r_46__11__sv2v_reg,r_46__10__sv2v_reg,r_46__9__sv2v_reg,
  r_46__8__sv2v_reg,r_46__7__sv2v_reg,r_46__6__sv2v_reg,r_46__5__sv2v_reg,
  r_46__4__sv2v_reg,r_46__3__sv2v_reg,r_46__2__sv2v_reg,r_46__1__sv2v_reg,r_46__0__sv2v_reg,
  r_47__15__sv2v_reg,r_47__14__sv2v_reg,r_47__13__sv2v_reg,r_47__12__sv2v_reg,
  r_47__11__sv2v_reg,r_47__10__sv2v_reg,r_47__9__sv2v_reg,r_47__8__sv2v_reg,
  r_47__7__sv2v_reg,r_47__6__sv2v_reg,r_47__5__sv2v_reg,r_47__4__sv2v_reg,r_47__3__sv2v_reg,
  r_47__2__sv2v_reg,r_47__1__sv2v_reg,r_47__0__sv2v_reg,r_48__15__sv2v_reg,
  r_48__14__sv2v_reg,r_48__13__sv2v_reg,r_48__12__sv2v_reg,r_48__11__sv2v_reg,
  r_48__10__sv2v_reg,r_48__9__sv2v_reg,r_48__8__sv2v_reg,r_48__7__sv2v_reg,r_48__6__sv2v_reg,
  r_48__5__sv2v_reg,r_48__4__sv2v_reg,r_48__3__sv2v_reg,r_48__2__sv2v_reg,
  r_48__1__sv2v_reg,r_48__0__sv2v_reg,r_49__15__sv2v_reg,r_49__14__sv2v_reg,r_49__13__sv2v_reg,
  r_49__12__sv2v_reg,r_49__11__sv2v_reg,r_49__10__sv2v_reg,r_49__9__sv2v_reg,
  r_49__8__sv2v_reg,r_49__7__sv2v_reg,r_49__6__sv2v_reg,r_49__5__sv2v_reg,
  r_49__4__sv2v_reg,r_49__3__sv2v_reg,r_49__2__sv2v_reg,r_49__1__sv2v_reg,r_49__0__sv2v_reg,
  r_50__15__sv2v_reg,r_50__14__sv2v_reg,r_50__13__sv2v_reg,r_50__12__sv2v_reg,
  r_50__11__sv2v_reg,r_50__10__sv2v_reg,r_50__9__sv2v_reg,r_50__8__sv2v_reg,
  r_50__7__sv2v_reg,r_50__6__sv2v_reg,r_50__5__sv2v_reg,r_50__4__sv2v_reg,r_50__3__sv2v_reg,
  r_50__2__sv2v_reg,r_50__1__sv2v_reg,r_50__0__sv2v_reg,r_51__15__sv2v_reg,
  r_51__14__sv2v_reg,r_51__13__sv2v_reg,r_51__12__sv2v_reg,r_51__11__sv2v_reg,
  r_51__10__sv2v_reg,r_51__9__sv2v_reg,r_51__8__sv2v_reg,r_51__7__sv2v_reg,r_51__6__sv2v_reg,
  r_51__5__sv2v_reg,r_51__4__sv2v_reg,r_51__3__sv2v_reg,r_51__2__sv2v_reg,
  r_51__1__sv2v_reg,r_51__0__sv2v_reg,r_52__15__sv2v_reg,r_52__14__sv2v_reg,
  r_52__13__sv2v_reg,r_52__12__sv2v_reg,r_52__11__sv2v_reg,r_52__10__sv2v_reg,r_52__9__sv2v_reg,
  r_52__8__sv2v_reg,r_52__7__sv2v_reg,r_52__6__sv2v_reg,r_52__5__sv2v_reg,
  r_52__4__sv2v_reg,r_52__3__sv2v_reg,r_52__2__sv2v_reg,r_52__1__sv2v_reg,r_52__0__sv2v_reg,
  r_53__15__sv2v_reg,r_53__14__sv2v_reg,r_53__13__sv2v_reg,r_53__12__sv2v_reg,
  r_53__11__sv2v_reg,r_53__10__sv2v_reg,r_53__9__sv2v_reg,r_53__8__sv2v_reg,
  r_53__7__sv2v_reg,r_53__6__sv2v_reg,r_53__5__sv2v_reg,r_53__4__sv2v_reg,r_53__3__sv2v_reg,
  r_53__2__sv2v_reg,r_53__1__sv2v_reg,r_53__0__sv2v_reg,r_54__15__sv2v_reg,
  r_54__14__sv2v_reg,r_54__13__sv2v_reg,r_54__12__sv2v_reg,r_54__11__sv2v_reg,
  r_54__10__sv2v_reg,r_54__9__sv2v_reg,r_54__8__sv2v_reg,r_54__7__sv2v_reg,r_54__6__sv2v_reg,
  r_54__5__sv2v_reg,r_54__4__sv2v_reg,r_54__3__sv2v_reg,r_54__2__sv2v_reg,
  r_54__1__sv2v_reg,r_54__0__sv2v_reg,r_55__15__sv2v_reg,r_55__14__sv2v_reg,
  r_55__13__sv2v_reg,r_55__12__sv2v_reg,r_55__11__sv2v_reg,r_55__10__sv2v_reg,r_55__9__sv2v_reg,
  r_55__8__sv2v_reg,r_55__7__sv2v_reg,r_55__6__sv2v_reg,r_55__5__sv2v_reg,
  r_55__4__sv2v_reg,r_55__3__sv2v_reg,r_55__2__sv2v_reg,r_55__1__sv2v_reg,r_55__0__sv2v_reg,
  r_56__15__sv2v_reg,r_56__14__sv2v_reg,r_56__13__sv2v_reg,r_56__12__sv2v_reg,
  r_56__11__sv2v_reg,r_56__10__sv2v_reg,r_56__9__sv2v_reg,r_56__8__sv2v_reg,
  r_56__7__sv2v_reg,r_56__6__sv2v_reg,r_56__5__sv2v_reg,r_56__4__sv2v_reg,r_56__3__sv2v_reg,
  r_56__2__sv2v_reg,r_56__1__sv2v_reg,r_56__0__sv2v_reg,r_57__15__sv2v_reg,
  r_57__14__sv2v_reg,r_57__13__sv2v_reg,r_57__12__sv2v_reg,r_57__11__sv2v_reg,
  r_57__10__sv2v_reg,r_57__9__sv2v_reg,r_57__8__sv2v_reg,r_57__7__sv2v_reg,r_57__6__sv2v_reg,
  r_57__5__sv2v_reg,r_57__4__sv2v_reg,r_57__3__sv2v_reg,r_57__2__sv2v_reg,
  r_57__1__sv2v_reg,r_57__0__sv2v_reg,r_58__15__sv2v_reg,r_58__14__sv2v_reg,
  r_58__13__sv2v_reg,r_58__12__sv2v_reg,r_58__11__sv2v_reg,r_58__10__sv2v_reg,r_58__9__sv2v_reg,
  r_58__8__sv2v_reg,r_58__7__sv2v_reg,r_58__6__sv2v_reg,r_58__5__sv2v_reg,
  r_58__4__sv2v_reg,r_58__3__sv2v_reg,r_58__2__sv2v_reg,r_58__1__sv2v_reg,
  r_58__0__sv2v_reg,r_59__15__sv2v_reg,r_59__14__sv2v_reg,r_59__13__sv2v_reg,r_59__12__sv2v_reg,
  r_59__11__sv2v_reg,r_59__10__sv2v_reg,r_59__9__sv2v_reg,r_59__8__sv2v_reg,
  r_59__7__sv2v_reg,r_59__6__sv2v_reg,r_59__5__sv2v_reg,r_59__4__sv2v_reg,
  r_59__3__sv2v_reg,r_59__2__sv2v_reg,r_59__1__sv2v_reg,r_59__0__sv2v_reg,r_60__15__sv2v_reg,
  r_60__14__sv2v_reg,r_60__13__sv2v_reg,r_60__12__sv2v_reg,r_60__11__sv2v_reg,
  r_60__10__sv2v_reg,r_60__9__sv2v_reg,r_60__8__sv2v_reg,r_60__7__sv2v_reg,
  r_60__6__sv2v_reg,r_60__5__sv2v_reg,r_60__4__sv2v_reg,r_60__3__sv2v_reg,r_60__2__sv2v_reg,
  r_60__1__sv2v_reg,r_60__0__sv2v_reg,r_61__15__sv2v_reg,r_61__14__sv2v_reg,
  r_61__13__sv2v_reg,r_61__12__sv2v_reg,r_61__11__sv2v_reg,r_61__10__sv2v_reg,
  r_61__9__sv2v_reg,r_61__8__sv2v_reg,r_61__7__sv2v_reg,r_61__6__sv2v_reg,r_61__5__sv2v_reg,
  r_61__4__sv2v_reg,r_61__3__sv2v_reg,r_61__2__sv2v_reg,r_61__1__sv2v_reg,
  r_61__0__sv2v_reg,r_62__15__sv2v_reg,r_62__14__sv2v_reg,r_62__13__sv2v_reg,r_62__12__sv2v_reg,
  r_62__11__sv2v_reg,r_62__10__sv2v_reg,r_62__9__sv2v_reg,r_62__8__sv2v_reg,
  r_62__7__sv2v_reg,r_62__6__sv2v_reg,r_62__5__sv2v_reg,r_62__4__sv2v_reg,
  r_62__3__sv2v_reg,r_62__2__sv2v_reg,r_62__1__sv2v_reg,r_62__0__sv2v_reg,r_63__15__sv2v_reg,
  r_63__14__sv2v_reg,r_63__13__sv2v_reg,r_63__12__sv2v_reg,r_63__11__sv2v_reg,
  r_63__10__sv2v_reg,r_63__9__sv2v_reg,r_63__8__sv2v_reg,r_63__7__sv2v_reg,
  r_63__6__sv2v_reg,r_63__5__sv2v_reg,r_63__4__sv2v_reg,r_63__3__sv2v_reg,r_63__2__sv2v_reg,
  r_63__1__sv2v_reg,r_63__0__sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;
  assign r_1__15_ = r_1__15__sv2v_reg;
  assign r_1__14_ = r_1__14__sv2v_reg;
  assign r_1__13_ = r_1__13__sv2v_reg;
  assign r_1__12_ = r_1__12__sv2v_reg;
  assign r_1__11_ = r_1__11__sv2v_reg;
  assign r_1__10_ = r_1__10__sv2v_reg;
  assign r_1__9_ = r_1__9__sv2v_reg;
  assign r_1__8_ = r_1__8__sv2v_reg;
  assign r_1__7_ = r_1__7__sv2v_reg;
  assign r_1__6_ = r_1__6__sv2v_reg;
  assign r_1__5_ = r_1__5__sv2v_reg;
  assign r_1__4_ = r_1__4__sv2v_reg;
  assign r_1__3_ = r_1__3__sv2v_reg;
  assign r_1__2_ = r_1__2__sv2v_reg;
  assign r_1__1_ = r_1__1__sv2v_reg;
  assign r_1__0_ = r_1__0__sv2v_reg;
  assign r_2__15_ = r_2__15__sv2v_reg;
  assign r_2__14_ = r_2__14__sv2v_reg;
  assign r_2__13_ = r_2__13__sv2v_reg;
  assign r_2__12_ = r_2__12__sv2v_reg;
  assign r_2__11_ = r_2__11__sv2v_reg;
  assign r_2__10_ = r_2__10__sv2v_reg;
  assign r_2__9_ = r_2__9__sv2v_reg;
  assign r_2__8_ = r_2__8__sv2v_reg;
  assign r_2__7_ = r_2__7__sv2v_reg;
  assign r_2__6_ = r_2__6__sv2v_reg;
  assign r_2__5_ = r_2__5__sv2v_reg;
  assign r_2__4_ = r_2__4__sv2v_reg;
  assign r_2__3_ = r_2__3__sv2v_reg;
  assign r_2__2_ = r_2__2__sv2v_reg;
  assign r_2__1_ = r_2__1__sv2v_reg;
  assign r_2__0_ = r_2__0__sv2v_reg;
  assign r_3__15_ = r_3__15__sv2v_reg;
  assign r_3__14_ = r_3__14__sv2v_reg;
  assign r_3__13_ = r_3__13__sv2v_reg;
  assign r_3__12_ = r_3__12__sv2v_reg;
  assign r_3__11_ = r_3__11__sv2v_reg;
  assign r_3__10_ = r_3__10__sv2v_reg;
  assign r_3__9_ = r_3__9__sv2v_reg;
  assign r_3__8_ = r_3__8__sv2v_reg;
  assign r_3__7_ = r_3__7__sv2v_reg;
  assign r_3__6_ = r_3__6__sv2v_reg;
  assign r_3__5_ = r_3__5__sv2v_reg;
  assign r_3__4_ = r_3__4__sv2v_reg;
  assign r_3__3_ = r_3__3__sv2v_reg;
  assign r_3__2_ = r_3__2__sv2v_reg;
  assign r_3__1_ = r_3__1__sv2v_reg;
  assign r_3__0_ = r_3__0__sv2v_reg;
  assign r_4__15_ = r_4__15__sv2v_reg;
  assign r_4__14_ = r_4__14__sv2v_reg;
  assign r_4__13_ = r_4__13__sv2v_reg;
  assign r_4__12_ = r_4__12__sv2v_reg;
  assign r_4__11_ = r_4__11__sv2v_reg;
  assign r_4__10_ = r_4__10__sv2v_reg;
  assign r_4__9_ = r_4__9__sv2v_reg;
  assign r_4__8_ = r_4__8__sv2v_reg;
  assign r_4__7_ = r_4__7__sv2v_reg;
  assign r_4__6_ = r_4__6__sv2v_reg;
  assign r_4__5_ = r_4__5__sv2v_reg;
  assign r_4__4_ = r_4__4__sv2v_reg;
  assign r_4__3_ = r_4__3__sv2v_reg;
  assign r_4__2_ = r_4__2__sv2v_reg;
  assign r_4__1_ = r_4__1__sv2v_reg;
  assign r_4__0_ = r_4__0__sv2v_reg;
  assign r_5__15_ = r_5__15__sv2v_reg;
  assign r_5__14_ = r_5__14__sv2v_reg;
  assign r_5__13_ = r_5__13__sv2v_reg;
  assign r_5__12_ = r_5__12__sv2v_reg;
  assign r_5__11_ = r_5__11__sv2v_reg;
  assign r_5__10_ = r_5__10__sv2v_reg;
  assign r_5__9_ = r_5__9__sv2v_reg;
  assign r_5__8_ = r_5__8__sv2v_reg;
  assign r_5__7_ = r_5__7__sv2v_reg;
  assign r_5__6_ = r_5__6__sv2v_reg;
  assign r_5__5_ = r_5__5__sv2v_reg;
  assign r_5__4_ = r_5__4__sv2v_reg;
  assign r_5__3_ = r_5__3__sv2v_reg;
  assign r_5__2_ = r_5__2__sv2v_reg;
  assign r_5__1_ = r_5__1__sv2v_reg;
  assign r_5__0_ = r_5__0__sv2v_reg;
  assign r_6__15_ = r_6__15__sv2v_reg;
  assign r_6__14_ = r_6__14__sv2v_reg;
  assign r_6__13_ = r_6__13__sv2v_reg;
  assign r_6__12_ = r_6__12__sv2v_reg;
  assign r_6__11_ = r_6__11__sv2v_reg;
  assign r_6__10_ = r_6__10__sv2v_reg;
  assign r_6__9_ = r_6__9__sv2v_reg;
  assign r_6__8_ = r_6__8__sv2v_reg;
  assign r_6__7_ = r_6__7__sv2v_reg;
  assign r_6__6_ = r_6__6__sv2v_reg;
  assign r_6__5_ = r_6__5__sv2v_reg;
  assign r_6__4_ = r_6__4__sv2v_reg;
  assign r_6__3_ = r_6__3__sv2v_reg;
  assign r_6__2_ = r_6__2__sv2v_reg;
  assign r_6__1_ = r_6__1__sv2v_reg;
  assign r_6__0_ = r_6__0__sv2v_reg;
  assign r_7__15_ = r_7__15__sv2v_reg;
  assign r_7__14_ = r_7__14__sv2v_reg;
  assign r_7__13_ = r_7__13__sv2v_reg;
  assign r_7__12_ = r_7__12__sv2v_reg;
  assign r_7__11_ = r_7__11__sv2v_reg;
  assign r_7__10_ = r_7__10__sv2v_reg;
  assign r_7__9_ = r_7__9__sv2v_reg;
  assign r_7__8_ = r_7__8__sv2v_reg;
  assign r_7__7_ = r_7__7__sv2v_reg;
  assign r_7__6_ = r_7__6__sv2v_reg;
  assign r_7__5_ = r_7__5__sv2v_reg;
  assign r_7__4_ = r_7__4__sv2v_reg;
  assign r_7__3_ = r_7__3__sv2v_reg;
  assign r_7__2_ = r_7__2__sv2v_reg;
  assign r_7__1_ = r_7__1__sv2v_reg;
  assign r_7__0_ = r_7__0__sv2v_reg;
  assign r_8__15_ = r_8__15__sv2v_reg;
  assign r_8__14_ = r_8__14__sv2v_reg;
  assign r_8__13_ = r_8__13__sv2v_reg;
  assign r_8__12_ = r_8__12__sv2v_reg;
  assign r_8__11_ = r_8__11__sv2v_reg;
  assign r_8__10_ = r_8__10__sv2v_reg;
  assign r_8__9_ = r_8__9__sv2v_reg;
  assign r_8__8_ = r_8__8__sv2v_reg;
  assign r_8__7_ = r_8__7__sv2v_reg;
  assign r_8__6_ = r_8__6__sv2v_reg;
  assign r_8__5_ = r_8__5__sv2v_reg;
  assign r_8__4_ = r_8__4__sv2v_reg;
  assign r_8__3_ = r_8__3__sv2v_reg;
  assign r_8__2_ = r_8__2__sv2v_reg;
  assign r_8__1_ = r_8__1__sv2v_reg;
  assign r_8__0_ = r_8__0__sv2v_reg;
  assign r_9__15_ = r_9__15__sv2v_reg;
  assign r_9__14_ = r_9__14__sv2v_reg;
  assign r_9__13_ = r_9__13__sv2v_reg;
  assign r_9__12_ = r_9__12__sv2v_reg;
  assign r_9__11_ = r_9__11__sv2v_reg;
  assign r_9__10_ = r_9__10__sv2v_reg;
  assign r_9__9_ = r_9__9__sv2v_reg;
  assign r_9__8_ = r_9__8__sv2v_reg;
  assign r_9__7_ = r_9__7__sv2v_reg;
  assign r_9__6_ = r_9__6__sv2v_reg;
  assign r_9__5_ = r_9__5__sv2v_reg;
  assign r_9__4_ = r_9__4__sv2v_reg;
  assign r_9__3_ = r_9__3__sv2v_reg;
  assign r_9__2_ = r_9__2__sv2v_reg;
  assign r_9__1_ = r_9__1__sv2v_reg;
  assign r_9__0_ = r_9__0__sv2v_reg;
  assign r_10__15_ = r_10__15__sv2v_reg;
  assign r_10__14_ = r_10__14__sv2v_reg;
  assign r_10__13_ = r_10__13__sv2v_reg;
  assign r_10__12_ = r_10__12__sv2v_reg;
  assign r_10__11_ = r_10__11__sv2v_reg;
  assign r_10__10_ = r_10__10__sv2v_reg;
  assign r_10__9_ = r_10__9__sv2v_reg;
  assign r_10__8_ = r_10__8__sv2v_reg;
  assign r_10__7_ = r_10__7__sv2v_reg;
  assign r_10__6_ = r_10__6__sv2v_reg;
  assign r_10__5_ = r_10__5__sv2v_reg;
  assign r_10__4_ = r_10__4__sv2v_reg;
  assign r_10__3_ = r_10__3__sv2v_reg;
  assign r_10__2_ = r_10__2__sv2v_reg;
  assign r_10__1_ = r_10__1__sv2v_reg;
  assign r_10__0_ = r_10__0__sv2v_reg;
  assign r_11__15_ = r_11__15__sv2v_reg;
  assign r_11__14_ = r_11__14__sv2v_reg;
  assign r_11__13_ = r_11__13__sv2v_reg;
  assign r_11__12_ = r_11__12__sv2v_reg;
  assign r_11__11_ = r_11__11__sv2v_reg;
  assign r_11__10_ = r_11__10__sv2v_reg;
  assign r_11__9_ = r_11__9__sv2v_reg;
  assign r_11__8_ = r_11__8__sv2v_reg;
  assign r_11__7_ = r_11__7__sv2v_reg;
  assign r_11__6_ = r_11__6__sv2v_reg;
  assign r_11__5_ = r_11__5__sv2v_reg;
  assign r_11__4_ = r_11__4__sv2v_reg;
  assign r_11__3_ = r_11__3__sv2v_reg;
  assign r_11__2_ = r_11__2__sv2v_reg;
  assign r_11__1_ = r_11__1__sv2v_reg;
  assign r_11__0_ = r_11__0__sv2v_reg;
  assign r_12__15_ = r_12__15__sv2v_reg;
  assign r_12__14_ = r_12__14__sv2v_reg;
  assign r_12__13_ = r_12__13__sv2v_reg;
  assign r_12__12_ = r_12__12__sv2v_reg;
  assign r_12__11_ = r_12__11__sv2v_reg;
  assign r_12__10_ = r_12__10__sv2v_reg;
  assign r_12__9_ = r_12__9__sv2v_reg;
  assign r_12__8_ = r_12__8__sv2v_reg;
  assign r_12__7_ = r_12__7__sv2v_reg;
  assign r_12__6_ = r_12__6__sv2v_reg;
  assign r_12__5_ = r_12__5__sv2v_reg;
  assign r_12__4_ = r_12__4__sv2v_reg;
  assign r_12__3_ = r_12__3__sv2v_reg;
  assign r_12__2_ = r_12__2__sv2v_reg;
  assign r_12__1_ = r_12__1__sv2v_reg;
  assign r_12__0_ = r_12__0__sv2v_reg;
  assign r_13__15_ = r_13__15__sv2v_reg;
  assign r_13__14_ = r_13__14__sv2v_reg;
  assign r_13__13_ = r_13__13__sv2v_reg;
  assign r_13__12_ = r_13__12__sv2v_reg;
  assign r_13__11_ = r_13__11__sv2v_reg;
  assign r_13__10_ = r_13__10__sv2v_reg;
  assign r_13__9_ = r_13__9__sv2v_reg;
  assign r_13__8_ = r_13__8__sv2v_reg;
  assign r_13__7_ = r_13__7__sv2v_reg;
  assign r_13__6_ = r_13__6__sv2v_reg;
  assign r_13__5_ = r_13__5__sv2v_reg;
  assign r_13__4_ = r_13__4__sv2v_reg;
  assign r_13__3_ = r_13__3__sv2v_reg;
  assign r_13__2_ = r_13__2__sv2v_reg;
  assign r_13__1_ = r_13__1__sv2v_reg;
  assign r_13__0_ = r_13__0__sv2v_reg;
  assign r_14__15_ = r_14__15__sv2v_reg;
  assign r_14__14_ = r_14__14__sv2v_reg;
  assign r_14__13_ = r_14__13__sv2v_reg;
  assign r_14__12_ = r_14__12__sv2v_reg;
  assign r_14__11_ = r_14__11__sv2v_reg;
  assign r_14__10_ = r_14__10__sv2v_reg;
  assign r_14__9_ = r_14__9__sv2v_reg;
  assign r_14__8_ = r_14__8__sv2v_reg;
  assign r_14__7_ = r_14__7__sv2v_reg;
  assign r_14__6_ = r_14__6__sv2v_reg;
  assign r_14__5_ = r_14__5__sv2v_reg;
  assign r_14__4_ = r_14__4__sv2v_reg;
  assign r_14__3_ = r_14__3__sv2v_reg;
  assign r_14__2_ = r_14__2__sv2v_reg;
  assign r_14__1_ = r_14__1__sv2v_reg;
  assign r_14__0_ = r_14__0__sv2v_reg;
  assign r_15__15_ = r_15__15__sv2v_reg;
  assign r_15__14_ = r_15__14__sv2v_reg;
  assign r_15__13_ = r_15__13__sv2v_reg;
  assign r_15__12_ = r_15__12__sv2v_reg;
  assign r_15__11_ = r_15__11__sv2v_reg;
  assign r_15__10_ = r_15__10__sv2v_reg;
  assign r_15__9_ = r_15__9__sv2v_reg;
  assign r_15__8_ = r_15__8__sv2v_reg;
  assign r_15__7_ = r_15__7__sv2v_reg;
  assign r_15__6_ = r_15__6__sv2v_reg;
  assign r_15__5_ = r_15__5__sv2v_reg;
  assign r_15__4_ = r_15__4__sv2v_reg;
  assign r_15__3_ = r_15__3__sv2v_reg;
  assign r_15__2_ = r_15__2__sv2v_reg;
  assign r_15__1_ = r_15__1__sv2v_reg;
  assign r_15__0_ = r_15__0__sv2v_reg;
  assign r_16__15_ = r_16__15__sv2v_reg;
  assign r_16__14_ = r_16__14__sv2v_reg;
  assign r_16__13_ = r_16__13__sv2v_reg;
  assign r_16__12_ = r_16__12__sv2v_reg;
  assign r_16__11_ = r_16__11__sv2v_reg;
  assign r_16__10_ = r_16__10__sv2v_reg;
  assign r_16__9_ = r_16__9__sv2v_reg;
  assign r_16__8_ = r_16__8__sv2v_reg;
  assign r_16__7_ = r_16__7__sv2v_reg;
  assign r_16__6_ = r_16__6__sv2v_reg;
  assign r_16__5_ = r_16__5__sv2v_reg;
  assign r_16__4_ = r_16__4__sv2v_reg;
  assign r_16__3_ = r_16__3__sv2v_reg;
  assign r_16__2_ = r_16__2__sv2v_reg;
  assign r_16__1_ = r_16__1__sv2v_reg;
  assign r_16__0_ = r_16__0__sv2v_reg;
  assign r_17__15_ = r_17__15__sv2v_reg;
  assign r_17__14_ = r_17__14__sv2v_reg;
  assign r_17__13_ = r_17__13__sv2v_reg;
  assign r_17__12_ = r_17__12__sv2v_reg;
  assign r_17__11_ = r_17__11__sv2v_reg;
  assign r_17__10_ = r_17__10__sv2v_reg;
  assign r_17__9_ = r_17__9__sv2v_reg;
  assign r_17__8_ = r_17__8__sv2v_reg;
  assign r_17__7_ = r_17__7__sv2v_reg;
  assign r_17__6_ = r_17__6__sv2v_reg;
  assign r_17__5_ = r_17__5__sv2v_reg;
  assign r_17__4_ = r_17__4__sv2v_reg;
  assign r_17__3_ = r_17__3__sv2v_reg;
  assign r_17__2_ = r_17__2__sv2v_reg;
  assign r_17__1_ = r_17__1__sv2v_reg;
  assign r_17__0_ = r_17__0__sv2v_reg;
  assign r_18__15_ = r_18__15__sv2v_reg;
  assign r_18__14_ = r_18__14__sv2v_reg;
  assign r_18__13_ = r_18__13__sv2v_reg;
  assign r_18__12_ = r_18__12__sv2v_reg;
  assign r_18__11_ = r_18__11__sv2v_reg;
  assign r_18__10_ = r_18__10__sv2v_reg;
  assign r_18__9_ = r_18__9__sv2v_reg;
  assign r_18__8_ = r_18__8__sv2v_reg;
  assign r_18__7_ = r_18__7__sv2v_reg;
  assign r_18__6_ = r_18__6__sv2v_reg;
  assign r_18__5_ = r_18__5__sv2v_reg;
  assign r_18__4_ = r_18__4__sv2v_reg;
  assign r_18__3_ = r_18__3__sv2v_reg;
  assign r_18__2_ = r_18__2__sv2v_reg;
  assign r_18__1_ = r_18__1__sv2v_reg;
  assign r_18__0_ = r_18__0__sv2v_reg;
  assign r_19__15_ = r_19__15__sv2v_reg;
  assign r_19__14_ = r_19__14__sv2v_reg;
  assign r_19__13_ = r_19__13__sv2v_reg;
  assign r_19__12_ = r_19__12__sv2v_reg;
  assign r_19__11_ = r_19__11__sv2v_reg;
  assign r_19__10_ = r_19__10__sv2v_reg;
  assign r_19__9_ = r_19__9__sv2v_reg;
  assign r_19__8_ = r_19__8__sv2v_reg;
  assign r_19__7_ = r_19__7__sv2v_reg;
  assign r_19__6_ = r_19__6__sv2v_reg;
  assign r_19__5_ = r_19__5__sv2v_reg;
  assign r_19__4_ = r_19__4__sv2v_reg;
  assign r_19__3_ = r_19__3__sv2v_reg;
  assign r_19__2_ = r_19__2__sv2v_reg;
  assign r_19__1_ = r_19__1__sv2v_reg;
  assign r_19__0_ = r_19__0__sv2v_reg;
  assign r_20__15_ = r_20__15__sv2v_reg;
  assign r_20__14_ = r_20__14__sv2v_reg;
  assign r_20__13_ = r_20__13__sv2v_reg;
  assign r_20__12_ = r_20__12__sv2v_reg;
  assign r_20__11_ = r_20__11__sv2v_reg;
  assign r_20__10_ = r_20__10__sv2v_reg;
  assign r_20__9_ = r_20__9__sv2v_reg;
  assign r_20__8_ = r_20__8__sv2v_reg;
  assign r_20__7_ = r_20__7__sv2v_reg;
  assign r_20__6_ = r_20__6__sv2v_reg;
  assign r_20__5_ = r_20__5__sv2v_reg;
  assign r_20__4_ = r_20__4__sv2v_reg;
  assign r_20__3_ = r_20__3__sv2v_reg;
  assign r_20__2_ = r_20__2__sv2v_reg;
  assign r_20__1_ = r_20__1__sv2v_reg;
  assign r_20__0_ = r_20__0__sv2v_reg;
  assign r_21__15_ = r_21__15__sv2v_reg;
  assign r_21__14_ = r_21__14__sv2v_reg;
  assign r_21__13_ = r_21__13__sv2v_reg;
  assign r_21__12_ = r_21__12__sv2v_reg;
  assign r_21__11_ = r_21__11__sv2v_reg;
  assign r_21__10_ = r_21__10__sv2v_reg;
  assign r_21__9_ = r_21__9__sv2v_reg;
  assign r_21__8_ = r_21__8__sv2v_reg;
  assign r_21__7_ = r_21__7__sv2v_reg;
  assign r_21__6_ = r_21__6__sv2v_reg;
  assign r_21__5_ = r_21__5__sv2v_reg;
  assign r_21__4_ = r_21__4__sv2v_reg;
  assign r_21__3_ = r_21__3__sv2v_reg;
  assign r_21__2_ = r_21__2__sv2v_reg;
  assign r_21__1_ = r_21__1__sv2v_reg;
  assign r_21__0_ = r_21__0__sv2v_reg;
  assign r_22__15_ = r_22__15__sv2v_reg;
  assign r_22__14_ = r_22__14__sv2v_reg;
  assign r_22__13_ = r_22__13__sv2v_reg;
  assign r_22__12_ = r_22__12__sv2v_reg;
  assign r_22__11_ = r_22__11__sv2v_reg;
  assign r_22__10_ = r_22__10__sv2v_reg;
  assign r_22__9_ = r_22__9__sv2v_reg;
  assign r_22__8_ = r_22__8__sv2v_reg;
  assign r_22__7_ = r_22__7__sv2v_reg;
  assign r_22__6_ = r_22__6__sv2v_reg;
  assign r_22__5_ = r_22__5__sv2v_reg;
  assign r_22__4_ = r_22__4__sv2v_reg;
  assign r_22__3_ = r_22__3__sv2v_reg;
  assign r_22__2_ = r_22__2__sv2v_reg;
  assign r_22__1_ = r_22__1__sv2v_reg;
  assign r_22__0_ = r_22__0__sv2v_reg;
  assign r_23__15_ = r_23__15__sv2v_reg;
  assign r_23__14_ = r_23__14__sv2v_reg;
  assign r_23__13_ = r_23__13__sv2v_reg;
  assign r_23__12_ = r_23__12__sv2v_reg;
  assign r_23__11_ = r_23__11__sv2v_reg;
  assign r_23__10_ = r_23__10__sv2v_reg;
  assign r_23__9_ = r_23__9__sv2v_reg;
  assign r_23__8_ = r_23__8__sv2v_reg;
  assign r_23__7_ = r_23__7__sv2v_reg;
  assign r_23__6_ = r_23__6__sv2v_reg;
  assign r_23__5_ = r_23__5__sv2v_reg;
  assign r_23__4_ = r_23__4__sv2v_reg;
  assign r_23__3_ = r_23__3__sv2v_reg;
  assign r_23__2_ = r_23__2__sv2v_reg;
  assign r_23__1_ = r_23__1__sv2v_reg;
  assign r_23__0_ = r_23__0__sv2v_reg;
  assign r_24__15_ = r_24__15__sv2v_reg;
  assign r_24__14_ = r_24__14__sv2v_reg;
  assign r_24__13_ = r_24__13__sv2v_reg;
  assign r_24__12_ = r_24__12__sv2v_reg;
  assign r_24__11_ = r_24__11__sv2v_reg;
  assign r_24__10_ = r_24__10__sv2v_reg;
  assign r_24__9_ = r_24__9__sv2v_reg;
  assign r_24__8_ = r_24__8__sv2v_reg;
  assign r_24__7_ = r_24__7__sv2v_reg;
  assign r_24__6_ = r_24__6__sv2v_reg;
  assign r_24__5_ = r_24__5__sv2v_reg;
  assign r_24__4_ = r_24__4__sv2v_reg;
  assign r_24__3_ = r_24__3__sv2v_reg;
  assign r_24__2_ = r_24__2__sv2v_reg;
  assign r_24__1_ = r_24__1__sv2v_reg;
  assign r_24__0_ = r_24__0__sv2v_reg;
  assign r_25__15_ = r_25__15__sv2v_reg;
  assign r_25__14_ = r_25__14__sv2v_reg;
  assign r_25__13_ = r_25__13__sv2v_reg;
  assign r_25__12_ = r_25__12__sv2v_reg;
  assign r_25__11_ = r_25__11__sv2v_reg;
  assign r_25__10_ = r_25__10__sv2v_reg;
  assign r_25__9_ = r_25__9__sv2v_reg;
  assign r_25__8_ = r_25__8__sv2v_reg;
  assign r_25__7_ = r_25__7__sv2v_reg;
  assign r_25__6_ = r_25__6__sv2v_reg;
  assign r_25__5_ = r_25__5__sv2v_reg;
  assign r_25__4_ = r_25__4__sv2v_reg;
  assign r_25__3_ = r_25__3__sv2v_reg;
  assign r_25__2_ = r_25__2__sv2v_reg;
  assign r_25__1_ = r_25__1__sv2v_reg;
  assign r_25__0_ = r_25__0__sv2v_reg;
  assign r_26__15_ = r_26__15__sv2v_reg;
  assign r_26__14_ = r_26__14__sv2v_reg;
  assign r_26__13_ = r_26__13__sv2v_reg;
  assign r_26__12_ = r_26__12__sv2v_reg;
  assign r_26__11_ = r_26__11__sv2v_reg;
  assign r_26__10_ = r_26__10__sv2v_reg;
  assign r_26__9_ = r_26__9__sv2v_reg;
  assign r_26__8_ = r_26__8__sv2v_reg;
  assign r_26__7_ = r_26__7__sv2v_reg;
  assign r_26__6_ = r_26__6__sv2v_reg;
  assign r_26__5_ = r_26__5__sv2v_reg;
  assign r_26__4_ = r_26__4__sv2v_reg;
  assign r_26__3_ = r_26__3__sv2v_reg;
  assign r_26__2_ = r_26__2__sv2v_reg;
  assign r_26__1_ = r_26__1__sv2v_reg;
  assign r_26__0_ = r_26__0__sv2v_reg;
  assign r_27__15_ = r_27__15__sv2v_reg;
  assign r_27__14_ = r_27__14__sv2v_reg;
  assign r_27__13_ = r_27__13__sv2v_reg;
  assign r_27__12_ = r_27__12__sv2v_reg;
  assign r_27__11_ = r_27__11__sv2v_reg;
  assign r_27__10_ = r_27__10__sv2v_reg;
  assign r_27__9_ = r_27__9__sv2v_reg;
  assign r_27__8_ = r_27__8__sv2v_reg;
  assign r_27__7_ = r_27__7__sv2v_reg;
  assign r_27__6_ = r_27__6__sv2v_reg;
  assign r_27__5_ = r_27__5__sv2v_reg;
  assign r_27__4_ = r_27__4__sv2v_reg;
  assign r_27__3_ = r_27__3__sv2v_reg;
  assign r_27__2_ = r_27__2__sv2v_reg;
  assign r_27__1_ = r_27__1__sv2v_reg;
  assign r_27__0_ = r_27__0__sv2v_reg;
  assign r_28__15_ = r_28__15__sv2v_reg;
  assign r_28__14_ = r_28__14__sv2v_reg;
  assign r_28__13_ = r_28__13__sv2v_reg;
  assign r_28__12_ = r_28__12__sv2v_reg;
  assign r_28__11_ = r_28__11__sv2v_reg;
  assign r_28__10_ = r_28__10__sv2v_reg;
  assign r_28__9_ = r_28__9__sv2v_reg;
  assign r_28__8_ = r_28__8__sv2v_reg;
  assign r_28__7_ = r_28__7__sv2v_reg;
  assign r_28__6_ = r_28__6__sv2v_reg;
  assign r_28__5_ = r_28__5__sv2v_reg;
  assign r_28__4_ = r_28__4__sv2v_reg;
  assign r_28__3_ = r_28__3__sv2v_reg;
  assign r_28__2_ = r_28__2__sv2v_reg;
  assign r_28__1_ = r_28__1__sv2v_reg;
  assign r_28__0_ = r_28__0__sv2v_reg;
  assign r_29__15_ = r_29__15__sv2v_reg;
  assign r_29__14_ = r_29__14__sv2v_reg;
  assign r_29__13_ = r_29__13__sv2v_reg;
  assign r_29__12_ = r_29__12__sv2v_reg;
  assign r_29__11_ = r_29__11__sv2v_reg;
  assign r_29__10_ = r_29__10__sv2v_reg;
  assign r_29__9_ = r_29__9__sv2v_reg;
  assign r_29__8_ = r_29__8__sv2v_reg;
  assign r_29__7_ = r_29__7__sv2v_reg;
  assign r_29__6_ = r_29__6__sv2v_reg;
  assign r_29__5_ = r_29__5__sv2v_reg;
  assign r_29__4_ = r_29__4__sv2v_reg;
  assign r_29__3_ = r_29__3__sv2v_reg;
  assign r_29__2_ = r_29__2__sv2v_reg;
  assign r_29__1_ = r_29__1__sv2v_reg;
  assign r_29__0_ = r_29__0__sv2v_reg;
  assign r_30__15_ = r_30__15__sv2v_reg;
  assign r_30__14_ = r_30__14__sv2v_reg;
  assign r_30__13_ = r_30__13__sv2v_reg;
  assign r_30__12_ = r_30__12__sv2v_reg;
  assign r_30__11_ = r_30__11__sv2v_reg;
  assign r_30__10_ = r_30__10__sv2v_reg;
  assign r_30__9_ = r_30__9__sv2v_reg;
  assign r_30__8_ = r_30__8__sv2v_reg;
  assign r_30__7_ = r_30__7__sv2v_reg;
  assign r_30__6_ = r_30__6__sv2v_reg;
  assign r_30__5_ = r_30__5__sv2v_reg;
  assign r_30__4_ = r_30__4__sv2v_reg;
  assign r_30__3_ = r_30__3__sv2v_reg;
  assign r_30__2_ = r_30__2__sv2v_reg;
  assign r_30__1_ = r_30__1__sv2v_reg;
  assign r_30__0_ = r_30__0__sv2v_reg;
  assign r_31__15_ = r_31__15__sv2v_reg;
  assign r_31__14_ = r_31__14__sv2v_reg;
  assign r_31__13_ = r_31__13__sv2v_reg;
  assign r_31__12_ = r_31__12__sv2v_reg;
  assign r_31__11_ = r_31__11__sv2v_reg;
  assign r_31__10_ = r_31__10__sv2v_reg;
  assign r_31__9_ = r_31__9__sv2v_reg;
  assign r_31__8_ = r_31__8__sv2v_reg;
  assign r_31__7_ = r_31__7__sv2v_reg;
  assign r_31__6_ = r_31__6__sv2v_reg;
  assign r_31__5_ = r_31__5__sv2v_reg;
  assign r_31__4_ = r_31__4__sv2v_reg;
  assign r_31__3_ = r_31__3__sv2v_reg;
  assign r_31__2_ = r_31__2__sv2v_reg;
  assign r_31__1_ = r_31__1__sv2v_reg;
  assign r_31__0_ = r_31__0__sv2v_reg;
  assign r_32__15_ = r_32__15__sv2v_reg;
  assign r_32__14_ = r_32__14__sv2v_reg;
  assign r_32__13_ = r_32__13__sv2v_reg;
  assign r_32__12_ = r_32__12__sv2v_reg;
  assign r_32__11_ = r_32__11__sv2v_reg;
  assign r_32__10_ = r_32__10__sv2v_reg;
  assign r_32__9_ = r_32__9__sv2v_reg;
  assign r_32__8_ = r_32__8__sv2v_reg;
  assign r_32__7_ = r_32__7__sv2v_reg;
  assign r_32__6_ = r_32__6__sv2v_reg;
  assign r_32__5_ = r_32__5__sv2v_reg;
  assign r_32__4_ = r_32__4__sv2v_reg;
  assign r_32__3_ = r_32__3__sv2v_reg;
  assign r_32__2_ = r_32__2__sv2v_reg;
  assign r_32__1_ = r_32__1__sv2v_reg;
  assign r_32__0_ = r_32__0__sv2v_reg;
  assign r_33__15_ = r_33__15__sv2v_reg;
  assign r_33__14_ = r_33__14__sv2v_reg;
  assign r_33__13_ = r_33__13__sv2v_reg;
  assign r_33__12_ = r_33__12__sv2v_reg;
  assign r_33__11_ = r_33__11__sv2v_reg;
  assign r_33__10_ = r_33__10__sv2v_reg;
  assign r_33__9_ = r_33__9__sv2v_reg;
  assign r_33__8_ = r_33__8__sv2v_reg;
  assign r_33__7_ = r_33__7__sv2v_reg;
  assign r_33__6_ = r_33__6__sv2v_reg;
  assign r_33__5_ = r_33__5__sv2v_reg;
  assign r_33__4_ = r_33__4__sv2v_reg;
  assign r_33__3_ = r_33__3__sv2v_reg;
  assign r_33__2_ = r_33__2__sv2v_reg;
  assign r_33__1_ = r_33__1__sv2v_reg;
  assign r_33__0_ = r_33__0__sv2v_reg;
  assign r_34__15_ = r_34__15__sv2v_reg;
  assign r_34__14_ = r_34__14__sv2v_reg;
  assign r_34__13_ = r_34__13__sv2v_reg;
  assign r_34__12_ = r_34__12__sv2v_reg;
  assign r_34__11_ = r_34__11__sv2v_reg;
  assign r_34__10_ = r_34__10__sv2v_reg;
  assign r_34__9_ = r_34__9__sv2v_reg;
  assign r_34__8_ = r_34__8__sv2v_reg;
  assign r_34__7_ = r_34__7__sv2v_reg;
  assign r_34__6_ = r_34__6__sv2v_reg;
  assign r_34__5_ = r_34__5__sv2v_reg;
  assign r_34__4_ = r_34__4__sv2v_reg;
  assign r_34__3_ = r_34__3__sv2v_reg;
  assign r_34__2_ = r_34__2__sv2v_reg;
  assign r_34__1_ = r_34__1__sv2v_reg;
  assign r_34__0_ = r_34__0__sv2v_reg;
  assign r_35__15_ = r_35__15__sv2v_reg;
  assign r_35__14_ = r_35__14__sv2v_reg;
  assign r_35__13_ = r_35__13__sv2v_reg;
  assign r_35__12_ = r_35__12__sv2v_reg;
  assign r_35__11_ = r_35__11__sv2v_reg;
  assign r_35__10_ = r_35__10__sv2v_reg;
  assign r_35__9_ = r_35__9__sv2v_reg;
  assign r_35__8_ = r_35__8__sv2v_reg;
  assign r_35__7_ = r_35__7__sv2v_reg;
  assign r_35__6_ = r_35__6__sv2v_reg;
  assign r_35__5_ = r_35__5__sv2v_reg;
  assign r_35__4_ = r_35__4__sv2v_reg;
  assign r_35__3_ = r_35__3__sv2v_reg;
  assign r_35__2_ = r_35__2__sv2v_reg;
  assign r_35__1_ = r_35__1__sv2v_reg;
  assign r_35__0_ = r_35__0__sv2v_reg;
  assign r_36__15_ = r_36__15__sv2v_reg;
  assign r_36__14_ = r_36__14__sv2v_reg;
  assign r_36__13_ = r_36__13__sv2v_reg;
  assign r_36__12_ = r_36__12__sv2v_reg;
  assign r_36__11_ = r_36__11__sv2v_reg;
  assign r_36__10_ = r_36__10__sv2v_reg;
  assign r_36__9_ = r_36__9__sv2v_reg;
  assign r_36__8_ = r_36__8__sv2v_reg;
  assign r_36__7_ = r_36__7__sv2v_reg;
  assign r_36__6_ = r_36__6__sv2v_reg;
  assign r_36__5_ = r_36__5__sv2v_reg;
  assign r_36__4_ = r_36__4__sv2v_reg;
  assign r_36__3_ = r_36__3__sv2v_reg;
  assign r_36__2_ = r_36__2__sv2v_reg;
  assign r_36__1_ = r_36__1__sv2v_reg;
  assign r_36__0_ = r_36__0__sv2v_reg;
  assign r_37__15_ = r_37__15__sv2v_reg;
  assign r_37__14_ = r_37__14__sv2v_reg;
  assign r_37__13_ = r_37__13__sv2v_reg;
  assign r_37__12_ = r_37__12__sv2v_reg;
  assign r_37__11_ = r_37__11__sv2v_reg;
  assign r_37__10_ = r_37__10__sv2v_reg;
  assign r_37__9_ = r_37__9__sv2v_reg;
  assign r_37__8_ = r_37__8__sv2v_reg;
  assign r_37__7_ = r_37__7__sv2v_reg;
  assign r_37__6_ = r_37__6__sv2v_reg;
  assign r_37__5_ = r_37__5__sv2v_reg;
  assign r_37__4_ = r_37__4__sv2v_reg;
  assign r_37__3_ = r_37__3__sv2v_reg;
  assign r_37__2_ = r_37__2__sv2v_reg;
  assign r_37__1_ = r_37__1__sv2v_reg;
  assign r_37__0_ = r_37__0__sv2v_reg;
  assign r_38__15_ = r_38__15__sv2v_reg;
  assign r_38__14_ = r_38__14__sv2v_reg;
  assign r_38__13_ = r_38__13__sv2v_reg;
  assign r_38__12_ = r_38__12__sv2v_reg;
  assign r_38__11_ = r_38__11__sv2v_reg;
  assign r_38__10_ = r_38__10__sv2v_reg;
  assign r_38__9_ = r_38__9__sv2v_reg;
  assign r_38__8_ = r_38__8__sv2v_reg;
  assign r_38__7_ = r_38__7__sv2v_reg;
  assign r_38__6_ = r_38__6__sv2v_reg;
  assign r_38__5_ = r_38__5__sv2v_reg;
  assign r_38__4_ = r_38__4__sv2v_reg;
  assign r_38__3_ = r_38__3__sv2v_reg;
  assign r_38__2_ = r_38__2__sv2v_reg;
  assign r_38__1_ = r_38__1__sv2v_reg;
  assign r_38__0_ = r_38__0__sv2v_reg;
  assign r_39__15_ = r_39__15__sv2v_reg;
  assign r_39__14_ = r_39__14__sv2v_reg;
  assign r_39__13_ = r_39__13__sv2v_reg;
  assign r_39__12_ = r_39__12__sv2v_reg;
  assign r_39__11_ = r_39__11__sv2v_reg;
  assign r_39__10_ = r_39__10__sv2v_reg;
  assign r_39__9_ = r_39__9__sv2v_reg;
  assign r_39__8_ = r_39__8__sv2v_reg;
  assign r_39__7_ = r_39__7__sv2v_reg;
  assign r_39__6_ = r_39__6__sv2v_reg;
  assign r_39__5_ = r_39__5__sv2v_reg;
  assign r_39__4_ = r_39__4__sv2v_reg;
  assign r_39__3_ = r_39__3__sv2v_reg;
  assign r_39__2_ = r_39__2__sv2v_reg;
  assign r_39__1_ = r_39__1__sv2v_reg;
  assign r_39__0_ = r_39__0__sv2v_reg;
  assign r_40__15_ = r_40__15__sv2v_reg;
  assign r_40__14_ = r_40__14__sv2v_reg;
  assign r_40__13_ = r_40__13__sv2v_reg;
  assign r_40__12_ = r_40__12__sv2v_reg;
  assign r_40__11_ = r_40__11__sv2v_reg;
  assign r_40__10_ = r_40__10__sv2v_reg;
  assign r_40__9_ = r_40__9__sv2v_reg;
  assign r_40__8_ = r_40__8__sv2v_reg;
  assign r_40__7_ = r_40__7__sv2v_reg;
  assign r_40__6_ = r_40__6__sv2v_reg;
  assign r_40__5_ = r_40__5__sv2v_reg;
  assign r_40__4_ = r_40__4__sv2v_reg;
  assign r_40__3_ = r_40__3__sv2v_reg;
  assign r_40__2_ = r_40__2__sv2v_reg;
  assign r_40__1_ = r_40__1__sv2v_reg;
  assign r_40__0_ = r_40__0__sv2v_reg;
  assign r_41__15_ = r_41__15__sv2v_reg;
  assign r_41__14_ = r_41__14__sv2v_reg;
  assign r_41__13_ = r_41__13__sv2v_reg;
  assign r_41__12_ = r_41__12__sv2v_reg;
  assign r_41__11_ = r_41__11__sv2v_reg;
  assign r_41__10_ = r_41__10__sv2v_reg;
  assign r_41__9_ = r_41__9__sv2v_reg;
  assign r_41__8_ = r_41__8__sv2v_reg;
  assign r_41__7_ = r_41__7__sv2v_reg;
  assign r_41__6_ = r_41__6__sv2v_reg;
  assign r_41__5_ = r_41__5__sv2v_reg;
  assign r_41__4_ = r_41__4__sv2v_reg;
  assign r_41__3_ = r_41__3__sv2v_reg;
  assign r_41__2_ = r_41__2__sv2v_reg;
  assign r_41__1_ = r_41__1__sv2v_reg;
  assign r_41__0_ = r_41__0__sv2v_reg;
  assign r_42__15_ = r_42__15__sv2v_reg;
  assign r_42__14_ = r_42__14__sv2v_reg;
  assign r_42__13_ = r_42__13__sv2v_reg;
  assign r_42__12_ = r_42__12__sv2v_reg;
  assign r_42__11_ = r_42__11__sv2v_reg;
  assign r_42__10_ = r_42__10__sv2v_reg;
  assign r_42__9_ = r_42__9__sv2v_reg;
  assign r_42__8_ = r_42__8__sv2v_reg;
  assign r_42__7_ = r_42__7__sv2v_reg;
  assign r_42__6_ = r_42__6__sv2v_reg;
  assign r_42__5_ = r_42__5__sv2v_reg;
  assign r_42__4_ = r_42__4__sv2v_reg;
  assign r_42__3_ = r_42__3__sv2v_reg;
  assign r_42__2_ = r_42__2__sv2v_reg;
  assign r_42__1_ = r_42__1__sv2v_reg;
  assign r_42__0_ = r_42__0__sv2v_reg;
  assign r_43__15_ = r_43__15__sv2v_reg;
  assign r_43__14_ = r_43__14__sv2v_reg;
  assign r_43__13_ = r_43__13__sv2v_reg;
  assign r_43__12_ = r_43__12__sv2v_reg;
  assign r_43__11_ = r_43__11__sv2v_reg;
  assign r_43__10_ = r_43__10__sv2v_reg;
  assign r_43__9_ = r_43__9__sv2v_reg;
  assign r_43__8_ = r_43__8__sv2v_reg;
  assign r_43__7_ = r_43__7__sv2v_reg;
  assign r_43__6_ = r_43__6__sv2v_reg;
  assign r_43__5_ = r_43__5__sv2v_reg;
  assign r_43__4_ = r_43__4__sv2v_reg;
  assign r_43__3_ = r_43__3__sv2v_reg;
  assign r_43__2_ = r_43__2__sv2v_reg;
  assign r_43__1_ = r_43__1__sv2v_reg;
  assign r_43__0_ = r_43__0__sv2v_reg;
  assign r_44__15_ = r_44__15__sv2v_reg;
  assign r_44__14_ = r_44__14__sv2v_reg;
  assign r_44__13_ = r_44__13__sv2v_reg;
  assign r_44__12_ = r_44__12__sv2v_reg;
  assign r_44__11_ = r_44__11__sv2v_reg;
  assign r_44__10_ = r_44__10__sv2v_reg;
  assign r_44__9_ = r_44__9__sv2v_reg;
  assign r_44__8_ = r_44__8__sv2v_reg;
  assign r_44__7_ = r_44__7__sv2v_reg;
  assign r_44__6_ = r_44__6__sv2v_reg;
  assign r_44__5_ = r_44__5__sv2v_reg;
  assign r_44__4_ = r_44__4__sv2v_reg;
  assign r_44__3_ = r_44__3__sv2v_reg;
  assign r_44__2_ = r_44__2__sv2v_reg;
  assign r_44__1_ = r_44__1__sv2v_reg;
  assign r_44__0_ = r_44__0__sv2v_reg;
  assign r_45__15_ = r_45__15__sv2v_reg;
  assign r_45__14_ = r_45__14__sv2v_reg;
  assign r_45__13_ = r_45__13__sv2v_reg;
  assign r_45__12_ = r_45__12__sv2v_reg;
  assign r_45__11_ = r_45__11__sv2v_reg;
  assign r_45__10_ = r_45__10__sv2v_reg;
  assign r_45__9_ = r_45__9__sv2v_reg;
  assign r_45__8_ = r_45__8__sv2v_reg;
  assign r_45__7_ = r_45__7__sv2v_reg;
  assign r_45__6_ = r_45__6__sv2v_reg;
  assign r_45__5_ = r_45__5__sv2v_reg;
  assign r_45__4_ = r_45__4__sv2v_reg;
  assign r_45__3_ = r_45__3__sv2v_reg;
  assign r_45__2_ = r_45__2__sv2v_reg;
  assign r_45__1_ = r_45__1__sv2v_reg;
  assign r_45__0_ = r_45__0__sv2v_reg;
  assign r_46__15_ = r_46__15__sv2v_reg;
  assign r_46__14_ = r_46__14__sv2v_reg;
  assign r_46__13_ = r_46__13__sv2v_reg;
  assign r_46__12_ = r_46__12__sv2v_reg;
  assign r_46__11_ = r_46__11__sv2v_reg;
  assign r_46__10_ = r_46__10__sv2v_reg;
  assign r_46__9_ = r_46__9__sv2v_reg;
  assign r_46__8_ = r_46__8__sv2v_reg;
  assign r_46__7_ = r_46__7__sv2v_reg;
  assign r_46__6_ = r_46__6__sv2v_reg;
  assign r_46__5_ = r_46__5__sv2v_reg;
  assign r_46__4_ = r_46__4__sv2v_reg;
  assign r_46__3_ = r_46__3__sv2v_reg;
  assign r_46__2_ = r_46__2__sv2v_reg;
  assign r_46__1_ = r_46__1__sv2v_reg;
  assign r_46__0_ = r_46__0__sv2v_reg;
  assign r_47__15_ = r_47__15__sv2v_reg;
  assign r_47__14_ = r_47__14__sv2v_reg;
  assign r_47__13_ = r_47__13__sv2v_reg;
  assign r_47__12_ = r_47__12__sv2v_reg;
  assign r_47__11_ = r_47__11__sv2v_reg;
  assign r_47__10_ = r_47__10__sv2v_reg;
  assign r_47__9_ = r_47__9__sv2v_reg;
  assign r_47__8_ = r_47__8__sv2v_reg;
  assign r_47__7_ = r_47__7__sv2v_reg;
  assign r_47__6_ = r_47__6__sv2v_reg;
  assign r_47__5_ = r_47__5__sv2v_reg;
  assign r_47__4_ = r_47__4__sv2v_reg;
  assign r_47__3_ = r_47__3__sv2v_reg;
  assign r_47__2_ = r_47__2__sv2v_reg;
  assign r_47__1_ = r_47__1__sv2v_reg;
  assign r_47__0_ = r_47__0__sv2v_reg;
  assign r_48__15_ = r_48__15__sv2v_reg;
  assign r_48__14_ = r_48__14__sv2v_reg;
  assign r_48__13_ = r_48__13__sv2v_reg;
  assign r_48__12_ = r_48__12__sv2v_reg;
  assign r_48__11_ = r_48__11__sv2v_reg;
  assign r_48__10_ = r_48__10__sv2v_reg;
  assign r_48__9_ = r_48__9__sv2v_reg;
  assign r_48__8_ = r_48__8__sv2v_reg;
  assign r_48__7_ = r_48__7__sv2v_reg;
  assign r_48__6_ = r_48__6__sv2v_reg;
  assign r_48__5_ = r_48__5__sv2v_reg;
  assign r_48__4_ = r_48__4__sv2v_reg;
  assign r_48__3_ = r_48__3__sv2v_reg;
  assign r_48__2_ = r_48__2__sv2v_reg;
  assign r_48__1_ = r_48__1__sv2v_reg;
  assign r_48__0_ = r_48__0__sv2v_reg;
  assign r_49__15_ = r_49__15__sv2v_reg;
  assign r_49__14_ = r_49__14__sv2v_reg;
  assign r_49__13_ = r_49__13__sv2v_reg;
  assign r_49__12_ = r_49__12__sv2v_reg;
  assign r_49__11_ = r_49__11__sv2v_reg;
  assign r_49__10_ = r_49__10__sv2v_reg;
  assign r_49__9_ = r_49__9__sv2v_reg;
  assign r_49__8_ = r_49__8__sv2v_reg;
  assign r_49__7_ = r_49__7__sv2v_reg;
  assign r_49__6_ = r_49__6__sv2v_reg;
  assign r_49__5_ = r_49__5__sv2v_reg;
  assign r_49__4_ = r_49__4__sv2v_reg;
  assign r_49__3_ = r_49__3__sv2v_reg;
  assign r_49__2_ = r_49__2__sv2v_reg;
  assign r_49__1_ = r_49__1__sv2v_reg;
  assign r_49__0_ = r_49__0__sv2v_reg;
  assign r_50__15_ = r_50__15__sv2v_reg;
  assign r_50__14_ = r_50__14__sv2v_reg;
  assign r_50__13_ = r_50__13__sv2v_reg;
  assign r_50__12_ = r_50__12__sv2v_reg;
  assign r_50__11_ = r_50__11__sv2v_reg;
  assign r_50__10_ = r_50__10__sv2v_reg;
  assign r_50__9_ = r_50__9__sv2v_reg;
  assign r_50__8_ = r_50__8__sv2v_reg;
  assign r_50__7_ = r_50__7__sv2v_reg;
  assign r_50__6_ = r_50__6__sv2v_reg;
  assign r_50__5_ = r_50__5__sv2v_reg;
  assign r_50__4_ = r_50__4__sv2v_reg;
  assign r_50__3_ = r_50__3__sv2v_reg;
  assign r_50__2_ = r_50__2__sv2v_reg;
  assign r_50__1_ = r_50__1__sv2v_reg;
  assign r_50__0_ = r_50__0__sv2v_reg;
  assign r_51__15_ = r_51__15__sv2v_reg;
  assign r_51__14_ = r_51__14__sv2v_reg;
  assign r_51__13_ = r_51__13__sv2v_reg;
  assign r_51__12_ = r_51__12__sv2v_reg;
  assign r_51__11_ = r_51__11__sv2v_reg;
  assign r_51__10_ = r_51__10__sv2v_reg;
  assign r_51__9_ = r_51__9__sv2v_reg;
  assign r_51__8_ = r_51__8__sv2v_reg;
  assign r_51__7_ = r_51__7__sv2v_reg;
  assign r_51__6_ = r_51__6__sv2v_reg;
  assign r_51__5_ = r_51__5__sv2v_reg;
  assign r_51__4_ = r_51__4__sv2v_reg;
  assign r_51__3_ = r_51__3__sv2v_reg;
  assign r_51__2_ = r_51__2__sv2v_reg;
  assign r_51__1_ = r_51__1__sv2v_reg;
  assign r_51__0_ = r_51__0__sv2v_reg;
  assign r_52__15_ = r_52__15__sv2v_reg;
  assign r_52__14_ = r_52__14__sv2v_reg;
  assign r_52__13_ = r_52__13__sv2v_reg;
  assign r_52__12_ = r_52__12__sv2v_reg;
  assign r_52__11_ = r_52__11__sv2v_reg;
  assign r_52__10_ = r_52__10__sv2v_reg;
  assign r_52__9_ = r_52__9__sv2v_reg;
  assign r_52__8_ = r_52__8__sv2v_reg;
  assign r_52__7_ = r_52__7__sv2v_reg;
  assign r_52__6_ = r_52__6__sv2v_reg;
  assign r_52__5_ = r_52__5__sv2v_reg;
  assign r_52__4_ = r_52__4__sv2v_reg;
  assign r_52__3_ = r_52__3__sv2v_reg;
  assign r_52__2_ = r_52__2__sv2v_reg;
  assign r_52__1_ = r_52__1__sv2v_reg;
  assign r_52__0_ = r_52__0__sv2v_reg;
  assign r_53__15_ = r_53__15__sv2v_reg;
  assign r_53__14_ = r_53__14__sv2v_reg;
  assign r_53__13_ = r_53__13__sv2v_reg;
  assign r_53__12_ = r_53__12__sv2v_reg;
  assign r_53__11_ = r_53__11__sv2v_reg;
  assign r_53__10_ = r_53__10__sv2v_reg;
  assign r_53__9_ = r_53__9__sv2v_reg;
  assign r_53__8_ = r_53__8__sv2v_reg;
  assign r_53__7_ = r_53__7__sv2v_reg;
  assign r_53__6_ = r_53__6__sv2v_reg;
  assign r_53__5_ = r_53__5__sv2v_reg;
  assign r_53__4_ = r_53__4__sv2v_reg;
  assign r_53__3_ = r_53__3__sv2v_reg;
  assign r_53__2_ = r_53__2__sv2v_reg;
  assign r_53__1_ = r_53__1__sv2v_reg;
  assign r_53__0_ = r_53__0__sv2v_reg;
  assign r_54__15_ = r_54__15__sv2v_reg;
  assign r_54__14_ = r_54__14__sv2v_reg;
  assign r_54__13_ = r_54__13__sv2v_reg;
  assign r_54__12_ = r_54__12__sv2v_reg;
  assign r_54__11_ = r_54__11__sv2v_reg;
  assign r_54__10_ = r_54__10__sv2v_reg;
  assign r_54__9_ = r_54__9__sv2v_reg;
  assign r_54__8_ = r_54__8__sv2v_reg;
  assign r_54__7_ = r_54__7__sv2v_reg;
  assign r_54__6_ = r_54__6__sv2v_reg;
  assign r_54__5_ = r_54__5__sv2v_reg;
  assign r_54__4_ = r_54__4__sv2v_reg;
  assign r_54__3_ = r_54__3__sv2v_reg;
  assign r_54__2_ = r_54__2__sv2v_reg;
  assign r_54__1_ = r_54__1__sv2v_reg;
  assign r_54__0_ = r_54__0__sv2v_reg;
  assign r_55__15_ = r_55__15__sv2v_reg;
  assign r_55__14_ = r_55__14__sv2v_reg;
  assign r_55__13_ = r_55__13__sv2v_reg;
  assign r_55__12_ = r_55__12__sv2v_reg;
  assign r_55__11_ = r_55__11__sv2v_reg;
  assign r_55__10_ = r_55__10__sv2v_reg;
  assign r_55__9_ = r_55__9__sv2v_reg;
  assign r_55__8_ = r_55__8__sv2v_reg;
  assign r_55__7_ = r_55__7__sv2v_reg;
  assign r_55__6_ = r_55__6__sv2v_reg;
  assign r_55__5_ = r_55__5__sv2v_reg;
  assign r_55__4_ = r_55__4__sv2v_reg;
  assign r_55__3_ = r_55__3__sv2v_reg;
  assign r_55__2_ = r_55__2__sv2v_reg;
  assign r_55__1_ = r_55__1__sv2v_reg;
  assign r_55__0_ = r_55__0__sv2v_reg;
  assign r_56__15_ = r_56__15__sv2v_reg;
  assign r_56__14_ = r_56__14__sv2v_reg;
  assign r_56__13_ = r_56__13__sv2v_reg;
  assign r_56__12_ = r_56__12__sv2v_reg;
  assign r_56__11_ = r_56__11__sv2v_reg;
  assign r_56__10_ = r_56__10__sv2v_reg;
  assign r_56__9_ = r_56__9__sv2v_reg;
  assign r_56__8_ = r_56__8__sv2v_reg;
  assign r_56__7_ = r_56__7__sv2v_reg;
  assign r_56__6_ = r_56__6__sv2v_reg;
  assign r_56__5_ = r_56__5__sv2v_reg;
  assign r_56__4_ = r_56__4__sv2v_reg;
  assign r_56__3_ = r_56__3__sv2v_reg;
  assign r_56__2_ = r_56__2__sv2v_reg;
  assign r_56__1_ = r_56__1__sv2v_reg;
  assign r_56__0_ = r_56__0__sv2v_reg;
  assign r_57__15_ = r_57__15__sv2v_reg;
  assign r_57__14_ = r_57__14__sv2v_reg;
  assign r_57__13_ = r_57__13__sv2v_reg;
  assign r_57__12_ = r_57__12__sv2v_reg;
  assign r_57__11_ = r_57__11__sv2v_reg;
  assign r_57__10_ = r_57__10__sv2v_reg;
  assign r_57__9_ = r_57__9__sv2v_reg;
  assign r_57__8_ = r_57__8__sv2v_reg;
  assign r_57__7_ = r_57__7__sv2v_reg;
  assign r_57__6_ = r_57__6__sv2v_reg;
  assign r_57__5_ = r_57__5__sv2v_reg;
  assign r_57__4_ = r_57__4__sv2v_reg;
  assign r_57__3_ = r_57__3__sv2v_reg;
  assign r_57__2_ = r_57__2__sv2v_reg;
  assign r_57__1_ = r_57__1__sv2v_reg;
  assign r_57__0_ = r_57__0__sv2v_reg;
  assign r_58__15_ = r_58__15__sv2v_reg;
  assign r_58__14_ = r_58__14__sv2v_reg;
  assign r_58__13_ = r_58__13__sv2v_reg;
  assign r_58__12_ = r_58__12__sv2v_reg;
  assign r_58__11_ = r_58__11__sv2v_reg;
  assign r_58__10_ = r_58__10__sv2v_reg;
  assign r_58__9_ = r_58__9__sv2v_reg;
  assign r_58__8_ = r_58__8__sv2v_reg;
  assign r_58__7_ = r_58__7__sv2v_reg;
  assign r_58__6_ = r_58__6__sv2v_reg;
  assign r_58__5_ = r_58__5__sv2v_reg;
  assign r_58__4_ = r_58__4__sv2v_reg;
  assign r_58__3_ = r_58__3__sv2v_reg;
  assign r_58__2_ = r_58__2__sv2v_reg;
  assign r_58__1_ = r_58__1__sv2v_reg;
  assign r_58__0_ = r_58__0__sv2v_reg;
  assign r_59__15_ = r_59__15__sv2v_reg;
  assign r_59__14_ = r_59__14__sv2v_reg;
  assign r_59__13_ = r_59__13__sv2v_reg;
  assign r_59__12_ = r_59__12__sv2v_reg;
  assign r_59__11_ = r_59__11__sv2v_reg;
  assign r_59__10_ = r_59__10__sv2v_reg;
  assign r_59__9_ = r_59__9__sv2v_reg;
  assign r_59__8_ = r_59__8__sv2v_reg;
  assign r_59__7_ = r_59__7__sv2v_reg;
  assign r_59__6_ = r_59__6__sv2v_reg;
  assign r_59__5_ = r_59__5__sv2v_reg;
  assign r_59__4_ = r_59__4__sv2v_reg;
  assign r_59__3_ = r_59__3__sv2v_reg;
  assign r_59__2_ = r_59__2__sv2v_reg;
  assign r_59__1_ = r_59__1__sv2v_reg;
  assign r_59__0_ = r_59__0__sv2v_reg;
  assign r_60__15_ = r_60__15__sv2v_reg;
  assign r_60__14_ = r_60__14__sv2v_reg;
  assign r_60__13_ = r_60__13__sv2v_reg;
  assign r_60__12_ = r_60__12__sv2v_reg;
  assign r_60__11_ = r_60__11__sv2v_reg;
  assign r_60__10_ = r_60__10__sv2v_reg;
  assign r_60__9_ = r_60__9__sv2v_reg;
  assign r_60__8_ = r_60__8__sv2v_reg;
  assign r_60__7_ = r_60__7__sv2v_reg;
  assign r_60__6_ = r_60__6__sv2v_reg;
  assign r_60__5_ = r_60__5__sv2v_reg;
  assign r_60__4_ = r_60__4__sv2v_reg;
  assign r_60__3_ = r_60__3__sv2v_reg;
  assign r_60__2_ = r_60__2__sv2v_reg;
  assign r_60__1_ = r_60__1__sv2v_reg;
  assign r_60__0_ = r_60__0__sv2v_reg;
  assign r_61__15_ = r_61__15__sv2v_reg;
  assign r_61__14_ = r_61__14__sv2v_reg;
  assign r_61__13_ = r_61__13__sv2v_reg;
  assign r_61__12_ = r_61__12__sv2v_reg;
  assign r_61__11_ = r_61__11__sv2v_reg;
  assign r_61__10_ = r_61__10__sv2v_reg;
  assign r_61__9_ = r_61__9__sv2v_reg;
  assign r_61__8_ = r_61__8__sv2v_reg;
  assign r_61__7_ = r_61__7__sv2v_reg;
  assign r_61__6_ = r_61__6__sv2v_reg;
  assign r_61__5_ = r_61__5__sv2v_reg;
  assign r_61__4_ = r_61__4__sv2v_reg;
  assign r_61__3_ = r_61__3__sv2v_reg;
  assign r_61__2_ = r_61__2__sv2v_reg;
  assign r_61__1_ = r_61__1__sv2v_reg;
  assign r_61__0_ = r_61__0__sv2v_reg;
  assign r_62__15_ = r_62__15__sv2v_reg;
  assign r_62__14_ = r_62__14__sv2v_reg;
  assign r_62__13_ = r_62__13__sv2v_reg;
  assign r_62__12_ = r_62__12__sv2v_reg;
  assign r_62__11_ = r_62__11__sv2v_reg;
  assign r_62__10_ = r_62__10__sv2v_reg;
  assign r_62__9_ = r_62__9__sv2v_reg;
  assign r_62__8_ = r_62__8__sv2v_reg;
  assign r_62__7_ = r_62__7__sv2v_reg;
  assign r_62__6_ = r_62__6__sv2v_reg;
  assign r_62__5_ = r_62__5__sv2v_reg;
  assign r_62__4_ = r_62__4__sv2v_reg;
  assign r_62__3_ = r_62__3__sv2v_reg;
  assign r_62__2_ = r_62__2__sv2v_reg;
  assign r_62__1_ = r_62__1__sv2v_reg;
  assign r_62__0_ = r_62__0__sv2v_reg;
  assign r_63__15_ = r_63__15__sv2v_reg;
  assign r_63__14_ = r_63__14__sv2v_reg;
  assign r_63__13_ = r_63__13__sv2v_reg;
  assign r_63__12_ = r_63__12__sv2v_reg;
  assign r_63__11_ = r_63__11__sv2v_reg;
  assign r_63__10_ = r_63__10__sv2v_reg;
  assign r_63__9_ = r_63__9__sv2v_reg;
  assign r_63__8_ = r_63__8__sv2v_reg;
  assign r_63__7_ = r_63__7__sv2v_reg;
  assign r_63__6_ = r_63__6__sv2v_reg;
  assign r_63__5_ = r_63__5__sv2v_reg;
  assign r_63__4_ = r_63__4__sv2v_reg;
  assign r_63__3_ = r_63__3__sv2v_reg;
  assign r_63__2_ = r_63__2__sv2v_reg;
  assign r_63__1_ = r_63__1__sv2v_reg;
  assign r_63__0_ = r_63__0__sv2v_reg;
  assign N126 = sel_i[1] & sel_i[0];
  assign N128 = N127 & N130;
  assign N131 = sel_i[3] & sel_i[2];
  assign N133 = N132 & N135;
  assign N136 = sel_i[5] & sel_i[4];
  assign N138 = N137 & N140;
  assign N141 = sel_i[7] & sel_i[6];
  assign N143 = N142 & N145;
  assign N146 = sel_i[9] & sel_i[8];
  assign N148 = N147 & N150;
  assign N151 = sel_i[11] & sel_i[10];
  assign N153 = N152 & N155;
  assign N156 = sel_i[13] & sel_i[12];
  assign N158 = N157 & N160;
  assign N161 = sel_i[15] & sel_i[14];
  assign N163 = N162 & N165;
  assign N166 = sel_i[17] & sel_i[16];
  assign N168 = N167 & N170;
  assign N171 = sel_i[19] & sel_i[18];
  assign N173 = N172 & N175;
  assign N176 = sel_i[21] & sel_i[20];
  assign N178 = N177 & N180;
  assign N181 = sel_i[23] & sel_i[22];
  assign N183 = N182 & N185;
  assign N186 = sel_i[25] & sel_i[24];
  assign N188 = N187 & N190;
  assign N191 = sel_i[27] & sel_i[26];
  assign N193 = N192 & N195;
  assign N196 = sel_i[29] & sel_i[28];
  assign N198 = N197 & N200;
  assign N201 = sel_i[31] & sel_i[30];
  assign N203 = N202 & N205;
  assign N206 = sel_i[33] & sel_i[32];
  assign N208 = N207 & N210;
  assign N211 = sel_i[35] & sel_i[34];
  assign N213 = N212 & N215;
  assign N216 = sel_i[37] & sel_i[36];
  assign N218 = N217 & N220;
  assign N221 = sel_i[39] & sel_i[38];
  assign N223 = N222 & N225;
  assign N226 = sel_i[41] & sel_i[40];
  assign N228 = N227 & N230;
  assign N231 = sel_i[43] & sel_i[42];
  assign N233 = N232 & N235;
  assign N236 = sel_i[45] & sel_i[44];
  assign N238 = N237 & N240;
  assign N241 = sel_i[47] & sel_i[46];
  assign N243 = N242 & N245;
  assign N246 = sel_i[49] & sel_i[48];
  assign N248 = N247 & N250;
  assign N251 = sel_i[51] & sel_i[50];
  assign N253 = N252 & N255;
  assign N256 = sel_i[53] & sel_i[52];
  assign N258 = N257 & N260;
  assign N261 = sel_i[55] & sel_i[54];
  assign N263 = N262 & N265;
  assign N266 = sel_i[57] & sel_i[56];
  assign N268 = N267 & N270;
  assign N271 = sel_i[59] & sel_i[58];
  assign N273 = N272 & N275;
  assign N276 = sel_i[61] & sel_i[60];
  assign N278 = N277 & N280;
  assign N281 = sel_i[63] & sel_i[62];
  assign N283 = N282 & N285;
  assign N286 = sel_i[65] & sel_i[64];
  assign N288 = N287 & N290;
  assign N291 = sel_i[67] & sel_i[66];
  assign N293 = N292 & N295;
  assign N296 = sel_i[69] & sel_i[68];
  assign N298 = N297 & N300;
  assign N301 = sel_i[71] & sel_i[70];
  assign N303 = N302 & N305;
  assign N306 = sel_i[73] & sel_i[72];
  assign N308 = N307 & N310;
  assign N311 = sel_i[75] & sel_i[74];
  assign N313 = N312 & N315;
  assign N316 = sel_i[77] & sel_i[76];
  assign N318 = N317 & N320;
  assign N321 = sel_i[79] & sel_i[78];
  assign N323 = N322 & N325;
  assign N326 = sel_i[81] & sel_i[80];
  assign N328 = N327 & N330;
  assign N331 = sel_i[83] & sel_i[82];
  assign N333 = N332 & N335;
  assign N336 = sel_i[85] & sel_i[84];
  assign N338 = N337 & N340;
  assign N341 = sel_i[87] & sel_i[86];
  assign N343 = N342 & N345;
  assign N346 = sel_i[89] & sel_i[88];
  assign N348 = N347 & N350;
  assign N351 = sel_i[91] & sel_i[90];
  assign N353 = N352 & N355;
  assign N356 = sel_i[93] & sel_i[92];
  assign N358 = N357 & N360;
  assign N361 = sel_i[95] & sel_i[94];
  assign N363 = N362 & N365;
  assign N366 = sel_i[97] & sel_i[96];
  assign N368 = N367 & N370;
  assign N371 = sel_i[99] & sel_i[98];
  assign N373 = N372 & N375;
  assign N376 = sel_i[101] & sel_i[100];
  assign N378 = N377 & N380;
  assign N381 = sel_i[103] & sel_i[102];
  assign N383 = N382 & N385;
  assign N386 = sel_i[105] & sel_i[104];
  assign N388 = N387 & N390;
  assign N391 = sel_i[107] & sel_i[106];
  assign N393 = N392 & N395;
  assign N396 = sel_i[109] & sel_i[108];
  assign N398 = N397 & N400;
  assign N401 = sel_i[111] & sel_i[110];
  assign N403 = N402 & N405;
  assign N406 = sel_i[113] & sel_i[112];
  assign N408 = N407 & N410;
  assign N411 = sel_i[115] & sel_i[114];
  assign N413 = N412 & N415;
  assign N416 = sel_i[117] & sel_i[116];
  assign N418 = N417 & N420;
  assign N421 = sel_i[119] & sel_i[118];
  assign N423 = N422 & N425;
  assign N426 = sel_i[121] & sel_i[120];
  assign N428 = N427 & N430;
  assign N431 = sel_i[123] & sel_i[122];
  assign N433 = N432 & N435;
  assign N436 = sel_i[125] & sel_i[124];
  assign N438 = N437 & N440;
  assign N442 = sel_i[127] | N441;
  assign N444 = sel_i[127] & sel_i[126];
  assign N446 = N445 & N441;
  assign N130 = ~sel_i[0];
  assign N135 = ~sel_i[2];
  assign N140 = ~sel_i[4];
  assign N145 = ~sel_i[6];
  assign N150 = ~sel_i[8];
  assign N155 = ~sel_i[10];
  assign N160 = ~sel_i[12];
  assign N165 = ~sel_i[14];
  assign N170 = ~sel_i[16];
  assign N175 = ~sel_i[18];
  assign N180 = ~sel_i[20];
  assign N185 = ~sel_i[22];
  assign N190 = ~sel_i[24];
  assign N195 = ~sel_i[26];
  assign N200 = ~sel_i[28];
  assign N205 = ~sel_i[30];
  assign N210 = ~sel_i[32];
  assign N215 = ~sel_i[34];
  assign N220 = ~sel_i[36];
  assign N225 = ~sel_i[38];
  assign N230 = ~sel_i[40];
  assign N235 = ~sel_i[42];
  assign N240 = ~sel_i[44];
  assign N245 = ~sel_i[46];
  assign N250 = ~sel_i[48];
  assign N255 = ~sel_i[50];
  assign N260 = ~sel_i[52];
  assign N265 = ~sel_i[54];
  assign N270 = ~sel_i[56];
  assign N275 = ~sel_i[58];
  assign N280 = ~sel_i[60];
  assign N285 = ~sel_i[62];
  assign N290 = ~sel_i[64];
  assign N295 = ~sel_i[66];
  assign N300 = ~sel_i[68];
  assign N305 = ~sel_i[70];
  assign N310 = ~sel_i[72];
  assign N315 = ~sel_i[74];
  assign N320 = ~sel_i[76];
  assign N325 = ~sel_i[78];
  assign N330 = ~sel_i[80];
  assign N335 = ~sel_i[82];
  assign N340 = ~sel_i[84];
  assign N345 = ~sel_i[86];
  assign N350 = ~sel_i[88];
  assign N355 = ~sel_i[90];
  assign N360 = ~sel_i[92];
  assign N365 = ~sel_i[94];
  assign N370 = ~sel_i[96];
  assign N375 = ~sel_i[98];
  assign N380 = ~sel_i[100];
  assign N385 = ~sel_i[102];
  assign N390 = ~sel_i[104];
  assign N395 = ~sel_i[106];
  assign N400 = ~sel_i[108];
  assign N405 = ~sel_i[110];
  assign N410 = ~sel_i[112];
  assign N415 = ~sel_i[114];
  assign N420 = ~sel_i[116];
  assign N425 = ~sel_i[118];
  assign N430 = ~sel_i[120];
  assign N435 = ~sel_i[122];
  assign N440 = ~sel_i[124];
  assign { r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ } = (N0)? { r_1__15_, r_1__14_, r_1__13_, r_1__12_, r_1__11_, r_1__10_, r_1__9_, r_1__8_, r_1__7_, r_1__6_, r_1__5_, r_1__4_, r_1__3_, r_1__2_, r_1__1_, r_1__0_ } : 
                                                                                                                                                                                                    (N1)? data_i : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = N130;
  assign { r_n_1__15_, r_n_1__14_, r_n_1__13_, r_n_1__12_, r_n_1__11_, r_n_1__10_, r_n_1__9_, r_n_1__8_, r_n_1__7_, r_n_1__6_, r_n_1__5_, r_n_1__4_, r_n_1__3_, r_n_1__2_, r_n_1__1_, r_n_1__0_ } = (N2)? { r_2__15_, r_2__14_, r_2__13_, r_2__12_, r_2__11_, r_2__10_, r_2__9_, r_2__8_, r_2__7_, r_2__6_, r_2__5_, r_2__4_, r_2__3_, r_2__2_, r_2__1_, r_2__0_ } : 
                                                                                                                                                                                                    (N3)? data_i : 1'b0;
  assign N2 = sel_i[2];
  assign N3 = N135;
  assign { r_n_2__15_, r_n_2__14_, r_n_2__13_, r_n_2__12_, r_n_2__11_, r_n_2__10_, r_n_2__9_, r_n_2__8_, r_n_2__7_, r_n_2__6_, r_n_2__5_, r_n_2__4_, r_n_2__3_, r_n_2__2_, r_n_2__1_, r_n_2__0_ } = (N4)? { r_3__15_, r_3__14_, r_3__13_, r_3__12_, r_3__11_, r_3__10_, r_3__9_, r_3__8_, r_3__7_, r_3__6_, r_3__5_, r_3__4_, r_3__3_, r_3__2_, r_3__1_, r_3__0_ } : 
                                                                                                                                                                                                    (N5)? data_i : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = N140;
  assign { r_n_3__15_, r_n_3__14_, r_n_3__13_, r_n_3__12_, r_n_3__11_, r_n_3__10_, r_n_3__9_, r_n_3__8_, r_n_3__7_, r_n_3__6_, r_n_3__5_, r_n_3__4_, r_n_3__3_, r_n_3__2_, r_n_3__1_, r_n_3__0_ } = (N6)? { r_4__15_, r_4__14_, r_4__13_, r_4__12_, r_4__11_, r_4__10_, r_4__9_, r_4__8_, r_4__7_, r_4__6_, r_4__5_, r_4__4_, r_4__3_, r_4__2_, r_4__1_, r_4__0_ } : 
                                                                                                                                                                                                    (N7)? data_i : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = N145;
  assign { r_n_4__15_, r_n_4__14_, r_n_4__13_, r_n_4__12_, r_n_4__11_, r_n_4__10_, r_n_4__9_, r_n_4__8_, r_n_4__7_, r_n_4__6_, r_n_4__5_, r_n_4__4_, r_n_4__3_, r_n_4__2_, r_n_4__1_, r_n_4__0_ } = (N8)? { r_5__15_, r_5__14_, r_5__13_, r_5__12_, r_5__11_, r_5__10_, r_5__9_, r_5__8_, r_5__7_, r_5__6_, r_5__5_, r_5__4_, r_5__3_, r_5__2_, r_5__1_, r_5__0_ } : 
                                                                                                                                                                                                    (N9)? data_i : 1'b0;
  assign N8 = sel_i[8];
  assign N9 = N150;
  assign { r_n_5__15_, r_n_5__14_, r_n_5__13_, r_n_5__12_, r_n_5__11_, r_n_5__10_, r_n_5__9_, r_n_5__8_, r_n_5__7_, r_n_5__6_, r_n_5__5_, r_n_5__4_, r_n_5__3_, r_n_5__2_, r_n_5__1_, r_n_5__0_ } = (N10)? { r_6__15_, r_6__14_, r_6__13_, r_6__12_, r_6__11_, r_6__10_, r_6__9_, r_6__8_, r_6__7_, r_6__6_, r_6__5_, r_6__4_, r_6__3_, r_6__2_, r_6__1_, r_6__0_ } : 
                                                                                                                                                                                                    (N11)? data_i : 1'b0;
  assign N10 = sel_i[10];
  assign N11 = N155;
  assign { r_n_6__15_, r_n_6__14_, r_n_6__13_, r_n_6__12_, r_n_6__11_, r_n_6__10_, r_n_6__9_, r_n_6__8_, r_n_6__7_, r_n_6__6_, r_n_6__5_, r_n_6__4_, r_n_6__3_, r_n_6__2_, r_n_6__1_, r_n_6__0_ } = (N12)? { r_7__15_, r_7__14_, r_7__13_, r_7__12_, r_7__11_, r_7__10_, r_7__9_, r_7__8_, r_7__7_, r_7__6_, r_7__5_, r_7__4_, r_7__3_, r_7__2_, r_7__1_, r_7__0_ } : 
                                                                                                                                                                                                    (N13)? data_i : 1'b0;
  assign N12 = sel_i[12];
  assign N13 = N160;
  assign { r_n_7__15_, r_n_7__14_, r_n_7__13_, r_n_7__12_, r_n_7__11_, r_n_7__10_, r_n_7__9_, r_n_7__8_, r_n_7__7_, r_n_7__6_, r_n_7__5_, r_n_7__4_, r_n_7__3_, r_n_7__2_, r_n_7__1_, r_n_7__0_ } = (N14)? { r_8__15_, r_8__14_, r_8__13_, r_8__12_, r_8__11_, r_8__10_, r_8__9_, r_8__8_, r_8__7_, r_8__6_, r_8__5_, r_8__4_, r_8__3_, r_8__2_, r_8__1_, r_8__0_ } : 
                                                                                                                                                                                                    (N15)? data_i : 1'b0;
  assign N14 = sel_i[14];
  assign N15 = N165;
  assign { r_n_8__15_, r_n_8__14_, r_n_8__13_, r_n_8__12_, r_n_8__11_, r_n_8__10_, r_n_8__9_, r_n_8__8_, r_n_8__7_, r_n_8__6_, r_n_8__5_, r_n_8__4_, r_n_8__3_, r_n_8__2_, r_n_8__1_, r_n_8__0_ } = (N16)? { r_9__15_, r_9__14_, r_9__13_, r_9__12_, r_9__11_, r_9__10_, r_9__9_, r_9__8_, r_9__7_, r_9__6_, r_9__5_, r_9__4_, r_9__3_, r_9__2_, r_9__1_, r_9__0_ } : 
                                                                                                                                                                                                    (N17)? data_i : 1'b0;
  assign N16 = sel_i[16];
  assign N17 = N170;
  assign { r_n_9__15_, r_n_9__14_, r_n_9__13_, r_n_9__12_, r_n_9__11_, r_n_9__10_, r_n_9__9_, r_n_9__8_, r_n_9__7_, r_n_9__6_, r_n_9__5_, r_n_9__4_, r_n_9__3_, r_n_9__2_, r_n_9__1_, r_n_9__0_ } = (N18)? { r_10__15_, r_10__14_, r_10__13_, r_10__12_, r_10__11_, r_10__10_, r_10__9_, r_10__8_, r_10__7_, r_10__6_, r_10__5_, r_10__4_, r_10__3_, r_10__2_, r_10__1_, r_10__0_ } : 
                                                                                                                                                                                                    (N19)? data_i : 1'b0;
  assign N18 = sel_i[18];
  assign N19 = N175;
  assign { r_n_10__15_, r_n_10__14_, r_n_10__13_, r_n_10__12_, r_n_10__11_, r_n_10__10_, r_n_10__9_, r_n_10__8_, r_n_10__7_, r_n_10__6_, r_n_10__5_, r_n_10__4_, r_n_10__3_, r_n_10__2_, r_n_10__1_, r_n_10__0_ } = (N20)? { r_11__15_, r_11__14_, r_11__13_, r_11__12_, r_11__11_, r_11__10_, r_11__9_, r_11__8_, r_11__7_, r_11__6_, r_11__5_, r_11__4_, r_11__3_, r_11__2_, r_11__1_, r_11__0_ } : 
                                                                                                                                                                                                                    (N21)? data_i : 1'b0;
  assign N20 = sel_i[20];
  assign N21 = N180;
  assign { r_n_11__15_, r_n_11__14_, r_n_11__13_, r_n_11__12_, r_n_11__11_, r_n_11__10_, r_n_11__9_, r_n_11__8_, r_n_11__7_, r_n_11__6_, r_n_11__5_, r_n_11__4_, r_n_11__3_, r_n_11__2_, r_n_11__1_, r_n_11__0_ } = (N22)? { r_12__15_, r_12__14_, r_12__13_, r_12__12_, r_12__11_, r_12__10_, r_12__9_, r_12__8_, r_12__7_, r_12__6_, r_12__5_, r_12__4_, r_12__3_, r_12__2_, r_12__1_, r_12__0_ } : 
                                                                                                                                                                                                                    (N23)? data_i : 1'b0;
  assign N22 = sel_i[22];
  assign N23 = N185;
  assign { r_n_12__15_, r_n_12__14_, r_n_12__13_, r_n_12__12_, r_n_12__11_, r_n_12__10_, r_n_12__9_, r_n_12__8_, r_n_12__7_, r_n_12__6_, r_n_12__5_, r_n_12__4_, r_n_12__3_, r_n_12__2_, r_n_12__1_, r_n_12__0_ } = (N24)? { r_13__15_, r_13__14_, r_13__13_, r_13__12_, r_13__11_, r_13__10_, r_13__9_, r_13__8_, r_13__7_, r_13__6_, r_13__5_, r_13__4_, r_13__3_, r_13__2_, r_13__1_, r_13__0_ } : 
                                                                                                                                                                                                                    (N25)? data_i : 1'b0;
  assign N24 = sel_i[24];
  assign N25 = N190;
  assign { r_n_13__15_, r_n_13__14_, r_n_13__13_, r_n_13__12_, r_n_13__11_, r_n_13__10_, r_n_13__9_, r_n_13__8_, r_n_13__7_, r_n_13__6_, r_n_13__5_, r_n_13__4_, r_n_13__3_, r_n_13__2_, r_n_13__1_, r_n_13__0_ } = (N26)? { r_14__15_, r_14__14_, r_14__13_, r_14__12_, r_14__11_, r_14__10_, r_14__9_, r_14__8_, r_14__7_, r_14__6_, r_14__5_, r_14__4_, r_14__3_, r_14__2_, r_14__1_, r_14__0_ } : 
                                                                                                                                                                                                                    (N27)? data_i : 1'b0;
  assign N26 = sel_i[26];
  assign N27 = N195;
  assign { r_n_14__15_, r_n_14__14_, r_n_14__13_, r_n_14__12_, r_n_14__11_, r_n_14__10_, r_n_14__9_, r_n_14__8_, r_n_14__7_, r_n_14__6_, r_n_14__5_, r_n_14__4_, r_n_14__3_, r_n_14__2_, r_n_14__1_, r_n_14__0_ } = (N28)? { r_15__15_, r_15__14_, r_15__13_, r_15__12_, r_15__11_, r_15__10_, r_15__9_, r_15__8_, r_15__7_, r_15__6_, r_15__5_, r_15__4_, r_15__3_, r_15__2_, r_15__1_, r_15__0_ } : 
                                                                                                                                                                                                                    (N29)? data_i : 1'b0;
  assign N28 = sel_i[28];
  assign N29 = N200;
  assign { r_n_15__15_, r_n_15__14_, r_n_15__13_, r_n_15__12_, r_n_15__11_, r_n_15__10_, r_n_15__9_, r_n_15__8_, r_n_15__7_, r_n_15__6_, r_n_15__5_, r_n_15__4_, r_n_15__3_, r_n_15__2_, r_n_15__1_, r_n_15__0_ } = (N30)? { r_16__15_, r_16__14_, r_16__13_, r_16__12_, r_16__11_, r_16__10_, r_16__9_, r_16__8_, r_16__7_, r_16__6_, r_16__5_, r_16__4_, r_16__3_, r_16__2_, r_16__1_, r_16__0_ } : 
                                                                                                                                                                                                                    (N31)? data_i : 1'b0;
  assign N30 = sel_i[30];
  assign N31 = N205;
  assign { r_n_16__15_, r_n_16__14_, r_n_16__13_, r_n_16__12_, r_n_16__11_, r_n_16__10_, r_n_16__9_, r_n_16__8_, r_n_16__7_, r_n_16__6_, r_n_16__5_, r_n_16__4_, r_n_16__3_, r_n_16__2_, r_n_16__1_, r_n_16__0_ } = (N32)? { r_17__15_, r_17__14_, r_17__13_, r_17__12_, r_17__11_, r_17__10_, r_17__9_, r_17__8_, r_17__7_, r_17__6_, r_17__5_, r_17__4_, r_17__3_, r_17__2_, r_17__1_, r_17__0_ } : 
                                                                                                                                                                                                                    (N33)? data_i : 1'b0;
  assign N32 = sel_i[32];
  assign N33 = N210;
  assign { r_n_17__15_, r_n_17__14_, r_n_17__13_, r_n_17__12_, r_n_17__11_, r_n_17__10_, r_n_17__9_, r_n_17__8_, r_n_17__7_, r_n_17__6_, r_n_17__5_, r_n_17__4_, r_n_17__3_, r_n_17__2_, r_n_17__1_, r_n_17__0_ } = (N34)? { r_18__15_, r_18__14_, r_18__13_, r_18__12_, r_18__11_, r_18__10_, r_18__9_, r_18__8_, r_18__7_, r_18__6_, r_18__5_, r_18__4_, r_18__3_, r_18__2_, r_18__1_, r_18__0_ } : 
                                                                                                                                                                                                                    (N35)? data_i : 1'b0;
  assign N34 = sel_i[34];
  assign N35 = N215;
  assign { r_n_18__15_, r_n_18__14_, r_n_18__13_, r_n_18__12_, r_n_18__11_, r_n_18__10_, r_n_18__9_, r_n_18__8_, r_n_18__7_, r_n_18__6_, r_n_18__5_, r_n_18__4_, r_n_18__3_, r_n_18__2_, r_n_18__1_, r_n_18__0_ } = (N36)? { r_19__15_, r_19__14_, r_19__13_, r_19__12_, r_19__11_, r_19__10_, r_19__9_, r_19__8_, r_19__7_, r_19__6_, r_19__5_, r_19__4_, r_19__3_, r_19__2_, r_19__1_, r_19__0_ } : 
                                                                                                                                                                                                                    (N37)? data_i : 1'b0;
  assign N36 = sel_i[36];
  assign N37 = N220;
  assign { r_n_19__15_, r_n_19__14_, r_n_19__13_, r_n_19__12_, r_n_19__11_, r_n_19__10_, r_n_19__9_, r_n_19__8_, r_n_19__7_, r_n_19__6_, r_n_19__5_, r_n_19__4_, r_n_19__3_, r_n_19__2_, r_n_19__1_, r_n_19__0_ } = (N38)? { r_20__15_, r_20__14_, r_20__13_, r_20__12_, r_20__11_, r_20__10_, r_20__9_, r_20__8_, r_20__7_, r_20__6_, r_20__5_, r_20__4_, r_20__3_, r_20__2_, r_20__1_, r_20__0_ } : 
                                                                                                                                                                                                                    (N39)? data_i : 1'b0;
  assign N38 = sel_i[38];
  assign N39 = N225;
  assign { r_n_20__15_, r_n_20__14_, r_n_20__13_, r_n_20__12_, r_n_20__11_, r_n_20__10_, r_n_20__9_, r_n_20__8_, r_n_20__7_, r_n_20__6_, r_n_20__5_, r_n_20__4_, r_n_20__3_, r_n_20__2_, r_n_20__1_, r_n_20__0_ } = (N40)? { r_21__15_, r_21__14_, r_21__13_, r_21__12_, r_21__11_, r_21__10_, r_21__9_, r_21__8_, r_21__7_, r_21__6_, r_21__5_, r_21__4_, r_21__3_, r_21__2_, r_21__1_, r_21__0_ } : 
                                                                                                                                                                                                                    (N41)? data_i : 1'b0;
  assign N40 = sel_i[40];
  assign N41 = N230;
  assign { r_n_21__15_, r_n_21__14_, r_n_21__13_, r_n_21__12_, r_n_21__11_, r_n_21__10_, r_n_21__9_, r_n_21__8_, r_n_21__7_, r_n_21__6_, r_n_21__5_, r_n_21__4_, r_n_21__3_, r_n_21__2_, r_n_21__1_, r_n_21__0_ } = (N42)? { r_22__15_, r_22__14_, r_22__13_, r_22__12_, r_22__11_, r_22__10_, r_22__9_, r_22__8_, r_22__7_, r_22__6_, r_22__5_, r_22__4_, r_22__3_, r_22__2_, r_22__1_, r_22__0_ } : 
                                                                                                                                                                                                                    (N43)? data_i : 1'b0;
  assign N42 = sel_i[42];
  assign N43 = N235;
  assign { r_n_22__15_, r_n_22__14_, r_n_22__13_, r_n_22__12_, r_n_22__11_, r_n_22__10_, r_n_22__9_, r_n_22__8_, r_n_22__7_, r_n_22__6_, r_n_22__5_, r_n_22__4_, r_n_22__3_, r_n_22__2_, r_n_22__1_, r_n_22__0_ } = (N44)? { r_23__15_, r_23__14_, r_23__13_, r_23__12_, r_23__11_, r_23__10_, r_23__9_, r_23__8_, r_23__7_, r_23__6_, r_23__5_, r_23__4_, r_23__3_, r_23__2_, r_23__1_, r_23__0_ } : 
                                                                                                                                                                                                                    (N45)? data_i : 1'b0;
  assign N44 = sel_i[44];
  assign N45 = N240;
  assign { r_n_23__15_, r_n_23__14_, r_n_23__13_, r_n_23__12_, r_n_23__11_, r_n_23__10_, r_n_23__9_, r_n_23__8_, r_n_23__7_, r_n_23__6_, r_n_23__5_, r_n_23__4_, r_n_23__3_, r_n_23__2_, r_n_23__1_, r_n_23__0_ } = (N46)? { r_24__15_, r_24__14_, r_24__13_, r_24__12_, r_24__11_, r_24__10_, r_24__9_, r_24__8_, r_24__7_, r_24__6_, r_24__5_, r_24__4_, r_24__3_, r_24__2_, r_24__1_, r_24__0_ } : 
                                                                                                                                                                                                                    (N47)? data_i : 1'b0;
  assign N46 = sel_i[46];
  assign N47 = N245;
  assign { r_n_24__15_, r_n_24__14_, r_n_24__13_, r_n_24__12_, r_n_24__11_, r_n_24__10_, r_n_24__9_, r_n_24__8_, r_n_24__7_, r_n_24__6_, r_n_24__5_, r_n_24__4_, r_n_24__3_, r_n_24__2_, r_n_24__1_, r_n_24__0_ } = (N48)? { r_25__15_, r_25__14_, r_25__13_, r_25__12_, r_25__11_, r_25__10_, r_25__9_, r_25__8_, r_25__7_, r_25__6_, r_25__5_, r_25__4_, r_25__3_, r_25__2_, r_25__1_, r_25__0_ } : 
                                                                                                                                                                                                                    (N49)? data_i : 1'b0;
  assign N48 = sel_i[48];
  assign N49 = N250;
  assign { r_n_25__15_, r_n_25__14_, r_n_25__13_, r_n_25__12_, r_n_25__11_, r_n_25__10_, r_n_25__9_, r_n_25__8_, r_n_25__7_, r_n_25__6_, r_n_25__5_, r_n_25__4_, r_n_25__3_, r_n_25__2_, r_n_25__1_, r_n_25__0_ } = (N50)? { r_26__15_, r_26__14_, r_26__13_, r_26__12_, r_26__11_, r_26__10_, r_26__9_, r_26__8_, r_26__7_, r_26__6_, r_26__5_, r_26__4_, r_26__3_, r_26__2_, r_26__1_, r_26__0_ } : 
                                                                                                                                                                                                                    (N51)? data_i : 1'b0;
  assign N50 = sel_i[50];
  assign N51 = N255;
  assign { r_n_26__15_, r_n_26__14_, r_n_26__13_, r_n_26__12_, r_n_26__11_, r_n_26__10_, r_n_26__9_, r_n_26__8_, r_n_26__7_, r_n_26__6_, r_n_26__5_, r_n_26__4_, r_n_26__3_, r_n_26__2_, r_n_26__1_, r_n_26__0_ } = (N52)? { r_27__15_, r_27__14_, r_27__13_, r_27__12_, r_27__11_, r_27__10_, r_27__9_, r_27__8_, r_27__7_, r_27__6_, r_27__5_, r_27__4_, r_27__3_, r_27__2_, r_27__1_, r_27__0_ } : 
                                                                                                                                                                                                                    (N53)? data_i : 1'b0;
  assign N52 = sel_i[52];
  assign N53 = N260;
  assign { r_n_27__15_, r_n_27__14_, r_n_27__13_, r_n_27__12_, r_n_27__11_, r_n_27__10_, r_n_27__9_, r_n_27__8_, r_n_27__7_, r_n_27__6_, r_n_27__5_, r_n_27__4_, r_n_27__3_, r_n_27__2_, r_n_27__1_, r_n_27__0_ } = (N54)? { r_28__15_, r_28__14_, r_28__13_, r_28__12_, r_28__11_, r_28__10_, r_28__9_, r_28__8_, r_28__7_, r_28__6_, r_28__5_, r_28__4_, r_28__3_, r_28__2_, r_28__1_, r_28__0_ } : 
                                                                                                                                                                                                                    (N55)? data_i : 1'b0;
  assign N54 = sel_i[54];
  assign N55 = N265;
  assign { r_n_28__15_, r_n_28__14_, r_n_28__13_, r_n_28__12_, r_n_28__11_, r_n_28__10_, r_n_28__9_, r_n_28__8_, r_n_28__7_, r_n_28__6_, r_n_28__5_, r_n_28__4_, r_n_28__3_, r_n_28__2_, r_n_28__1_, r_n_28__0_ } = (N56)? { r_29__15_, r_29__14_, r_29__13_, r_29__12_, r_29__11_, r_29__10_, r_29__9_, r_29__8_, r_29__7_, r_29__6_, r_29__5_, r_29__4_, r_29__3_, r_29__2_, r_29__1_, r_29__0_ } : 
                                                                                                                                                                                                                    (N57)? data_i : 1'b0;
  assign N56 = sel_i[56];
  assign N57 = N270;
  assign { r_n_29__15_, r_n_29__14_, r_n_29__13_, r_n_29__12_, r_n_29__11_, r_n_29__10_, r_n_29__9_, r_n_29__8_, r_n_29__7_, r_n_29__6_, r_n_29__5_, r_n_29__4_, r_n_29__3_, r_n_29__2_, r_n_29__1_, r_n_29__0_ } = (N58)? { r_30__15_, r_30__14_, r_30__13_, r_30__12_, r_30__11_, r_30__10_, r_30__9_, r_30__8_, r_30__7_, r_30__6_, r_30__5_, r_30__4_, r_30__3_, r_30__2_, r_30__1_, r_30__0_ } : 
                                                                                                                                                                                                                    (N59)? data_i : 1'b0;
  assign N58 = sel_i[58];
  assign N59 = N275;
  assign { r_n_30__15_, r_n_30__14_, r_n_30__13_, r_n_30__12_, r_n_30__11_, r_n_30__10_, r_n_30__9_, r_n_30__8_, r_n_30__7_, r_n_30__6_, r_n_30__5_, r_n_30__4_, r_n_30__3_, r_n_30__2_, r_n_30__1_, r_n_30__0_ } = (N60)? { r_31__15_, r_31__14_, r_31__13_, r_31__12_, r_31__11_, r_31__10_, r_31__9_, r_31__8_, r_31__7_, r_31__6_, r_31__5_, r_31__4_, r_31__3_, r_31__2_, r_31__1_, r_31__0_ } : 
                                                                                                                                                                                                                    (N61)? data_i : 1'b0;
  assign N60 = sel_i[60];
  assign N61 = N280;
  assign { r_n_31__15_, r_n_31__14_, r_n_31__13_, r_n_31__12_, r_n_31__11_, r_n_31__10_, r_n_31__9_, r_n_31__8_, r_n_31__7_, r_n_31__6_, r_n_31__5_, r_n_31__4_, r_n_31__3_, r_n_31__2_, r_n_31__1_, r_n_31__0_ } = (N62)? { r_32__15_, r_32__14_, r_32__13_, r_32__12_, r_32__11_, r_32__10_, r_32__9_, r_32__8_, r_32__7_, r_32__6_, r_32__5_, r_32__4_, r_32__3_, r_32__2_, r_32__1_, r_32__0_ } : 
                                                                                                                                                                                                                    (N63)? data_i : 1'b0;
  assign N62 = sel_i[62];
  assign N63 = N285;
  assign { r_n_32__15_, r_n_32__14_, r_n_32__13_, r_n_32__12_, r_n_32__11_, r_n_32__10_, r_n_32__9_, r_n_32__8_, r_n_32__7_, r_n_32__6_, r_n_32__5_, r_n_32__4_, r_n_32__3_, r_n_32__2_, r_n_32__1_, r_n_32__0_ } = (N64)? { r_33__15_, r_33__14_, r_33__13_, r_33__12_, r_33__11_, r_33__10_, r_33__9_, r_33__8_, r_33__7_, r_33__6_, r_33__5_, r_33__4_, r_33__3_, r_33__2_, r_33__1_, r_33__0_ } : 
                                                                                                                                                                                                                    (N65)? data_i : 1'b0;
  assign N64 = sel_i[64];
  assign N65 = N290;
  assign { r_n_33__15_, r_n_33__14_, r_n_33__13_, r_n_33__12_, r_n_33__11_, r_n_33__10_, r_n_33__9_, r_n_33__8_, r_n_33__7_, r_n_33__6_, r_n_33__5_, r_n_33__4_, r_n_33__3_, r_n_33__2_, r_n_33__1_, r_n_33__0_ } = (N66)? { r_34__15_, r_34__14_, r_34__13_, r_34__12_, r_34__11_, r_34__10_, r_34__9_, r_34__8_, r_34__7_, r_34__6_, r_34__5_, r_34__4_, r_34__3_, r_34__2_, r_34__1_, r_34__0_ } : 
                                                                                                                                                                                                                    (N67)? data_i : 1'b0;
  assign N66 = sel_i[66];
  assign N67 = N295;
  assign { r_n_34__15_, r_n_34__14_, r_n_34__13_, r_n_34__12_, r_n_34__11_, r_n_34__10_, r_n_34__9_, r_n_34__8_, r_n_34__7_, r_n_34__6_, r_n_34__5_, r_n_34__4_, r_n_34__3_, r_n_34__2_, r_n_34__1_, r_n_34__0_ } = (N68)? { r_35__15_, r_35__14_, r_35__13_, r_35__12_, r_35__11_, r_35__10_, r_35__9_, r_35__8_, r_35__7_, r_35__6_, r_35__5_, r_35__4_, r_35__3_, r_35__2_, r_35__1_, r_35__0_ } : 
                                                                                                                                                                                                                    (N69)? data_i : 1'b0;
  assign N68 = sel_i[68];
  assign N69 = N300;
  assign { r_n_35__15_, r_n_35__14_, r_n_35__13_, r_n_35__12_, r_n_35__11_, r_n_35__10_, r_n_35__9_, r_n_35__8_, r_n_35__7_, r_n_35__6_, r_n_35__5_, r_n_35__4_, r_n_35__3_, r_n_35__2_, r_n_35__1_, r_n_35__0_ } = (N70)? { r_36__15_, r_36__14_, r_36__13_, r_36__12_, r_36__11_, r_36__10_, r_36__9_, r_36__8_, r_36__7_, r_36__6_, r_36__5_, r_36__4_, r_36__3_, r_36__2_, r_36__1_, r_36__0_ } : 
                                                                                                                                                                                                                    (N71)? data_i : 1'b0;
  assign N70 = sel_i[70];
  assign N71 = N305;
  assign { r_n_36__15_, r_n_36__14_, r_n_36__13_, r_n_36__12_, r_n_36__11_, r_n_36__10_, r_n_36__9_, r_n_36__8_, r_n_36__7_, r_n_36__6_, r_n_36__5_, r_n_36__4_, r_n_36__3_, r_n_36__2_, r_n_36__1_, r_n_36__0_ } = (N72)? { r_37__15_, r_37__14_, r_37__13_, r_37__12_, r_37__11_, r_37__10_, r_37__9_, r_37__8_, r_37__7_, r_37__6_, r_37__5_, r_37__4_, r_37__3_, r_37__2_, r_37__1_, r_37__0_ } : 
                                                                                                                                                                                                                    (N73)? data_i : 1'b0;
  assign N72 = sel_i[72];
  assign N73 = N310;
  assign { r_n_37__15_, r_n_37__14_, r_n_37__13_, r_n_37__12_, r_n_37__11_, r_n_37__10_, r_n_37__9_, r_n_37__8_, r_n_37__7_, r_n_37__6_, r_n_37__5_, r_n_37__4_, r_n_37__3_, r_n_37__2_, r_n_37__1_, r_n_37__0_ } = (N74)? { r_38__15_, r_38__14_, r_38__13_, r_38__12_, r_38__11_, r_38__10_, r_38__9_, r_38__8_, r_38__7_, r_38__6_, r_38__5_, r_38__4_, r_38__3_, r_38__2_, r_38__1_, r_38__0_ } : 
                                                                                                                                                                                                                    (N75)? data_i : 1'b0;
  assign N74 = sel_i[74];
  assign N75 = N315;
  assign { r_n_38__15_, r_n_38__14_, r_n_38__13_, r_n_38__12_, r_n_38__11_, r_n_38__10_, r_n_38__9_, r_n_38__8_, r_n_38__7_, r_n_38__6_, r_n_38__5_, r_n_38__4_, r_n_38__3_, r_n_38__2_, r_n_38__1_, r_n_38__0_ } = (N76)? { r_39__15_, r_39__14_, r_39__13_, r_39__12_, r_39__11_, r_39__10_, r_39__9_, r_39__8_, r_39__7_, r_39__6_, r_39__5_, r_39__4_, r_39__3_, r_39__2_, r_39__1_, r_39__0_ } : 
                                                                                                                                                                                                                    (N77)? data_i : 1'b0;
  assign N76 = sel_i[76];
  assign N77 = N320;
  assign { r_n_39__15_, r_n_39__14_, r_n_39__13_, r_n_39__12_, r_n_39__11_, r_n_39__10_, r_n_39__9_, r_n_39__8_, r_n_39__7_, r_n_39__6_, r_n_39__5_, r_n_39__4_, r_n_39__3_, r_n_39__2_, r_n_39__1_, r_n_39__0_ } = (N78)? { r_40__15_, r_40__14_, r_40__13_, r_40__12_, r_40__11_, r_40__10_, r_40__9_, r_40__8_, r_40__7_, r_40__6_, r_40__5_, r_40__4_, r_40__3_, r_40__2_, r_40__1_, r_40__0_ } : 
                                                                                                                                                                                                                    (N79)? data_i : 1'b0;
  assign N78 = sel_i[78];
  assign N79 = N325;
  assign { r_n_40__15_, r_n_40__14_, r_n_40__13_, r_n_40__12_, r_n_40__11_, r_n_40__10_, r_n_40__9_, r_n_40__8_, r_n_40__7_, r_n_40__6_, r_n_40__5_, r_n_40__4_, r_n_40__3_, r_n_40__2_, r_n_40__1_, r_n_40__0_ } = (N80)? { r_41__15_, r_41__14_, r_41__13_, r_41__12_, r_41__11_, r_41__10_, r_41__9_, r_41__8_, r_41__7_, r_41__6_, r_41__5_, r_41__4_, r_41__3_, r_41__2_, r_41__1_, r_41__0_ } : 
                                                                                                                                                                                                                    (N81)? data_i : 1'b0;
  assign N80 = sel_i[80];
  assign N81 = N330;
  assign { r_n_41__15_, r_n_41__14_, r_n_41__13_, r_n_41__12_, r_n_41__11_, r_n_41__10_, r_n_41__9_, r_n_41__8_, r_n_41__7_, r_n_41__6_, r_n_41__5_, r_n_41__4_, r_n_41__3_, r_n_41__2_, r_n_41__1_, r_n_41__0_ } = (N82)? { r_42__15_, r_42__14_, r_42__13_, r_42__12_, r_42__11_, r_42__10_, r_42__9_, r_42__8_, r_42__7_, r_42__6_, r_42__5_, r_42__4_, r_42__3_, r_42__2_, r_42__1_, r_42__0_ } : 
                                                                                                                                                                                                                    (N83)? data_i : 1'b0;
  assign N82 = sel_i[82];
  assign N83 = N335;
  assign { r_n_42__15_, r_n_42__14_, r_n_42__13_, r_n_42__12_, r_n_42__11_, r_n_42__10_, r_n_42__9_, r_n_42__8_, r_n_42__7_, r_n_42__6_, r_n_42__5_, r_n_42__4_, r_n_42__3_, r_n_42__2_, r_n_42__1_, r_n_42__0_ } = (N84)? { r_43__15_, r_43__14_, r_43__13_, r_43__12_, r_43__11_, r_43__10_, r_43__9_, r_43__8_, r_43__7_, r_43__6_, r_43__5_, r_43__4_, r_43__3_, r_43__2_, r_43__1_, r_43__0_ } : 
                                                                                                                                                                                                                    (N85)? data_i : 1'b0;
  assign N84 = sel_i[84];
  assign N85 = N340;
  assign { r_n_43__15_, r_n_43__14_, r_n_43__13_, r_n_43__12_, r_n_43__11_, r_n_43__10_, r_n_43__9_, r_n_43__8_, r_n_43__7_, r_n_43__6_, r_n_43__5_, r_n_43__4_, r_n_43__3_, r_n_43__2_, r_n_43__1_, r_n_43__0_ } = (N86)? { r_44__15_, r_44__14_, r_44__13_, r_44__12_, r_44__11_, r_44__10_, r_44__9_, r_44__8_, r_44__7_, r_44__6_, r_44__5_, r_44__4_, r_44__3_, r_44__2_, r_44__1_, r_44__0_ } : 
                                                                                                                                                                                                                    (N87)? data_i : 1'b0;
  assign N86 = sel_i[86];
  assign N87 = N345;
  assign { r_n_44__15_, r_n_44__14_, r_n_44__13_, r_n_44__12_, r_n_44__11_, r_n_44__10_, r_n_44__9_, r_n_44__8_, r_n_44__7_, r_n_44__6_, r_n_44__5_, r_n_44__4_, r_n_44__3_, r_n_44__2_, r_n_44__1_, r_n_44__0_ } = (N88)? { r_45__15_, r_45__14_, r_45__13_, r_45__12_, r_45__11_, r_45__10_, r_45__9_, r_45__8_, r_45__7_, r_45__6_, r_45__5_, r_45__4_, r_45__3_, r_45__2_, r_45__1_, r_45__0_ } : 
                                                                                                                                                                                                                    (N89)? data_i : 1'b0;
  assign N88 = sel_i[88];
  assign N89 = N350;
  assign { r_n_45__15_, r_n_45__14_, r_n_45__13_, r_n_45__12_, r_n_45__11_, r_n_45__10_, r_n_45__9_, r_n_45__8_, r_n_45__7_, r_n_45__6_, r_n_45__5_, r_n_45__4_, r_n_45__3_, r_n_45__2_, r_n_45__1_, r_n_45__0_ } = (N90)? { r_46__15_, r_46__14_, r_46__13_, r_46__12_, r_46__11_, r_46__10_, r_46__9_, r_46__8_, r_46__7_, r_46__6_, r_46__5_, r_46__4_, r_46__3_, r_46__2_, r_46__1_, r_46__0_ } : 
                                                                                                                                                                                                                    (N91)? data_i : 1'b0;
  assign N90 = sel_i[90];
  assign N91 = N355;
  assign { r_n_46__15_, r_n_46__14_, r_n_46__13_, r_n_46__12_, r_n_46__11_, r_n_46__10_, r_n_46__9_, r_n_46__8_, r_n_46__7_, r_n_46__6_, r_n_46__5_, r_n_46__4_, r_n_46__3_, r_n_46__2_, r_n_46__1_, r_n_46__0_ } = (N92)? { r_47__15_, r_47__14_, r_47__13_, r_47__12_, r_47__11_, r_47__10_, r_47__9_, r_47__8_, r_47__7_, r_47__6_, r_47__5_, r_47__4_, r_47__3_, r_47__2_, r_47__1_, r_47__0_ } : 
                                                                                                                                                                                                                    (N93)? data_i : 1'b0;
  assign N92 = sel_i[92];
  assign N93 = N360;
  assign { r_n_47__15_, r_n_47__14_, r_n_47__13_, r_n_47__12_, r_n_47__11_, r_n_47__10_, r_n_47__9_, r_n_47__8_, r_n_47__7_, r_n_47__6_, r_n_47__5_, r_n_47__4_, r_n_47__3_, r_n_47__2_, r_n_47__1_, r_n_47__0_ } = (N94)? { r_48__15_, r_48__14_, r_48__13_, r_48__12_, r_48__11_, r_48__10_, r_48__9_, r_48__8_, r_48__7_, r_48__6_, r_48__5_, r_48__4_, r_48__3_, r_48__2_, r_48__1_, r_48__0_ } : 
                                                                                                                                                                                                                    (N95)? data_i : 1'b0;
  assign N94 = sel_i[94];
  assign N95 = N365;
  assign { r_n_48__15_, r_n_48__14_, r_n_48__13_, r_n_48__12_, r_n_48__11_, r_n_48__10_, r_n_48__9_, r_n_48__8_, r_n_48__7_, r_n_48__6_, r_n_48__5_, r_n_48__4_, r_n_48__3_, r_n_48__2_, r_n_48__1_, r_n_48__0_ } = (N96)? { r_49__15_, r_49__14_, r_49__13_, r_49__12_, r_49__11_, r_49__10_, r_49__9_, r_49__8_, r_49__7_, r_49__6_, r_49__5_, r_49__4_, r_49__3_, r_49__2_, r_49__1_, r_49__0_ } : 
                                                                                                                                                                                                                    (N97)? data_i : 1'b0;
  assign N96 = sel_i[96];
  assign N97 = N370;
  assign { r_n_49__15_, r_n_49__14_, r_n_49__13_, r_n_49__12_, r_n_49__11_, r_n_49__10_, r_n_49__9_, r_n_49__8_, r_n_49__7_, r_n_49__6_, r_n_49__5_, r_n_49__4_, r_n_49__3_, r_n_49__2_, r_n_49__1_, r_n_49__0_ } = (N98)? { r_50__15_, r_50__14_, r_50__13_, r_50__12_, r_50__11_, r_50__10_, r_50__9_, r_50__8_, r_50__7_, r_50__6_, r_50__5_, r_50__4_, r_50__3_, r_50__2_, r_50__1_, r_50__0_ } : 
                                                                                                                                                                                                                    (N99)? data_i : 1'b0;
  assign N98 = sel_i[98];
  assign N99 = N375;
  assign { r_n_50__15_, r_n_50__14_, r_n_50__13_, r_n_50__12_, r_n_50__11_, r_n_50__10_, r_n_50__9_, r_n_50__8_, r_n_50__7_, r_n_50__6_, r_n_50__5_, r_n_50__4_, r_n_50__3_, r_n_50__2_, r_n_50__1_, r_n_50__0_ } = (N100)? { r_51__15_, r_51__14_, r_51__13_, r_51__12_, r_51__11_, r_51__10_, r_51__9_, r_51__8_, r_51__7_, r_51__6_, r_51__5_, r_51__4_, r_51__3_, r_51__2_, r_51__1_, r_51__0_ } : 
                                                                                                                                                                                                                    (N101)? data_i : 1'b0;
  assign N100 = sel_i[100];
  assign N101 = N380;
  assign { r_n_51__15_, r_n_51__14_, r_n_51__13_, r_n_51__12_, r_n_51__11_, r_n_51__10_, r_n_51__9_, r_n_51__8_, r_n_51__7_, r_n_51__6_, r_n_51__5_, r_n_51__4_, r_n_51__3_, r_n_51__2_, r_n_51__1_, r_n_51__0_ } = (N102)? { r_52__15_, r_52__14_, r_52__13_, r_52__12_, r_52__11_, r_52__10_, r_52__9_, r_52__8_, r_52__7_, r_52__6_, r_52__5_, r_52__4_, r_52__3_, r_52__2_, r_52__1_, r_52__0_ } : 
                                                                                                                                                                                                                    (N103)? data_i : 1'b0;
  assign N102 = sel_i[102];
  assign N103 = N385;
  assign { r_n_52__15_, r_n_52__14_, r_n_52__13_, r_n_52__12_, r_n_52__11_, r_n_52__10_, r_n_52__9_, r_n_52__8_, r_n_52__7_, r_n_52__6_, r_n_52__5_, r_n_52__4_, r_n_52__3_, r_n_52__2_, r_n_52__1_, r_n_52__0_ } = (N104)? { r_53__15_, r_53__14_, r_53__13_, r_53__12_, r_53__11_, r_53__10_, r_53__9_, r_53__8_, r_53__7_, r_53__6_, r_53__5_, r_53__4_, r_53__3_, r_53__2_, r_53__1_, r_53__0_ } : 
                                                                                                                                                                                                                    (N105)? data_i : 1'b0;
  assign N104 = sel_i[104];
  assign N105 = N390;
  assign { r_n_53__15_, r_n_53__14_, r_n_53__13_, r_n_53__12_, r_n_53__11_, r_n_53__10_, r_n_53__9_, r_n_53__8_, r_n_53__7_, r_n_53__6_, r_n_53__5_, r_n_53__4_, r_n_53__3_, r_n_53__2_, r_n_53__1_, r_n_53__0_ } = (N106)? { r_54__15_, r_54__14_, r_54__13_, r_54__12_, r_54__11_, r_54__10_, r_54__9_, r_54__8_, r_54__7_, r_54__6_, r_54__5_, r_54__4_, r_54__3_, r_54__2_, r_54__1_, r_54__0_ } : 
                                                                                                                                                                                                                    (N107)? data_i : 1'b0;
  assign N106 = sel_i[106];
  assign N107 = N395;
  assign { r_n_54__15_, r_n_54__14_, r_n_54__13_, r_n_54__12_, r_n_54__11_, r_n_54__10_, r_n_54__9_, r_n_54__8_, r_n_54__7_, r_n_54__6_, r_n_54__5_, r_n_54__4_, r_n_54__3_, r_n_54__2_, r_n_54__1_, r_n_54__0_ } = (N108)? { r_55__15_, r_55__14_, r_55__13_, r_55__12_, r_55__11_, r_55__10_, r_55__9_, r_55__8_, r_55__7_, r_55__6_, r_55__5_, r_55__4_, r_55__3_, r_55__2_, r_55__1_, r_55__0_ } : 
                                                                                                                                                                                                                    (N109)? data_i : 1'b0;
  assign N108 = sel_i[108];
  assign N109 = N400;
  assign { r_n_55__15_, r_n_55__14_, r_n_55__13_, r_n_55__12_, r_n_55__11_, r_n_55__10_, r_n_55__9_, r_n_55__8_, r_n_55__7_, r_n_55__6_, r_n_55__5_, r_n_55__4_, r_n_55__3_, r_n_55__2_, r_n_55__1_, r_n_55__0_ } = (N110)? { r_56__15_, r_56__14_, r_56__13_, r_56__12_, r_56__11_, r_56__10_, r_56__9_, r_56__8_, r_56__7_, r_56__6_, r_56__5_, r_56__4_, r_56__3_, r_56__2_, r_56__1_, r_56__0_ } : 
                                                                                                                                                                                                                    (N111)? data_i : 1'b0;
  assign N110 = sel_i[110];
  assign N111 = N405;
  assign { r_n_56__15_, r_n_56__14_, r_n_56__13_, r_n_56__12_, r_n_56__11_, r_n_56__10_, r_n_56__9_, r_n_56__8_, r_n_56__7_, r_n_56__6_, r_n_56__5_, r_n_56__4_, r_n_56__3_, r_n_56__2_, r_n_56__1_, r_n_56__0_ } = (N112)? { r_57__15_, r_57__14_, r_57__13_, r_57__12_, r_57__11_, r_57__10_, r_57__9_, r_57__8_, r_57__7_, r_57__6_, r_57__5_, r_57__4_, r_57__3_, r_57__2_, r_57__1_, r_57__0_ } : 
                                                                                                                                                                                                                    (N113)? data_i : 1'b0;
  assign N112 = sel_i[112];
  assign N113 = N410;
  assign { r_n_57__15_, r_n_57__14_, r_n_57__13_, r_n_57__12_, r_n_57__11_, r_n_57__10_, r_n_57__9_, r_n_57__8_, r_n_57__7_, r_n_57__6_, r_n_57__5_, r_n_57__4_, r_n_57__3_, r_n_57__2_, r_n_57__1_, r_n_57__0_ } = (N114)? { r_58__15_, r_58__14_, r_58__13_, r_58__12_, r_58__11_, r_58__10_, r_58__9_, r_58__8_, r_58__7_, r_58__6_, r_58__5_, r_58__4_, r_58__3_, r_58__2_, r_58__1_, r_58__0_ } : 
                                                                                                                                                                                                                    (N115)? data_i : 1'b0;
  assign N114 = sel_i[114];
  assign N115 = N415;
  assign { r_n_58__15_, r_n_58__14_, r_n_58__13_, r_n_58__12_, r_n_58__11_, r_n_58__10_, r_n_58__9_, r_n_58__8_, r_n_58__7_, r_n_58__6_, r_n_58__5_, r_n_58__4_, r_n_58__3_, r_n_58__2_, r_n_58__1_, r_n_58__0_ } = (N116)? { r_59__15_, r_59__14_, r_59__13_, r_59__12_, r_59__11_, r_59__10_, r_59__9_, r_59__8_, r_59__7_, r_59__6_, r_59__5_, r_59__4_, r_59__3_, r_59__2_, r_59__1_, r_59__0_ } : 
                                                                                                                                                                                                                    (N117)? data_i : 1'b0;
  assign N116 = sel_i[116];
  assign N117 = N420;
  assign { r_n_59__15_, r_n_59__14_, r_n_59__13_, r_n_59__12_, r_n_59__11_, r_n_59__10_, r_n_59__9_, r_n_59__8_, r_n_59__7_, r_n_59__6_, r_n_59__5_, r_n_59__4_, r_n_59__3_, r_n_59__2_, r_n_59__1_, r_n_59__0_ } = (N118)? { r_60__15_, r_60__14_, r_60__13_, r_60__12_, r_60__11_, r_60__10_, r_60__9_, r_60__8_, r_60__7_, r_60__6_, r_60__5_, r_60__4_, r_60__3_, r_60__2_, r_60__1_, r_60__0_ } : 
                                                                                                                                                                                                                    (N119)? data_i : 1'b0;
  assign N118 = sel_i[118];
  assign N119 = N425;
  assign { r_n_60__15_, r_n_60__14_, r_n_60__13_, r_n_60__12_, r_n_60__11_, r_n_60__10_, r_n_60__9_, r_n_60__8_, r_n_60__7_, r_n_60__6_, r_n_60__5_, r_n_60__4_, r_n_60__3_, r_n_60__2_, r_n_60__1_, r_n_60__0_ } = (N120)? { r_61__15_, r_61__14_, r_61__13_, r_61__12_, r_61__11_, r_61__10_, r_61__9_, r_61__8_, r_61__7_, r_61__6_, r_61__5_, r_61__4_, r_61__3_, r_61__2_, r_61__1_, r_61__0_ } : 
                                                                                                                                                                                                                    (N121)? data_i : 1'b0;
  assign N120 = sel_i[120];
  assign N121 = N430;
  assign { r_n_61__15_, r_n_61__14_, r_n_61__13_, r_n_61__12_, r_n_61__11_, r_n_61__10_, r_n_61__9_, r_n_61__8_, r_n_61__7_, r_n_61__6_, r_n_61__5_, r_n_61__4_, r_n_61__3_, r_n_61__2_, r_n_61__1_, r_n_61__0_ } = (N122)? { r_62__15_, r_62__14_, r_62__13_, r_62__12_, r_62__11_, r_62__10_, r_62__9_, r_62__8_, r_62__7_, r_62__6_, r_62__5_, r_62__4_, r_62__3_, r_62__2_, r_62__1_, r_62__0_ } : 
                                                                                                                                                                                                                    (N123)? data_i : 1'b0;
  assign N122 = sel_i[122];
  assign N123 = N435;
  assign { r_n_62__15_, r_n_62__14_, r_n_62__13_, r_n_62__12_, r_n_62__11_, r_n_62__10_, r_n_62__9_, r_n_62__8_, r_n_62__7_, r_n_62__6_, r_n_62__5_, r_n_62__4_, r_n_62__3_, r_n_62__2_, r_n_62__1_, r_n_62__0_ } = (N124)? { r_63__15_, r_63__14_, r_63__13_, r_63__12_, r_63__11_, r_63__10_, r_63__9_, r_63__8_, r_63__7_, r_63__6_, r_63__5_, r_63__4_, r_63__3_, r_63__2_, r_63__1_, r_63__0_ } : 
                                                                                                                                                                                                                    (N125)? data_i : 1'b0;
  assign N124 = sel_i[124];
  assign N125 = N440;
  assign N127 = ~sel_i[1];
  assign N129 = N126 | N128;
  assign N132 = ~sel_i[3];
  assign N134 = N131 | N133;
  assign N137 = ~sel_i[5];
  assign N139 = N136 | N138;
  assign N142 = ~sel_i[7];
  assign N144 = N141 | N143;
  assign N147 = ~sel_i[9];
  assign N149 = N146 | N148;
  assign N152 = ~sel_i[11];
  assign N154 = N151 | N153;
  assign N157 = ~sel_i[13];
  assign N159 = N156 | N158;
  assign N162 = ~sel_i[15];
  assign N164 = N161 | N163;
  assign N167 = ~sel_i[17];
  assign N169 = N166 | N168;
  assign N172 = ~sel_i[19];
  assign N174 = N171 | N173;
  assign N177 = ~sel_i[21];
  assign N179 = N176 | N178;
  assign N182 = ~sel_i[23];
  assign N184 = N181 | N183;
  assign N187 = ~sel_i[25];
  assign N189 = N186 | N188;
  assign N192 = ~sel_i[27];
  assign N194 = N191 | N193;
  assign N197 = ~sel_i[29];
  assign N199 = N196 | N198;
  assign N202 = ~sel_i[31];
  assign N204 = N201 | N203;
  assign N207 = ~sel_i[33];
  assign N209 = N206 | N208;
  assign N212 = ~sel_i[35];
  assign N214 = N211 | N213;
  assign N217 = ~sel_i[37];
  assign N219 = N216 | N218;
  assign N222 = ~sel_i[39];
  assign N224 = N221 | N223;
  assign N227 = ~sel_i[41];
  assign N229 = N226 | N228;
  assign N232 = ~sel_i[43];
  assign N234 = N231 | N233;
  assign N237 = ~sel_i[45];
  assign N239 = N236 | N238;
  assign N242 = ~sel_i[47];
  assign N244 = N241 | N243;
  assign N247 = ~sel_i[49];
  assign N249 = N246 | N248;
  assign N252 = ~sel_i[51];
  assign N254 = N251 | N253;
  assign N257 = ~sel_i[53];
  assign N259 = N256 | N258;
  assign N262 = ~sel_i[55];
  assign N264 = N261 | N263;
  assign N267 = ~sel_i[57];
  assign N269 = N266 | N268;
  assign N272 = ~sel_i[59];
  assign N274 = N271 | N273;
  assign N277 = ~sel_i[61];
  assign N279 = N276 | N278;
  assign N282 = ~sel_i[63];
  assign N284 = N281 | N283;
  assign N287 = ~sel_i[65];
  assign N289 = N286 | N288;
  assign N292 = ~sel_i[67];
  assign N294 = N291 | N293;
  assign N297 = ~sel_i[69];
  assign N299 = N296 | N298;
  assign N302 = ~sel_i[71];
  assign N304 = N301 | N303;
  assign N307 = ~sel_i[73];
  assign N309 = N306 | N308;
  assign N312 = ~sel_i[75];
  assign N314 = N311 | N313;
  assign N317 = ~sel_i[77];
  assign N319 = N316 | N318;
  assign N322 = ~sel_i[79];
  assign N324 = N321 | N323;
  assign N327 = ~sel_i[81];
  assign N329 = N326 | N328;
  assign N332 = ~sel_i[83];
  assign N334 = N331 | N333;
  assign N337 = ~sel_i[85];
  assign N339 = N336 | N338;
  assign N342 = ~sel_i[87];
  assign N344 = N341 | N343;
  assign N347 = ~sel_i[89];
  assign N349 = N346 | N348;
  assign N352 = ~sel_i[91];
  assign N354 = N351 | N353;
  assign N357 = ~sel_i[93];
  assign N359 = N356 | N358;
  assign N362 = ~sel_i[95];
  assign N364 = N361 | N363;
  assign N367 = ~sel_i[97];
  assign N369 = N366 | N368;
  assign N372 = ~sel_i[99];
  assign N374 = N371 | N373;
  assign N377 = ~sel_i[101];
  assign N379 = N376 | N378;
  assign N382 = ~sel_i[103];
  assign N384 = N381 | N383;
  assign N387 = ~sel_i[105];
  assign N389 = N386 | N388;
  assign N392 = ~sel_i[107];
  assign N394 = N391 | N393;
  assign N397 = ~sel_i[109];
  assign N399 = N396 | N398;
  assign N402 = ~sel_i[111];
  assign N404 = N401 | N403;
  assign N407 = ~sel_i[113];
  assign N409 = N406 | N408;
  assign N412 = ~sel_i[115];
  assign N414 = N411 | N413;
  assign N417 = ~sel_i[117];
  assign N419 = N416 | N418;
  assign N422 = ~sel_i[119];
  assign N424 = N421 | N423;
  assign N427 = ~sel_i[121];
  assign N429 = N426 | N428;
  assign N432 = ~sel_i[123];
  assign N434 = N431 | N433;
  assign N437 = ~sel_i[125];
  assign N439 = N436 | N438;
  assign N441 = ~sel_i[126];
  assign N443 = ~N442;
  assign N445 = ~sel_i[127];
  assign N447 = N444 | N446;
  assign N448 = ~N129;
  assign N449 = ~N134;
  assign N450 = ~N139;
  assign N451 = ~N144;
  assign N452 = ~N149;
  assign N453 = ~N154;
  assign N454 = ~N159;
  assign N455 = ~N164;
  assign N456 = ~N169;
  assign N457 = ~N174;
  assign N458 = ~N179;
  assign N459 = ~N184;
  assign N460 = ~N189;
  assign N461 = ~N194;
  assign N462 = ~N199;
  assign N463 = ~N204;
  assign N464 = ~N209;
  assign N465 = ~N214;
  assign N466 = ~N219;
  assign N467 = ~N224;
  assign N468 = ~N229;
  assign N469 = ~N234;
  assign N470 = ~N239;
  assign N471 = ~N244;
  assign N472 = ~N249;
  assign N473 = ~N254;
  assign N474 = ~N259;
  assign N475 = ~N264;
  assign N476 = ~N269;
  assign N477 = ~N274;
  assign N478 = ~N279;
  assign N479 = ~N284;
  assign N480 = ~N289;
  assign N481 = ~N294;
  assign N482 = ~N299;
  assign N483 = ~N304;
  assign N484 = ~N309;
  assign N485 = ~N314;
  assign N486 = ~N319;
  assign N487 = ~N324;
  assign N488 = ~N329;
  assign N489 = ~N334;
  assign N490 = ~N339;
  assign N491 = ~N344;
  assign N492 = ~N349;
  assign N493 = ~N354;
  assign N494 = ~N359;
  assign N495 = ~N364;
  assign N496 = ~N369;
  assign N497 = ~N374;
  assign N498 = ~N379;
  assign N499 = ~N384;
  assign N500 = ~N389;
  assign N501 = ~N394;
  assign N502 = ~N399;
  assign N503 = ~N404;
  assign N504 = ~N409;
  assign N505 = ~N414;
  assign N506 = ~N419;
  assign N507 = ~N424;
  assign N508 = ~N429;
  assign N509 = ~N434;
  assign N510 = ~N439;
  assign N511 = ~N447;

  always @(posedge clk_i) begin
    if(N448) begin
      data_o_15_sv2v_reg <= r_n_0__15_;
      data_o_14_sv2v_reg <= r_n_0__14_;
      data_o_13_sv2v_reg <= r_n_0__13_;
      data_o_12_sv2v_reg <= r_n_0__12_;
      data_o_11_sv2v_reg <= r_n_0__11_;
      data_o_10_sv2v_reg <= r_n_0__10_;
      data_o_9_sv2v_reg <= r_n_0__9_;
      data_o_8_sv2v_reg <= r_n_0__8_;
      data_o_7_sv2v_reg <= r_n_0__7_;
      data_o_6_sv2v_reg <= r_n_0__6_;
      data_o_5_sv2v_reg <= r_n_0__5_;
      data_o_4_sv2v_reg <= r_n_0__4_;
      data_o_3_sv2v_reg <= r_n_0__3_;
      data_o_2_sv2v_reg <= r_n_0__2_;
      data_o_1_sv2v_reg <= r_n_0__1_;
      data_o_0_sv2v_reg <= r_n_0__0_;
    end 
    if(N449) begin
      r_1__15__sv2v_reg <= r_n_1__15_;
      r_1__14__sv2v_reg <= r_n_1__14_;
      r_1__13__sv2v_reg <= r_n_1__13_;
      r_1__12__sv2v_reg <= r_n_1__12_;
      r_1__11__sv2v_reg <= r_n_1__11_;
      r_1__10__sv2v_reg <= r_n_1__10_;
      r_1__9__sv2v_reg <= r_n_1__9_;
      r_1__8__sv2v_reg <= r_n_1__8_;
      r_1__7__sv2v_reg <= r_n_1__7_;
      r_1__6__sv2v_reg <= r_n_1__6_;
      r_1__5__sv2v_reg <= r_n_1__5_;
      r_1__4__sv2v_reg <= r_n_1__4_;
      r_1__3__sv2v_reg <= r_n_1__3_;
      r_1__2__sv2v_reg <= r_n_1__2_;
      r_1__1__sv2v_reg <= r_n_1__1_;
      r_1__0__sv2v_reg <= r_n_1__0_;
    end 
    if(N450) begin
      r_2__15__sv2v_reg <= r_n_2__15_;
      r_2__14__sv2v_reg <= r_n_2__14_;
      r_2__13__sv2v_reg <= r_n_2__13_;
      r_2__12__sv2v_reg <= r_n_2__12_;
      r_2__11__sv2v_reg <= r_n_2__11_;
      r_2__10__sv2v_reg <= r_n_2__10_;
      r_2__9__sv2v_reg <= r_n_2__9_;
      r_2__8__sv2v_reg <= r_n_2__8_;
      r_2__7__sv2v_reg <= r_n_2__7_;
      r_2__6__sv2v_reg <= r_n_2__6_;
      r_2__5__sv2v_reg <= r_n_2__5_;
      r_2__4__sv2v_reg <= r_n_2__4_;
      r_2__3__sv2v_reg <= r_n_2__3_;
      r_2__2__sv2v_reg <= r_n_2__2_;
      r_2__1__sv2v_reg <= r_n_2__1_;
      r_2__0__sv2v_reg <= r_n_2__0_;
    end 
    if(N451) begin
      r_3__15__sv2v_reg <= r_n_3__15_;
      r_3__14__sv2v_reg <= r_n_3__14_;
      r_3__13__sv2v_reg <= r_n_3__13_;
      r_3__12__sv2v_reg <= r_n_3__12_;
      r_3__11__sv2v_reg <= r_n_3__11_;
      r_3__10__sv2v_reg <= r_n_3__10_;
      r_3__9__sv2v_reg <= r_n_3__9_;
      r_3__8__sv2v_reg <= r_n_3__8_;
      r_3__7__sv2v_reg <= r_n_3__7_;
      r_3__6__sv2v_reg <= r_n_3__6_;
      r_3__5__sv2v_reg <= r_n_3__5_;
      r_3__4__sv2v_reg <= r_n_3__4_;
      r_3__3__sv2v_reg <= r_n_3__3_;
      r_3__2__sv2v_reg <= r_n_3__2_;
      r_3__1__sv2v_reg <= r_n_3__1_;
      r_3__0__sv2v_reg <= r_n_3__0_;
    end 
    if(N452) begin
      r_4__15__sv2v_reg <= r_n_4__15_;
      r_4__14__sv2v_reg <= r_n_4__14_;
      r_4__13__sv2v_reg <= r_n_4__13_;
      r_4__12__sv2v_reg <= r_n_4__12_;
      r_4__11__sv2v_reg <= r_n_4__11_;
      r_4__10__sv2v_reg <= r_n_4__10_;
      r_4__9__sv2v_reg <= r_n_4__9_;
      r_4__8__sv2v_reg <= r_n_4__8_;
      r_4__7__sv2v_reg <= r_n_4__7_;
      r_4__6__sv2v_reg <= r_n_4__6_;
      r_4__5__sv2v_reg <= r_n_4__5_;
      r_4__4__sv2v_reg <= r_n_4__4_;
      r_4__3__sv2v_reg <= r_n_4__3_;
      r_4__2__sv2v_reg <= r_n_4__2_;
      r_4__1__sv2v_reg <= r_n_4__1_;
      r_4__0__sv2v_reg <= r_n_4__0_;
    end 
    if(N453) begin
      r_5__15__sv2v_reg <= r_n_5__15_;
      r_5__14__sv2v_reg <= r_n_5__14_;
      r_5__13__sv2v_reg <= r_n_5__13_;
      r_5__12__sv2v_reg <= r_n_5__12_;
      r_5__11__sv2v_reg <= r_n_5__11_;
      r_5__10__sv2v_reg <= r_n_5__10_;
      r_5__9__sv2v_reg <= r_n_5__9_;
      r_5__8__sv2v_reg <= r_n_5__8_;
      r_5__7__sv2v_reg <= r_n_5__7_;
      r_5__6__sv2v_reg <= r_n_5__6_;
      r_5__5__sv2v_reg <= r_n_5__5_;
      r_5__4__sv2v_reg <= r_n_5__4_;
      r_5__3__sv2v_reg <= r_n_5__3_;
      r_5__2__sv2v_reg <= r_n_5__2_;
      r_5__1__sv2v_reg <= r_n_5__1_;
      r_5__0__sv2v_reg <= r_n_5__0_;
    end 
    if(N454) begin
      r_6__15__sv2v_reg <= r_n_6__15_;
      r_6__14__sv2v_reg <= r_n_6__14_;
      r_6__13__sv2v_reg <= r_n_6__13_;
      r_6__12__sv2v_reg <= r_n_6__12_;
      r_6__11__sv2v_reg <= r_n_6__11_;
      r_6__10__sv2v_reg <= r_n_6__10_;
      r_6__9__sv2v_reg <= r_n_6__9_;
      r_6__8__sv2v_reg <= r_n_6__8_;
      r_6__7__sv2v_reg <= r_n_6__7_;
      r_6__6__sv2v_reg <= r_n_6__6_;
      r_6__5__sv2v_reg <= r_n_6__5_;
      r_6__4__sv2v_reg <= r_n_6__4_;
      r_6__3__sv2v_reg <= r_n_6__3_;
      r_6__2__sv2v_reg <= r_n_6__2_;
      r_6__1__sv2v_reg <= r_n_6__1_;
      r_6__0__sv2v_reg <= r_n_6__0_;
    end 
    if(N455) begin
      r_7__15__sv2v_reg <= r_n_7__15_;
      r_7__14__sv2v_reg <= r_n_7__14_;
      r_7__13__sv2v_reg <= r_n_7__13_;
      r_7__12__sv2v_reg <= r_n_7__12_;
      r_7__11__sv2v_reg <= r_n_7__11_;
      r_7__10__sv2v_reg <= r_n_7__10_;
      r_7__9__sv2v_reg <= r_n_7__9_;
      r_7__8__sv2v_reg <= r_n_7__8_;
      r_7__7__sv2v_reg <= r_n_7__7_;
      r_7__6__sv2v_reg <= r_n_7__6_;
      r_7__5__sv2v_reg <= r_n_7__5_;
      r_7__4__sv2v_reg <= r_n_7__4_;
      r_7__3__sv2v_reg <= r_n_7__3_;
      r_7__2__sv2v_reg <= r_n_7__2_;
      r_7__1__sv2v_reg <= r_n_7__1_;
      r_7__0__sv2v_reg <= r_n_7__0_;
    end 
    if(N456) begin
      r_8__15__sv2v_reg <= r_n_8__15_;
      r_8__14__sv2v_reg <= r_n_8__14_;
      r_8__13__sv2v_reg <= r_n_8__13_;
      r_8__12__sv2v_reg <= r_n_8__12_;
      r_8__11__sv2v_reg <= r_n_8__11_;
      r_8__10__sv2v_reg <= r_n_8__10_;
      r_8__9__sv2v_reg <= r_n_8__9_;
      r_8__8__sv2v_reg <= r_n_8__8_;
      r_8__7__sv2v_reg <= r_n_8__7_;
      r_8__6__sv2v_reg <= r_n_8__6_;
      r_8__5__sv2v_reg <= r_n_8__5_;
      r_8__4__sv2v_reg <= r_n_8__4_;
      r_8__3__sv2v_reg <= r_n_8__3_;
      r_8__2__sv2v_reg <= r_n_8__2_;
      r_8__1__sv2v_reg <= r_n_8__1_;
      r_8__0__sv2v_reg <= r_n_8__0_;
    end 
    if(N457) begin
      r_9__15__sv2v_reg <= r_n_9__15_;
      r_9__14__sv2v_reg <= r_n_9__14_;
      r_9__13__sv2v_reg <= r_n_9__13_;
      r_9__12__sv2v_reg <= r_n_9__12_;
      r_9__11__sv2v_reg <= r_n_9__11_;
      r_9__10__sv2v_reg <= r_n_9__10_;
      r_9__9__sv2v_reg <= r_n_9__9_;
      r_9__8__sv2v_reg <= r_n_9__8_;
      r_9__7__sv2v_reg <= r_n_9__7_;
      r_9__6__sv2v_reg <= r_n_9__6_;
      r_9__5__sv2v_reg <= r_n_9__5_;
      r_9__4__sv2v_reg <= r_n_9__4_;
      r_9__3__sv2v_reg <= r_n_9__3_;
      r_9__2__sv2v_reg <= r_n_9__2_;
      r_9__1__sv2v_reg <= r_n_9__1_;
      r_9__0__sv2v_reg <= r_n_9__0_;
    end 
    if(N458) begin
      r_10__15__sv2v_reg <= r_n_10__15_;
      r_10__14__sv2v_reg <= r_n_10__14_;
      r_10__13__sv2v_reg <= r_n_10__13_;
      r_10__12__sv2v_reg <= r_n_10__12_;
      r_10__11__sv2v_reg <= r_n_10__11_;
      r_10__10__sv2v_reg <= r_n_10__10_;
      r_10__9__sv2v_reg <= r_n_10__9_;
      r_10__8__sv2v_reg <= r_n_10__8_;
      r_10__7__sv2v_reg <= r_n_10__7_;
      r_10__6__sv2v_reg <= r_n_10__6_;
      r_10__5__sv2v_reg <= r_n_10__5_;
      r_10__4__sv2v_reg <= r_n_10__4_;
      r_10__3__sv2v_reg <= r_n_10__3_;
      r_10__2__sv2v_reg <= r_n_10__2_;
      r_10__1__sv2v_reg <= r_n_10__1_;
      r_10__0__sv2v_reg <= r_n_10__0_;
    end 
    if(N459) begin
      r_11__15__sv2v_reg <= r_n_11__15_;
      r_11__14__sv2v_reg <= r_n_11__14_;
      r_11__13__sv2v_reg <= r_n_11__13_;
      r_11__12__sv2v_reg <= r_n_11__12_;
      r_11__11__sv2v_reg <= r_n_11__11_;
      r_11__10__sv2v_reg <= r_n_11__10_;
      r_11__9__sv2v_reg <= r_n_11__9_;
      r_11__8__sv2v_reg <= r_n_11__8_;
      r_11__7__sv2v_reg <= r_n_11__7_;
      r_11__6__sv2v_reg <= r_n_11__6_;
      r_11__5__sv2v_reg <= r_n_11__5_;
      r_11__4__sv2v_reg <= r_n_11__4_;
      r_11__3__sv2v_reg <= r_n_11__3_;
      r_11__2__sv2v_reg <= r_n_11__2_;
      r_11__1__sv2v_reg <= r_n_11__1_;
      r_11__0__sv2v_reg <= r_n_11__0_;
    end 
    if(N460) begin
      r_12__15__sv2v_reg <= r_n_12__15_;
      r_12__14__sv2v_reg <= r_n_12__14_;
      r_12__13__sv2v_reg <= r_n_12__13_;
      r_12__12__sv2v_reg <= r_n_12__12_;
      r_12__11__sv2v_reg <= r_n_12__11_;
      r_12__10__sv2v_reg <= r_n_12__10_;
      r_12__9__sv2v_reg <= r_n_12__9_;
      r_12__8__sv2v_reg <= r_n_12__8_;
      r_12__7__sv2v_reg <= r_n_12__7_;
      r_12__6__sv2v_reg <= r_n_12__6_;
      r_12__5__sv2v_reg <= r_n_12__5_;
      r_12__4__sv2v_reg <= r_n_12__4_;
      r_12__3__sv2v_reg <= r_n_12__3_;
      r_12__2__sv2v_reg <= r_n_12__2_;
      r_12__1__sv2v_reg <= r_n_12__1_;
      r_12__0__sv2v_reg <= r_n_12__0_;
    end 
    if(N461) begin
      r_13__15__sv2v_reg <= r_n_13__15_;
      r_13__14__sv2v_reg <= r_n_13__14_;
      r_13__13__sv2v_reg <= r_n_13__13_;
      r_13__12__sv2v_reg <= r_n_13__12_;
      r_13__11__sv2v_reg <= r_n_13__11_;
      r_13__10__sv2v_reg <= r_n_13__10_;
      r_13__9__sv2v_reg <= r_n_13__9_;
      r_13__8__sv2v_reg <= r_n_13__8_;
      r_13__7__sv2v_reg <= r_n_13__7_;
      r_13__6__sv2v_reg <= r_n_13__6_;
      r_13__5__sv2v_reg <= r_n_13__5_;
      r_13__4__sv2v_reg <= r_n_13__4_;
      r_13__3__sv2v_reg <= r_n_13__3_;
      r_13__2__sv2v_reg <= r_n_13__2_;
      r_13__1__sv2v_reg <= r_n_13__1_;
      r_13__0__sv2v_reg <= r_n_13__0_;
    end 
    if(N462) begin
      r_14__15__sv2v_reg <= r_n_14__15_;
      r_14__14__sv2v_reg <= r_n_14__14_;
      r_14__13__sv2v_reg <= r_n_14__13_;
      r_14__12__sv2v_reg <= r_n_14__12_;
      r_14__11__sv2v_reg <= r_n_14__11_;
      r_14__10__sv2v_reg <= r_n_14__10_;
      r_14__9__sv2v_reg <= r_n_14__9_;
      r_14__8__sv2v_reg <= r_n_14__8_;
      r_14__7__sv2v_reg <= r_n_14__7_;
      r_14__6__sv2v_reg <= r_n_14__6_;
      r_14__5__sv2v_reg <= r_n_14__5_;
      r_14__4__sv2v_reg <= r_n_14__4_;
      r_14__3__sv2v_reg <= r_n_14__3_;
      r_14__2__sv2v_reg <= r_n_14__2_;
      r_14__1__sv2v_reg <= r_n_14__1_;
      r_14__0__sv2v_reg <= r_n_14__0_;
    end 
    if(N463) begin
      r_15__15__sv2v_reg <= r_n_15__15_;
      r_15__14__sv2v_reg <= r_n_15__14_;
      r_15__13__sv2v_reg <= r_n_15__13_;
      r_15__12__sv2v_reg <= r_n_15__12_;
      r_15__11__sv2v_reg <= r_n_15__11_;
      r_15__10__sv2v_reg <= r_n_15__10_;
      r_15__9__sv2v_reg <= r_n_15__9_;
      r_15__8__sv2v_reg <= r_n_15__8_;
      r_15__7__sv2v_reg <= r_n_15__7_;
      r_15__6__sv2v_reg <= r_n_15__6_;
      r_15__5__sv2v_reg <= r_n_15__5_;
      r_15__4__sv2v_reg <= r_n_15__4_;
      r_15__3__sv2v_reg <= r_n_15__3_;
      r_15__2__sv2v_reg <= r_n_15__2_;
      r_15__1__sv2v_reg <= r_n_15__1_;
      r_15__0__sv2v_reg <= r_n_15__0_;
    end 
    if(N464) begin
      r_16__15__sv2v_reg <= r_n_16__15_;
      r_16__14__sv2v_reg <= r_n_16__14_;
      r_16__13__sv2v_reg <= r_n_16__13_;
      r_16__12__sv2v_reg <= r_n_16__12_;
      r_16__11__sv2v_reg <= r_n_16__11_;
      r_16__10__sv2v_reg <= r_n_16__10_;
      r_16__9__sv2v_reg <= r_n_16__9_;
      r_16__8__sv2v_reg <= r_n_16__8_;
      r_16__7__sv2v_reg <= r_n_16__7_;
      r_16__6__sv2v_reg <= r_n_16__6_;
      r_16__5__sv2v_reg <= r_n_16__5_;
      r_16__4__sv2v_reg <= r_n_16__4_;
      r_16__3__sv2v_reg <= r_n_16__3_;
      r_16__2__sv2v_reg <= r_n_16__2_;
      r_16__1__sv2v_reg <= r_n_16__1_;
      r_16__0__sv2v_reg <= r_n_16__0_;
    end 
    if(N465) begin
      r_17__15__sv2v_reg <= r_n_17__15_;
      r_17__14__sv2v_reg <= r_n_17__14_;
      r_17__13__sv2v_reg <= r_n_17__13_;
      r_17__12__sv2v_reg <= r_n_17__12_;
      r_17__11__sv2v_reg <= r_n_17__11_;
      r_17__10__sv2v_reg <= r_n_17__10_;
      r_17__9__sv2v_reg <= r_n_17__9_;
      r_17__8__sv2v_reg <= r_n_17__8_;
      r_17__7__sv2v_reg <= r_n_17__7_;
      r_17__6__sv2v_reg <= r_n_17__6_;
      r_17__5__sv2v_reg <= r_n_17__5_;
      r_17__4__sv2v_reg <= r_n_17__4_;
      r_17__3__sv2v_reg <= r_n_17__3_;
      r_17__2__sv2v_reg <= r_n_17__2_;
      r_17__1__sv2v_reg <= r_n_17__1_;
      r_17__0__sv2v_reg <= r_n_17__0_;
    end 
    if(N466) begin
      r_18__15__sv2v_reg <= r_n_18__15_;
      r_18__14__sv2v_reg <= r_n_18__14_;
      r_18__13__sv2v_reg <= r_n_18__13_;
      r_18__12__sv2v_reg <= r_n_18__12_;
      r_18__11__sv2v_reg <= r_n_18__11_;
      r_18__10__sv2v_reg <= r_n_18__10_;
      r_18__9__sv2v_reg <= r_n_18__9_;
      r_18__8__sv2v_reg <= r_n_18__8_;
      r_18__7__sv2v_reg <= r_n_18__7_;
      r_18__6__sv2v_reg <= r_n_18__6_;
      r_18__5__sv2v_reg <= r_n_18__5_;
      r_18__4__sv2v_reg <= r_n_18__4_;
      r_18__3__sv2v_reg <= r_n_18__3_;
      r_18__2__sv2v_reg <= r_n_18__2_;
      r_18__1__sv2v_reg <= r_n_18__1_;
      r_18__0__sv2v_reg <= r_n_18__0_;
    end 
    if(N467) begin
      r_19__15__sv2v_reg <= r_n_19__15_;
      r_19__14__sv2v_reg <= r_n_19__14_;
      r_19__13__sv2v_reg <= r_n_19__13_;
      r_19__12__sv2v_reg <= r_n_19__12_;
      r_19__11__sv2v_reg <= r_n_19__11_;
      r_19__10__sv2v_reg <= r_n_19__10_;
      r_19__9__sv2v_reg <= r_n_19__9_;
      r_19__8__sv2v_reg <= r_n_19__8_;
      r_19__7__sv2v_reg <= r_n_19__7_;
      r_19__6__sv2v_reg <= r_n_19__6_;
      r_19__5__sv2v_reg <= r_n_19__5_;
      r_19__4__sv2v_reg <= r_n_19__4_;
      r_19__3__sv2v_reg <= r_n_19__3_;
      r_19__2__sv2v_reg <= r_n_19__2_;
      r_19__1__sv2v_reg <= r_n_19__1_;
      r_19__0__sv2v_reg <= r_n_19__0_;
    end 
    if(N468) begin
      r_20__15__sv2v_reg <= r_n_20__15_;
      r_20__14__sv2v_reg <= r_n_20__14_;
      r_20__13__sv2v_reg <= r_n_20__13_;
      r_20__12__sv2v_reg <= r_n_20__12_;
      r_20__11__sv2v_reg <= r_n_20__11_;
      r_20__10__sv2v_reg <= r_n_20__10_;
      r_20__9__sv2v_reg <= r_n_20__9_;
      r_20__8__sv2v_reg <= r_n_20__8_;
      r_20__7__sv2v_reg <= r_n_20__7_;
      r_20__6__sv2v_reg <= r_n_20__6_;
      r_20__5__sv2v_reg <= r_n_20__5_;
      r_20__4__sv2v_reg <= r_n_20__4_;
      r_20__3__sv2v_reg <= r_n_20__3_;
      r_20__2__sv2v_reg <= r_n_20__2_;
      r_20__1__sv2v_reg <= r_n_20__1_;
      r_20__0__sv2v_reg <= r_n_20__0_;
    end 
    if(N469) begin
      r_21__15__sv2v_reg <= r_n_21__15_;
      r_21__14__sv2v_reg <= r_n_21__14_;
      r_21__13__sv2v_reg <= r_n_21__13_;
      r_21__12__sv2v_reg <= r_n_21__12_;
      r_21__11__sv2v_reg <= r_n_21__11_;
      r_21__10__sv2v_reg <= r_n_21__10_;
      r_21__9__sv2v_reg <= r_n_21__9_;
      r_21__8__sv2v_reg <= r_n_21__8_;
      r_21__7__sv2v_reg <= r_n_21__7_;
      r_21__6__sv2v_reg <= r_n_21__6_;
      r_21__5__sv2v_reg <= r_n_21__5_;
      r_21__4__sv2v_reg <= r_n_21__4_;
      r_21__3__sv2v_reg <= r_n_21__3_;
      r_21__2__sv2v_reg <= r_n_21__2_;
      r_21__1__sv2v_reg <= r_n_21__1_;
      r_21__0__sv2v_reg <= r_n_21__0_;
    end 
    if(N470) begin
      r_22__15__sv2v_reg <= r_n_22__15_;
      r_22__14__sv2v_reg <= r_n_22__14_;
      r_22__13__sv2v_reg <= r_n_22__13_;
      r_22__12__sv2v_reg <= r_n_22__12_;
      r_22__11__sv2v_reg <= r_n_22__11_;
      r_22__10__sv2v_reg <= r_n_22__10_;
      r_22__9__sv2v_reg <= r_n_22__9_;
      r_22__8__sv2v_reg <= r_n_22__8_;
      r_22__7__sv2v_reg <= r_n_22__7_;
      r_22__6__sv2v_reg <= r_n_22__6_;
      r_22__5__sv2v_reg <= r_n_22__5_;
      r_22__4__sv2v_reg <= r_n_22__4_;
      r_22__3__sv2v_reg <= r_n_22__3_;
      r_22__2__sv2v_reg <= r_n_22__2_;
      r_22__1__sv2v_reg <= r_n_22__1_;
      r_22__0__sv2v_reg <= r_n_22__0_;
    end 
    if(N471) begin
      r_23__15__sv2v_reg <= r_n_23__15_;
      r_23__14__sv2v_reg <= r_n_23__14_;
      r_23__13__sv2v_reg <= r_n_23__13_;
      r_23__12__sv2v_reg <= r_n_23__12_;
      r_23__11__sv2v_reg <= r_n_23__11_;
      r_23__10__sv2v_reg <= r_n_23__10_;
      r_23__9__sv2v_reg <= r_n_23__9_;
      r_23__8__sv2v_reg <= r_n_23__8_;
      r_23__7__sv2v_reg <= r_n_23__7_;
      r_23__6__sv2v_reg <= r_n_23__6_;
      r_23__5__sv2v_reg <= r_n_23__5_;
      r_23__4__sv2v_reg <= r_n_23__4_;
      r_23__3__sv2v_reg <= r_n_23__3_;
      r_23__2__sv2v_reg <= r_n_23__2_;
      r_23__1__sv2v_reg <= r_n_23__1_;
      r_23__0__sv2v_reg <= r_n_23__0_;
    end 
    if(N472) begin
      r_24__15__sv2v_reg <= r_n_24__15_;
      r_24__14__sv2v_reg <= r_n_24__14_;
      r_24__13__sv2v_reg <= r_n_24__13_;
      r_24__12__sv2v_reg <= r_n_24__12_;
      r_24__11__sv2v_reg <= r_n_24__11_;
      r_24__10__sv2v_reg <= r_n_24__10_;
      r_24__9__sv2v_reg <= r_n_24__9_;
      r_24__8__sv2v_reg <= r_n_24__8_;
      r_24__7__sv2v_reg <= r_n_24__7_;
      r_24__6__sv2v_reg <= r_n_24__6_;
      r_24__5__sv2v_reg <= r_n_24__5_;
      r_24__4__sv2v_reg <= r_n_24__4_;
      r_24__3__sv2v_reg <= r_n_24__3_;
      r_24__2__sv2v_reg <= r_n_24__2_;
      r_24__1__sv2v_reg <= r_n_24__1_;
      r_24__0__sv2v_reg <= r_n_24__0_;
    end 
    if(N473) begin
      r_25__15__sv2v_reg <= r_n_25__15_;
      r_25__14__sv2v_reg <= r_n_25__14_;
      r_25__13__sv2v_reg <= r_n_25__13_;
      r_25__12__sv2v_reg <= r_n_25__12_;
      r_25__11__sv2v_reg <= r_n_25__11_;
      r_25__10__sv2v_reg <= r_n_25__10_;
      r_25__9__sv2v_reg <= r_n_25__9_;
      r_25__8__sv2v_reg <= r_n_25__8_;
      r_25__7__sv2v_reg <= r_n_25__7_;
      r_25__6__sv2v_reg <= r_n_25__6_;
      r_25__5__sv2v_reg <= r_n_25__5_;
      r_25__4__sv2v_reg <= r_n_25__4_;
      r_25__3__sv2v_reg <= r_n_25__3_;
      r_25__2__sv2v_reg <= r_n_25__2_;
      r_25__1__sv2v_reg <= r_n_25__1_;
      r_25__0__sv2v_reg <= r_n_25__0_;
    end 
    if(N474) begin
      r_26__15__sv2v_reg <= r_n_26__15_;
      r_26__14__sv2v_reg <= r_n_26__14_;
      r_26__13__sv2v_reg <= r_n_26__13_;
      r_26__12__sv2v_reg <= r_n_26__12_;
      r_26__11__sv2v_reg <= r_n_26__11_;
      r_26__10__sv2v_reg <= r_n_26__10_;
      r_26__9__sv2v_reg <= r_n_26__9_;
      r_26__8__sv2v_reg <= r_n_26__8_;
      r_26__7__sv2v_reg <= r_n_26__7_;
      r_26__6__sv2v_reg <= r_n_26__6_;
      r_26__5__sv2v_reg <= r_n_26__5_;
      r_26__4__sv2v_reg <= r_n_26__4_;
      r_26__3__sv2v_reg <= r_n_26__3_;
      r_26__2__sv2v_reg <= r_n_26__2_;
      r_26__1__sv2v_reg <= r_n_26__1_;
      r_26__0__sv2v_reg <= r_n_26__0_;
    end 
    if(N475) begin
      r_27__15__sv2v_reg <= r_n_27__15_;
      r_27__14__sv2v_reg <= r_n_27__14_;
      r_27__13__sv2v_reg <= r_n_27__13_;
      r_27__12__sv2v_reg <= r_n_27__12_;
      r_27__11__sv2v_reg <= r_n_27__11_;
      r_27__10__sv2v_reg <= r_n_27__10_;
      r_27__9__sv2v_reg <= r_n_27__9_;
      r_27__8__sv2v_reg <= r_n_27__8_;
      r_27__7__sv2v_reg <= r_n_27__7_;
      r_27__6__sv2v_reg <= r_n_27__6_;
      r_27__5__sv2v_reg <= r_n_27__5_;
      r_27__4__sv2v_reg <= r_n_27__4_;
      r_27__3__sv2v_reg <= r_n_27__3_;
      r_27__2__sv2v_reg <= r_n_27__2_;
      r_27__1__sv2v_reg <= r_n_27__1_;
      r_27__0__sv2v_reg <= r_n_27__0_;
    end 
    if(N476) begin
      r_28__15__sv2v_reg <= r_n_28__15_;
      r_28__14__sv2v_reg <= r_n_28__14_;
      r_28__13__sv2v_reg <= r_n_28__13_;
      r_28__12__sv2v_reg <= r_n_28__12_;
      r_28__11__sv2v_reg <= r_n_28__11_;
      r_28__10__sv2v_reg <= r_n_28__10_;
      r_28__9__sv2v_reg <= r_n_28__9_;
      r_28__8__sv2v_reg <= r_n_28__8_;
      r_28__7__sv2v_reg <= r_n_28__7_;
      r_28__6__sv2v_reg <= r_n_28__6_;
      r_28__5__sv2v_reg <= r_n_28__5_;
      r_28__4__sv2v_reg <= r_n_28__4_;
      r_28__3__sv2v_reg <= r_n_28__3_;
      r_28__2__sv2v_reg <= r_n_28__2_;
      r_28__1__sv2v_reg <= r_n_28__1_;
      r_28__0__sv2v_reg <= r_n_28__0_;
    end 
    if(N477) begin
      r_29__15__sv2v_reg <= r_n_29__15_;
      r_29__14__sv2v_reg <= r_n_29__14_;
      r_29__13__sv2v_reg <= r_n_29__13_;
      r_29__12__sv2v_reg <= r_n_29__12_;
      r_29__11__sv2v_reg <= r_n_29__11_;
      r_29__10__sv2v_reg <= r_n_29__10_;
      r_29__9__sv2v_reg <= r_n_29__9_;
      r_29__8__sv2v_reg <= r_n_29__8_;
      r_29__7__sv2v_reg <= r_n_29__7_;
      r_29__6__sv2v_reg <= r_n_29__6_;
      r_29__5__sv2v_reg <= r_n_29__5_;
      r_29__4__sv2v_reg <= r_n_29__4_;
      r_29__3__sv2v_reg <= r_n_29__3_;
      r_29__2__sv2v_reg <= r_n_29__2_;
      r_29__1__sv2v_reg <= r_n_29__1_;
      r_29__0__sv2v_reg <= r_n_29__0_;
    end 
    if(N478) begin
      r_30__15__sv2v_reg <= r_n_30__15_;
      r_30__14__sv2v_reg <= r_n_30__14_;
      r_30__13__sv2v_reg <= r_n_30__13_;
      r_30__12__sv2v_reg <= r_n_30__12_;
      r_30__11__sv2v_reg <= r_n_30__11_;
      r_30__10__sv2v_reg <= r_n_30__10_;
      r_30__9__sv2v_reg <= r_n_30__9_;
      r_30__8__sv2v_reg <= r_n_30__8_;
      r_30__7__sv2v_reg <= r_n_30__7_;
      r_30__6__sv2v_reg <= r_n_30__6_;
      r_30__5__sv2v_reg <= r_n_30__5_;
      r_30__4__sv2v_reg <= r_n_30__4_;
      r_30__3__sv2v_reg <= r_n_30__3_;
      r_30__2__sv2v_reg <= r_n_30__2_;
      r_30__1__sv2v_reg <= r_n_30__1_;
      r_30__0__sv2v_reg <= r_n_30__0_;
    end 
    if(N479) begin
      r_31__15__sv2v_reg <= r_n_31__15_;
      r_31__14__sv2v_reg <= r_n_31__14_;
      r_31__13__sv2v_reg <= r_n_31__13_;
      r_31__12__sv2v_reg <= r_n_31__12_;
      r_31__11__sv2v_reg <= r_n_31__11_;
      r_31__10__sv2v_reg <= r_n_31__10_;
      r_31__9__sv2v_reg <= r_n_31__9_;
      r_31__8__sv2v_reg <= r_n_31__8_;
      r_31__7__sv2v_reg <= r_n_31__7_;
      r_31__6__sv2v_reg <= r_n_31__6_;
      r_31__5__sv2v_reg <= r_n_31__5_;
      r_31__4__sv2v_reg <= r_n_31__4_;
      r_31__3__sv2v_reg <= r_n_31__3_;
      r_31__2__sv2v_reg <= r_n_31__2_;
      r_31__1__sv2v_reg <= r_n_31__1_;
      r_31__0__sv2v_reg <= r_n_31__0_;
    end 
    if(N480) begin
      r_32__15__sv2v_reg <= r_n_32__15_;
      r_32__14__sv2v_reg <= r_n_32__14_;
      r_32__13__sv2v_reg <= r_n_32__13_;
      r_32__12__sv2v_reg <= r_n_32__12_;
      r_32__11__sv2v_reg <= r_n_32__11_;
      r_32__10__sv2v_reg <= r_n_32__10_;
      r_32__9__sv2v_reg <= r_n_32__9_;
      r_32__8__sv2v_reg <= r_n_32__8_;
      r_32__7__sv2v_reg <= r_n_32__7_;
      r_32__6__sv2v_reg <= r_n_32__6_;
      r_32__5__sv2v_reg <= r_n_32__5_;
      r_32__4__sv2v_reg <= r_n_32__4_;
      r_32__3__sv2v_reg <= r_n_32__3_;
      r_32__2__sv2v_reg <= r_n_32__2_;
      r_32__1__sv2v_reg <= r_n_32__1_;
      r_32__0__sv2v_reg <= r_n_32__0_;
    end 
    if(N481) begin
      r_33__15__sv2v_reg <= r_n_33__15_;
      r_33__14__sv2v_reg <= r_n_33__14_;
      r_33__13__sv2v_reg <= r_n_33__13_;
      r_33__12__sv2v_reg <= r_n_33__12_;
      r_33__11__sv2v_reg <= r_n_33__11_;
      r_33__10__sv2v_reg <= r_n_33__10_;
      r_33__9__sv2v_reg <= r_n_33__9_;
      r_33__8__sv2v_reg <= r_n_33__8_;
      r_33__7__sv2v_reg <= r_n_33__7_;
      r_33__6__sv2v_reg <= r_n_33__6_;
      r_33__5__sv2v_reg <= r_n_33__5_;
      r_33__4__sv2v_reg <= r_n_33__4_;
      r_33__3__sv2v_reg <= r_n_33__3_;
      r_33__2__sv2v_reg <= r_n_33__2_;
      r_33__1__sv2v_reg <= r_n_33__1_;
      r_33__0__sv2v_reg <= r_n_33__0_;
    end 
    if(N482) begin
      r_34__15__sv2v_reg <= r_n_34__15_;
      r_34__14__sv2v_reg <= r_n_34__14_;
      r_34__13__sv2v_reg <= r_n_34__13_;
      r_34__12__sv2v_reg <= r_n_34__12_;
      r_34__11__sv2v_reg <= r_n_34__11_;
      r_34__10__sv2v_reg <= r_n_34__10_;
      r_34__9__sv2v_reg <= r_n_34__9_;
      r_34__8__sv2v_reg <= r_n_34__8_;
      r_34__7__sv2v_reg <= r_n_34__7_;
      r_34__6__sv2v_reg <= r_n_34__6_;
      r_34__5__sv2v_reg <= r_n_34__5_;
      r_34__4__sv2v_reg <= r_n_34__4_;
      r_34__3__sv2v_reg <= r_n_34__3_;
      r_34__2__sv2v_reg <= r_n_34__2_;
      r_34__1__sv2v_reg <= r_n_34__1_;
      r_34__0__sv2v_reg <= r_n_34__0_;
    end 
    if(N483) begin
      r_35__15__sv2v_reg <= r_n_35__15_;
      r_35__14__sv2v_reg <= r_n_35__14_;
      r_35__13__sv2v_reg <= r_n_35__13_;
      r_35__12__sv2v_reg <= r_n_35__12_;
      r_35__11__sv2v_reg <= r_n_35__11_;
      r_35__10__sv2v_reg <= r_n_35__10_;
      r_35__9__sv2v_reg <= r_n_35__9_;
      r_35__8__sv2v_reg <= r_n_35__8_;
      r_35__7__sv2v_reg <= r_n_35__7_;
      r_35__6__sv2v_reg <= r_n_35__6_;
      r_35__5__sv2v_reg <= r_n_35__5_;
      r_35__4__sv2v_reg <= r_n_35__4_;
      r_35__3__sv2v_reg <= r_n_35__3_;
      r_35__2__sv2v_reg <= r_n_35__2_;
      r_35__1__sv2v_reg <= r_n_35__1_;
      r_35__0__sv2v_reg <= r_n_35__0_;
    end 
    if(N484) begin
      r_36__15__sv2v_reg <= r_n_36__15_;
      r_36__14__sv2v_reg <= r_n_36__14_;
      r_36__13__sv2v_reg <= r_n_36__13_;
      r_36__12__sv2v_reg <= r_n_36__12_;
      r_36__11__sv2v_reg <= r_n_36__11_;
      r_36__10__sv2v_reg <= r_n_36__10_;
      r_36__9__sv2v_reg <= r_n_36__9_;
      r_36__8__sv2v_reg <= r_n_36__8_;
      r_36__7__sv2v_reg <= r_n_36__7_;
      r_36__6__sv2v_reg <= r_n_36__6_;
      r_36__5__sv2v_reg <= r_n_36__5_;
      r_36__4__sv2v_reg <= r_n_36__4_;
      r_36__3__sv2v_reg <= r_n_36__3_;
      r_36__2__sv2v_reg <= r_n_36__2_;
      r_36__1__sv2v_reg <= r_n_36__1_;
      r_36__0__sv2v_reg <= r_n_36__0_;
    end 
    if(N485) begin
      r_37__15__sv2v_reg <= r_n_37__15_;
      r_37__14__sv2v_reg <= r_n_37__14_;
      r_37__13__sv2v_reg <= r_n_37__13_;
      r_37__12__sv2v_reg <= r_n_37__12_;
      r_37__11__sv2v_reg <= r_n_37__11_;
      r_37__10__sv2v_reg <= r_n_37__10_;
      r_37__9__sv2v_reg <= r_n_37__9_;
      r_37__8__sv2v_reg <= r_n_37__8_;
      r_37__7__sv2v_reg <= r_n_37__7_;
      r_37__6__sv2v_reg <= r_n_37__6_;
      r_37__5__sv2v_reg <= r_n_37__5_;
      r_37__4__sv2v_reg <= r_n_37__4_;
      r_37__3__sv2v_reg <= r_n_37__3_;
      r_37__2__sv2v_reg <= r_n_37__2_;
      r_37__1__sv2v_reg <= r_n_37__1_;
      r_37__0__sv2v_reg <= r_n_37__0_;
    end 
    if(N486) begin
      r_38__15__sv2v_reg <= r_n_38__15_;
      r_38__14__sv2v_reg <= r_n_38__14_;
      r_38__13__sv2v_reg <= r_n_38__13_;
      r_38__12__sv2v_reg <= r_n_38__12_;
      r_38__11__sv2v_reg <= r_n_38__11_;
      r_38__10__sv2v_reg <= r_n_38__10_;
      r_38__9__sv2v_reg <= r_n_38__9_;
      r_38__8__sv2v_reg <= r_n_38__8_;
      r_38__7__sv2v_reg <= r_n_38__7_;
      r_38__6__sv2v_reg <= r_n_38__6_;
      r_38__5__sv2v_reg <= r_n_38__5_;
      r_38__4__sv2v_reg <= r_n_38__4_;
      r_38__3__sv2v_reg <= r_n_38__3_;
      r_38__2__sv2v_reg <= r_n_38__2_;
      r_38__1__sv2v_reg <= r_n_38__1_;
      r_38__0__sv2v_reg <= r_n_38__0_;
    end 
    if(N487) begin
      r_39__15__sv2v_reg <= r_n_39__15_;
      r_39__14__sv2v_reg <= r_n_39__14_;
      r_39__13__sv2v_reg <= r_n_39__13_;
      r_39__12__sv2v_reg <= r_n_39__12_;
      r_39__11__sv2v_reg <= r_n_39__11_;
      r_39__10__sv2v_reg <= r_n_39__10_;
      r_39__9__sv2v_reg <= r_n_39__9_;
      r_39__8__sv2v_reg <= r_n_39__8_;
      r_39__7__sv2v_reg <= r_n_39__7_;
      r_39__6__sv2v_reg <= r_n_39__6_;
      r_39__5__sv2v_reg <= r_n_39__5_;
      r_39__4__sv2v_reg <= r_n_39__4_;
      r_39__3__sv2v_reg <= r_n_39__3_;
      r_39__2__sv2v_reg <= r_n_39__2_;
      r_39__1__sv2v_reg <= r_n_39__1_;
      r_39__0__sv2v_reg <= r_n_39__0_;
    end 
    if(N488) begin
      r_40__15__sv2v_reg <= r_n_40__15_;
      r_40__14__sv2v_reg <= r_n_40__14_;
      r_40__13__sv2v_reg <= r_n_40__13_;
      r_40__12__sv2v_reg <= r_n_40__12_;
      r_40__11__sv2v_reg <= r_n_40__11_;
      r_40__10__sv2v_reg <= r_n_40__10_;
      r_40__9__sv2v_reg <= r_n_40__9_;
      r_40__8__sv2v_reg <= r_n_40__8_;
      r_40__7__sv2v_reg <= r_n_40__7_;
      r_40__6__sv2v_reg <= r_n_40__6_;
      r_40__5__sv2v_reg <= r_n_40__5_;
      r_40__4__sv2v_reg <= r_n_40__4_;
      r_40__3__sv2v_reg <= r_n_40__3_;
      r_40__2__sv2v_reg <= r_n_40__2_;
      r_40__1__sv2v_reg <= r_n_40__1_;
      r_40__0__sv2v_reg <= r_n_40__0_;
    end 
    if(N489) begin
      r_41__15__sv2v_reg <= r_n_41__15_;
      r_41__14__sv2v_reg <= r_n_41__14_;
      r_41__13__sv2v_reg <= r_n_41__13_;
      r_41__12__sv2v_reg <= r_n_41__12_;
      r_41__11__sv2v_reg <= r_n_41__11_;
      r_41__10__sv2v_reg <= r_n_41__10_;
      r_41__9__sv2v_reg <= r_n_41__9_;
      r_41__8__sv2v_reg <= r_n_41__8_;
      r_41__7__sv2v_reg <= r_n_41__7_;
      r_41__6__sv2v_reg <= r_n_41__6_;
      r_41__5__sv2v_reg <= r_n_41__5_;
      r_41__4__sv2v_reg <= r_n_41__4_;
      r_41__3__sv2v_reg <= r_n_41__3_;
      r_41__2__sv2v_reg <= r_n_41__2_;
      r_41__1__sv2v_reg <= r_n_41__1_;
      r_41__0__sv2v_reg <= r_n_41__0_;
    end 
    if(N490) begin
      r_42__15__sv2v_reg <= r_n_42__15_;
      r_42__14__sv2v_reg <= r_n_42__14_;
      r_42__13__sv2v_reg <= r_n_42__13_;
      r_42__12__sv2v_reg <= r_n_42__12_;
      r_42__11__sv2v_reg <= r_n_42__11_;
      r_42__10__sv2v_reg <= r_n_42__10_;
      r_42__9__sv2v_reg <= r_n_42__9_;
      r_42__8__sv2v_reg <= r_n_42__8_;
      r_42__7__sv2v_reg <= r_n_42__7_;
      r_42__6__sv2v_reg <= r_n_42__6_;
      r_42__5__sv2v_reg <= r_n_42__5_;
      r_42__4__sv2v_reg <= r_n_42__4_;
      r_42__3__sv2v_reg <= r_n_42__3_;
      r_42__2__sv2v_reg <= r_n_42__2_;
      r_42__1__sv2v_reg <= r_n_42__1_;
      r_42__0__sv2v_reg <= r_n_42__0_;
    end 
    if(N491) begin
      r_43__15__sv2v_reg <= r_n_43__15_;
      r_43__14__sv2v_reg <= r_n_43__14_;
      r_43__13__sv2v_reg <= r_n_43__13_;
      r_43__12__sv2v_reg <= r_n_43__12_;
      r_43__11__sv2v_reg <= r_n_43__11_;
      r_43__10__sv2v_reg <= r_n_43__10_;
      r_43__9__sv2v_reg <= r_n_43__9_;
      r_43__8__sv2v_reg <= r_n_43__8_;
      r_43__7__sv2v_reg <= r_n_43__7_;
      r_43__6__sv2v_reg <= r_n_43__6_;
      r_43__5__sv2v_reg <= r_n_43__5_;
      r_43__4__sv2v_reg <= r_n_43__4_;
      r_43__3__sv2v_reg <= r_n_43__3_;
      r_43__2__sv2v_reg <= r_n_43__2_;
      r_43__1__sv2v_reg <= r_n_43__1_;
      r_43__0__sv2v_reg <= r_n_43__0_;
    end 
    if(N492) begin
      r_44__15__sv2v_reg <= r_n_44__15_;
      r_44__14__sv2v_reg <= r_n_44__14_;
      r_44__13__sv2v_reg <= r_n_44__13_;
      r_44__12__sv2v_reg <= r_n_44__12_;
      r_44__11__sv2v_reg <= r_n_44__11_;
      r_44__10__sv2v_reg <= r_n_44__10_;
      r_44__9__sv2v_reg <= r_n_44__9_;
      r_44__8__sv2v_reg <= r_n_44__8_;
      r_44__7__sv2v_reg <= r_n_44__7_;
      r_44__6__sv2v_reg <= r_n_44__6_;
      r_44__5__sv2v_reg <= r_n_44__5_;
      r_44__4__sv2v_reg <= r_n_44__4_;
      r_44__3__sv2v_reg <= r_n_44__3_;
      r_44__2__sv2v_reg <= r_n_44__2_;
      r_44__1__sv2v_reg <= r_n_44__1_;
      r_44__0__sv2v_reg <= r_n_44__0_;
    end 
    if(N493) begin
      r_45__15__sv2v_reg <= r_n_45__15_;
      r_45__14__sv2v_reg <= r_n_45__14_;
      r_45__13__sv2v_reg <= r_n_45__13_;
      r_45__12__sv2v_reg <= r_n_45__12_;
      r_45__11__sv2v_reg <= r_n_45__11_;
      r_45__10__sv2v_reg <= r_n_45__10_;
      r_45__9__sv2v_reg <= r_n_45__9_;
      r_45__8__sv2v_reg <= r_n_45__8_;
      r_45__7__sv2v_reg <= r_n_45__7_;
      r_45__6__sv2v_reg <= r_n_45__6_;
      r_45__5__sv2v_reg <= r_n_45__5_;
      r_45__4__sv2v_reg <= r_n_45__4_;
      r_45__3__sv2v_reg <= r_n_45__3_;
      r_45__2__sv2v_reg <= r_n_45__2_;
      r_45__1__sv2v_reg <= r_n_45__1_;
      r_45__0__sv2v_reg <= r_n_45__0_;
    end 
    if(N494) begin
      r_46__15__sv2v_reg <= r_n_46__15_;
      r_46__14__sv2v_reg <= r_n_46__14_;
      r_46__13__sv2v_reg <= r_n_46__13_;
      r_46__12__sv2v_reg <= r_n_46__12_;
      r_46__11__sv2v_reg <= r_n_46__11_;
      r_46__10__sv2v_reg <= r_n_46__10_;
      r_46__9__sv2v_reg <= r_n_46__9_;
      r_46__8__sv2v_reg <= r_n_46__8_;
      r_46__7__sv2v_reg <= r_n_46__7_;
      r_46__6__sv2v_reg <= r_n_46__6_;
      r_46__5__sv2v_reg <= r_n_46__5_;
      r_46__4__sv2v_reg <= r_n_46__4_;
      r_46__3__sv2v_reg <= r_n_46__3_;
      r_46__2__sv2v_reg <= r_n_46__2_;
      r_46__1__sv2v_reg <= r_n_46__1_;
      r_46__0__sv2v_reg <= r_n_46__0_;
    end 
    if(N495) begin
      r_47__15__sv2v_reg <= r_n_47__15_;
      r_47__14__sv2v_reg <= r_n_47__14_;
      r_47__13__sv2v_reg <= r_n_47__13_;
      r_47__12__sv2v_reg <= r_n_47__12_;
      r_47__11__sv2v_reg <= r_n_47__11_;
      r_47__10__sv2v_reg <= r_n_47__10_;
      r_47__9__sv2v_reg <= r_n_47__9_;
      r_47__8__sv2v_reg <= r_n_47__8_;
      r_47__7__sv2v_reg <= r_n_47__7_;
      r_47__6__sv2v_reg <= r_n_47__6_;
      r_47__5__sv2v_reg <= r_n_47__5_;
      r_47__4__sv2v_reg <= r_n_47__4_;
      r_47__3__sv2v_reg <= r_n_47__3_;
      r_47__2__sv2v_reg <= r_n_47__2_;
      r_47__1__sv2v_reg <= r_n_47__1_;
      r_47__0__sv2v_reg <= r_n_47__0_;
    end 
    if(N496) begin
      r_48__15__sv2v_reg <= r_n_48__15_;
      r_48__14__sv2v_reg <= r_n_48__14_;
      r_48__13__sv2v_reg <= r_n_48__13_;
      r_48__12__sv2v_reg <= r_n_48__12_;
      r_48__11__sv2v_reg <= r_n_48__11_;
      r_48__10__sv2v_reg <= r_n_48__10_;
      r_48__9__sv2v_reg <= r_n_48__9_;
      r_48__8__sv2v_reg <= r_n_48__8_;
      r_48__7__sv2v_reg <= r_n_48__7_;
      r_48__6__sv2v_reg <= r_n_48__6_;
      r_48__5__sv2v_reg <= r_n_48__5_;
      r_48__4__sv2v_reg <= r_n_48__4_;
      r_48__3__sv2v_reg <= r_n_48__3_;
      r_48__2__sv2v_reg <= r_n_48__2_;
      r_48__1__sv2v_reg <= r_n_48__1_;
      r_48__0__sv2v_reg <= r_n_48__0_;
    end 
    if(N497) begin
      r_49__15__sv2v_reg <= r_n_49__15_;
      r_49__14__sv2v_reg <= r_n_49__14_;
      r_49__13__sv2v_reg <= r_n_49__13_;
      r_49__12__sv2v_reg <= r_n_49__12_;
      r_49__11__sv2v_reg <= r_n_49__11_;
      r_49__10__sv2v_reg <= r_n_49__10_;
      r_49__9__sv2v_reg <= r_n_49__9_;
      r_49__8__sv2v_reg <= r_n_49__8_;
      r_49__7__sv2v_reg <= r_n_49__7_;
      r_49__6__sv2v_reg <= r_n_49__6_;
      r_49__5__sv2v_reg <= r_n_49__5_;
      r_49__4__sv2v_reg <= r_n_49__4_;
      r_49__3__sv2v_reg <= r_n_49__3_;
      r_49__2__sv2v_reg <= r_n_49__2_;
      r_49__1__sv2v_reg <= r_n_49__1_;
      r_49__0__sv2v_reg <= r_n_49__0_;
    end 
    if(N498) begin
      r_50__15__sv2v_reg <= r_n_50__15_;
      r_50__14__sv2v_reg <= r_n_50__14_;
      r_50__13__sv2v_reg <= r_n_50__13_;
      r_50__12__sv2v_reg <= r_n_50__12_;
      r_50__11__sv2v_reg <= r_n_50__11_;
      r_50__10__sv2v_reg <= r_n_50__10_;
      r_50__9__sv2v_reg <= r_n_50__9_;
      r_50__8__sv2v_reg <= r_n_50__8_;
      r_50__7__sv2v_reg <= r_n_50__7_;
      r_50__6__sv2v_reg <= r_n_50__6_;
      r_50__5__sv2v_reg <= r_n_50__5_;
      r_50__4__sv2v_reg <= r_n_50__4_;
      r_50__3__sv2v_reg <= r_n_50__3_;
      r_50__2__sv2v_reg <= r_n_50__2_;
      r_50__1__sv2v_reg <= r_n_50__1_;
      r_50__0__sv2v_reg <= r_n_50__0_;
    end 
    if(N499) begin
      r_51__15__sv2v_reg <= r_n_51__15_;
      r_51__14__sv2v_reg <= r_n_51__14_;
      r_51__13__sv2v_reg <= r_n_51__13_;
      r_51__12__sv2v_reg <= r_n_51__12_;
      r_51__11__sv2v_reg <= r_n_51__11_;
      r_51__10__sv2v_reg <= r_n_51__10_;
      r_51__9__sv2v_reg <= r_n_51__9_;
      r_51__8__sv2v_reg <= r_n_51__8_;
      r_51__7__sv2v_reg <= r_n_51__7_;
      r_51__6__sv2v_reg <= r_n_51__6_;
      r_51__5__sv2v_reg <= r_n_51__5_;
      r_51__4__sv2v_reg <= r_n_51__4_;
      r_51__3__sv2v_reg <= r_n_51__3_;
      r_51__2__sv2v_reg <= r_n_51__2_;
      r_51__1__sv2v_reg <= r_n_51__1_;
      r_51__0__sv2v_reg <= r_n_51__0_;
    end 
    if(N500) begin
      r_52__15__sv2v_reg <= r_n_52__15_;
      r_52__14__sv2v_reg <= r_n_52__14_;
      r_52__13__sv2v_reg <= r_n_52__13_;
      r_52__12__sv2v_reg <= r_n_52__12_;
      r_52__11__sv2v_reg <= r_n_52__11_;
      r_52__10__sv2v_reg <= r_n_52__10_;
      r_52__9__sv2v_reg <= r_n_52__9_;
      r_52__8__sv2v_reg <= r_n_52__8_;
      r_52__7__sv2v_reg <= r_n_52__7_;
      r_52__6__sv2v_reg <= r_n_52__6_;
      r_52__5__sv2v_reg <= r_n_52__5_;
      r_52__4__sv2v_reg <= r_n_52__4_;
      r_52__3__sv2v_reg <= r_n_52__3_;
      r_52__2__sv2v_reg <= r_n_52__2_;
      r_52__1__sv2v_reg <= r_n_52__1_;
      r_52__0__sv2v_reg <= r_n_52__0_;
    end 
    if(N501) begin
      r_53__15__sv2v_reg <= r_n_53__15_;
      r_53__14__sv2v_reg <= r_n_53__14_;
      r_53__13__sv2v_reg <= r_n_53__13_;
      r_53__12__sv2v_reg <= r_n_53__12_;
      r_53__11__sv2v_reg <= r_n_53__11_;
      r_53__10__sv2v_reg <= r_n_53__10_;
      r_53__9__sv2v_reg <= r_n_53__9_;
      r_53__8__sv2v_reg <= r_n_53__8_;
      r_53__7__sv2v_reg <= r_n_53__7_;
      r_53__6__sv2v_reg <= r_n_53__6_;
      r_53__5__sv2v_reg <= r_n_53__5_;
      r_53__4__sv2v_reg <= r_n_53__4_;
      r_53__3__sv2v_reg <= r_n_53__3_;
      r_53__2__sv2v_reg <= r_n_53__2_;
      r_53__1__sv2v_reg <= r_n_53__1_;
      r_53__0__sv2v_reg <= r_n_53__0_;
    end 
    if(N502) begin
      r_54__15__sv2v_reg <= r_n_54__15_;
      r_54__14__sv2v_reg <= r_n_54__14_;
      r_54__13__sv2v_reg <= r_n_54__13_;
      r_54__12__sv2v_reg <= r_n_54__12_;
      r_54__11__sv2v_reg <= r_n_54__11_;
      r_54__10__sv2v_reg <= r_n_54__10_;
      r_54__9__sv2v_reg <= r_n_54__9_;
      r_54__8__sv2v_reg <= r_n_54__8_;
      r_54__7__sv2v_reg <= r_n_54__7_;
      r_54__6__sv2v_reg <= r_n_54__6_;
      r_54__5__sv2v_reg <= r_n_54__5_;
      r_54__4__sv2v_reg <= r_n_54__4_;
      r_54__3__sv2v_reg <= r_n_54__3_;
      r_54__2__sv2v_reg <= r_n_54__2_;
      r_54__1__sv2v_reg <= r_n_54__1_;
      r_54__0__sv2v_reg <= r_n_54__0_;
    end 
    if(N503) begin
      r_55__15__sv2v_reg <= r_n_55__15_;
      r_55__14__sv2v_reg <= r_n_55__14_;
      r_55__13__sv2v_reg <= r_n_55__13_;
      r_55__12__sv2v_reg <= r_n_55__12_;
      r_55__11__sv2v_reg <= r_n_55__11_;
      r_55__10__sv2v_reg <= r_n_55__10_;
      r_55__9__sv2v_reg <= r_n_55__9_;
      r_55__8__sv2v_reg <= r_n_55__8_;
      r_55__7__sv2v_reg <= r_n_55__7_;
      r_55__6__sv2v_reg <= r_n_55__6_;
      r_55__5__sv2v_reg <= r_n_55__5_;
      r_55__4__sv2v_reg <= r_n_55__4_;
      r_55__3__sv2v_reg <= r_n_55__3_;
      r_55__2__sv2v_reg <= r_n_55__2_;
      r_55__1__sv2v_reg <= r_n_55__1_;
      r_55__0__sv2v_reg <= r_n_55__0_;
    end 
    if(N504) begin
      r_56__15__sv2v_reg <= r_n_56__15_;
      r_56__14__sv2v_reg <= r_n_56__14_;
      r_56__13__sv2v_reg <= r_n_56__13_;
      r_56__12__sv2v_reg <= r_n_56__12_;
      r_56__11__sv2v_reg <= r_n_56__11_;
      r_56__10__sv2v_reg <= r_n_56__10_;
      r_56__9__sv2v_reg <= r_n_56__9_;
      r_56__8__sv2v_reg <= r_n_56__8_;
      r_56__7__sv2v_reg <= r_n_56__7_;
      r_56__6__sv2v_reg <= r_n_56__6_;
      r_56__5__sv2v_reg <= r_n_56__5_;
      r_56__4__sv2v_reg <= r_n_56__4_;
      r_56__3__sv2v_reg <= r_n_56__3_;
      r_56__2__sv2v_reg <= r_n_56__2_;
      r_56__1__sv2v_reg <= r_n_56__1_;
      r_56__0__sv2v_reg <= r_n_56__0_;
    end 
    if(N505) begin
      r_57__15__sv2v_reg <= r_n_57__15_;
      r_57__14__sv2v_reg <= r_n_57__14_;
      r_57__13__sv2v_reg <= r_n_57__13_;
      r_57__12__sv2v_reg <= r_n_57__12_;
      r_57__11__sv2v_reg <= r_n_57__11_;
      r_57__10__sv2v_reg <= r_n_57__10_;
      r_57__9__sv2v_reg <= r_n_57__9_;
      r_57__8__sv2v_reg <= r_n_57__8_;
      r_57__7__sv2v_reg <= r_n_57__7_;
      r_57__6__sv2v_reg <= r_n_57__6_;
      r_57__5__sv2v_reg <= r_n_57__5_;
      r_57__4__sv2v_reg <= r_n_57__4_;
      r_57__3__sv2v_reg <= r_n_57__3_;
      r_57__2__sv2v_reg <= r_n_57__2_;
      r_57__1__sv2v_reg <= r_n_57__1_;
      r_57__0__sv2v_reg <= r_n_57__0_;
    end 
    if(N506) begin
      r_58__15__sv2v_reg <= r_n_58__15_;
      r_58__14__sv2v_reg <= r_n_58__14_;
      r_58__13__sv2v_reg <= r_n_58__13_;
      r_58__12__sv2v_reg <= r_n_58__12_;
      r_58__11__sv2v_reg <= r_n_58__11_;
      r_58__10__sv2v_reg <= r_n_58__10_;
      r_58__9__sv2v_reg <= r_n_58__9_;
      r_58__8__sv2v_reg <= r_n_58__8_;
      r_58__7__sv2v_reg <= r_n_58__7_;
      r_58__6__sv2v_reg <= r_n_58__6_;
      r_58__5__sv2v_reg <= r_n_58__5_;
      r_58__4__sv2v_reg <= r_n_58__4_;
      r_58__3__sv2v_reg <= r_n_58__3_;
      r_58__2__sv2v_reg <= r_n_58__2_;
      r_58__1__sv2v_reg <= r_n_58__1_;
      r_58__0__sv2v_reg <= r_n_58__0_;
    end 
    if(N507) begin
      r_59__15__sv2v_reg <= r_n_59__15_;
      r_59__14__sv2v_reg <= r_n_59__14_;
      r_59__13__sv2v_reg <= r_n_59__13_;
      r_59__12__sv2v_reg <= r_n_59__12_;
      r_59__11__sv2v_reg <= r_n_59__11_;
      r_59__10__sv2v_reg <= r_n_59__10_;
      r_59__9__sv2v_reg <= r_n_59__9_;
      r_59__8__sv2v_reg <= r_n_59__8_;
      r_59__7__sv2v_reg <= r_n_59__7_;
      r_59__6__sv2v_reg <= r_n_59__6_;
      r_59__5__sv2v_reg <= r_n_59__5_;
      r_59__4__sv2v_reg <= r_n_59__4_;
      r_59__3__sv2v_reg <= r_n_59__3_;
      r_59__2__sv2v_reg <= r_n_59__2_;
      r_59__1__sv2v_reg <= r_n_59__1_;
      r_59__0__sv2v_reg <= r_n_59__0_;
    end 
    if(N508) begin
      r_60__15__sv2v_reg <= r_n_60__15_;
      r_60__14__sv2v_reg <= r_n_60__14_;
      r_60__13__sv2v_reg <= r_n_60__13_;
      r_60__12__sv2v_reg <= r_n_60__12_;
      r_60__11__sv2v_reg <= r_n_60__11_;
      r_60__10__sv2v_reg <= r_n_60__10_;
      r_60__9__sv2v_reg <= r_n_60__9_;
      r_60__8__sv2v_reg <= r_n_60__8_;
      r_60__7__sv2v_reg <= r_n_60__7_;
      r_60__6__sv2v_reg <= r_n_60__6_;
      r_60__5__sv2v_reg <= r_n_60__5_;
      r_60__4__sv2v_reg <= r_n_60__4_;
      r_60__3__sv2v_reg <= r_n_60__3_;
      r_60__2__sv2v_reg <= r_n_60__2_;
      r_60__1__sv2v_reg <= r_n_60__1_;
      r_60__0__sv2v_reg <= r_n_60__0_;
    end 
    if(N509) begin
      r_61__15__sv2v_reg <= r_n_61__15_;
      r_61__14__sv2v_reg <= r_n_61__14_;
      r_61__13__sv2v_reg <= r_n_61__13_;
      r_61__12__sv2v_reg <= r_n_61__12_;
      r_61__11__sv2v_reg <= r_n_61__11_;
      r_61__10__sv2v_reg <= r_n_61__10_;
      r_61__9__sv2v_reg <= r_n_61__9_;
      r_61__8__sv2v_reg <= r_n_61__8_;
      r_61__7__sv2v_reg <= r_n_61__7_;
      r_61__6__sv2v_reg <= r_n_61__6_;
      r_61__5__sv2v_reg <= r_n_61__5_;
      r_61__4__sv2v_reg <= r_n_61__4_;
      r_61__3__sv2v_reg <= r_n_61__3_;
      r_61__2__sv2v_reg <= r_n_61__2_;
      r_61__1__sv2v_reg <= r_n_61__1_;
      r_61__0__sv2v_reg <= r_n_61__0_;
    end 
    if(N510) begin
      r_62__15__sv2v_reg <= r_n_62__15_;
      r_62__14__sv2v_reg <= r_n_62__14_;
      r_62__13__sv2v_reg <= r_n_62__13_;
      r_62__12__sv2v_reg <= r_n_62__12_;
      r_62__11__sv2v_reg <= r_n_62__11_;
      r_62__10__sv2v_reg <= r_n_62__10_;
      r_62__9__sv2v_reg <= r_n_62__9_;
      r_62__8__sv2v_reg <= r_n_62__8_;
      r_62__7__sv2v_reg <= r_n_62__7_;
      r_62__6__sv2v_reg <= r_n_62__6_;
      r_62__5__sv2v_reg <= r_n_62__5_;
      r_62__4__sv2v_reg <= r_n_62__4_;
      r_62__3__sv2v_reg <= r_n_62__3_;
      r_62__2__sv2v_reg <= r_n_62__2_;
      r_62__1__sv2v_reg <= r_n_62__1_;
      r_62__0__sv2v_reg <= r_n_62__0_;
    end 
    if(N443) begin
      r_63__15__sv2v_reg <= 1'b0;
      r_63__14__sv2v_reg <= 1'b0;
      r_63__13__sv2v_reg <= 1'b0;
      r_63__12__sv2v_reg <= 1'b0;
      r_63__11__sv2v_reg <= 1'b0;
      r_63__10__sv2v_reg <= 1'b0;
      r_63__9__sv2v_reg <= 1'b0;
      r_63__8__sv2v_reg <= 1'b0;
      r_63__7__sv2v_reg <= 1'b0;
      r_63__6__sv2v_reg <= 1'b0;
      r_63__5__sv2v_reg <= 1'b0;
      r_63__4__sv2v_reg <= 1'b0;
      r_63__3__sv2v_reg <= 1'b0;
      r_63__2__sv2v_reg <= 1'b0;
      r_63__1__sv2v_reg <= 1'b0;
      r_63__0__sv2v_reg <= 1'b0;
    end else if(N511) begin
      r_63__15__sv2v_reg <= data_i[15];
      r_63__14__sv2v_reg <= data_i[14];
      r_63__13__sv2v_reg <= data_i[13];
      r_63__12__sv2v_reg <= data_i[12];
      r_63__11__sv2v_reg <= data_i[11];
      r_63__10__sv2v_reg <= data_i[10];
      r_63__9__sv2v_reg <= data_i[9];
      r_63__8__sv2v_reg <= data_i[8];
      r_63__7__sv2v_reg <= data_i[7];
      r_63__6__sv2v_reg <= data_i[6];
      r_63__5__sv2v_reg <= data_i[5];
      r_63__4__sv2v_reg <= data_i[4];
      r_63__3__sv2v_reg <= data_i[3];
      r_63__2__sv2v_reg <= data_i[2];
      r_63__1__sv2v_reg <= data_i[1];
      r_63__0__sv2v_reg <= data_i[0];
    end 
  end


endmodule

