

module top
(
  L_clk_i,
  L_reset_i,
  L_en_o,
  L_v_o,
  L_data_o,
  L_ready_i,
  L_v_i,
  L_data_i,
  L_yumi_o,
  R_clk_i,
  R_reset_i,
  R_en_i,
  R_v_i,
  R_data_i,
  R_ready_o,
  R_v_o,
  R_data_o,
  R_yumi_i
);

  output [49:0] L_data_o;
  input [49:0] L_data_i;
  input [49:0] R_data_i;
  output [49:0] R_data_o;
  input L_clk_i;
  input L_reset_i;
  input L_ready_i;
  input L_v_i;
  input R_clk_i;
  input R_reset_i;
  input R_en_i;
  input R_v_i;
  input R_yumi_i;
  output L_en_o;
  output L_v_o;
  output L_yumi_o;
  output R_ready_o;
  output R_v_o;

  bsg_fsb_node_async_buffer
  wrapper
  (
    .L_data_o(L_data_o),
    .L_data_i(L_data_i),
    .R_data_i(R_data_i),
    .R_data_o(R_data_o),
    .L_clk_i(L_clk_i),
    .L_reset_i(L_reset_i),
    .L_ready_i(L_ready_i),
    .L_v_i(L_v_i),
    .R_clk_i(R_clk_i),
    .R_reset_i(R_reset_i),
    .R_en_i(R_en_i),
    .R_v_i(R_v_i),
    .R_yumi_i(R_yumi_i),
    .L_en_o(L_en_o),
    .L_v_o(L_v_o),
    .L_yumi_o(L_yumi_o),
    .R_ready_o(R_ready_o),
    .R_v_o(R_v_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p50_els_p64_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [49:0] w_data_i;
  input [5:0] r_addr_i;
  output [49:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [49:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294;
  reg [3199:0] mem;
  assign r_data_o[49] = (N76)? mem[49] : 
                        (N78)? mem[99] : 
                        (N80)? mem[149] : 
                        (N82)? mem[199] : 
                        (N84)? mem[249] : 
                        (N86)? mem[299] : 
                        (N88)? mem[349] : 
                        (N90)? mem[399] : 
                        (N92)? mem[449] : 
                        (N94)? mem[499] : 
                        (N96)? mem[549] : 
                        (N98)? mem[599] : 
                        (N100)? mem[649] : 
                        (N102)? mem[699] : 
                        (N104)? mem[749] : 
                        (N106)? mem[799] : 
                        (N108)? mem[849] : 
                        (N110)? mem[899] : 
                        (N112)? mem[949] : 
                        (N114)? mem[999] : 
                        (N116)? mem[1049] : 
                        (N118)? mem[1099] : 
                        (N120)? mem[1149] : 
                        (N122)? mem[1199] : 
                        (N124)? mem[1249] : 
                        (N126)? mem[1299] : 
                        (N128)? mem[1349] : 
                        (N130)? mem[1399] : 
                        (N132)? mem[1449] : 
                        (N134)? mem[1499] : 
                        (N136)? mem[1549] : 
                        (N138)? mem[1599] : 
                        (N77)? mem[1649] : 
                        (N79)? mem[1699] : 
                        (N81)? mem[1749] : 
                        (N83)? mem[1799] : 
                        (N85)? mem[1849] : 
                        (N87)? mem[1899] : 
                        (N89)? mem[1949] : 
                        (N91)? mem[1999] : 
                        (N93)? mem[2049] : 
                        (N95)? mem[2099] : 
                        (N97)? mem[2149] : 
                        (N99)? mem[2199] : 
                        (N101)? mem[2249] : 
                        (N103)? mem[2299] : 
                        (N105)? mem[2349] : 
                        (N107)? mem[2399] : 
                        (N109)? mem[2449] : 
                        (N111)? mem[2499] : 
                        (N113)? mem[2549] : 
                        (N115)? mem[2599] : 
                        (N117)? mem[2649] : 
                        (N119)? mem[2699] : 
                        (N121)? mem[2749] : 
                        (N123)? mem[2799] : 
                        (N125)? mem[2849] : 
                        (N127)? mem[2899] : 
                        (N129)? mem[2949] : 
                        (N131)? mem[2999] : 
                        (N133)? mem[3049] : 
                        (N135)? mem[3099] : 
                        (N137)? mem[3149] : 
                        (N139)? mem[3199] : 1'b0;
  assign r_data_o[48] = (N76)? mem[48] : 
                        (N78)? mem[98] : 
                        (N80)? mem[148] : 
                        (N82)? mem[198] : 
                        (N84)? mem[248] : 
                        (N86)? mem[298] : 
                        (N88)? mem[348] : 
                        (N90)? mem[398] : 
                        (N92)? mem[448] : 
                        (N94)? mem[498] : 
                        (N96)? mem[548] : 
                        (N98)? mem[598] : 
                        (N100)? mem[648] : 
                        (N102)? mem[698] : 
                        (N104)? mem[748] : 
                        (N106)? mem[798] : 
                        (N108)? mem[848] : 
                        (N110)? mem[898] : 
                        (N112)? mem[948] : 
                        (N114)? mem[998] : 
                        (N116)? mem[1048] : 
                        (N118)? mem[1098] : 
                        (N120)? mem[1148] : 
                        (N122)? mem[1198] : 
                        (N124)? mem[1248] : 
                        (N126)? mem[1298] : 
                        (N128)? mem[1348] : 
                        (N130)? mem[1398] : 
                        (N132)? mem[1448] : 
                        (N134)? mem[1498] : 
                        (N136)? mem[1548] : 
                        (N138)? mem[1598] : 
                        (N77)? mem[1648] : 
                        (N79)? mem[1698] : 
                        (N81)? mem[1748] : 
                        (N83)? mem[1798] : 
                        (N85)? mem[1848] : 
                        (N87)? mem[1898] : 
                        (N89)? mem[1948] : 
                        (N91)? mem[1998] : 
                        (N93)? mem[2048] : 
                        (N95)? mem[2098] : 
                        (N97)? mem[2148] : 
                        (N99)? mem[2198] : 
                        (N101)? mem[2248] : 
                        (N103)? mem[2298] : 
                        (N105)? mem[2348] : 
                        (N107)? mem[2398] : 
                        (N109)? mem[2448] : 
                        (N111)? mem[2498] : 
                        (N113)? mem[2548] : 
                        (N115)? mem[2598] : 
                        (N117)? mem[2648] : 
                        (N119)? mem[2698] : 
                        (N121)? mem[2748] : 
                        (N123)? mem[2798] : 
                        (N125)? mem[2848] : 
                        (N127)? mem[2898] : 
                        (N129)? mem[2948] : 
                        (N131)? mem[2998] : 
                        (N133)? mem[3048] : 
                        (N135)? mem[3098] : 
                        (N137)? mem[3148] : 
                        (N139)? mem[3198] : 1'b0;
  assign r_data_o[47] = (N76)? mem[47] : 
                        (N78)? mem[97] : 
                        (N80)? mem[147] : 
                        (N82)? mem[197] : 
                        (N84)? mem[247] : 
                        (N86)? mem[297] : 
                        (N88)? mem[347] : 
                        (N90)? mem[397] : 
                        (N92)? mem[447] : 
                        (N94)? mem[497] : 
                        (N96)? mem[547] : 
                        (N98)? mem[597] : 
                        (N100)? mem[647] : 
                        (N102)? mem[697] : 
                        (N104)? mem[747] : 
                        (N106)? mem[797] : 
                        (N108)? mem[847] : 
                        (N110)? mem[897] : 
                        (N112)? mem[947] : 
                        (N114)? mem[997] : 
                        (N116)? mem[1047] : 
                        (N118)? mem[1097] : 
                        (N120)? mem[1147] : 
                        (N122)? mem[1197] : 
                        (N124)? mem[1247] : 
                        (N126)? mem[1297] : 
                        (N128)? mem[1347] : 
                        (N130)? mem[1397] : 
                        (N132)? mem[1447] : 
                        (N134)? mem[1497] : 
                        (N136)? mem[1547] : 
                        (N138)? mem[1597] : 
                        (N77)? mem[1647] : 
                        (N79)? mem[1697] : 
                        (N81)? mem[1747] : 
                        (N83)? mem[1797] : 
                        (N85)? mem[1847] : 
                        (N87)? mem[1897] : 
                        (N89)? mem[1947] : 
                        (N91)? mem[1997] : 
                        (N93)? mem[2047] : 
                        (N95)? mem[2097] : 
                        (N97)? mem[2147] : 
                        (N99)? mem[2197] : 
                        (N101)? mem[2247] : 
                        (N103)? mem[2297] : 
                        (N105)? mem[2347] : 
                        (N107)? mem[2397] : 
                        (N109)? mem[2447] : 
                        (N111)? mem[2497] : 
                        (N113)? mem[2547] : 
                        (N115)? mem[2597] : 
                        (N117)? mem[2647] : 
                        (N119)? mem[2697] : 
                        (N121)? mem[2747] : 
                        (N123)? mem[2797] : 
                        (N125)? mem[2847] : 
                        (N127)? mem[2897] : 
                        (N129)? mem[2947] : 
                        (N131)? mem[2997] : 
                        (N133)? mem[3047] : 
                        (N135)? mem[3097] : 
                        (N137)? mem[3147] : 
                        (N139)? mem[3197] : 1'b0;
  assign r_data_o[46] = (N76)? mem[46] : 
                        (N78)? mem[96] : 
                        (N80)? mem[146] : 
                        (N82)? mem[196] : 
                        (N84)? mem[246] : 
                        (N86)? mem[296] : 
                        (N88)? mem[346] : 
                        (N90)? mem[396] : 
                        (N92)? mem[446] : 
                        (N94)? mem[496] : 
                        (N96)? mem[546] : 
                        (N98)? mem[596] : 
                        (N100)? mem[646] : 
                        (N102)? mem[696] : 
                        (N104)? mem[746] : 
                        (N106)? mem[796] : 
                        (N108)? mem[846] : 
                        (N110)? mem[896] : 
                        (N112)? mem[946] : 
                        (N114)? mem[996] : 
                        (N116)? mem[1046] : 
                        (N118)? mem[1096] : 
                        (N120)? mem[1146] : 
                        (N122)? mem[1196] : 
                        (N124)? mem[1246] : 
                        (N126)? mem[1296] : 
                        (N128)? mem[1346] : 
                        (N130)? mem[1396] : 
                        (N132)? mem[1446] : 
                        (N134)? mem[1496] : 
                        (N136)? mem[1546] : 
                        (N138)? mem[1596] : 
                        (N77)? mem[1646] : 
                        (N79)? mem[1696] : 
                        (N81)? mem[1746] : 
                        (N83)? mem[1796] : 
                        (N85)? mem[1846] : 
                        (N87)? mem[1896] : 
                        (N89)? mem[1946] : 
                        (N91)? mem[1996] : 
                        (N93)? mem[2046] : 
                        (N95)? mem[2096] : 
                        (N97)? mem[2146] : 
                        (N99)? mem[2196] : 
                        (N101)? mem[2246] : 
                        (N103)? mem[2296] : 
                        (N105)? mem[2346] : 
                        (N107)? mem[2396] : 
                        (N109)? mem[2446] : 
                        (N111)? mem[2496] : 
                        (N113)? mem[2546] : 
                        (N115)? mem[2596] : 
                        (N117)? mem[2646] : 
                        (N119)? mem[2696] : 
                        (N121)? mem[2746] : 
                        (N123)? mem[2796] : 
                        (N125)? mem[2846] : 
                        (N127)? mem[2896] : 
                        (N129)? mem[2946] : 
                        (N131)? mem[2996] : 
                        (N133)? mem[3046] : 
                        (N135)? mem[3096] : 
                        (N137)? mem[3146] : 
                        (N139)? mem[3196] : 1'b0;
  assign r_data_o[45] = (N76)? mem[45] : 
                        (N78)? mem[95] : 
                        (N80)? mem[145] : 
                        (N82)? mem[195] : 
                        (N84)? mem[245] : 
                        (N86)? mem[295] : 
                        (N88)? mem[345] : 
                        (N90)? mem[395] : 
                        (N92)? mem[445] : 
                        (N94)? mem[495] : 
                        (N96)? mem[545] : 
                        (N98)? mem[595] : 
                        (N100)? mem[645] : 
                        (N102)? mem[695] : 
                        (N104)? mem[745] : 
                        (N106)? mem[795] : 
                        (N108)? mem[845] : 
                        (N110)? mem[895] : 
                        (N112)? mem[945] : 
                        (N114)? mem[995] : 
                        (N116)? mem[1045] : 
                        (N118)? mem[1095] : 
                        (N120)? mem[1145] : 
                        (N122)? mem[1195] : 
                        (N124)? mem[1245] : 
                        (N126)? mem[1295] : 
                        (N128)? mem[1345] : 
                        (N130)? mem[1395] : 
                        (N132)? mem[1445] : 
                        (N134)? mem[1495] : 
                        (N136)? mem[1545] : 
                        (N138)? mem[1595] : 
                        (N77)? mem[1645] : 
                        (N79)? mem[1695] : 
                        (N81)? mem[1745] : 
                        (N83)? mem[1795] : 
                        (N85)? mem[1845] : 
                        (N87)? mem[1895] : 
                        (N89)? mem[1945] : 
                        (N91)? mem[1995] : 
                        (N93)? mem[2045] : 
                        (N95)? mem[2095] : 
                        (N97)? mem[2145] : 
                        (N99)? mem[2195] : 
                        (N101)? mem[2245] : 
                        (N103)? mem[2295] : 
                        (N105)? mem[2345] : 
                        (N107)? mem[2395] : 
                        (N109)? mem[2445] : 
                        (N111)? mem[2495] : 
                        (N113)? mem[2545] : 
                        (N115)? mem[2595] : 
                        (N117)? mem[2645] : 
                        (N119)? mem[2695] : 
                        (N121)? mem[2745] : 
                        (N123)? mem[2795] : 
                        (N125)? mem[2845] : 
                        (N127)? mem[2895] : 
                        (N129)? mem[2945] : 
                        (N131)? mem[2995] : 
                        (N133)? mem[3045] : 
                        (N135)? mem[3095] : 
                        (N137)? mem[3145] : 
                        (N139)? mem[3195] : 1'b0;
  assign r_data_o[44] = (N76)? mem[44] : 
                        (N78)? mem[94] : 
                        (N80)? mem[144] : 
                        (N82)? mem[194] : 
                        (N84)? mem[244] : 
                        (N86)? mem[294] : 
                        (N88)? mem[344] : 
                        (N90)? mem[394] : 
                        (N92)? mem[444] : 
                        (N94)? mem[494] : 
                        (N96)? mem[544] : 
                        (N98)? mem[594] : 
                        (N100)? mem[644] : 
                        (N102)? mem[694] : 
                        (N104)? mem[744] : 
                        (N106)? mem[794] : 
                        (N108)? mem[844] : 
                        (N110)? mem[894] : 
                        (N112)? mem[944] : 
                        (N114)? mem[994] : 
                        (N116)? mem[1044] : 
                        (N118)? mem[1094] : 
                        (N120)? mem[1144] : 
                        (N122)? mem[1194] : 
                        (N124)? mem[1244] : 
                        (N126)? mem[1294] : 
                        (N128)? mem[1344] : 
                        (N130)? mem[1394] : 
                        (N132)? mem[1444] : 
                        (N134)? mem[1494] : 
                        (N136)? mem[1544] : 
                        (N138)? mem[1594] : 
                        (N77)? mem[1644] : 
                        (N79)? mem[1694] : 
                        (N81)? mem[1744] : 
                        (N83)? mem[1794] : 
                        (N85)? mem[1844] : 
                        (N87)? mem[1894] : 
                        (N89)? mem[1944] : 
                        (N91)? mem[1994] : 
                        (N93)? mem[2044] : 
                        (N95)? mem[2094] : 
                        (N97)? mem[2144] : 
                        (N99)? mem[2194] : 
                        (N101)? mem[2244] : 
                        (N103)? mem[2294] : 
                        (N105)? mem[2344] : 
                        (N107)? mem[2394] : 
                        (N109)? mem[2444] : 
                        (N111)? mem[2494] : 
                        (N113)? mem[2544] : 
                        (N115)? mem[2594] : 
                        (N117)? mem[2644] : 
                        (N119)? mem[2694] : 
                        (N121)? mem[2744] : 
                        (N123)? mem[2794] : 
                        (N125)? mem[2844] : 
                        (N127)? mem[2894] : 
                        (N129)? mem[2944] : 
                        (N131)? mem[2994] : 
                        (N133)? mem[3044] : 
                        (N135)? mem[3094] : 
                        (N137)? mem[3144] : 
                        (N139)? mem[3194] : 1'b0;
  assign r_data_o[43] = (N76)? mem[43] : 
                        (N78)? mem[93] : 
                        (N80)? mem[143] : 
                        (N82)? mem[193] : 
                        (N84)? mem[243] : 
                        (N86)? mem[293] : 
                        (N88)? mem[343] : 
                        (N90)? mem[393] : 
                        (N92)? mem[443] : 
                        (N94)? mem[493] : 
                        (N96)? mem[543] : 
                        (N98)? mem[593] : 
                        (N100)? mem[643] : 
                        (N102)? mem[693] : 
                        (N104)? mem[743] : 
                        (N106)? mem[793] : 
                        (N108)? mem[843] : 
                        (N110)? mem[893] : 
                        (N112)? mem[943] : 
                        (N114)? mem[993] : 
                        (N116)? mem[1043] : 
                        (N118)? mem[1093] : 
                        (N120)? mem[1143] : 
                        (N122)? mem[1193] : 
                        (N124)? mem[1243] : 
                        (N126)? mem[1293] : 
                        (N128)? mem[1343] : 
                        (N130)? mem[1393] : 
                        (N132)? mem[1443] : 
                        (N134)? mem[1493] : 
                        (N136)? mem[1543] : 
                        (N138)? mem[1593] : 
                        (N77)? mem[1643] : 
                        (N79)? mem[1693] : 
                        (N81)? mem[1743] : 
                        (N83)? mem[1793] : 
                        (N85)? mem[1843] : 
                        (N87)? mem[1893] : 
                        (N89)? mem[1943] : 
                        (N91)? mem[1993] : 
                        (N93)? mem[2043] : 
                        (N95)? mem[2093] : 
                        (N97)? mem[2143] : 
                        (N99)? mem[2193] : 
                        (N101)? mem[2243] : 
                        (N103)? mem[2293] : 
                        (N105)? mem[2343] : 
                        (N107)? mem[2393] : 
                        (N109)? mem[2443] : 
                        (N111)? mem[2493] : 
                        (N113)? mem[2543] : 
                        (N115)? mem[2593] : 
                        (N117)? mem[2643] : 
                        (N119)? mem[2693] : 
                        (N121)? mem[2743] : 
                        (N123)? mem[2793] : 
                        (N125)? mem[2843] : 
                        (N127)? mem[2893] : 
                        (N129)? mem[2943] : 
                        (N131)? mem[2993] : 
                        (N133)? mem[3043] : 
                        (N135)? mem[3093] : 
                        (N137)? mem[3143] : 
                        (N139)? mem[3193] : 1'b0;
  assign r_data_o[42] = (N76)? mem[42] : 
                        (N78)? mem[92] : 
                        (N80)? mem[142] : 
                        (N82)? mem[192] : 
                        (N84)? mem[242] : 
                        (N86)? mem[292] : 
                        (N88)? mem[342] : 
                        (N90)? mem[392] : 
                        (N92)? mem[442] : 
                        (N94)? mem[492] : 
                        (N96)? mem[542] : 
                        (N98)? mem[592] : 
                        (N100)? mem[642] : 
                        (N102)? mem[692] : 
                        (N104)? mem[742] : 
                        (N106)? mem[792] : 
                        (N108)? mem[842] : 
                        (N110)? mem[892] : 
                        (N112)? mem[942] : 
                        (N114)? mem[992] : 
                        (N116)? mem[1042] : 
                        (N118)? mem[1092] : 
                        (N120)? mem[1142] : 
                        (N122)? mem[1192] : 
                        (N124)? mem[1242] : 
                        (N126)? mem[1292] : 
                        (N128)? mem[1342] : 
                        (N130)? mem[1392] : 
                        (N132)? mem[1442] : 
                        (N134)? mem[1492] : 
                        (N136)? mem[1542] : 
                        (N138)? mem[1592] : 
                        (N77)? mem[1642] : 
                        (N79)? mem[1692] : 
                        (N81)? mem[1742] : 
                        (N83)? mem[1792] : 
                        (N85)? mem[1842] : 
                        (N87)? mem[1892] : 
                        (N89)? mem[1942] : 
                        (N91)? mem[1992] : 
                        (N93)? mem[2042] : 
                        (N95)? mem[2092] : 
                        (N97)? mem[2142] : 
                        (N99)? mem[2192] : 
                        (N101)? mem[2242] : 
                        (N103)? mem[2292] : 
                        (N105)? mem[2342] : 
                        (N107)? mem[2392] : 
                        (N109)? mem[2442] : 
                        (N111)? mem[2492] : 
                        (N113)? mem[2542] : 
                        (N115)? mem[2592] : 
                        (N117)? mem[2642] : 
                        (N119)? mem[2692] : 
                        (N121)? mem[2742] : 
                        (N123)? mem[2792] : 
                        (N125)? mem[2842] : 
                        (N127)? mem[2892] : 
                        (N129)? mem[2942] : 
                        (N131)? mem[2992] : 
                        (N133)? mem[3042] : 
                        (N135)? mem[3092] : 
                        (N137)? mem[3142] : 
                        (N139)? mem[3192] : 1'b0;
  assign r_data_o[41] = (N76)? mem[41] : 
                        (N78)? mem[91] : 
                        (N80)? mem[141] : 
                        (N82)? mem[191] : 
                        (N84)? mem[241] : 
                        (N86)? mem[291] : 
                        (N88)? mem[341] : 
                        (N90)? mem[391] : 
                        (N92)? mem[441] : 
                        (N94)? mem[491] : 
                        (N96)? mem[541] : 
                        (N98)? mem[591] : 
                        (N100)? mem[641] : 
                        (N102)? mem[691] : 
                        (N104)? mem[741] : 
                        (N106)? mem[791] : 
                        (N108)? mem[841] : 
                        (N110)? mem[891] : 
                        (N112)? mem[941] : 
                        (N114)? mem[991] : 
                        (N116)? mem[1041] : 
                        (N118)? mem[1091] : 
                        (N120)? mem[1141] : 
                        (N122)? mem[1191] : 
                        (N124)? mem[1241] : 
                        (N126)? mem[1291] : 
                        (N128)? mem[1341] : 
                        (N130)? mem[1391] : 
                        (N132)? mem[1441] : 
                        (N134)? mem[1491] : 
                        (N136)? mem[1541] : 
                        (N138)? mem[1591] : 
                        (N77)? mem[1641] : 
                        (N79)? mem[1691] : 
                        (N81)? mem[1741] : 
                        (N83)? mem[1791] : 
                        (N85)? mem[1841] : 
                        (N87)? mem[1891] : 
                        (N89)? mem[1941] : 
                        (N91)? mem[1991] : 
                        (N93)? mem[2041] : 
                        (N95)? mem[2091] : 
                        (N97)? mem[2141] : 
                        (N99)? mem[2191] : 
                        (N101)? mem[2241] : 
                        (N103)? mem[2291] : 
                        (N105)? mem[2341] : 
                        (N107)? mem[2391] : 
                        (N109)? mem[2441] : 
                        (N111)? mem[2491] : 
                        (N113)? mem[2541] : 
                        (N115)? mem[2591] : 
                        (N117)? mem[2641] : 
                        (N119)? mem[2691] : 
                        (N121)? mem[2741] : 
                        (N123)? mem[2791] : 
                        (N125)? mem[2841] : 
                        (N127)? mem[2891] : 
                        (N129)? mem[2941] : 
                        (N131)? mem[2991] : 
                        (N133)? mem[3041] : 
                        (N135)? mem[3091] : 
                        (N137)? mem[3141] : 
                        (N139)? mem[3191] : 1'b0;
  assign r_data_o[40] = (N76)? mem[40] : 
                        (N78)? mem[90] : 
                        (N80)? mem[140] : 
                        (N82)? mem[190] : 
                        (N84)? mem[240] : 
                        (N86)? mem[290] : 
                        (N88)? mem[340] : 
                        (N90)? mem[390] : 
                        (N92)? mem[440] : 
                        (N94)? mem[490] : 
                        (N96)? mem[540] : 
                        (N98)? mem[590] : 
                        (N100)? mem[640] : 
                        (N102)? mem[690] : 
                        (N104)? mem[740] : 
                        (N106)? mem[790] : 
                        (N108)? mem[840] : 
                        (N110)? mem[890] : 
                        (N112)? mem[940] : 
                        (N114)? mem[990] : 
                        (N116)? mem[1040] : 
                        (N118)? mem[1090] : 
                        (N120)? mem[1140] : 
                        (N122)? mem[1190] : 
                        (N124)? mem[1240] : 
                        (N126)? mem[1290] : 
                        (N128)? mem[1340] : 
                        (N130)? mem[1390] : 
                        (N132)? mem[1440] : 
                        (N134)? mem[1490] : 
                        (N136)? mem[1540] : 
                        (N138)? mem[1590] : 
                        (N77)? mem[1640] : 
                        (N79)? mem[1690] : 
                        (N81)? mem[1740] : 
                        (N83)? mem[1790] : 
                        (N85)? mem[1840] : 
                        (N87)? mem[1890] : 
                        (N89)? mem[1940] : 
                        (N91)? mem[1990] : 
                        (N93)? mem[2040] : 
                        (N95)? mem[2090] : 
                        (N97)? mem[2140] : 
                        (N99)? mem[2190] : 
                        (N101)? mem[2240] : 
                        (N103)? mem[2290] : 
                        (N105)? mem[2340] : 
                        (N107)? mem[2390] : 
                        (N109)? mem[2440] : 
                        (N111)? mem[2490] : 
                        (N113)? mem[2540] : 
                        (N115)? mem[2590] : 
                        (N117)? mem[2640] : 
                        (N119)? mem[2690] : 
                        (N121)? mem[2740] : 
                        (N123)? mem[2790] : 
                        (N125)? mem[2840] : 
                        (N127)? mem[2890] : 
                        (N129)? mem[2940] : 
                        (N131)? mem[2990] : 
                        (N133)? mem[3040] : 
                        (N135)? mem[3090] : 
                        (N137)? mem[3140] : 
                        (N139)? mem[3190] : 1'b0;
  assign r_data_o[39] = (N76)? mem[39] : 
                        (N78)? mem[89] : 
                        (N80)? mem[139] : 
                        (N82)? mem[189] : 
                        (N84)? mem[239] : 
                        (N86)? mem[289] : 
                        (N88)? mem[339] : 
                        (N90)? mem[389] : 
                        (N92)? mem[439] : 
                        (N94)? mem[489] : 
                        (N96)? mem[539] : 
                        (N98)? mem[589] : 
                        (N100)? mem[639] : 
                        (N102)? mem[689] : 
                        (N104)? mem[739] : 
                        (N106)? mem[789] : 
                        (N108)? mem[839] : 
                        (N110)? mem[889] : 
                        (N112)? mem[939] : 
                        (N114)? mem[989] : 
                        (N116)? mem[1039] : 
                        (N118)? mem[1089] : 
                        (N120)? mem[1139] : 
                        (N122)? mem[1189] : 
                        (N124)? mem[1239] : 
                        (N126)? mem[1289] : 
                        (N128)? mem[1339] : 
                        (N130)? mem[1389] : 
                        (N132)? mem[1439] : 
                        (N134)? mem[1489] : 
                        (N136)? mem[1539] : 
                        (N138)? mem[1589] : 
                        (N77)? mem[1639] : 
                        (N79)? mem[1689] : 
                        (N81)? mem[1739] : 
                        (N83)? mem[1789] : 
                        (N85)? mem[1839] : 
                        (N87)? mem[1889] : 
                        (N89)? mem[1939] : 
                        (N91)? mem[1989] : 
                        (N93)? mem[2039] : 
                        (N95)? mem[2089] : 
                        (N97)? mem[2139] : 
                        (N99)? mem[2189] : 
                        (N101)? mem[2239] : 
                        (N103)? mem[2289] : 
                        (N105)? mem[2339] : 
                        (N107)? mem[2389] : 
                        (N109)? mem[2439] : 
                        (N111)? mem[2489] : 
                        (N113)? mem[2539] : 
                        (N115)? mem[2589] : 
                        (N117)? mem[2639] : 
                        (N119)? mem[2689] : 
                        (N121)? mem[2739] : 
                        (N123)? mem[2789] : 
                        (N125)? mem[2839] : 
                        (N127)? mem[2889] : 
                        (N129)? mem[2939] : 
                        (N131)? mem[2989] : 
                        (N133)? mem[3039] : 
                        (N135)? mem[3089] : 
                        (N137)? mem[3139] : 
                        (N139)? mem[3189] : 1'b0;
  assign r_data_o[38] = (N76)? mem[38] : 
                        (N78)? mem[88] : 
                        (N80)? mem[138] : 
                        (N82)? mem[188] : 
                        (N84)? mem[238] : 
                        (N86)? mem[288] : 
                        (N88)? mem[338] : 
                        (N90)? mem[388] : 
                        (N92)? mem[438] : 
                        (N94)? mem[488] : 
                        (N96)? mem[538] : 
                        (N98)? mem[588] : 
                        (N100)? mem[638] : 
                        (N102)? mem[688] : 
                        (N104)? mem[738] : 
                        (N106)? mem[788] : 
                        (N108)? mem[838] : 
                        (N110)? mem[888] : 
                        (N112)? mem[938] : 
                        (N114)? mem[988] : 
                        (N116)? mem[1038] : 
                        (N118)? mem[1088] : 
                        (N120)? mem[1138] : 
                        (N122)? mem[1188] : 
                        (N124)? mem[1238] : 
                        (N126)? mem[1288] : 
                        (N128)? mem[1338] : 
                        (N130)? mem[1388] : 
                        (N132)? mem[1438] : 
                        (N134)? mem[1488] : 
                        (N136)? mem[1538] : 
                        (N138)? mem[1588] : 
                        (N77)? mem[1638] : 
                        (N79)? mem[1688] : 
                        (N81)? mem[1738] : 
                        (N83)? mem[1788] : 
                        (N85)? mem[1838] : 
                        (N87)? mem[1888] : 
                        (N89)? mem[1938] : 
                        (N91)? mem[1988] : 
                        (N93)? mem[2038] : 
                        (N95)? mem[2088] : 
                        (N97)? mem[2138] : 
                        (N99)? mem[2188] : 
                        (N101)? mem[2238] : 
                        (N103)? mem[2288] : 
                        (N105)? mem[2338] : 
                        (N107)? mem[2388] : 
                        (N109)? mem[2438] : 
                        (N111)? mem[2488] : 
                        (N113)? mem[2538] : 
                        (N115)? mem[2588] : 
                        (N117)? mem[2638] : 
                        (N119)? mem[2688] : 
                        (N121)? mem[2738] : 
                        (N123)? mem[2788] : 
                        (N125)? mem[2838] : 
                        (N127)? mem[2888] : 
                        (N129)? mem[2938] : 
                        (N131)? mem[2988] : 
                        (N133)? mem[3038] : 
                        (N135)? mem[3088] : 
                        (N137)? mem[3138] : 
                        (N139)? mem[3188] : 1'b0;
  assign r_data_o[37] = (N76)? mem[37] : 
                        (N78)? mem[87] : 
                        (N80)? mem[137] : 
                        (N82)? mem[187] : 
                        (N84)? mem[237] : 
                        (N86)? mem[287] : 
                        (N88)? mem[337] : 
                        (N90)? mem[387] : 
                        (N92)? mem[437] : 
                        (N94)? mem[487] : 
                        (N96)? mem[537] : 
                        (N98)? mem[587] : 
                        (N100)? mem[637] : 
                        (N102)? mem[687] : 
                        (N104)? mem[737] : 
                        (N106)? mem[787] : 
                        (N108)? mem[837] : 
                        (N110)? mem[887] : 
                        (N112)? mem[937] : 
                        (N114)? mem[987] : 
                        (N116)? mem[1037] : 
                        (N118)? mem[1087] : 
                        (N120)? mem[1137] : 
                        (N122)? mem[1187] : 
                        (N124)? mem[1237] : 
                        (N126)? mem[1287] : 
                        (N128)? mem[1337] : 
                        (N130)? mem[1387] : 
                        (N132)? mem[1437] : 
                        (N134)? mem[1487] : 
                        (N136)? mem[1537] : 
                        (N138)? mem[1587] : 
                        (N77)? mem[1637] : 
                        (N79)? mem[1687] : 
                        (N81)? mem[1737] : 
                        (N83)? mem[1787] : 
                        (N85)? mem[1837] : 
                        (N87)? mem[1887] : 
                        (N89)? mem[1937] : 
                        (N91)? mem[1987] : 
                        (N93)? mem[2037] : 
                        (N95)? mem[2087] : 
                        (N97)? mem[2137] : 
                        (N99)? mem[2187] : 
                        (N101)? mem[2237] : 
                        (N103)? mem[2287] : 
                        (N105)? mem[2337] : 
                        (N107)? mem[2387] : 
                        (N109)? mem[2437] : 
                        (N111)? mem[2487] : 
                        (N113)? mem[2537] : 
                        (N115)? mem[2587] : 
                        (N117)? mem[2637] : 
                        (N119)? mem[2687] : 
                        (N121)? mem[2737] : 
                        (N123)? mem[2787] : 
                        (N125)? mem[2837] : 
                        (N127)? mem[2887] : 
                        (N129)? mem[2937] : 
                        (N131)? mem[2987] : 
                        (N133)? mem[3037] : 
                        (N135)? mem[3087] : 
                        (N137)? mem[3137] : 
                        (N139)? mem[3187] : 1'b0;
  assign r_data_o[36] = (N76)? mem[36] : 
                        (N78)? mem[86] : 
                        (N80)? mem[136] : 
                        (N82)? mem[186] : 
                        (N84)? mem[236] : 
                        (N86)? mem[286] : 
                        (N88)? mem[336] : 
                        (N90)? mem[386] : 
                        (N92)? mem[436] : 
                        (N94)? mem[486] : 
                        (N96)? mem[536] : 
                        (N98)? mem[586] : 
                        (N100)? mem[636] : 
                        (N102)? mem[686] : 
                        (N104)? mem[736] : 
                        (N106)? mem[786] : 
                        (N108)? mem[836] : 
                        (N110)? mem[886] : 
                        (N112)? mem[936] : 
                        (N114)? mem[986] : 
                        (N116)? mem[1036] : 
                        (N118)? mem[1086] : 
                        (N120)? mem[1136] : 
                        (N122)? mem[1186] : 
                        (N124)? mem[1236] : 
                        (N126)? mem[1286] : 
                        (N128)? mem[1336] : 
                        (N130)? mem[1386] : 
                        (N132)? mem[1436] : 
                        (N134)? mem[1486] : 
                        (N136)? mem[1536] : 
                        (N138)? mem[1586] : 
                        (N77)? mem[1636] : 
                        (N79)? mem[1686] : 
                        (N81)? mem[1736] : 
                        (N83)? mem[1786] : 
                        (N85)? mem[1836] : 
                        (N87)? mem[1886] : 
                        (N89)? mem[1936] : 
                        (N91)? mem[1986] : 
                        (N93)? mem[2036] : 
                        (N95)? mem[2086] : 
                        (N97)? mem[2136] : 
                        (N99)? mem[2186] : 
                        (N101)? mem[2236] : 
                        (N103)? mem[2286] : 
                        (N105)? mem[2336] : 
                        (N107)? mem[2386] : 
                        (N109)? mem[2436] : 
                        (N111)? mem[2486] : 
                        (N113)? mem[2536] : 
                        (N115)? mem[2586] : 
                        (N117)? mem[2636] : 
                        (N119)? mem[2686] : 
                        (N121)? mem[2736] : 
                        (N123)? mem[2786] : 
                        (N125)? mem[2836] : 
                        (N127)? mem[2886] : 
                        (N129)? mem[2936] : 
                        (N131)? mem[2986] : 
                        (N133)? mem[3036] : 
                        (N135)? mem[3086] : 
                        (N137)? mem[3136] : 
                        (N139)? mem[3186] : 1'b0;
  assign r_data_o[35] = (N76)? mem[35] : 
                        (N78)? mem[85] : 
                        (N80)? mem[135] : 
                        (N82)? mem[185] : 
                        (N84)? mem[235] : 
                        (N86)? mem[285] : 
                        (N88)? mem[335] : 
                        (N90)? mem[385] : 
                        (N92)? mem[435] : 
                        (N94)? mem[485] : 
                        (N96)? mem[535] : 
                        (N98)? mem[585] : 
                        (N100)? mem[635] : 
                        (N102)? mem[685] : 
                        (N104)? mem[735] : 
                        (N106)? mem[785] : 
                        (N108)? mem[835] : 
                        (N110)? mem[885] : 
                        (N112)? mem[935] : 
                        (N114)? mem[985] : 
                        (N116)? mem[1035] : 
                        (N118)? mem[1085] : 
                        (N120)? mem[1135] : 
                        (N122)? mem[1185] : 
                        (N124)? mem[1235] : 
                        (N126)? mem[1285] : 
                        (N128)? mem[1335] : 
                        (N130)? mem[1385] : 
                        (N132)? mem[1435] : 
                        (N134)? mem[1485] : 
                        (N136)? mem[1535] : 
                        (N138)? mem[1585] : 
                        (N77)? mem[1635] : 
                        (N79)? mem[1685] : 
                        (N81)? mem[1735] : 
                        (N83)? mem[1785] : 
                        (N85)? mem[1835] : 
                        (N87)? mem[1885] : 
                        (N89)? mem[1935] : 
                        (N91)? mem[1985] : 
                        (N93)? mem[2035] : 
                        (N95)? mem[2085] : 
                        (N97)? mem[2135] : 
                        (N99)? mem[2185] : 
                        (N101)? mem[2235] : 
                        (N103)? mem[2285] : 
                        (N105)? mem[2335] : 
                        (N107)? mem[2385] : 
                        (N109)? mem[2435] : 
                        (N111)? mem[2485] : 
                        (N113)? mem[2535] : 
                        (N115)? mem[2585] : 
                        (N117)? mem[2635] : 
                        (N119)? mem[2685] : 
                        (N121)? mem[2735] : 
                        (N123)? mem[2785] : 
                        (N125)? mem[2835] : 
                        (N127)? mem[2885] : 
                        (N129)? mem[2935] : 
                        (N131)? mem[2985] : 
                        (N133)? mem[3035] : 
                        (N135)? mem[3085] : 
                        (N137)? mem[3135] : 
                        (N139)? mem[3185] : 1'b0;
  assign r_data_o[34] = (N76)? mem[34] : 
                        (N78)? mem[84] : 
                        (N80)? mem[134] : 
                        (N82)? mem[184] : 
                        (N84)? mem[234] : 
                        (N86)? mem[284] : 
                        (N88)? mem[334] : 
                        (N90)? mem[384] : 
                        (N92)? mem[434] : 
                        (N94)? mem[484] : 
                        (N96)? mem[534] : 
                        (N98)? mem[584] : 
                        (N100)? mem[634] : 
                        (N102)? mem[684] : 
                        (N104)? mem[734] : 
                        (N106)? mem[784] : 
                        (N108)? mem[834] : 
                        (N110)? mem[884] : 
                        (N112)? mem[934] : 
                        (N114)? mem[984] : 
                        (N116)? mem[1034] : 
                        (N118)? mem[1084] : 
                        (N120)? mem[1134] : 
                        (N122)? mem[1184] : 
                        (N124)? mem[1234] : 
                        (N126)? mem[1284] : 
                        (N128)? mem[1334] : 
                        (N130)? mem[1384] : 
                        (N132)? mem[1434] : 
                        (N134)? mem[1484] : 
                        (N136)? mem[1534] : 
                        (N138)? mem[1584] : 
                        (N77)? mem[1634] : 
                        (N79)? mem[1684] : 
                        (N81)? mem[1734] : 
                        (N83)? mem[1784] : 
                        (N85)? mem[1834] : 
                        (N87)? mem[1884] : 
                        (N89)? mem[1934] : 
                        (N91)? mem[1984] : 
                        (N93)? mem[2034] : 
                        (N95)? mem[2084] : 
                        (N97)? mem[2134] : 
                        (N99)? mem[2184] : 
                        (N101)? mem[2234] : 
                        (N103)? mem[2284] : 
                        (N105)? mem[2334] : 
                        (N107)? mem[2384] : 
                        (N109)? mem[2434] : 
                        (N111)? mem[2484] : 
                        (N113)? mem[2534] : 
                        (N115)? mem[2584] : 
                        (N117)? mem[2634] : 
                        (N119)? mem[2684] : 
                        (N121)? mem[2734] : 
                        (N123)? mem[2784] : 
                        (N125)? mem[2834] : 
                        (N127)? mem[2884] : 
                        (N129)? mem[2934] : 
                        (N131)? mem[2984] : 
                        (N133)? mem[3034] : 
                        (N135)? mem[3084] : 
                        (N137)? mem[3134] : 
                        (N139)? mem[3184] : 1'b0;
  assign r_data_o[33] = (N76)? mem[33] : 
                        (N78)? mem[83] : 
                        (N80)? mem[133] : 
                        (N82)? mem[183] : 
                        (N84)? mem[233] : 
                        (N86)? mem[283] : 
                        (N88)? mem[333] : 
                        (N90)? mem[383] : 
                        (N92)? mem[433] : 
                        (N94)? mem[483] : 
                        (N96)? mem[533] : 
                        (N98)? mem[583] : 
                        (N100)? mem[633] : 
                        (N102)? mem[683] : 
                        (N104)? mem[733] : 
                        (N106)? mem[783] : 
                        (N108)? mem[833] : 
                        (N110)? mem[883] : 
                        (N112)? mem[933] : 
                        (N114)? mem[983] : 
                        (N116)? mem[1033] : 
                        (N118)? mem[1083] : 
                        (N120)? mem[1133] : 
                        (N122)? mem[1183] : 
                        (N124)? mem[1233] : 
                        (N126)? mem[1283] : 
                        (N128)? mem[1333] : 
                        (N130)? mem[1383] : 
                        (N132)? mem[1433] : 
                        (N134)? mem[1483] : 
                        (N136)? mem[1533] : 
                        (N138)? mem[1583] : 
                        (N77)? mem[1633] : 
                        (N79)? mem[1683] : 
                        (N81)? mem[1733] : 
                        (N83)? mem[1783] : 
                        (N85)? mem[1833] : 
                        (N87)? mem[1883] : 
                        (N89)? mem[1933] : 
                        (N91)? mem[1983] : 
                        (N93)? mem[2033] : 
                        (N95)? mem[2083] : 
                        (N97)? mem[2133] : 
                        (N99)? mem[2183] : 
                        (N101)? mem[2233] : 
                        (N103)? mem[2283] : 
                        (N105)? mem[2333] : 
                        (N107)? mem[2383] : 
                        (N109)? mem[2433] : 
                        (N111)? mem[2483] : 
                        (N113)? mem[2533] : 
                        (N115)? mem[2583] : 
                        (N117)? mem[2633] : 
                        (N119)? mem[2683] : 
                        (N121)? mem[2733] : 
                        (N123)? mem[2783] : 
                        (N125)? mem[2833] : 
                        (N127)? mem[2883] : 
                        (N129)? mem[2933] : 
                        (N131)? mem[2983] : 
                        (N133)? mem[3033] : 
                        (N135)? mem[3083] : 
                        (N137)? mem[3133] : 
                        (N139)? mem[3183] : 1'b0;
  assign r_data_o[32] = (N76)? mem[32] : 
                        (N78)? mem[82] : 
                        (N80)? mem[132] : 
                        (N82)? mem[182] : 
                        (N84)? mem[232] : 
                        (N86)? mem[282] : 
                        (N88)? mem[332] : 
                        (N90)? mem[382] : 
                        (N92)? mem[432] : 
                        (N94)? mem[482] : 
                        (N96)? mem[532] : 
                        (N98)? mem[582] : 
                        (N100)? mem[632] : 
                        (N102)? mem[682] : 
                        (N104)? mem[732] : 
                        (N106)? mem[782] : 
                        (N108)? mem[832] : 
                        (N110)? mem[882] : 
                        (N112)? mem[932] : 
                        (N114)? mem[982] : 
                        (N116)? mem[1032] : 
                        (N118)? mem[1082] : 
                        (N120)? mem[1132] : 
                        (N122)? mem[1182] : 
                        (N124)? mem[1232] : 
                        (N126)? mem[1282] : 
                        (N128)? mem[1332] : 
                        (N130)? mem[1382] : 
                        (N132)? mem[1432] : 
                        (N134)? mem[1482] : 
                        (N136)? mem[1532] : 
                        (N138)? mem[1582] : 
                        (N77)? mem[1632] : 
                        (N79)? mem[1682] : 
                        (N81)? mem[1732] : 
                        (N83)? mem[1782] : 
                        (N85)? mem[1832] : 
                        (N87)? mem[1882] : 
                        (N89)? mem[1932] : 
                        (N91)? mem[1982] : 
                        (N93)? mem[2032] : 
                        (N95)? mem[2082] : 
                        (N97)? mem[2132] : 
                        (N99)? mem[2182] : 
                        (N101)? mem[2232] : 
                        (N103)? mem[2282] : 
                        (N105)? mem[2332] : 
                        (N107)? mem[2382] : 
                        (N109)? mem[2432] : 
                        (N111)? mem[2482] : 
                        (N113)? mem[2532] : 
                        (N115)? mem[2582] : 
                        (N117)? mem[2632] : 
                        (N119)? mem[2682] : 
                        (N121)? mem[2732] : 
                        (N123)? mem[2782] : 
                        (N125)? mem[2832] : 
                        (N127)? mem[2882] : 
                        (N129)? mem[2932] : 
                        (N131)? mem[2982] : 
                        (N133)? mem[3032] : 
                        (N135)? mem[3082] : 
                        (N137)? mem[3132] : 
                        (N139)? mem[3182] : 1'b0;
  assign r_data_o[31] = (N76)? mem[31] : 
                        (N78)? mem[81] : 
                        (N80)? mem[131] : 
                        (N82)? mem[181] : 
                        (N84)? mem[231] : 
                        (N86)? mem[281] : 
                        (N88)? mem[331] : 
                        (N90)? mem[381] : 
                        (N92)? mem[431] : 
                        (N94)? mem[481] : 
                        (N96)? mem[531] : 
                        (N98)? mem[581] : 
                        (N100)? mem[631] : 
                        (N102)? mem[681] : 
                        (N104)? mem[731] : 
                        (N106)? mem[781] : 
                        (N108)? mem[831] : 
                        (N110)? mem[881] : 
                        (N112)? mem[931] : 
                        (N114)? mem[981] : 
                        (N116)? mem[1031] : 
                        (N118)? mem[1081] : 
                        (N120)? mem[1131] : 
                        (N122)? mem[1181] : 
                        (N124)? mem[1231] : 
                        (N126)? mem[1281] : 
                        (N128)? mem[1331] : 
                        (N130)? mem[1381] : 
                        (N132)? mem[1431] : 
                        (N134)? mem[1481] : 
                        (N136)? mem[1531] : 
                        (N138)? mem[1581] : 
                        (N77)? mem[1631] : 
                        (N79)? mem[1681] : 
                        (N81)? mem[1731] : 
                        (N83)? mem[1781] : 
                        (N85)? mem[1831] : 
                        (N87)? mem[1881] : 
                        (N89)? mem[1931] : 
                        (N91)? mem[1981] : 
                        (N93)? mem[2031] : 
                        (N95)? mem[2081] : 
                        (N97)? mem[2131] : 
                        (N99)? mem[2181] : 
                        (N101)? mem[2231] : 
                        (N103)? mem[2281] : 
                        (N105)? mem[2331] : 
                        (N107)? mem[2381] : 
                        (N109)? mem[2431] : 
                        (N111)? mem[2481] : 
                        (N113)? mem[2531] : 
                        (N115)? mem[2581] : 
                        (N117)? mem[2631] : 
                        (N119)? mem[2681] : 
                        (N121)? mem[2731] : 
                        (N123)? mem[2781] : 
                        (N125)? mem[2831] : 
                        (N127)? mem[2881] : 
                        (N129)? mem[2931] : 
                        (N131)? mem[2981] : 
                        (N133)? mem[3031] : 
                        (N135)? mem[3081] : 
                        (N137)? mem[3131] : 
                        (N139)? mem[3181] : 1'b0;
  assign r_data_o[30] = (N76)? mem[30] : 
                        (N78)? mem[80] : 
                        (N80)? mem[130] : 
                        (N82)? mem[180] : 
                        (N84)? mem[230] : 
                        (N86)? mem[280] : 
                        (N88)? mem[330] : 
                        (N90)? mem[380] : 
                        (N92)? mem[430] : 
                        (N94)? mem[480] : 
                        (N96)? mem[530] : 
                        (N98)? mem[580] : 
                        (N100)? mem[630] : 
                        (N102)? mem[680] : 
                        (N104)? mem[730] : 
                        (N106)? mem[780] : 
                        (N108)? mem[830] : 
                        (N110)? mem[880] : 
                        (N112)? mem[930] : 
                        (N114)? mem[980] : 
                        (N116)? mem[1030] : 
                        (N118)? mem[1080] : 
                        (N120)? mem[1130] : 
                        (N122)? mem[1180] : 
                        (N124)? mem[1230] : 
                        (N126)? mem[1280] : 
                        (N128)? mem[1330] : 
                        (N130)? mem[1380] : 
                        (N132)? mem[1430] : 
                        (N134)? mem[1480] : 
                        (N136)? mem[1530] : 
                        (N138)? mem[1580] : 
                        (N77)? mem[1630] : 
                        (N79)? mem[1680] : 
                        (N81)? mem[1730] : 
                        (N83)? mem[1780] : 
                        (N85)? mem[1830] : 
                        (N87)? mem[1880] : 
                        (N89)? mem[1930] : 
                        (N91)? mem[1980] : 
                        (N93)? mem[2030] : 
                        (N95)? mem[2080] : 
                        (N97)? mem[2130] : 
                        (N99)? mem[2180] : 
                        (N101)? mem[2230] : 
                        (N103)? mem[2280] : 
                        (N105)? mem[2330] : 
                        (N107)? mem[2380] : 
                        (N109)? mem[2430] : 
                        (N111)? mem[2480] : 
                        (N113)? mem[2530] : 
                        (N115)? mem[2580] : 
                        (N117)? mem[2630] : 
                        (N119)? mem[2680] : 
                        (N121)? mem[2730] : 
                        (N123)? mem[2780] : 
                        (N125)? mem[2830] : 
                        (N127)? mem[2880] : 
                        (N129)? mem[2930] : 
                        (N131)? mem[2980] : 
                        (N133)? mem[3030] : 
                        (N135)? mem[3080] : 
                        (N137)? mem[3130] : 
                        (N139)? mem[3180] : 1'b0;
  assign r_data_o[29] = (N76)? mem[29] : 
                        (N78)? mem[79] : 
                        (N80)? mem[129] : 
                        (N82)? mem[179] : 
                        (N84)? mem[229] : 
                        (N86)? mem[279] : 
                        (N88)? mem[329] : 
                        (N90)? mem[379] : 
                        (N92)? mem[429] : 
                        (N94)? mem[479] : 
                        (N96)? mem[529] : 
                        (N98)? mem[579] : 
                        (N100)? mem[629] : 
                        (N102)? mem[679] : 
                        (N104)? mem[729] : 
                        (N106)? mem[779] : 
                        (N108)? mem[829] : 
                        (N110)? mem[879] : 
                        (N112)? mem[929] : 
                        (N114)? mem[979] : 
                        (N116)? mem[1029] : 
                        (N118)? mem[1079] : 
                        (N120)? mem[1129] : 
                        (N122)? mem[1179] : 
                        (N124)? mem[1229] : 
                        (N126)? mem[1279] : 
                        (N128)? mem[1329] : 
                        (N130)? mem[1379] : 
                        (N132)? mem[1429] : 
                        (N134)? mem[1479] : 
                        (N136)? mem[1529] : 
                        (N138)? mem[1579] : 
                        (N77)? mem[1629] : 
                        (N79)? mem[1679] : 
                        (N81)? mem[1729] : 
                        (N83)? mem[1779] : 
                        (N85)? mem[1829] : 
                        (N87)? mem[1879] : 
                        (N89)? mem[1929] : 
                        (N91)? mem[1979] : 
                        (N93)? mem[2029] : 
                        (N95)? mem[2079] : 
                        (N97)? mem[2129] : 
                        (N99)? mem[2179] : 
                        (N101)? mem[2229] : 
                        (N103)? mem[2279] : 
                        (N105)? mem[2329] : 
                        (N107)? mem[2379] : 
                        (N109)? mem[2429] : 
                        (N111)? mem[2479] : 
                        (N113)? mem[2529] : 
                        (N115)? mem[2579] : 
                        (N117)? mem[2629] : 
                        (N119)? mem[2679] : 
                        (N121)? mem[2729] : 
                        (N123)? mem[2779] : 
                        (N125)? mem[2829] : 
                        (N127)? mem[2879] : 
                        (N129)? mem[2929] : 
                        (N131)? mem[2979] : 
                        (N133)? mem[3029] : 
                        (N135)? mem[3079] : 
                        (N137)? mem[3129] : 
                        (N139)? mem[3179] : 1'b0;
  assign r_data_o[28] = (N76)? mem[28] : 
                        (N78)? mem[78] : 
                        (N80)? mem[128] : 
                        (N82)? mem[178] : 
                        (N84)? mem[228] : 
                        (N86)? mem[278] : 
                        (N88)? mem[328] : 
                        (N90)? mem[378] : 
                        (N92)? mem[428] : 
                        (N94)? mem[478] : 
                        (N96)? mem[528] : 
                        (N98)? mem[578] : 
                        (N100)? mem[628] : 
                        (N102)? mem[678] : 
                        (N104)? mem[728] : 
                        (N106)? mem[778] : 
                        (N108)? mem[828] : 
                        (N110)? mem[878] : 
                        (N112)? mem[928] : 
                        (N114)? mem[978] : 
                        (N116)? mem[1028] : 
                        (N118)? mem[1078] : 
                        (N120)? mem[1128] : 
                        (N122)? mem[1178] : 
                        (N124)? mem[1228] : 
                        (N126)? mem[1278] : 
                        (N128)? mem[1328] : 
                        (N130)? mem[1378] : 
                        (N132)? mem[1428] : 
                        (N134)? mem[1478] : 
                        (N136)? mem[1528] : 
                        (N138)? mem[1578] : 
                        (N77)? mem[1628] : 
                        (N79)? mem[1678] : 
                        (N81)? mem[1728] : 
                        (N83)? mem[1778] : 
                        (N85)? mem[1828] : 
                        (N87)? mem[1878] : 
                        (N89)? mem[1928] : 
                        (N91)? mem[1978] : 
                        (N93)? mem[2028] : 
                        (N95)? mem[2078] : 
                        (N97)? mem[2128] : 
                        (N99)? mem[2178] : 
                        (N101)? mem[2228] : 
                        (N103)? mem[2278] : 
                        (N105)? mem[2328] : 
                        (N107)? mem[2378] : 
                        (N109)? mem[2428] : 
                        (N111)? mem[2478] : 
                        (N113)? mem[2528] : 
                        (N115)? mem[2578] : 
                        (N117)? mem[2628] : 
                        (N119)? mem[2678] : 
                        (N121)? mem[2728] : 
                        (N123)? mem[2778] : 
                        (N125)? mem[2828] : 
                        (N127)? mem[2878] : 
                        (N129)? mem[2928] : 
                        (N131)? mem[2978] : 
                        (N133)? mem[3028] : 
                        (N135)? mem[3078] : 
                        (N137)? mem[3128] : 
                        (N139)? mem[3178] : 1'b0;
  assign r_data_o[27] = (N76)? mem[27] : 
                        (N78)? mem[77] : 
                        (N80)? mem[127] : 
                        (N82)? mem[177] : 
                        (N84)? mem[227] : 
                        (N86)? mem[277] : 
                        (N88)? mem[327] : 
                        (N90)? mem[377] : 
                        (N92)? mem[427] : 
                        (N94)? mem[477] : 
                        (N96)? mem[527] : 
                        (N98)? mem[577] : 
                        (N100)? mem[627] : 
                        (N102)? mem[677] : 
                        (N104)? mem[727] : 
                        (N106)? mem[777] : 
                        (N108)? mem[827] : 
                        (N110)? mem[877] : 
                        (N112)? mem[927] : 
                        (N114)? mem[977] : 
                        (N116)? mem[1027] : 
                        (N118)? mem[1077] : 
                        (N120)? mem[1127] : 
                        (N122)? mem[1177] : 
                        (N124)? mem[1227] : 
                        (N126)? mem[1277] : 
                        (N128)? mem[1327] : 
                        (N130)? mem[1377] : 
                        (N132)? mem[1427] : 
                        (N134)? mem[1477] : 
                        (N136)? mem[1527] : 
                        (N138)? mem[1577] : 
                        (N77)? mem[1627] : 
                        (N79)? mem[1677] : 
                        (N81)? mem[1727] : 
                        (N83)? mem[1777] : 
                        (N85)? mem[1827] : 
                        (N87)? mem[1877] : 
                        (N89)? mem[1927] : 
                        (N91)? mem[1977] : 
                        (N93)? mem[2027] : 
                        (N95)? mem[2077] : 
                        (N97)? mem[2127] : 
                        (N99)? mem[2177] : 
                        (N101)? mem[2227] : 
                        (N103)? mem[2277] : 
                        (N105)? mem[2327] : 
                        (N107)? mem[2377] : 
                        (N109)? mem[2427] : 
                        (N111)? mem[2477] : 
                        (N113)? mem[2527] : 
                        (N115)? mem[2577] : 
                        (N117)? mem[2627] : 
                        (N119)? mem[2677] : 
                        (N121)? mem[2727] : 
                        (N123)? mem[2777] : 
                        (N125)? mem[2827] : 
                        (N127)? mem[2877] : 
                        (N129)? mem[2927] : 
                        (N131)? mem[2977] : 
                        (N133)? mem[3027] : 
                        (N135)? mem[3077] : 
                        (N137)? mem[3127] : 
                        (N139)? mem[3177] : 1'b0;
  assign r_data_o[26] = (N76)? mem[26] : 
                        (N78)? mem[76] : 
                        (N80)? mem[126] : 
                        (N82)? mem[176] : 
                        (N84)? mem[226] : 
                        (N86)? mem[276] : 
                        (N88)? mem[326] : 
                        (N90)? mem[376] : 
                        (N92)? mem[426] : 
                        (N94)? mem[476] : 
                        (N96)? mem[526] : 
                        (N98)? mem[576] : 
                        (N100)? mem[626] : 
                        (N102)? mem[676] : 
                        (N104)? mem[726] : 
                        (N106)? mem[776] : 
                        (N108)? mem[826] : 
                        (N110)? mem[876] : 
                        (N112)? mem[926] : 
                        (N114)? mem[976] : 
                        (N116)? mem[1026] : 
                        (N118)? mem[1076] : 
                        (N120)? mem[1126] : 
                        (N122)? mem[1176] : 
                        (N124)? mem[1226] : 
                        (N126)? mem[1276] : 
                        (N128)? mem[1326] : 
                        (N130)? mem[1376] : 
                        (N132)? mem[1426] : 
                        (N134)? mem[1476] : 
                        (N136)? mem[1526] : 
                        (N138)? mem[1576] : 
                        (N77)? mem[1626] : 
                        (N79)? mem[1676] : 
                        (N81)? mem[1726] : 
                        (N83)? mem[1776] : 
                        (N85)? mem[1826] : 
                        (N87)? mem[1876] : 
                        (N89)? mem[1926] : 
                        (N91)? mem[1976] : 
                        (N93)? mem[2026] : 
                        (N95)? mem[2076] : 
                        (N97)? mem[2126] : 
                        (N99)? mem[2176] : 
                        (N101)? mem[2226] : 
                        (N103)? mem[2276] : 
                        (N105)? mem[2326] : 
                        (N107)? mem[2376] : 
                        (N109)? mem[2426] : 
                        (N111)? mem[2476] : 
                        (N113)? mem[2526] : 
                        (N115)? mem[2576] : 
                        (N117)? mem[2626] : 
                        (N119)? mem[2676] : 
                        (N121)? mem[2726] : 
                        (N123)? mem[2776] : 
                        (N125)? mem[2826] : 
                        (N127)? mem[2876] : 
                        (N129)? mem[2926] : 
                        (N131)? mem[2976] : 
                        (N133)? mem[3026] : 
                        (N135)? mem[3076] : 
                        (N137)? mem[3126] : 
                        (N139)? mem[3176] : 1'b0;
  assign r_data_o[25] = (N76)? mem[25] : 
                        (N78)? mem[75] : 
                        (N80)? mem[125] : 
                        (N82)? mem[175] : 
                        (N84)? mem[225] : 
                        (N86)? mem[275] : 
                        (N88)? mem[325] : 
                        (N90)? mem[375] : 
                        (N92)? mem[425] : 
                        (N94)? mem[475] : 
                        (N96)? mem[525] : 
                        (N98)? mem[575] : 
                        (N100)? mem[625] : 
                        (N102)? mem[675] : 
                        (N104)? mem[725] : 
                        (N106)? mem[775] : 
                        (N108)? mem[825] : 
                        (N110)? mem[875] : 
                        (N112)? mem[925] : 
                        (N114)? mem[975] : 
                        (N116)? mem[1025] : 
                        (N118)? mem[1075] : 
                        (N120)? mem[1125] : 
                        (N122)? mem[1175] : 
                        (N124)? mem[1225] : 
                        (N126)? mem[1275] : 
                        (N128)? mem[1325] : 
                        (N130)? mem[1375] : 
                        (N132)? mem[1425] : 
                        (N134)? mem[1475] : 
                        (N136)? mem[1525] : 
                        (N138)? mem[1575] : 
                        (N77)? mem[1625] : 
                        (N79)? mem[1675] : 
                        (N81)? mem[1725] : 
                        (N83)? mem[1775] : 
                        (N85)? mem[1825] : 
                        (N87)? mem[1875] : 
                        (N89)? mem[1925] : 
                        (N91)? mem[1975] : 
                        (N93)? mem[2025] : 
                        (N95)? mem[2075] : 
                        (N97)? mem[2125] : 
                        (N99)? mem[2175] : 
                        (N101)? mem[2225] : 
                        (N103)? mem[2275] : 
                        (N105)? mem[2325] : 
                        (N107)? mem[2375] : 
                        (N109)? mem[2425] : 
                        (N111)? mem[2475] : 
                        (N113)? mem[2525] : 
                        (N115)? mem[2575] : 
                        (N117)? mem[2625] : 
                        (N119)? mem[2675] : 
                        (N121)? mem[2725] : 
                        (N123)? mem[2775] : 
                        (N125)? mem[2825] : 
                        (N127)? mem[2875] : 
                        (N129)? mem[2925] : 
                        (N131)? mem[2975] : 
                        (N133)? mem[3025] : 
                        (N135)? mem[3075] : 
                        (N137)? mem[3125] : 
                        (N139)? mem[3175] : 1'b0;
  assign r_data_o[24] = (N76)? mem[24] : 
                        (N78)? mem[74] : 
                        (N80)? mem[124] : 
                        (N82)? mem[174] : 
                        (N84)? mem[224] : 
                        (N86)? mem[274] : 
                        (N88)? mem[324] : 
                        (N90)? mem[374] : 
                        (N92)? mem[424] : 
                        (N94)? mem[474] : 
                        (N96)? mem[524] : 
                        (N98)? mem[574] : 
                        (N100)? mem[624] : 
                        (N102)? mem[674] : 
                        (N104)? mem[724] : 
                        (N106)? mem[774] : 
                        (N108)? mem[824] : 
                        (N110)? mem[874] : 
                        (N112)? mem[924] : 
                        (N114)? mem[974] : 
                        (N116)? mem[1024] : 
                        (N118)? mem[1074] : 
                        (N120)? mem[1124] : 
                        (N122)? mem[1174] : 
                        (N124)? mem[1224] : 
                        (N126)? mem[1274] : 
                        (N128)? mem[1324] : 
                        (N130)? mem[1374] : 
                        (N132)? mem[1424] : 
                        (N134)? mem[1474] : 
                        (N136)? mem[1524] : 
                        (N138)? mem[1574] : 
                        (N77)? mem[1624] : 
                        (N79)? mem[1674] : 
                        (N81)? mem[1724] : 
                        (N83)? mem[1774] : 
                        (N85)? mem[1824] : 
                        (N87)? mem[1874] : 
                        (N89)? mem[1924] : 
                        (N91)? mem[1974] : 
                        (N93)? mem[2024] : 
                        (N95)? mem[2074] : 
                        (N97)? mem[2124] : 
                        (N99)? mem[2174] : 
                        (N101)? mem[2224] : 
                        (N103)? mem[2274] : 
                        (N105)? mem[2324] : 
                        (N107)? mem[2374] : 
                        (N109)? mem[2424] : 
                        (N111)? mem[2474] : 
                        (N113)? mem[2524] : 
                        (N115)? mem[2574] : 
                        (N117)? mem[2624] : 
                        (N119)? mem[2674] : 
                        (N121)? mem[2724] : 
                        (N123)? mem[2774] : 
                        (N125)? mem[2824] : 
                        (N127)? mem[2874] : 
                        (N129)? mem[2924] : 
                        (N131)? mem[2974] : 
                        (N133)? mem[3024] : 
                        (N135)? mem[3074] : 
                        (N137)? mem[3124] : 
                        (N139)? mem[3174] : 1'b0;
  assign r_data_o[23] = (N76)? mem[23] : 
                        (N78)? mem[73] : 
                        (N80)? mem[123] : 
                        (N82)? mem[173] : 
                        (N84)? mem[223] : 
                        (N86)? mem[273] : 
                        (N88)? mem[323] : 
                        (N90)? mem[373] : 
                        (N92)? mem[423] : 
                        (N94)? mem[473] : 
                        (N96)? mem[523] : 
                        (N98)? mem[573] : 
                        (N100)? mem[623] : 
                        (N102)? mem[673] : 
                        (N104)? mem[723] : 
                        (N106)? mem[773] : 
                        (N108)? mem[823] : 
                        (N110)? mem[873] : 
                        (N112)? mem[923] : 
                        (N114)? mem[973] : 
                        (N116)? mem[1023] : 
                        (N118)? mem[1073] : 
                        (N120)? mem[1123] : 
                        (N122)? mem[1173] : 
                        (N124)? mem[1223] : 
                        (N126)? mem[1273] : 
                        (N128)? mem[1323] : 
                        (N130)? mem[1373] : 
                        (N132)? mem[1423] : 
                        (N134)? mem[1473] : 
                        (N136)? mem[1523] : 
                        (N138)? mem[1573] : 
                        (N77)? mem[1623] : 
                        (N79)? mem[1673] : 
                        (N81)? mem[1723] : 
                        (N83)? mem[1773] : 
                        (N85)? mem[1823] : 
                        (N87)? mem[1873] : 
                        (N89)? mem[1923] : 
                        (N91)? mem[1973] : 
                        (N93)? mem[2023] : 
                        (N95)? mem[2073] : 
                        (N97)? mem[2123] : 
                        (N99)? mem[2173] : 
                        (N101)? mem[2223] : 
                        (N103)? mem[2273] : 
                        (N105)? mem[2323] : 
                        (N107)? mem[2373] : 
                        (N109)? mem[2423] : 
                        (N111)? mem[2473] : 
                        (N113)? mem[2523] : 
                        (N115)? mem[2573] : 
                        (N117)? mem[2623] : 
                        (N119)? mem[2673] : 
                        (N121)? mem[2723] : 
                        (N123)? mem[2773] : 
                        (N125)? mem[2823] : 
                        (N127)? mem[2873] : 
                        (N129)? mem[2923] : 
                        (N131)? mem[2973] : 
                        (N133)? mem[3023] : 
                        (N135)? mem[3073] : 
                        (N137)? mem[3123] : 
                        (N139)? mem[3173] : 1'b0;
  assign r_data_o[22] = (N76)? mem[22] : 
                        (N78)? mem[72] : 
                        (N80)? mem[122] : 
                        (N82)? mem[172] : 
                        (N84)? mem[222] : 
                        (N86)? mem[272] : 
                        (N88)? mem[322] : 
                        (N90)? mem[372] : 
                        (N92)? mem[422] : 
                        (N94)? mem[472] : 
                        (N96)? mem[522] : 
                        (N98)? mem[572] : 
                        (N100)? mem[622] : 
                        (N102)? mem[672] : 
                        (N104)? mem[722] : 
                        (N106)? mem[772] : 
                        (N108)? mem[822] : 
                        (N110)? mem[872] : 
                        (N112)? mem[922] : 
                        (N114)? mem[972] : 
                        (N116)? mem[1022] : 
                        (N118)? mem[1072] : 
                        (N120)? mem[1122] : 
                        (N122)? mem[1172] : 
                        (N124)? mem[1222] : 
                        (N126)? mem[1272] : 
                        (N128)? mem[1322] : 
                        (N130)? mem[1372] : 
                        (N132)? mem[1422] : 
                        (N134)? mem[1472] : 
                        (N136)? mem[1522] : 
                        (N138)? mem[1572] : 
                        (N77)? mem[1622] : 
                        (N79)? mem[1672] : 
                        (N81)? mem[1722] : 
                        (N83)? mem[1772] : 
                        (N85)? mem[1822] : 
                        (N87)? mem[1872] : 
                        (N89)? mem[1922] : 
                        (N91)? mem[1972] : 
                        (N93)? mem[2022] : 
                        (N95)? mem[2072] : 
                        (N97)? mem[2122] : 
                        (N99)? mem[2172] : 
                        (N101)? mem[2222] : 
                        (N103)? mem[2272] : 
                        (N105)? mem[2322] : 
                        (N107)? mem[2372] : 
                        (N109)? mem[2422] : 
                        (N111)? mem[2472] : 
                        (N113)? mem[2522] : 
                        (N115)? mem[2572] : 
                        (N117)? mem[2622] : 
                        (N119)? mem[2672] : 
                        (N121)? mem[2722] : 
                        (N123)? mem[2772] : 
                        (N125)? mem[2822] : 
                        (N127)? mem[2872] : 
                        (N129)? mem[2922] : 
                        (N131)? mem[2972] : 
                        (N133)? mem[3022] : 
                        (N135)? mem[3072] : 
                        (N137)? mem[3122] : 
                        (N139)? mem[3172] : 1'b0;
  assign r_data_o[21] = (N76)? mem[21] : 
                        (N78)? mem[71] : 
                        (N80)? mem[121] : 
                        (N82)? mem[171] : 
                        (N84)? mem[221] : 
                        (N86)? mem[271] : 
                        (N88)? mem[321] : 
                        (N90)? mem[371] : 
                        (N92)? mem[421] : 
                        (N94)? mem[471] : 
                        (N96)? mem[521] : 
                        (N98)? mem[571] : 
                        (N100)? mem[621] : 
                        (N102)? mem[671] : 
                        (N104)? mem[721] : 
                        (N106)? mem[771] : 
                        (N108)? mem[821] : 
                        (N110)? mem[871] : 
                        (N112)? mem[921] : 
                        (N114)? mem[971] : 
                        (N116)? mem[1021] : 
                        (N118)? mem[1071] : 
                        (N120)? mem[1121] : 
                        (N122)? mem[1171] : 
                        (N124)? mem[1221] : 
                        (N126)? mem[1271] : 
                        (N128)? mem[1321] : 
                        (N130)? mem[1371] : 
                        (N132)? mem[1421] : 
                        (N134)? mem[1471] : 
                        (N136)? mem[1521] : 
                        (N138)? mem[1571] : 
                        (N77)? mem[1621] : 
                        (N79)? mem[1671] : 
                        (N81)? mem[1721] : 
                        (N83)? mem[1771] : 
                        (N85)? mem[1821] : 
                        (N87)? mem[1871] : 
                        (N89)? mem[1921] : 
                        (N91)? mem[1971] : 
                        (N93)? mem[2021] : 
                        (N95)? mem[2071] : 
                        (N97)? mem[2121] : 
                        (N99)? mem[2171] : 
                        (N101)? mem[2221] : 
                        (N103)? mem[2271] : 
                        (N105)? mem[2321] : 
                        (N107)? mem[2371] : 
                        (N109)? mem[2421] : 
                        (N111)? mem[2471] : 
                        (N113)? mem[2521] : 
                        (N115)? mem[2571] : 
                        (N117)? mem[2621] : 
                        (N119)? mem[2671] : 
                        (N121)? mem[2721] : 
                        (N123)? mem[2771] : 
                        (N125)? mem[2821] : 
                        (N127)? mem[2871] : 
                        (N129)? mem[2921] : 
                        (N131)? mem[2971] : 
                        (N133)? mem[3021] : 
                        (N135)? mem[3071] : 
                        (N137)? mem[3121] : 
                        (N139)? mem[3171] : 1'b0;
  assign r_data_o[20] = (N76)? mem[20] : 
                        (N78)? mem[70] : 
                        (N80)? mem[120] : 
                        (N82)? mem[170] : 
                        (N84)? mem[220] : 
                        (N86)? mem[270] : 
                        (N88)? mem[320] : 
                        (N90)? mem[370] : 
                        (N92)? mem[420] : 
                        (N94)? mem[470] : 
                        (N96)? mem[520] : 
                        (N98)? mem[570] : 
                        (N100)? mem[620] : 
                        (N102)? mem[670] : 
                        (N104)? mem[720] : 
                        (N106)? mem[770] : 
                        (N108)? mem[820] : 
                        (N110)? mem[870] : 
                        (N112)? mem[920] : 
                        (N114)? mem[970] : 
                        (N116)? mem[1020] : 
                        (N118)? mem[1070] : 
                        (N120)? mem[1120] : 
                        (N122)? mem[1170] : 
                        (N124)? mem[1220] : 
                        (N126)? mem[1270] : 
                        (N128)? mem[1320] : 
                        (N130)? mem[1370] : 
                        (N132)? mem[1420] : 
                        (N134)? mem[1470] : 
                        (N136)? mem[1520] : 
                        (N138)? mem[1570] : 
                        (N77)? mem[1620] : 
                        (N79)? mem[1670] : 
                        (N81)? mem[1720] : 
                        (N83)? mem[1770] : 
                        (N85)? mem[1820] : 
                        (N87)? mem[1870] : 
                        (N89)? mem[1920] : 
                        (N91)? mem[1970] : 
                        (N93)? mem[2020] : 
                        (N95)? mem[2070] : 
                        (N97)? mem[2120] : 
                        (N99)? mem[2170] : 
                        (N101)? mem[2220] : 
                        (N103)? mem[2270] : 
                        (N105)? mem[2320] : 
                        (N107)? mem[2370] : 
                        (N109)? mem[2420] : 
                        (N111)? mem[2470] : 
                        (N113)? mem[2520] : 
                        (N115)? mem[2570] : 
                        (N117)? mem[2620] : 
                        (N119)? mem[2670] : 
                        (N121)? mem[2720] : 
                        (N123)? mem[2770] : 
                        (N125)? mem[2820] : 
                        (N127)? mem[2870] : 
                        (N129)? mem[2920] : 
                        (N131)? mem[2970] : 
                        (N133)? mem[3020] : 
                        (N135)? mem[3070] : 
                        (N137)? mem[3120] : 
                        (N139)? mem[3170] : 1'b0;
  assign r_data_o[19] = (N76)? mem[19] : 
                        (N78)? mem[69] : 
                        (N80)? mem[119] : 
                        (N82)? mem[169] : 
                        (N84)? mem[219] : 
                        (N86)? mem[269] : 
                        (N88)? mem[319] : 
                        (N90)? mem[369] : 
                        (N92)? mem[419] : 
                        (N94)? mem[469] : 
                        (N96)? mem[519] : 
                        (N98)? mem[569] : 
                        (N100)? mem[619] : 
                        (N102)? mem[669] : 
                        (N104)? mem[719] : 
                        (N106)? mem[769] : 
                        (N108)? mem[819] : 
                        (N110)? mem[869] : 
                        (N112)? mem[919] : 
                        (N114)? mem[969] : 
                        (N116)? mem[1019] : 
                        (N118)? mem[1069] : 
                        (N120)? mem[1119] : 
                        (N122)? mem[1169] : 
                        (N124)? mem[1219] : 
                        (N126)? mem[1269] : 
                        (N128)? mem[1319] : 
                        (N130)? mem[1369] : 
                        (N132)? mem[1419] : 
                        (N134)? mem[1469] : 
                        (N136)? mem[1519] : 
                        (N138)? mem[1569] : 
                        (N77)? mem[1619] : 
                        (N79)? mem[1669] : 
                        (N81)? mem[1719] : 
                        (N83)? mem[1769] : 
                        (N85)? mem[1819] : 
                        (N87)? mem[1869] : 
                        (N89)? mem[1919] : 
                        (N91)? mem[1969] : 
                        (N93)? mem[2019] : 
                        (N95)? mem[2069] : 
                        (N97)? mem[2119] : 
                        (N99)? mem[2169] : 
                        (N101)? mem[2219] : 
                        (N103)? mem[2269] : 
                        (N105)? mem[2319] : 
                        (N107)? mem[2369] : 
                        (N109)? mem[2419] : 
                        (N111)? mem[2469] : 
                        (N113)? mem[2519] : 
                        (N115)? mem[2569] : 
                        (N117)? mem[2619] : 
                        (N119)? mem[2669] : 
                        (N121)? mem[2719] : 
                        (N123)? mem[2769] : 
                        (N125)? mem[2819] : 
                        (N127)? mem[2869] : 
                        (N129)? mem[2919] : 
                        (N131)? mem[2969] : 
                        (N133)? mem[3019] : 
                        (N135)? mem[3069] : 
                        (N137)? mem[3119] : 
                        (N139)? mem[3169] : 1'b0;
  assign r_data_o[18] = (N76)? mem[18] : 
                        (N78)? mem[68] : 
                        (N80)? mem[118] : 
                        (N82)? mem[168] : 
                        (N84)? mem[218] : 
                        (N86)? mem[268] : 
                        (N88)? mem[318] : 
                        (N90)? mem[368] : 
                        (N92)? mem[418] : 
                        (N94)? mem[468] : 
                        (N96)? mem[518] : 
                        (N98)? mem[568] : 
                        (N100)? mem[618] : 
                        (N102)? mem[668] : 
                        (N104)? mem[718] : 
                        (N106)? mem[768] : 
                        (N108)? mem[818] : 
                        (N110)? mem[868] : 
                        (N112)? mem[918] : 
                        (N114)? mem[968] : 
                        (N116)? mem[1018] : 
                        (N118)? mem[1068] : 
                        (N120)? mem[1118] : 
                        (N122)? mem[1168] : 
                        (N124)? mem[1218] : 
                        (N126)? mem[1268] : 
                        (N128)? mem[1318] : 
                        (N130)? mem[1368] : 
                        (N132)? mem[1418] : 
                        (N134)? mem[1468] : 
                        (N136)? mem[1518] : 
                        (N138)? mem[1568] : 
                        (N77)? mem[1618] : 
                        (N79)? mem[1668] : 
                        (N81)? mem[1718] : 
                        (N83)? mem[1768] : 
                        (N85)? mem[1818] : 
                        (N87)? mem[1868] : 
                        (N89)? mem[1918] : 
                        (N91)? mem[1968] : 
                        (N93)? mem[2018] : 
                        (N95)? mem[2068] : 
                        (N97)? mem[2118] : 
                        (N99)? mem[2168] : 
                        (N101)? mem[2218] : 
                        (N103)? mem[2268] : 
                        (N105)? mem[2318] : 
                        (N107)? mem[2368] : 
                        (N109)? mem[2418] : 
                        (N111)? mem[2468] : 
                        (N113)? mem[2518] : 
                        (N115)? mem[2568] : 
                        (N117)? mem[2618] : 
                        (N119)? mem[2668] : 
                        (N121)? mem[2718] : 
                        (N123)? mem[2768] : 
                        (N125)? mem[2818] : 
                        (N127)? mem[2868] : 
                        (N129)? mem[2918] : 
                        (N131)? mem[2968] : 
                        (N133)? mem[3018] : 
                        (N135)? mem[3068] : 
                        (N137)? mem[3118] : 
                        (N139)? mem[3168] : 1'b0;
  assign r_data_o[17] = (N76)? mem[17] : 
                        (N78)? mem[67] : 
                        (N80)? mem[117] : 
                        (N82)? mem[167] : 
                        (N84)? mem[217] : 
                        (N86)? mem[267] : 
                        (N88)? mem[317] : 
                        (N90)? mem[367] : 
                        (N92)? mem[417] : 
                        (N94)? mem[467] : 
                        (N96)? mem[517] : 
                        (N98)? mem[567] : 
                        (N100)? mem[617] : 
                        (N102)? mem[667] : 
                        (N104)? mem[717] : 
                        (N106)? mem[767] : 
                        (N108)? mem[817] : 
                        (N110)? mem[867] : 
                        (N112)? mem[917] : 
                        (N114)? mem[967] : 
                        (N116)? mem[1017] : 
                        (N118)? mem[1067] : 
                        (N120)? mem[1117] : 
                        (N122)? mem[1167] : 
                        (N124)? mem[1217] : 
                        (N126)? mem[1267] : 
                        (N128)? mem[1317] : 
                        (N130)? mem[1367] : 
                        (N132)? mem[1417] : 
                        (N134)? mem[1467] : 
                        (N136)? mem[1517] : 
                        (N138)? mem[1567] : 
                        (N77)? mem[1617] : 
                        (N79)? mem[1667] : 
                        (N81)? mem[1717] : 
                        (N83)? mem[1767] : 
                        (N85)? mem[1817] : 
                        (N87)? mem[1867] : 
                        (N89)? mem[1917] : 
                        (N91)? mem[1967] : 
                        (N93)? mem[2017] : 
                        (N95)? mem[2067] : 
                        (N97)? mem[2117] : 
                        (N99)? mem[2167] : 
                        (N101)? mem[2217] : 
                        (N103)? mem[2267] : 
                        (N105)? mem[2317] : 
                        (N107)? mem[2367] : 
                        (N109)? mem[2417] : 
                        (N111)? mem[2467] : 
                        (N113)? mem[2517] : 
                        (N115)? mem[2567] : 
                        (N117)? mem[2617] : 
                        (N119)? mem[2667] : 
                        (N121)? mem[2717] : 
                        (N123)? mem[2767] : 
                        (N125)? mem[2817] : 
                        (N127)? mem[2867] : 
                        (N129)? mem[2917] : 
                        (N131)? mem[2967] : 
                        (N133)? mem[3017] : 
                        (N135)? mem[3067] : 
                        (N137)? mem[3117] : 
                        (N139)? mem[3167] : 1'b0;
  assign r_data_o[16] = (N76)? mem[16] : 
                        (N78)? mem[66] : 
                        (N80)? mem[116] : 
                        (N82)? mem[166] : 
                        (N84)? mem[216] : 
                        (N86)? mem[266] : 
                        (N88)? mem[316] : 
                        (N90)? mem[366] : 
                        (N92)? mem[416] : 
                        (N94)? mem[466] : 
                        (N96)? mem[516] : 
                        (N98)? mem[566] : 
                        (N100)? mem[616] : 
                        (N102)? mem[666] : 
                        (N104)? mem[716] : 
                        (N106)? mem[766] : 
                        (N108)? mem[816] : 
                        (N110)? mem[866] : 
                        (N112)? mem[916] : 
                        (N114)? mem[966] : 
                        (N116)? mem[1016] : 
                        (N118)? mem[1066] : 
                        (N120)? mem[1116] : 
                        (N122)? mem[1166] : 
                        (N124)? mem[1216] : 
                        (N126)? mem[1266] : 
                        (N128)? mem[1316] : 
                        (N130)? mem[1366] : 
                        (N132)? mem[1416] : 
                        (N134)? mem[1466] : 
                        (N136)? mem[1516] : 
                        (N138)? mem[1566] : 
                        (N77)? mem[1616] : 
                        (N79)? mem[1666] : 
                        (N81)? mem[1716] : 
                        (N83)? mem[1766] : 
                        (N85)? mem[1816] : 
                        (N87)? mem[1866] : 
                        (N89)? mem[1916] : 
                        (N91)? mem[1966] : 
                        (N93)? mem[2016] : 
                        (N95)? mem[2066] : 
                        (N97)? mem[2116] : 
                        (N99)? mem[2166] : 
                        (N101)? mem[2216] : 
                        (N103)? mem[2266] : 
                        (N105)? mem[2316] : 
                        (N107)? mem[2366] : 
                        (N109)? mem[2416] : 
                        (N111)? mem[2466] : 
                        (N113)? mem[2516] : 
                        (N115)? mem[2566] : 
                        (N117)? mem[2616] : 
                        (N119)? mem[2666] : 
                        (N121)? mem[2716] : 
                        (N123)? mem[2766] : 
                        (N125)? mem[2816] : 
                        (N127)? mem[2866] : 
                        (N129)? mem[2916] : 
                        (N131)? mem[2966] : 
                        (N133)? mem[3016] : 
                        (N135)? mem[3066] : 
                        (N137)? mem[3116] : 
                        (N139)? mem[3166] : 1'b0;
  assign r_data_o[15] = (N76)? mem[15] : 
                        (N78)? mem[65] : 
                        (N80)? mem[115] : 
                        (N82)? mem[165] : 
                        (N84)? mem[215] : 
                        (N86)? mem[265] : 
                        (N88)? mem[315] : 
                        (N90)? mem[365] : 
                        (N92)? mem[415] : 
                        (N94)? mem[465] : 
                        (N96)? mem[515] : 
                        (N98)? mem[565] : 
                        (N100)? mem[615] : 
                        (N102)? mem[665] : 
                        (N104)? mem[715] : 
                        (N106)? mem[765] : 
                        (N108)? mem[815] : 
                        (N110)? mem[865] : 
                        (N112)? mem[915] : 
                        (N114)? mem[965] : 
                        (N116)? mem[1015] : 
                        (N118)? mem[1065] : 
                        (N120)? mem[1115] : 
                        (N122)? mem[1165] : 
                        (N124)? mem[1215] : 
                        (N126)? mem[1265] : 
                        (N128)? mem[1315] : 
                        (N130)? mem[1365] : 
                        (N132)? mem[1415] : 
                        (N134)? mem[1465] : 
                        (N136)? mem[1515] : 
                        (N138)? mem[1565] : 
                        (N77)? mem[1615] : 
                        (N79)? mem[1665] : 
                        (N81)? mem[1715] : 
                        (N83)? mem[1765] : 
                        (N85)? mem[1815] : 
                        (N87)? mem[1865] : 
                        (N89)? mem[1915] : 
                        (N91)? mem[1965] : 
                        (N93)? mem[2015] : 
                        (N95)? mem[2065] : 
                        (N97)? mem[2115] : 
                        (N99)? mem[2165] : 
                        (N101)? mem[2215] : 
                        (N103)? mem[2265] : 
                        (N105)? mem[2315] : 
                        (N107)? mem[2365] : 
                        (N109)? mem[2415] : 
                        (N111)? mem[2465] : 
                        (N113)? mem[2515] : 
                        (N115)? mem[2565] : 
                        (N117)? mem[2615] : 
                        (N119)? mem[2665] : 
                        (N121)? mem[2715] : 
                        (N123)? mem[2765] : 
                        (N125)? mem[2815] : 
                        (N127)? mem[2865] : 
                        (N129)? mem[2915] : 
                        (N131)? mem[2965] : 
                        (N133)? mem[3015] : 
                        (N135)? mem[3065] : 
                        (N137)? mem[3115] : 
                        (N139)? mem[3165] : 1'b0;
  assign r_data_o[14] = (N76)? mem[14] : 
                        (N78)? mem[64] : 
                        (N80)? mem[114] : 
                        (N82)? mem[164] : 
                        (N84)? mem[214] : 
                        (N86)? mem[264] : 
                        (N88)? mem[314] : 
                        (N90)? mem[364] : 
                        (N92)? mem[414] : 
                        (N94)? mem[464] : 
                        (N96)? mem[514] : 
                        (N98)? mem[564] : 
                        (N100)? mem[614] : 
                        (N102)? mem[664] : 
                        (N104)? mem[714] : 
                        (N106)? mem[764] : 
                        (N108)? mem[814] : 
                        (N110)? mem[864] : 
                        (N112)? mem[914] : 
                        (N114)? mem[964] : 
                        (N116)? mem[1014] : 
                        (N118)? mem[1064] : 
                        (N120)? mem[1114] : 
                        (N122)? mem[1164] : 
                        (N124)? mem[1214] : 
                        (N126)? mem[1264] : 
                        (N128)? mem[1314] : 
                        (N130)? mem[1364] : 
                        (N132)? mem[1414] : 
                        (N134)? mem[1464] : 
                        (N136)? mem[1514] : 
                        (N138)? mem[1564] : 
                        (N77)? mem[1614] : 
                        (N79)? mem[1664] : 
                        (N81)? mem[1714] : 
                        (N83)? mem[1764] : 
                        (N85)? mem[1814] : 
                        (N87)? mem[1864] : 
                        (N89)? mem[1914] : 
                        (N91)? mem[1964] : 
                        (N93)? mem[2014] : 
                        (N95)? mem[2064] : 
                        (N97)? mem[2114] : 
                        (N99)? mem[2164] : 
                        (N101)? mem[2214] : 
                        (N103)? mem[2264] : 
                        (N105)? mem[2314] : 
                        (N107)? mem[2364] : 
                        (N109)? mem[2414] : 
                        (N111)? mem[2464] : 
                        (N113)? mem[2514] : 
                        (N115)? mem[2564] : 
                        (N117)? mem[2614] : 
                        (N119)? mem[2664] : 
                        (N121)? mem[2714] : 
                        (N123)? mem[2764] : 
                        (N125)? mem[2814] : 
                        (N127)? mem[2864] : 
                        (N129)? mem[2914] : 
                        (N131)? mem[2964] : 
                        (N133)? mem[3014] : 
                        (N135)? mem[3064] : 
                        (N137)? mem[3114] : 
                        (N139)? mem[3164] : 1'b0;
  assign r_data_o[13] = (N76)? mem[13] : 
                        (N78)? mem[63] : 
                        (N80)? mem[113] : 
                        (N82)? mem[163] : 
                        (N84)? mem[213] : 
                        (N86)? mem[263] : 
                        (N88)? mem[313] : 
                        (N90)? mem[363] : 
                        (N92)? mem[413] : 
                        (N94)? mem[463] : 
                        (N96)? mem[513] : 
                        (N98)? mem[563] : 
                        (N100)? mem[613] : 
                        (N102)? mem[663] : 
                        (N104)? mem[713] : 
                        (N106)? mem[763] : 
                        (N108)? mem[813] : 
                        (N110)? mem[863] : 
                        (N112)? mem[913] : 
                        (N114)? mem[963] : 
                        (N116)? mem[1013] : 
                        (N118)? mem[1063] : 
                        (N120)? mem[1113] : 
                        (N122)? mem[1163] : 
                        (N124)? mem[1213] : 
                        (N126)? mem[1263] : 
                        (N128)? mem[1313] : 
                        (N130)? mem[1363] : 
                        (N132)? mem[1413] : 
                        (N134)? mem[1463] : 
                        (N136)? mem[1513] : 
                        (N138)? mem[1563] : 
                        (N77)? mem[1613] : 
                        (N79)? mem[1663] : 
                        (N81)? mem[1713] : 
                        (N83)? mem[1763] : 
                        (N85)? mem[1813] : 
                        (N87)? mem[1863] : 
                        (N89)? mem[1913] : 
                        (N91)? mem[1963] : 
                        (N93)? mem[2013] : 
                        (N95)? mem[2063] : 
                        (N97)? mem[2113] : 
                        (N99)? mem[2163] : 
                        (N101)? mem[2213] : 
                        (N103)? mem[2263] : 
                        (N105)? mem[2313] : 
                        (N107)? mem[2363] : 
                        (N109)? mem[2413] : 
                        (N111)? mem[2463] : 
                        (N113)? mem[2513] : 
                        (N115)? mem[2563] : 
                        (N117)? mem[2613] : 
                        (N119)? mem[2663] : 
                        (N121)? mem[2713] : 
                        (N123)? mem[2763] : 
                        (N125)? mem[2813] : 
                        (N127)? mem[2863] : 
                        (N129)? mem[2913] : 
                        (N131)? mem[2963] : 
                        (N133)? mem[3013] : 
                        (N135)? mem[3063] : 
                        (N137)? mem[3113] : 
                        (N139)? mem[3163] : 1'b0;
  assign r_data_o[12] = (N76)? mem[12] : 
                        (N78)? mem[62] : 
                        (N80)? mem[112] : 
                        (N82)? mem[162] : 
                        (N84)? mem[212] : 
                        (N86)? mem[262] : 
                        (N88)? mem[312] : 
                        (N90)? mem[362] : 
                        (N92)? mem[412] : 
                        (N94)? mem[462] : 
                        (N96)? mem[512] : 
                        (N98)? mem[562] : 
                        (N100)? mem[612] : 
                        (N102)? mem[662] : 
                        (N104)? mem[712] : 
                        (N106)? mem[762] : 
                        (N108)? mem[812] : 
                        (N110)? mem[862] : 
                        (N112)? mem[912] : 
                        (N114)? mem[962] : 
                        (N116)? mem[1012] : 
                        (N118)? mem[1062] : 
                        (N120)? mem[1112] : 
                        (N122)? mem[1162] : 
                        (N124)? mem[1212] : 
                        (N126)? mem[1262] : 
                        (N128)? mem[1312] : 
                        (N130)? mem[1362] : 
                        (N132)? mem[1412] : 
                        (N134)? mem[1462] : 
                        (N136)? mem[1512] : 
                        (N138)? mem[1562] : 
                        (N77)? mem[1612] : 
                        (N79)? mem[1662] : 
                        (N81)? mem[1712] : 
                        (N83)? mem[1762] : 
                        (N85)? mem[1812] : 
                        (N87)? mem[1862] : 
                        (N89)? mem[1912] : 
                        (N91)? mem[1962] : 
                        (N93)? mem[2012] : 
                        (N95)? mem[2062] : 
                        (N97)? mem[2112] : 
                        (N99)? mem[2162] : 
                        (N101)? mem[2212] : 
                        (N103)? mem[2262] : 
                        (N105)? mem[2312] : 
                        (N107)? mem[2362] : 
                        (N109)? mem[2412] : 
                        (N111)? mem[2462] : 
                        (N113)? mem[2512] : 
                        (N115)? mem[2562] : 
                        (N117)? mem[2612] : 
                        (N119)? mem[2662] : 
                        (N121)? mem[2712] : 
                        (N123)? mem[2762] : 
                        (N125)? mem[2812] : 
                        (N127)? mem[2862] : 
                        (N129)? mem[2912] : 
                        (N131)? mem[2962] : 
                        (N133)? mem[3012] : 
                        (N135)? mem[3062] : 
                        (N137)? mem[3112] : 
                        (N139)? mem[3162] : 1'b0;
  assign r_data_o[11] = (N76)? mem[11] : 
                        (N78)? mem[61] : 
                        (N80)? mem[111] : 
                        (N82)? mem[161] : 
                        (N84)? mem[211] : 
                        (N86)? mem[261] : 
                        (N88)? mem[311] : 
                        (N90)? mem[361] : 
                        (N92)? mem[411] : 
                        (N94)? mem[461] : 
                        (N96)? mem[511] : 
                        (N98)? mem[561] : 
                        (N100)? mem[611] : 
                        (N102)? mem[661] : 
                        (N104)? mem[711] : 
                        (N106)? mem[761] : 
                        (N108)? mem[811] : 
                        (N110)? mem[861] : 
                        (N112)? mem[911] : 
                        (N114)? mem[961] : 
                        (N116)? mem[1011] : 
                        (N118)? mem[1061] : 
                        (N120)? mem[1111] : 
                        (N122)? mem[1161] : 
                        (N124)? mem[1211] : 
                        (N126)? mem[1261] : 
                        (N128)? mem[1311] : 
                        (N130)? mem[1361] : 
                        (N132)? mem[1411] : 
                        (N134)? mem[1461] : 
                        (N136)? mem[1511] : 
                        (N138)? mem[1561] : 
                        (N77)? mem[1611] : 
                        (N79)? mem[1661] : 
                        (N81)? mem[1711] : 
                        (N83)? mem[1761] : 
                        (N85)? mem[1811] : 
                        (N87)? mem[1861] : 
                        (N89)? mem[1911] : 
                        (N91)? mem[1961] : 
                        (N93)? mem[2011] : 
                        (N95)? mem[2061] : 
                        (N97)? mem[2111] : 
                        (N99)? mem[2161] : 
                        (N101)? mem[2211] : 
                        (N103)? mem[2261] : 
                        (N105)? mem[2311] : 
                        (N107)? mem[2361] : 
                        (N109)? mem[2411] : 
                        (N111)? mem[2461] : 
                        (N113)? mem[2511] : 
                        (N115)? mem[2561] : 
                        (N117)? mem[2611] : 
                        (N119)? mem[2661] : 
                        (N121)? mem[2711] : 
                        (N123)? mem[2761] : 
                        (N125)? mem[2811] : 
                        (N127)? mem[2861] : 
                        (N129)? mem[2911] : 
                        (N131)? mem[2961] : 
                        (N133)? mem[3011] : 
                        (N135)? mem[3061] : 
                        (N137)? mem[3111] : 
                        (N139)? mem[3161] : 1'b0;
  assign r_data_o[10] = (N76)? mem[10] : 
                        (N78)? mem[60] : 
                        (N80)? mem[110] : 
                        (N82)? mem[160] : 
                        (N84)? mem[210] : 
                        (N86)? mem[260] : 
                        (N88)? mem[310] : 
                        (N90)? mem[360] : 
                        (N92)? mem[410] : 
                        (N94)? mem[460] : 
                        (N96)? mem[510] : 
                        (N98)? mem[560] : 
                        (N100)? mem[610] : 
                        (N102)? mem[660] : 
                        (N104)? mem[710] : 
                        (N106)? mem[760] : 
                        (N108)? mem[810] : 
                        (N110)? mem[860] : 
                        (N112)? mem[910] : 
                        (N114)? mem[960] : 
                        (N116)? mem[1010] : 
                        (N118)? mem[1060] : 
                        (N120)? mem[1110] : 
                        (N122)? mem[1160] : 
                        (N124)? mem[1210] : 
                        (N126)? mem[1260] : 
                        (N128)? mem[1310] : 
                        (N130)? mem[1360] : 
                        (N132)? mem[1410] : 
                        (N134)? mem[1460] : 
                        (N136)? mem[1510] : 
                        (N138)? mem[1560] : 
                        (N77)? mem[1610] : 
                        (N79)? mem[1660] : 
                        (N81)? mem[1710] : 
                        (N83)? mem[1760] : 
                        (N85)? mem[1810] : 
                        (N87)? mem[1860] : 
                        (N89)? mem[1910] : 
                        (N91)? mem[1960] : 
                        (N93)? mem[2010] : 
                        (N95)? mem[2060] : 
                        (N97)? mem[2110] : 
                        (N99)? mem[2160] : 
                        (N101)? mem[2210] : 
                        (N103)? mem[2260] : 
                        (N105)? mem[2310] : 
                        (N107)? mem[2360] : 
                        (N109)? mem[2410] : 
                        (N111)? mem[2460] : 
                        (N113)? mem[2510] : 
                        (N115)? mem[2560] : 
                        (N117)? mem[2610] : 
                        (N119)? mem[2660] : 
                        (N121)? mem[2710] : 
                        (N123)? mem[2760] : 
                        (N125)? mem[2810] : 
                        (N127)? mem[2860] : 
                        (N129)? mem[2910] : 
                        (N131)? mem[2960] : 
                        (N133)? mem[3010] : 
                        (N135)? mem[3060] : 
                        (N137)? mem[3110] : 
                        (N139)? mem[3160] : 1'b0;
  assign r_data_o[9] = (N76)? mem[9] : 
                       (N78)? mem[59] : 
                       (N80)? mem[109] : 
                       (N82)? mem[159] : 
                       (N84)? mem[209] : 
                       (N86)? mem[259] : 
                       (N88)? mem[309] : 
                       (N90)? mem[359] : 
                       (N92)? mem[409] : 
                       (N94)? mem[459] : 
                       (N96)? mem[509] : 
                       (N98)? mem[559] : 
                       (N100)? mem[609] : 
                       (N102)? mem[659] : 
                       (N104)? mem[709] : 
                       (N106)? mem[759] : 
                       (N108)? mem[809] : 
                       (N110)? mem[859] : 
                       (N112)? mem[909] : 
                       (N114)? mem[959] : 
                       (N116)? mem[1009] : 
                       (N118)? mem[1059] : 
                       (N120)? mem[1109] : 
                       (N122)? mem[1159] : 
                       (N124)? mem[1209] : 
                       (N126)? mem[1259] : 
                       (N128)? mem[1309] : 
                       (N130)? mem[1359] : 
                       (N132)? mem[1409] : 
                       (N134)? mem[1459] : 
                       (N136)? mem[1509] : 
                       (N138)? mem[1559] : 
                       (N77)? mem[1609] : 
                       (N79)? mem[1659] : 
                       (N81)? mem[1709] : 
                       (N83)? mem[1759] : 
                       (N85)? mem[1809] : 
                       (N87)? mem[1859] : 
                       (N89)? mem[1909] : 
                       (N91)? mem[1959] : 
                       (N93)? mem[2009] : 
                       (N95)? mem[2059] : 
                       (N97)? mem[2109] : 
                       (N99)? mem[2159] : 
                       (N101)? mem[2209] : 
                       (N103)? mem[2259] : 
                       (N105)? mem[2309] : 
                       (N107)? mem[2359] : 
                       (N109)? mem[2409] : 
                       (N111)? mem[2459] : 
                       (N113)? mem[2509] : 
                       (N115)? mem[2559] : 
                       (N117)? mem[2609] : 
                       (N119)? mem[2659] : 
                       (N121)? mem[2709] : 
                       (N123)? mem[2759] : 
                       (N125)? mem[2809] : 
                       (N127)? mem[2859] : 
                       (N129)? mem[2909] : 
                       (N131)? mem[2959] : 
                       (N133)? mem[3009] : 
                       (N135)? mem[3059] : 
                       (N137)? mem[3109] : 
                       (N139)? mem[3159] : 1'b0;
  assign r_data_o[8] = (N76)? mem[8] : 
                       (N78)? mem[58] : 
                       (N80)? mem[108] : 
                       (N82)? mem[158] : 
                       (N84)? mem[208] : 
                       (N86)? mem[258] : 
                       (N88)? mem[308] : 
                       (N90)? mem[358] : 
                       (N92)? mem[408] : 
                       (N94)? mem[458] : 
                       (N96)? mem[508] : 
                       (N98)? mem[558] : 
                       (N100)? mem[608] : 
                       (N102)? mem[658] : 
                       (N104)? mem[708] : 
                       (N106)? mem[758] : 
                       (N108)? mem[808] : 
                       (N110)? mem[858] : 
                       (N112)? mem[908] : 
                       (N114)? mem[958] : 
                       (N116)? mem[1008] : 
                       (N118)? mem[1058] : 
                       (N120)? mem[1108] : 
                       (N122)? mem[1158] : 
                       (N124)? mem[1208] : 
                       (N126)? mem[1258] : 
                       (N128)? mem[1308] : 
                       (N130)? mem[1358] : 
                       (N132)? mem[1408] : 
                       (N134)? mem[1458] : 
                       (N136)? mem[1508] : 
                       (N138)? mem[1558] : 
                       (N77)? mem[1608] : 
                       (N79)? mem[1658] : 
                       (N81)? mem[1708] : 
                       (N83)? mem[1758] : 
                       (N85)? mem[1808] : 
                       (N87)? mem[1858] : 
                       (N89)? mem[1908] : 
                       (N91)? mem[1958] : 
                       (N93)? mem[2008] : 
                       (N95)? mem[2058] : 
                       (N97)? mem[2108] : 
                       (N99)? mem[2158] : 
                       (N101)? mem[2208] : 
                       (N103)? mem[2258] : 
                       (N105)? mem[2308] : 
                       (N107)? mem[2358] : 
                       (N109)? mem[2408] : 
                       (N111)? mem[2458] : 
                       (N113)? mem[2508] : 
                       (N115)? mem[2558] : 
                       (N117)? mem[2608] : 
                       (N119)? mem[2658] : 
                       (N121)? mem[2708] : 
                       (N123)? mem[2758] : 
                       (N125)? mem[2808] : 
                       (N127)? mem[2858] : 
                       (N129)? mem[2908] : 
                       (N131)? mem[2958] : 
                       (N133)? mem[3008] : 
                       (N135)? mem[3058] : 
                       (N137)? mem[3108] : 
                       (N139)? mem[3158] : 1'b0;
  assign r_data_o[7] = (N76)? mem[7] : 
                       (N78)? mem[57] : 
                       (N80)? mem[107] : 
                       (N82)? mem[157] : 
                       (N84)? mem[207] : 
                       (N86)? mem[257] : 
                       (N88)? mem[307] : 
                       (N90)? mem[357] : 
                       (N92)? mem[407] : 
                       (N94)? mem[457] : 
                       (N96)? mem[507] : 
                       (N98)? mem[557] : 
                       (N100)? mem[607] : 
                       (N102)? mem[657] : 
                       (N104)? mem[707] : 
                       (N106)? mem[757] : 
                       (N108)? mem[807] : 
                       (N110)? mem[857] : 
                       (N112)? mem[907] : 
                       (N114)? mem[957] : 
                       (N116)? mem[1007] : 
                       (N118)? mem[1057] : 
                       (N120)? mem[1107] : 
                       (N122)? mem[1157] : 
                       (N124)? mem[1207] : 
                       (N126)? mem[1257] : 
                       (N128)? mem[1307] : 
                       (N130)? mem[1357] : 
                       (N132)? mem[1407] : 
                       (N134)? mem[1457] : 
                       (N136)? mem[1507] : 
                       (N138)? mem[1557] : 
                       (N77)? mem[1607] : 
                       (N79)? mem[1657] : 
                       (N81)? mem[1707] : 
                       (N83)? mem[1757] : 
                       (N85)? mem[1807] : 
                       (N87)? mem[1857] : 
                       (N89)? mem[1907] : 
                       (N91)? mem[1957] : 
                       (N93)? mem[2007] : 
                       (N95)? mem[2057] : 
                       (N97)? mem[2107] : 
                       (N99)? mem[2157] : 
                       (N101)? mem[2207] : 
                       (N103)? mem[2257] : 
                       (N105)? mem[2307] : 
                       (N107)? mem[2357] : 
                       (N109)? mem[2407] : 
                       (N111)? mem[2457] : 
                       (N113)? mem[2507] : 
                       (N115)? mem[2557] : 
                       (N117)? mem[2607] : 
                       (N119)? mem[2657] : 
                       (N121)? mem[2707] : 
                       (N123)? mem[2757] : 
                       (N125)? mem[2807] : 
                       (N127)? mem[2857] : 
                       (N129)? mem[2907] : 
                       (N131)? mem[2957] : 
                       (N133)? mem[3007] : 
                       (N135)? mem[3057] : 
                       (N137)? mem[3107] : 
                       (N139)? mem[3157] : 1'b0;
  assign r_data_o[6] = (N76)? mem[6] : 
                       (N78)? mem[56] : 
                       (N80)? mem[106] : 
                       (N82)? mem[156] : 
                       (N84)? mem[206] : 
                       (N86)? mem[256] : 
                       (N88)? mem[306] : 
                       (N90)? mem[356] : 
                       (N92)? mem[406] : 
                       (N94)? mem[456] : 
                       (N96)? mem[506] : 
                       (N98)? mem[556] : 
                       (N100)? mem[606] : 
                       (N102)? mem[656] : 
                       (N104)? mem[706] : 
                       (N106)? mem[756] : 
                       (N108)? mem[806] : 
                       (N110)? mem[856] : 
                       (N112)? mem[906] : 
                       (N114)? mem[956] : 
                       (N116)? mem[1006] : 
                       (N118)? mem[1056] : 
                       (N120)? mem[1106] : 
                       (N122)? mem[1156] : 
                       (N124)? mem[1206] : 
                       (N126)? mem[1256] : 
                       (N128)? mem[1306] : 
                       (N130)? mem[1356] : 
                       (N132)? mem[1406] : 
                       (N134)? mem[1456] : 
                       (N136)? mem[1506] : 
                       (N138)? mem[1556] : 
                       (N77)? mem[1606] : 
                       (N79)? mem[1656] : 
                       (N81)? mem[1706] : 
                       (N83)? mem[1756] : 
                       (N85)? mem[1806] : 
                       (N87)? mem[1856] : 
                       (N89)? mem[1906] : 
                       (N91)? mem[1956] : 
                       (N93)? mem[2006] : 
                       (N95)? mem[2056] : 
                       (N97)? mem[2106] : 
                       (N99)? mem[2156] : 
                       (N101)? mem[2206] : 
                       (N103)? mem[2256] : 
                       (N105)? mem[2306] : 
                       (N107)? mem[2356] : 
                       (N109)? mem[2406] : 
                       (N111)? mem[2456] : 
                       (N113)? mem[2506] : 
                       (N115)? mem[2556] : 
                       (N117)? mem[2606] : 
                       (N119)? mem[2656] : 
                       (N121)? mem[2706] : 
                       (N123)? mem[2756] : 
                       (N125)? mem[2806] : 
                       (N127)? mem[2856] : 
                       (N129)? mem[2906] : 
                       (N131)? mem[2956] : 
                       (N133)? mem[3006] : 
                       (N135)? mem[3056] : 
                       (N137)? mem[3106] : 
                       (N139)? mem[3156] : 1'b0;
  assign r_data_o[5] = (N76)? mem[5] : 
                       (N78)? mem[55] : 
                       (N80)? mem[105] : 
                       (N82)? mem[155] : 
                       (N84)? mem[205] : 
                       (N86)? mem[255] : 
                       (N88)? mem[305] : 
                       (N90)? mem[355] : 
                       (N92)? mem[405] : 
                       (N94)? mem[455] : 
                       (N96)? mem[505] : 
                       (N98)? mem[555] : 
                       (N100)? mem[605] : 
                       (N102)? mem[655] : 
                       (N104)? mem[705] : 
                       (N106)? mem[755] : 
                       (N108)? mem[805] : 
                       (N110)? mem[855] : 
                       (N112)? mem[905] : 
                       (N114)? mem[955] : 
                       (N116)? mem[1005] : 
                       (N118)? mem[1055] : 
                       (N120)? mem[1105] : 
                       (N122)? mem[1155] : 
                       (N124)? mem[1205] : 
                       (N126)? mem[1255] : 
                       (N128)? mem[1305] : 
                       (N130)? mem[1355] : 
                       (N132)? mem[1405] : 
                       (N134)? mem[1455] : 
                       (N136)? mem[1505] : 
                       (N138)? mem[1555] : 
                       (N77)? mem[1605] : 
                       (N79)? mem[1655] : 
                       (N81)? mem[1705] : 
                       (N83)? mem[1755] : 
                       (N85)? mem[1805] : 
                       (N87)? mem[1855] : 
                       (N89)? mem[1905] : 
                       (N91)? mem[1955] : 
                       (N93)? mem[2005] : 
                       (N95)? mem[2055] : 
                       (N97)? mem[2105] : 
                       (N99)? mem[2155] : 
                       (N101)? mem[2205] : 
                       (N103)? mem[2255] : 
                       (N105)? mem[2305] : 
                       (N107)? mem[2355] : 
                       (N109)? mem[2405] : 
                       (N111)? mem[2455] : 
                       (N113)? mem[2505] : 
                       (N115)? mem[2555] : 
                       (N117)? mem[2605] : 
                       (N119)? mem[2655] : 
                       (N121)? mem[2705] : 
                       (N123)? mem[2755] : 
                       (N125)? mem[2805] : 
                       (N127)? mem[2855] : 
                       (N129)? mem[2905] : 
                       (N131)? mem[2955] : 
                       (N133)? mem[3005] : 
                       (N135)? mem[3055] : 
                       (N137)? mem[3105] : 
                       (N139)? mem[3155] : 1'b0;
  assign r_data_o[4] = (N76)? mem[4] : 
                       (N78)? mem[54] : 
                       (N80)? mem[104] : 
                       (N82)? mem[154] : 
                       (N84)? mem[204] : 
                       (N86)? mem[254] : 
                       (N88)? mem[304] : 
                       (N90)? mem[354] : 
                       (N92)? mem[404] : 
                       (N94)? mem[454] : 
                       (N96)? mem[504] : 
                       (N98)? mem[554] : 
                       (N100)? mem[604] : 
                       (N102)? mem[654] : 
                       (N104)? mem[704] : 
                       (N106)? mem[754] : 
                       (N108)? mem[804] : 
                       (N110)? mem[854] : 
                       (N112)? mem[904] : 
                       (N114)? mem[954] : 
                       (N116)? mem[1004] : 
                       (N118)? mem[1054] : 
                       (N120)? mem[1104] : 
                       (N122)? mem[1154] : 
                       (N124)? mem[1204] : 
                       (N126)? mem[1254] : 
                       (N128)? mem[1304] : 
                       (N130)? mem[1354] : 
                       (N132)? mem[1404] : 
                       (N134)? mem[1454] : 
                       (N136)? mem[1504] : 
                       (N138)? mem[1554] : 
                       (N77)? mem[1604] : 
                       (N79)? mem[1654] : 
                       (N81)? mem[1704] : 
                       (N83)? mem[1754] : 
                       (N85)? mem[1804] : 
                       (N87)? mem[1854] : 
                       (N89)? mem[1904] : 
                       (N91)? mem[1954] : 
                       (N93)? mem[2004] : 
                       (N95)? mem[2054] : 
                       (N97)? mem[2104] : 
                       (N99)? mem[2154] : 
                       (N101)? mem[2204] : 
                       (N103)? mem[2254] : 
                       (N105)? mem[2304] : 
                       (N107)? mem[2354] : 
                       (N109)? mem[2404] : 
                       (N111)? mem[2454] : 
                       (N113)? mem[2504] : 
                       (N115)? mem[2554] : 
                       (N117)? mem[2604] : 
                       (N119)? mem[2654] : 
                       (N121)? mem[2704] : 
                       (N123)? mem[2754] : 
                       (N125)? mem[2804] : 
                       (N127)? mem[2854] : 
                       (N129)? mem[2904] : 
                       (N131)? mem[2954] : 
                       (N133)? mem[3004] : 
                       (N135)? mem[3054] : 
                       (N137)? mem[3104] : 
                       (N139)? mem[3154] : 1'b0;
  assign r_data_o[3] = (N76)? mem[3] : 
                       (N78)? mem[53] : 
                       (N80)? mem[103] : 
                       (N82)? mem[153] : 
                       (N84)? mem[203] : 
                       (N86)? mem[253] : 
                       (N88)? mem[303] : 
                       (N90)? mem[353] : 
                       (N92)? mem[403] : 
                       (N94)? mem[453] : 
                       (N96)? mem[503] : 
                       (N98)? mem[553] : 
                       (N100)? mem[603] : 
                       (N102)? mem[653] : 
                       (N104)? mem[703] : 
                       (N106)? mem[753] : 
                       (N108)? mem[803] : 
                       (N110)? mem[853] : 
                       (N112)? mem[903] : 
                       (N114)? mem[953] : 
                       (N116)? mem[1003] : 
                       (N118)? mem[1053] : 
                       (N120)? mem[1103] : 
                       (N122)? mem[1153] : 
                       (N124)? mem[1203] : 
                       (N126)? mem[1253] : 
                       (N128)? mem[1303] : 
                       (N130)? mem[1353] : 
                       (N132)? mem[1403] : 
                       (N134)? mem[1453] : 
                       (N136)? mem[1503] : 
                       (N138)? mem[1553] : 
                       (N77)? mem[1603] : 
                       (N79)? mem[1653] : 
                       (N81)? mem[1703] : 
                       (N83)? mem[1753] : 
                       (N85)? mem[1803] : 
                       (N87)? mem[1853] : 
                       (N89)? mem[1903] : 
                       (N91)? mem[1953] : 
                       (N93)? mem[2003] : 
                       (N95)? mem[2053] : 
                       (N97)? mem[2103] : 
                       (N99)? mem[2153] : 
                       (N101)? mem[2203] : 
                       (N103)? mem[2253] : 
                       (N105)? mem[2303] : 
                       (N107)? mem[2353] : 
                       (N109)? mem[2403] : 
                       (N111)? mem[2453] : 
                       (N113)? mem[2503] : 
                       (N115)? mem[2553] : 
                       (N117)? mem[2603] : 
                       (N119)? mem[2653] : 
                       (N121)? mem[2703] : 
                       (N123)? mem[2753] : 
                       (N125)? mem[2803] : 
                       (N127)? mem[2853] : 
                       (N129)? mem[2903] : 
                       (N131)? mem[2953] : 
                       (N133)? mem[3003] : 
                       (N135)? mem[3053] : 
                       (N137)? mem[3103] : 
                       (N139)? mem[3153] : 1'b0;
  assign r_data_o[2] = (N76)? mem[2] : 
                       (N78)? mem[52] : 
                       (N80)? mem[102] : 
                       (N82)? mem[152] : 
                       (N84)? mem[202] : 
                       (N86)? mem[252] : 
                       (N88)? mem[302] : 
                       (N90)? mem[352] : 
                       (N92)? mem[402] : 
                       (N94)? mem[452] : 
                       (N96)? mem[502] : 
                       (N98)? mem[552] : 
                       (N100)? mem[602] : 
                       (N102)? mem[652] : 
                       (N104)? mem[702] : 
                       (N106)? mem[752] : 
                       (N108)? mem[802] : 
                       (N110)? mem[852] : 
                       (N112)? mem[902] : 
                       (N114)? mem[952] : 
                       (N116)? mem[1002] : 
                       (N118)? mem[1052] : 
                       (N120)? mem[1102] : 
                       (N122)? mem[1152] : 
                       (N124)? mem[1202] : 
                       (N126)? mem[1252] : 
                       (N128)? mem[1302] : 
                       (N130)? mem[1352] : 
                       (N132)? mem[1402] : 
                       (N134)? mem[1452] : 
                       (N136)? mem[1502] : 
                       (N138)? mem[1552] : 
                       (N77)? mem[1602] : 
                       (N79)? mem[1652] : 
                       (N81)? mem[1702] : 
                       (N83)? mem[1752] : 
                       (N85)? mem[1802] : 
                       (N87)? mem[1852] : 
                       (N89)? mem[1902] : 
                       (N91)? mem[1952] : 
                       (N93)? mem[2002] : 
                       (N95)? mem[2052] : 
                       (N97)? mem[2102] : 
                       (N99)? mem[2152] : 
                       (N101)? mem[2202] : 
                       (N103)? mem[2252] : 
                       (N105)? mem[2302] : 
                       (N107)? mem[2352] : 
                       (N109)? mem[2402] : 
                       (N111)? mem[2452] : 
                       (N113)? mem[2502] : 
                       (N115)? mem[2552] : 
                       (N117)? mem[2602] : 
                       (N119)? mem[2652] : 
                       (N121)? mem[2702] : 
                       (N123)? mem[2752] : 
                       (N125)? mem[2802] : 
                       (N127)? mem[2852] : 
                       (N129)? mem[2902] : 
                       (N131)? mem[2952] : 
                       (N133)? mem[3002] : 
                       (N135)? mem[3052] : 
                       (N137)? mem[3102] : 
                       (N139)? mem[3152] : 1'b0;
  assign r_data_o[1] = (N76)? mem[1] : 
                       (N78)? mem[51] : 
                       (N80)? mem[101] : 
                       (N82)? mem[151] : 
                       (N84)? mem[201] : 
                       (N86)? mem[251] : 
                       (N88)? mem[301] : 
                       (N90)? mem[351] : 
                       (N92)? mem[401] : 
                       (N94)? mem[451] : 
                       (N96)? mem[501] : 
                       (N98)? mem[551] : 
                       (N100)? mem[601] : 
                       (N102)? mem[651] : 
                       (N104)? mem[701] : 
                       (N106)? mem[751] : 
                       (N108)? mem[801] : 
                       (N110)? mem[851] : 
                       (N112)? mem[901] : 
                       (N114)? mem[951] : 
                       (N116)? mem[1001] : 
                       (N118)? mem[1051] : 
                       (N120)? mem[1101] : 
                       (N122)? mem[1151] : 
                       (N124)? mem[1201] : 
                       (N126)? mem[1251] : 
                       (N128)? mem[1301] : 
                       (N130)? mem[1351] : 
                       (N132)? mem[1401] : 
                       (N134)? mem[1451] : 
                       (N136)? mem[1501] : 
                       (N138)? mem[1551] : 
                       (N77)? mem[1601] : 
                       (N79)? mem[1651] : 
                       (N81)? mem[1701] : 
                       (N83)? mem[1751] : 
                       (N85)? mem[1801] : 
                       (N87)? mem[1851] : 
                       (N89)? mem[1901] : 
                       (N91)? mem[1951] : 
                       (N93)? mem[2001] : 
                       (N95)? mem[2051] : 
                       (N97)? mem[2101] : 
                       (N99)? mem[2151] : 
                       (N101)? mem[2201] : 
                       (N103)? mem[2251] : 
                       (N105)? mem[2301] : 
                       (N107)? mem[2351] : 
                       (N109)? mem[2401] : 
                       (N111)? mem[2451] : 
                       (N113)? mem[2501] : 
                       (N115)? mem[2551] : 
                       (N117)? mem[2601] : 
                       (N119)? mem[2651] : 
                       (N121)? mem[2701] : 
                       (N123)? mem[2751] : 
                       (N125)? mem[2801] : 
                       (N127)? mem[2851] : 
                       (N129)? mem[2901] : 
                       (N131)? mem[2951] : 
                       (N133)? mem[3001] : 
                       (N135)? mem[3051] : 
                       (N137)? mem[3101] : 
                       (N139)? mem[3151] : 1'b0;
  assign r_data_o[0] = (N76)? mem[0] : 
                       (N78)? mem[50] : 
                       (N80)? mem[100] : 
                       (N82)? mem[150] : 
                       (N84)? mem[200] : 
                       (N86)? mem[250] : 
                       (N88)? mem[300] : 
                       (N90)? mem[350] : 
                       (N92)? mem[400] : 
                       (N94)? mem[450] : 
                       (N96)? mem[500] : 
                       (N98)? mem[550] : 
                       (N100)? mem[600] : 
                       (N102)? mem[650] : 
                       (N104)? mem[700] : 
                       (N106)? mem[750] : 
                       (N108)? mem[800] : 
                       (N110)? mem[850] : 
                       (N112)? mem[900] : 
                       (N114)? mem[950] : 
                       (N116)? mem[1000] : 
                       (N118)? mem[1050] : 
                       (N120)? mem[1100] : 
                       (N122)? mem[1150] : 
                       (N124)? mem[1200] : 
                       (N126)? mem[1250] : 
                       (N128)? mem[1300] : 
                       (N130)? mem[1350] : 
                       (N132)? mem[1400] : 
                       (N134)? mem[1450] : 
                       (N136)? mem[1500] : 
                       (N138)? mem[1550] : 
                       (N77)? mem[1600] : 
                       (N79)? mem[1650] : 
                       (N81)? mem[1700] : 
                       (N83)? mem[1750] : 
                       (N85)? mem[1800] : 
                       (N87)? mem[1850] : 
                       (N89)? mem[1900] : 
                       (N91)? mem[1950] : 
                       (N93)? mem[2000] : 
                       (N95)? mem[2050] : 
                       (N97)? mem[2100] : 
                       (N99)? mem[2150] : 
                       (N101)? mem[2200] : 
                       (N103)? mem[2250] : 
                       (N105)? mem[2300] : 
                       (N107)? mem[2350] : 
                       (N109)? mem[2400] : 
                       (N111)? mem[2450] : 
                       (N113)? mem[2500] : 
                       (N115)? mem[2550] : 
                       (N117)? mem[2600] : 
                       (N119)? mem[2650] : 
                       (N121)? mem[2700] : 
                       (N123)? mem[2750] : 
                       (N125)? mem[2800] : 
                       (N127)? mem[2850] : 
                       (N129)? mem[2900] : 
                       (N131)? mem[2950] : 
                       (N133)? mem[3000] : 
                       (N135)? mem[3050] : 
                       (N137)? mem[3100] : 
                       (N139)? mem[3150] : 1'b0;
  assign N269 = ~w_addr_i[5];
  assign N270 = w_addr_i[3] & w_addr_i[4];
  assign N271 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N272 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N273 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N274 = w_addr_i[5] & N270;
  assign N275 = w_addr_i[5] & N271;
  assign N276 = w_addr_i[5] & N272;
  assign N277 = w_addr_i[5] & N273;
  assign N278 = N269 & N270;
  assign N279 = N269 & N271;
  assign N280 = N269 & N272;
  assign N281 = N269 & N273;
  assign N282 = ~w_addr_i[2];
  assign N283 = w_addr_i[0] & w_addr_i[1];
  assign N284 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N285 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N286 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N287 = w_addr_i[2] & N283;
  assign N288 = w_addr_i[2] & N284;
  assign N289 = w_addr_i[2] & N285;
  assign N290 = w_addr_i[2] & N286;
  assign N291 = N282 & N283;
  assign N292 = N282 & N284;
  assign N293 = N282 & N285;
  assign N294 = N282 & N286;
  assign N204 = N274 & N287;
  assign N203 = N274 & N288;
  assign N202 = N274 & N289;
  assign N201 = N274 & N290;
  assign N200 = N274 & N291;
  assign N199 = N274 & N292;
  assign N198 = N274 & N293;
  assign N197 = N274 & N294;
  assign N196 = N275 & N287;
  assign N195 = N275 & N288;
  assign N194 = N275 & N289;
  assign N193 = N275 & N290;
  assign N192 = N275 & N291;
  assign N191 = N275 & N292;
  assign N190 = N275 & N293;
  assign N189 = N275 & N294;
  assign N188 = N276 & N287;
  assign N187 = N276 & N288;
  assign N186 = N276 & N289;
  assign N185 = N276 & N290;
  assign N184 = N276 & N291;
  assign N183 = N276 & N292;
  assign N182 = N276 & N293;
  assign N181 = N276 & N294;
  assign N180 = N277 & N287;
  assign N179 = N277 & N288;
  assign N178 = N277 & N289;
  assign N177 = N277 & N290;
  assign N176 = N277 & N291;
  assign N175 = N277 & N292;
  assign N174 = N277 & N293;
  assign N173 = N277 & N294;
  assign N172 = N278 & N287;
  assign N171 = N278 & N288;
  assign N170 = N278 & N289;
  assign N169 = N278 & N290;
  assign N168 = N278 & N291;
  assign N167 = N278 & N292;
  assign N166 = N278 & N293;
  assign N165 = N278 & N294;
  assign N164 = N279 & N287;
  assign N163 = N279 & N288;
  assign N162 = N279 & N289;
  assign N161 = N279 & N290;
  assign N160 = N279 & N291;
  assign N159 = N279 & N292;
  assign N158 = N279 & N293;
  assign N157 = N279 & N294;
  assign N156 = N280 & N287;
  assign N155 = N280 & N288;
  assign N154 = N280 & N289;
  assign N153 = N280 & N290;
  assign N152 = N280 & N291;
  assign N151 = N280 & N292;
  assign N150 = N280 & N293;
  assign N149 = N280 & N294;
  assign N148 = N281 & N287;
  assign N147 = N281 & N288;
  assign N146 = N281 & N289;
  assign N145 = N281 & N290;
  assign N144 = N281 & N291;
  assign N143 = N281 & N292;
  assign N142 = N281 & N293;
  assign N141 = N281 & N294;
  assign { N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205 } = (N8)? { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~r_addr_i[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r_addr_i[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r_addr_i[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r_addr_i[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r_addr_i[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r_addr_i[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r_addr_i[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r_addr_i[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r_addr_i[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r_addr_i[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r_addr_i[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r_addr_i[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r_addr_i[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r_addr_i[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r_addr_i[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r_addr_i[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r_addr_i[4];
  assign N75 = ~r_addr_i[5];
  assign N76 = N43 & N75;
  assign N77 = N43 & r_addr_i[5];
  assign N78 = N45 & N75;
  assign N79 = N45 & r_addr_i[5];
  assign N80 = N47 & N75;
  assign N81 = N47 & r_addr_i[5];
  assign N82 = N49 & N75;
  assign N83 = N49 & r_addr_i[5];
  assign N84 = N51 & N75;
  assign N85 = N51 & r_addr_i[5];
  assign N86 = N53 & N75;
  assign N87 = N53 & r_addr_i[5];
  assign N88 = N55 & N75;
  assign N89 = N55 & r_addr_i[5];
  assign N90 = N57 & N75;
  assign N91 = N57 & r_addr_i[5];
  assign N92 = N59 & N75;
  assign N93 = N59 & r_addr_i[5];
  assign N94 = N61 & N75;
  assign N95 = N61 & r_addr_i[5];
  assign N96 = N63 & N75;
  assign N97 = N63 & r_addr_i[5];
  assign N98 = N65 & N75;
  assign N99 = N65 & r_addr_i[5];
  assign N100 = N67 & N75;
  assign N101 = N67 & r_addr_i[5];
  assign N102 = N69 & N75;
  assign N103 = N69 & r_addr_i[5];
  assign N104 = N71 & N75;
  assign N105 = N71 & r_addr_i[5];
  assign N106 = N73 & N75;
  assign N107 = N73 & r_addr_i[5];
  assign N108 = N44 & N75;
  assign N109 = N44 & r_addr_i[5];
  assign N110 = N46 & N75;
  assign N111 = N46 & r_addr_i[5];
  assign N112 = N48 & N75;
  assign N113 = N48 & r_addr_i[5];
  assign N114 = N50 & N75;
  assign N115 = N50 & r_addr_i[5];
  assign N116 = N52 & N75;
  assign N117 = N52 & r_addr_i[5];
  assign N118 = N54 & N75;
  assign N119 = N54 & r_addr_i[5];
  assign N120 = N56 & N75;
  assign N121 = N56 & r_addr_i[5];
  assign N122 = N58 & N75;
  assign N123 = N58 & r_addr_i[5];
  assign N124 = N60 & N75;
  assign N125 = N60 & r_addr_i[5];
  assign N126 = N62 & N75;
  assign N127 = N62 & r_addr_i[5];
  assign N128 = N64 & N75;
  assign N129 = N64 & r_addr_i[5];
  assign N130 = N66 & N75;
  assign N131 = N66 & r_addr_i[5];
  assign N132 = N68 & N75;
  assign N133 = N68 & r_addr_i[5];
  assign N134 = N70 & N75;
  assign N135 = N70 & r_addr_i[5];
  assign N136 = N72 & N75;
  assign N137 = N72 & r_addr_i[5];
  assign N138 = N74 & N75;
  assign N139 = N74 & r_addr_i[5];
  assign N140 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N268) begin
      { mem[3199:3150] } <= { w_data_i[49:0] };
    end 
    if(N267) begin
      { mem[3149:3100] } <= { w_data_i[49:0] };
    end 
    if(N266) begin
      { mem[3099:3050] } <= { w_data_i[49:0] };
    end 
    if(N265) begin
      { mem[3049:3000] } <= { w_data_i[49:0] };
    end 
    if(N264) begin
      { mem[2999:2950] } <= { w_data_i[49:0] };
    end 
    if(N263) begin
      { mem[2949:2900] } <= { w_data_i[49:0] };
    end 
    if(N262) begin
      { mem[2899:2850] } <= { w_data_i[49:0] };
    end 
    if(N261) begin
      { mem[2849:2800] } <= { w_data_i[49:0] };
    end 
    if(N260) begin
      { mem[2799:2750] } <= { w_data_i[49:0] };
    end 
    if(N259) begin
      { mem[2749:2700] } <= { w_data_i[49:0] };
    end 
    if(N258) begin
      { mem[2699:2650] } <= { w_data_i[49:0] };
    end 
    if(N257) begin
      { mem[2649:2600] } <= { w_data_i[49:0] };
    end 
    if(N256) begin
      { mem[2599:2550] } <= { w_data_i[49:0] };
    end 
    if(N255) begin
      { mem[2549:2500] } <= { w_data_i[49:0] };
    end 
    if(N254) begin
      { mem[2499:2450] } <= { w_data_i[49:0] };
    end 
    if(N253) begin
      { mem[2449:2400] } <= { w_data_i[49:0] };
    end 
    if(N252) begin
      { mem[2399:2350] } <= { w_data_i[49:0] };
    end 
    if(N251) begin
      { mem[2349:2300] } <= { w_data_i[49:0] };
    end 
    if(N250) begin
      { mem[2299:2250] } <= { w_data_i[49:0] };
    end 
    if(N249) begin
      { mem[2249:2200] } <= { w_data_i[49:0] };
    end 
    if(N248) begin
      { mem[2199:2150] } <= { w_data_i[49:0] };
    end 
    if(N247) begin
      { mem[2149:2100] } <= { w_data_i[49:0] };
    end 
    if(N246) begin
      { mem[2099:2050] } <= { w_data_i[49:0] };
    end 
    if(N245) begin
      { mem[2049:2000] } <= { w_data_i[49:0] };
    end 
    if(N244) begin
      { mem[1999:1950] } <= { w_data_i[49:0] };
    end 
    if(N243) begin
      { mem[1949:1900] } <= { w_data_i[49:0] };
    end 
    if(N242) begin
      { mem[1899:1850] } <= { w_data_i[49:0] };
    end 
    if(N241) begin
      { mem[1849:1800] } <= { w_data_i[49:0] };
    end 
    if(N240) begin
      { mem[1799:1750] } <= { w_data_i[49:0] };
    end 
    if(N239) begin
      { mem[1749:1700] } <= { w_data_i[49:0] };
    end 
    if(N238) begin
      { mem[1699:1650] } <= { w_data_i[49:0] };
    end 
    if(N237) begin
      { mem[1649:1600] } <= { w_data_i[49:0] };
    end 
    if(N236) begin
      { mem[1599:1550] } <= { w_data_i[49:0] };
    end 
    if(N235) begin
      { mem[1549:1500] } <= { w_data_i[49:0] };
    end 
    if(N234) begin
      { mem[1499:1450] } <= { w_data_i[49:0] };
    end 
    if(N233) begin
      { mem[1449:1400] } <= { w_data_i[49:0] };
    end 
    if(N232) begin
      { mem[1399:1350] } <= { w_data_i[49:0] };
    end 
    if(N231) begin
      { mem[1349:1300] } <= { w_data_i[49:0] };
    end 
    if(N230) begin
      { mem[1299:1250] } <= { w_data_i[49:0] };
    end 
    if(N229) begin
      { mem[1249:1200] } <= { w_data_i[49:0] };
    end 
    if(N228) begin
      { mem[1199:1150] } <= { w_data_i[49:0] };
    end 
    if(N227) begin
      { mem[1149:1100] } <= { w_data_i[49:0] };
    end 
    if(N226) begin
      { mem[1099:1050] } <= { w_data_i[49:0] };
    end 
    if(N225) begin
      { mem[1049:1000] } <= { w_data_i[49:0] };
    end 
    if(N224) begin
      { mem[999:950] } <= { w_data_i[49:0] };
    end 
    if(N223) begin
      { mem[949:900] } <= { w_data_i[49:0] };
    end 
    if(N222) begin
      { mem[899:850] } <= { w_data_i[49:0] };
    end 
    if(N221) begin
      { mem[849:800] } <= { w_data_i[49:0] };
    end 
    if(N220) begin
      { mem[799:750] } <= { w_data_i[49:0] };
    end 
    if(N219) begin
      { mem[749:700] } <= { w_data_i[49:0] };
    end 
    if(N218) begin
      { mem[699:650] } <= { w_data_i[49:0] };
    end 
    if(N217) begin
      { mem[649:600] } <= { w_data_i[49:0] };
    end 
    if(N216) begin
      { mem[599:550] } <= { w_data_i[49:0] };
    end 
    if(N215) begin
      { mem[549:500] } <= { w_data_i[49:0] };
    end 
    if(N214) begin
      { mem[499:450] } <= { w_data_i[49:0] };
    end 
    if(N213) begin
      { mem[449:400] } <= { w_data_i[49:0] };
    end 
    if(N212) begin
      { mem[399:350] } <= { w_data_i[49:0] };
    end 
    if(N211) begin
      { mem[349:300] } <= { w_data_i[49:0] };
    end 
    if(N210) begin
      { mem[299:250] } <= { w_data_i[49:0] };
    end 
    if(N209) begin
      { mem[249:200] } <= { w_data_i[49:0] };
    end 
    if(N208) begin
      { mem[199:150] } <= { w_data_i[49:0] };
    end 
    if(N207) begin
      { mem[149:100] } <= { w_data_i[49:0] };
    end 
    if(N206) begin
      { mem[99:50] } <= { w_data_i[49:0] };
    end 
    if(N205) begin
      { mem[49:0] } <= { w_data_i[49:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p50_els_p64_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [49:0] w_data_i;
  input [5:0] r_addr_i;
  output [49:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [49:0] r_data_o;

  bsg_mem_1r1w_synth_width_p50_els_p64_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_launch_sync_sync_posedge_7_unit
(
  iclk_i,
  iclk_reset_i,
  oclk_i,
  iclk_data_i,
  iclk_data_o,
  oclk_data_o
);

  input [6:0] iclk_data_i;
  output [6:0] iclk_data_o;
  output [6:0] oclk_data_o;
  input iclk_i;
  input iclk_reset_i;
  input oclk_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  reg [6:0] iclk_data_o,bsg_SYNC_1_r,oclk_data_o;
  assign { N9, N8, N7, N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N1)? iclk_data_i : 1'b0;
  assign N0 = iclk_reset_i;
  assign N1 = N2;
  assign N2 = ~iclk_reset_i;

  always @(posedge iclk_i) begin
    if(1'b1) begin
      { iclk_data_o[6:0] } <= { N9, N8, N7, N6, N5, N4, N3 };
    end 
  end


  always @(posedge oclk_i) begin
    if(1'b1) begin
      { bsg_SYNC_1_r[6:0] } <= { iclk_data_o[6:0] };
      { oclk_data_o[6:0] } <= { bsg_SYNC_1_r[6:0] };
    end 
  end


endmodule



module bsg_launch_sync_sync_width_p7_use_negedge_for_launch_p0_use_async_reset_p0
(
  iclk_i,
  iclk_reset_i,
  oclk_i,
  iclk_data_i,
  iclk_data_o,
  oclk_data_o
);

  input [6:0] iclk_data_i;
  output [6:0] iclk_data_o;
  output [6:0] oclk_data_o;
  input iclk_i;
  input iclk_reset_i;
  input oclk_i;
  wire [6:0] iclk_data_o,oclk_data_o;

  bsg_launch_sync_sync_posedge_7_unit
  sync_p_z_blss
  (
    .iclk_i(iclk_i),
    .iclk_reset_i(iclk_reset_i),
    .oclk_i(oclk_i),
    .iclk_data_i(iclk_data_i),
    .iclk_data_o(iclk_data_o),
    .oclk_data_o(oclk_data_o)
  );


endmodule



module bsg_async_ptr_gray_lg_size_p7
(
  w_clk_i,
  w_reset_i,
  w_inc_i,
  r_clk_i,
  w_ptr_binary_r_o,
  w_ptr_gray_r_o,
  w_ptr_gray_r_rsync_o
);

  output [6:0] w_ptr_binary_r_o;
  output [6:0] w_ptr_gray_r_o;
  output [6:0] w_ptr_gray_r_rsync_o;
  input w_clk_i;
  input w_reset_i;
  input w_inc_i;
  input r_clk_i;
  wire [6:0] w_ptr_gray_r_o,w_ptr_gray_r_rsync_o,w_ptr_p2,w_ptr_gray_n;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  reg [6:0] w_ptr_p1_r,w_ptr_binary_r_o;

  bsg_launch_sync_sync_width_p7_use_negedge_for_launch_p0_use_async_reset_p0
  ptr_sync
  (
    .iclk_i(w_clk_i),
    .iclk_reset_i(w_reset_i),
    .oclk_i(r_clk_i),
    .iclk_data_i(w_ptr_gray_n),
    .iclk_data_o(w_ptr_gray_r_o),
    .oclk_data_o(w_ptr_gray_r_rsync_o)
  );

  assign w_ptr_p2 = w_ptr_p1_r + 1'b1;
  assign w_ptr_gray_n = (N0)? { w_ptr_p1_r[6:6], N3, N4, N5, N6, N7, N8 } : 
                        (N1)? w_ptr_gray_r_o : 1'b0;
  assign N0 = w_inc_i;
  assign N1 = N2;
  assign N2 = ~w_inc_i;
  assign N3 = w_ptr_p1_r[6] ^ w_ptr_p1_r[5];
  assign N4 = w_ptr_p1_r[5] ^ w_ptr_p1_r[4];
  assign N5 = w_ptr_p1_r[4] ^ w_ptr_p1_r[3];
  assign N6 = w_ptr_p1_r[3] ^ w_ptr_p1_r[2];
  assign N7 = w_ptr_p1_r[2] ^ w_ptr_p1_r[1];
  assign N8 = w_ptr_p1_r[1] ^ w_ptr_p1_r[0];

  always @(posedge w_clk_i) begin
    if(w_reset_i) begin
      { w_ptr_p1_r[6:0] } <= { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 };
      { w_ptr_binary_r_o[6:0] } <= { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
    end else if(w_inc_i) begin
      { w_ptr_p1_r[6:0] } <= { w_ptr_p2[6:0] };
      { w_ptr_binary_r_o[6:0] } <= { w_ptr_p1_r[6:0] };
    end 
  end


endmodule



module bsg_async_fifo_lg_size_p6_width_p50
(
  w_clk_i,
  w_reset_i,
  w_enq_i,
  w_data_i,
  w_full_o,
  r_clk_i,
  r_reset_i,
  r_deq_i,
  r_data_o,
  r_valid_o
);

  input [49:0] w_data_i;
  output [49:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_enq_i;
  input r_clk_i;
  input r_reset_i;
  input r_deq_i;
  output w_full_o;
  output r_valid_o;
  wire [49:0] r_data_o;
  wire w_full_o,r_valid_o,N0,N1;
  wire [6:0] w_ptr_binary_r,r_ptr_binary_r,w_ptr_gray_r,w_ptr_gray_r_rsync,r_ptr_gray_r,
  r_ptr_gray_r_wsync;

  bsg_mem_1r1w_width_p50_els_p64_read_write_same_addr_p0
  MSYNC_1r1w
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_enq_i),
    .w_addr_i(w_ptr_binary_r[5:0]),
    .w_data_i(w_data_i),
    .r_v_i(r_valid_o),
    .r_addr_i(r_ptr_binary_r[5:0]),
    .r_data_o(r_data_o)
  );


  bsg_async_ptr_gray_lg_size_p7
  bapg_wr
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_inc_i(w_enq_i),
    .r_clk_i(r_clk_i),
    .w_ptr_binary_r_o(w_ptr_binary_r),
    .w_ptr_gray_r_o(w_ptr_gray_r),
    .w_ptr_gray_r_rsync_o(w_ptr_gray_r_rsync)
  );


  bsg_async_ptr_gray_lg_size_p7
  bapg_rd
  (
    .w_clk_i(r_clk_i),
    .w_reset_i(r_reset_i),
    .w_inc_i(r_deq_i),
    .r_clk_i(w_clk_i),
    .w_ptr_binary_r_o(r_ptr_binary_r),
    .w_ptr_gray_r_o(r_ptr_gray_r),
    .w_ptr_gray_r_rsync_o(r_ptr_gray_r_wsync)
  );

  assign r_valid_o = r_ptr_gray_r != w_ptr_gray_r_rsync;
  assign w_full_o = w_ptr_gray_r == { N0, N1, r_ptr_gray_r_wsync[4:0] };
  assign N0 = ~r_ptr_gray_r_wsync[6];
  assign N1 = ~r_ptr_gray_r_wsync[5];

endmodule



module bsg_sync_sync_1_unit
(
  oclk_i,
  iclk_data_i,
  oclk_data_o
);

  input [0:0] iclk_data_i;
  output [0:0] oclk_data_o;
  input oclk_i;
  reg [0:0] bsg_SYNC_1_r,oclk_data_o;

  always @(posedge oclk_i) begin
    if(1'b1) begin
      { bsg_SYNC_1_r[0:0] } <= { iclk_data_i[0:0] };
      { oclk_data_o[0:0] } <= { bsg_SYNC_1_r[0:0] };
    end 
  end


endmodule



module bsg_sync_sync_width_p1
(
  oclk_i,
  iclk_data_i,
  oclk_data_o
);

  input [0:0] iclk_data_i;
  output [0:0] oclk_data_o;
  input oclk_i;
  wire [0:0] oclk_data_o;

  bsg_sync_sync_1_unit
  z_bss
  (
    .oclk_i(oclk_i),
    .iclk_data_i(iclk_data_i[0]),
    .oclk_data_o(oclk_data_o[0])
  );


endmodule



module bsg_fsb_node_async_buffer
(
  L_clk_i,
  L_reset_i,
  L_en_o,
  L_v_o,
  L_data_o,
  L_ready_i,
  L_v_i,
  L_data_i,
  L_yumi_o,
  R_clk_i,
  R_reset_i,
  R_en_i,
  R_v_i,
  R_data_i,
  R_ready_o,
  R_v_o,
  R_data_o,
  R_yumi_i
);

  output [49:0] L_data_o;
  input [49:0] L_data_i;
  input [49:0] R_data_i;
  output [49:0] R_data_o;
  input L_clk_i;
  input L_reset_i;
  input L_ready_i;
  input L_v_i;
  input R_clk_i;
  input R_reset_i;
  input R_en_i;
  input R_v_i;
  input R_yumi_i;
  output L_en_o;
  output L_v_o;
  output L_yumi_o;
  output R_ready_o;
  output R_v_o;
  wire [49:0] L_data_o,R_data_o;
  wire L_en_o,L_v_o,L_yumi_o,R_ready_o,R_v_o,R_w_full_lo,n_0_net_,n_1_net_,L_w_full_lo,
  N0,N1;

  bsg_async_fifo_lg_size_p6_width_p50
  r2l_fifo
  (
    .w_clk_i(R_clk_i),
    .w_reset_i(R_reset_i),
    .w_enq_i(n_0_net_),
    .w_data_i(R_data_i),
    .w_full_o(R_w_full_lo),
    .r_clk_i(L_clk_i),
    .r_reset_i(L_reset_i),
    .r_deq_i(n_1_net_),
    .r_data_o(L_data_o),
    .r_valid_o(L_v_o)
  );


  bsg_async_fifo_lg_size_p6_width_p50
  l2r_fifo
  (
    .w_clk_i(L_clk_i),
    .w_reset_i(L_reset_i),
    .w_enq_i(L_yumi_o),
    .w_data_i(L_data_i),
    .w_full_o(L_w_full_lo),
    .r_clk_i(R_clk_i),
    .r_reset_i(R_reset_i),
    .r_deq_i(R_yumi_i),
    .r_data_o(R_data_o),
    .r_valid_o(R_v_o)
  );


  bsg_sync_sync_width_p1
  fsb_en_sync
  (
    .oclk_i(L_clk_i),
    .iclk_data_i(R_en_i),
    .oclk_data_o(L_en_o)
  );

  assign R_ready_o = ~R_w_full_lo;
  assign n_1_net_ = L_v_o & L_ready_i;
  assign n_0_net_ = N0 & R_v_i;
  assign N0 = ~R_w_full_lo;
  assign L_yumi_o = N1 & L_v_i;
  assign N1 = ~L_w_full_lo;

endmodule

