

module top
(
  i,
  shamt_i,
  sticky_o
);

  input [63:0] i;
  input [6:0] shamt_i;
  output sticky_o;

  bsg_fpu_sticky
  wrapper
  (
    .i(i),
    .shamt_i(shamt_i),
    .sticky_o(sticky_o)
  );


endmodule



module bsg_scan_width_p64_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [63:0] i;
  output [63:0] o;
  wire [63:0] o;
  wire t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,t_5__11_,
  t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,t_5__1_,
  t_5__0_,t_4__63_,t_4__62_,t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,
  t_4__55_,t_4__54_,t_4__53_,t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,
  t_4__46_,t_4__45_,t_4__44_,t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,
  t_4__37_,t_4__36_,t_4__35_,t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,
  t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,
  t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,
  t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,
  t_4__1_,t_4__0_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,
  t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,
  t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,
  t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,
  t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,
  t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,
  t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,
  t_3__2_,t_3__1_,t_3__0_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,
  t_2__57_,t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,
  t_2__48_,t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,
  t_2__39_,t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,
  t_2__30_,t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__63_,t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,
  t_1__57_,t_1__56_,t_1__55_,t_1__54_,t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,
  t_1__48_,t_1__47_,t_1__46_,t_1__45_,t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,
  t_1__39_,t_1__38_,t_1__37_,t_1__36_,t_1__35_,t_1__34_,t_1__33_,t_1__32_,
  t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,
  t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,
  t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,
  t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__63_ = i[0] | 1'b0;
  assign t_1__62_ = i[1] | i[0];
  assign t_1__61_ = i[2] | i[1];
  assign t_1__60_ = i[3] | i[2];
  assign t_1__59_ = i[4] | i[3];
  assign t_1__58_ = i[5] | i[4];
  assign t_1__57_ = i[6] | i[5];
  assign t_1__56_ = i[7] | i[6];
  assign t_1__55_ = i[8] | i[7];
  assign t_1__54_ = i[9] | i[8];
  assign t_1__53_ = i[10] | i[9];
  assign t_1__52_ = i[11] | i[10];
  assign t_1__51_ = i[12] | i[11];
  assign t_1__50_ = i[13] | i[12];
  assign t_1__49_ = i[14] | i[13];
  assign t_1__48_ = i[15] | i[14];
  assign t_1__47_ = i[16] | i[15];
  assign t_1__46_ = i[17] | i[16];
  assign t_1__45_ = i[18] | i[17];
  assign t_1__44_ = i[19] | i[18];
  assign t_1__43_ = i[20] | i[19];
  assign t_1__42_ = i[21] | i[20];
  assign t_1__41_ = i[22] | i[21];
  assign t_1__40_ = i[23] | i[22];
  assign t_1__39_ = i[24] | i[23];
  assign t_1__38_ = i[25] | i[24];
  assign t_1__37_ = i[26] | i[25];
  assign t_1__36_ = i[27] | i[26];
  assign t_1__35_ = i[28] | i[27];
  assign t_1__34_ = i[29] | i[28];
  assign t_1__33_ = i[30] | i[29];
  assign t_1__32_ = i[31] | i[30];
  assign t_1__31_ = i[32] | i[31];
  assign t_1__30_ = i[33] | i[32];
  assign t_1__29_ = i[34] | i[33];
  assign t_1__28_ = i[35] | i[34];
  assign t_1__27_ = i[36] | i[35];
  assign t_1__26_ = i[37] | i[36];
  assign t_1__25_ = i[38] | i[37];
  assign t_1__24_ = i[39] | i[38];
  assign t_1__23_ = i[40] | i[39];
  assign t_1__22_ = i[41] | i[40];
  assign t_1__21_ = i[42] | i[41];
  assign t_1__20_ = i[43] | i[42];
  assign t_1__19_ = i[44] | i[43];
  assign t_1__18_ = i[45] | i[44];
  assign t_1__17_ = i[46] | i[45];
  assign t_1__16_ = i[47] | i[46];
  assign t_1__15_ = i[48] | i[47];
  assign t_1__14_ = i[49] | i[48];
  assign t_1__13_ = i[50] | i[49];
  assign t_1__12_ = i[51] | i[50];
  assign t_1__11_ = i[52] | i[51];
  assign t_1__10_ = i[53] | i[52];
  assign t_1__9_ = i[54] | i[53];
  assign t_1__8_ = i[55] | i[54];
  assign t_1__7_ = i[56] | i[55];
  assign t_1__6_ = i[57] | i[56];
  assign t_1__5_ = i[58] | i[57];
  assign t_1__4_ = i[59] | i[58];
  assign t_1__3_ = i[60] | i[59];
  assign t_1__2_ = i[61] | i[60];
  assign t_1__1_ = i[62] | i[61];
  assign t_1__0_ = i[63] | i[62];
  assign t_2__63_ = t_1__63_ | 1'b0;
  assign t_2__62_ = t_1__62_ | 1'b0;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__63_ = t_2__63_ | 1'b0;
  assign t_3__62_ = t_2__62_ | 1'b0;
  assign t_3__61_ = t_2__61_ | 1'b0;
  assign t_3__60_ = t_2__60_ | 1'b0;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__63_ = t_3__63_ | 1'b0;
  assign t_4__62_ = t_3__62_ | 1'b0;
  assign t_4__61_ = t_3__61_ | 1'b0;
  assign t_4__60_ = t_3__60_ | 1'b0;
  assign t_4__59_ = t_3__59_ | 1'b0;
  assign t_4__58_ = t_3__58_ | 1'b0;
  assign t_4__57_ = t_3__57_ | 1'b0;
  assign t_4__56_ = t_3__56_ | 1'b0;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__63_ = t_4__63_ | 1'b0;
  assign t_5__62_ = t_4__62_ | 1'b0;
  assign t_5__61_ = t_4__61_ | 1'b0;
  assign t_5__60_ = t_4__60_ | 1'b0;
  assign t_5__59_ = t_4__59_ | 1'b0;
  assign t_5__58_ = t_4__58_ | 1'b0;
  assign t_5__57_ = t_4__57_ | 1'b0;
  assign t_5__56_ = t_4__56_ | 1'b0;
  assign t_5__55_ = t_4__55_ | 1'b0;
  assign t_5__54_ = t_4__54_ | 1'b0;
  assign t_5__53_ = t_4__53_ | 1'b0;
  assign t_5__52_ = t_4__52_ | 1'b0;
  assign t_5__51_ = t_4__51_ | 1'b0;
  assign t_5__50_ = t_4__50_ | 1'b0;
  assign t_5__49_ = t_4__49_ | 1'b0;
  assign t_5__48_ = t_4__48_ | 1'b0;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign o[0] = t_5__63_ | 1'b0;
  assign o[1] = t_5__62_ | 1'b0;
  assign o[2] = t_5__61_ | 1'b0;
  assign o[3] = t_5__60_ | 1'b0;
  assign o[4] = t_5__59_ | 1'b0;
  assign o[5] = t_5__58_ | 1'b0;
  assign o[6] = t_5__57_ | 1'b0;
  assign o[7] = t_5__56_ | 1'b0;
  assign o[8] = t_5__55_ | 1'b0;
  assign o[9] = t_5__54_ | 1'b0;
  assign o[10] = t_5__53_ | 1'b0;
  assign o[11] = t_5__52_ | 1'b0;
  assign o[12] = t_5__51_ | 1'b0;
  assign o[13] = t_5__50_ | 1'b0;
  assign o[14] = t_5__49_ | 1'b0;
  assign o[15] = t_5__48_ | 1'b0;
  assign o[16] = t_5__47_ | 1'b0;
  assign o[17] = t_5__46_ | 1'b0;
  assign o[18] = t_5__45_ | 1'b0;
  assign o[19] = t_5__44_ | 1'b0;
  assign o[20] = t_5__43_ | 1'b0;
  assign o[21] = t_5__42_ | 1'b0;
  assign o[22] = t_5__41_ | 1'b0;
  assign o[23] = t_5__40_ | 1'b0;
  assign o[24] = t_5__39_ | 1'b0;
  assign o[25] = t_5__38_ | 1'b0;
  assign o[26] = t_5__37_ | 1'b0;
  assign o[27] = t_5__36_ | 1'b0;
  assign o[28] = t_5__35_ | 1'b0;
  assign o[29] = t_5__34_ | 1'b0;
  assign o[30] = t_5__33_ | 1'b0;
  assign o[31] = t_5__32_ | 1'b0;
  assign o[32] = t_5__31_ | t_5__63_;
  assign o[33] = t_5__30_ | t_5__62_;
  assign o[34] = t_5__29_ | t_5__61_;
  assign o[35] = t_5__28_ | t_5__60_;
  assign o[36] = t_5__27_ | t_5__59_;
  assign o[37] = t_5__26_ | t_5__58_;
  assign o[38] = t_5__25_ | t_5__57_;
  assign o[39] = t_5__24_ | t_5__56_;
  assign o[40] = t_5__23_ | t_5__55_;
  assign o[41] = t_5__22_ | t_5__54_;
  assign o[42] = t_5__21_ | t_5__53_;
  assign o[43] = t_5__20_ | t_5__52_;
  assign o[44] = t_5__19_ | t_5__51_;
  assign o[45] = t_5__18_ | t_5__50_;
  assign o[46] = t_5__17_ | t_5__49_;
  assign o[47] = t_5__16_ | t_5__48_;
  assign o[48] = t_5__15_ | t_5__47_;
  assign o[49] = t_5__14_ | t_5__46_;
  assign o[50] = t_5__13_ | t_5__45_;
  assign o[51] = t_5__12_ | t_5__44_;
  assign o[52] = t_5__11_ | t_5__43_;
  assign o[53] = t_5__10_ | t_5__42_;
  assign o[54] = t_5__9_ | t_5__41_;
  assign o[55] = t_5__8_ | t_5__40_;
  assign o[56] = t_5__7_ | t_5__39_;
  assign o[57] = t_5__6_ | t_5__38_;
  assign o[58] = t_5__5_ | t_5__37_;
  assign o[59] = t_5__4_ | t_5__36_;
  assign o[60] = t_5__3_ | t_5__35_;
  assign o[61] = t_5__2_ | t_5__34_;
  assign o[62] = t_5__1_ | t_5__33_;
  assign o[63] = t_5__0_ | t_5__32_;

endmodule



module bsg_fpu_sticky
(
  i,
  shamt_i,
  sticky_o
);

  input [63:0] i;
  input [6:0] shamt_i;
  output sticky_o;
  wire sticky_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582;
  wire [63:0] scan_out;

  bsg_scan_width_p64_or_p1_lo_to_hi_p1
  scan0
  (
    .i(i),
    .o(scan_out)
  );

  assign N516 = shamt_i > { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign N0 = N5 & N6;
  assign N1 = N0 & N7;
  assign N2 = N1 & N8;
  assign N3 = N2 & N9;
  assign N4 = N3 & N10;
  assign N518 = N4 & N11;
  assign N5 = ~shamt_i[6];
  assign N6 = ~shamt_i[5];
  assign N7 = ~shamt_i[4];
  assign N8 = ~shamt_i[3];
  assign N9 = ~shamt_i[2];
  assign N10 = ~shamt_i[0];
  assign N11 = ~shamt_i[1];
  assign N12 = N16 & N17;
  assign N13 = N12 & N18;
  assign N14 = N13 & N19;
  assign N15 = N14 & shamt_i[0];
  assign N519 = N15 & N20;
  assign N16 = ~shamt_i[5];
  assign N17 = ~shamt_i[4];
  assign N18 = ~shamt_i[3];
  assign N19 = ~shamt_i[2];
  assign N20 = ~shamt_i[1];
  assign N21 = N25 & N26;
  assign N22 = N21 & N27;
  assign N23 = N22 & N28;
  assign N24 = N23 & N29;
  assign N520 = N24 & shamt_i[1];
  assign N25 = ~shamt_i[5];
  assign N26 = ~shamt_i[4];
  assign N27 = ~shamt_i[3];
  assign N28 = ~shamt_i[2];
  assign N29 = ~shamt_i[0];
  assign N30 = N34 & N35;
  assign N31 = N30 & N36;
  assign N32 = N31 & N37;
  assign N33 = N32 & shamt_i[0];
  assign N521 = N33 & shamt_i[1];
  assign N34 = ~shamt_i[5];
  assign N35 = ~shamt_i[4];
  assign N36 = ~shamt_i[3];
  assign N37 = ~shamt_i[2];
  assign N38 = N42 & N43;
  assign N39 = N38 & N44;
  assign N40 = N39 & shamt_i[2];
  assign N41 = N40 & N45;
  assign N522 = N41 & N46;
  assign N42 = ~shamt_i[5];
  assign N43 = ~shamt_i[4];
  assign N44 = ~shamt_i[3];
  assign N45 = ~shamt_i[0];
  assign N46 = ~shamt_i[1];
  assign N47 = N51 & N52;
  assign N48 = N47 & N53;
  assign N49 = N48 & shamt_i[2];
  assign N50 = N49 & shamt_i[0];
  assign N523 = N50 & N54;
  assign N51 = ~shamt_i[5];
  assign N52 = ~shamt_i[4];
  assign N53 = ~shamt_i[3];
  assign N54 = ~shamt_i[1];
  assign N55 = N59 & N60;
  assign N56 = N55 & N61;
  assign N57 = N56 & shamt_i[2];
  assign N58 = N57 & N62;
  assign N524 = N58 & shamt_i[1];
  assign N59 = ~shamt_i[5];
  assign N60 = ~shamt_i[4];
  assign N61 = ~shamt_i[3];
  assign N62 = ~shamt_i[0];
  assign N63 = N67 & N68;
  assign N64 = N63 & N69;
  assign N65 = N64 & shamt_i[2];
  assign N66 = N65 & shamt_i[0];
  assign N525 = N66 & shamt_i[1];
  assign N67 = ~shamt_i[5];
  assign N68 = ~shamt_i[4];
  assign N69 = ~shamt_i[3];
  assign N70 = N74 & N75;
  assign N71 = N70 & shamt_i[3];
  assign N72 = N71 & N76;
  assign N73 = N72 & N77;
  assign N526 = N73 & N78;
  assign N74 = ~shamt_i[5];
  assign N75 = ~shamt_i[4];
  assign N76 = ~shamt_i[2];
  assign N77 = ~shamt_i[0];
  assign N78 = ~shamt_i[1];
  assign N79 = N83 & N84;
  assign N80 = N79 & shamt_i[3];
  assign N81 = N80 & N85;
  assign N82 = N81 & shamt_i[0];
  assign N527 = N82 & N86;
  assign N83 = ~shamt_i[5];
  assign N84 = ~shamt_i[4];
  assign N85 = ~shamt_i[2];
  assign N86 = ~shamt_i[1];
  assign N87 = N91 & N92;
  assign N88 = N87 & shamt_i[3];
  assign N89 = N88 & N93;
  assign N90 = N89 & N94;
  assign N528 = N90 & shamt_i[1];
  assign N91 = ~shamt_i[5];
  assign N92 = ~shamt_i[4];
  assign N93 = ~shamt_i[2];
  assign N94 = ~shamt_i[0];
  assign N95 = N99 & N100;
  assign N96 = N95 & shamt_i[3];
  assign N97 = N96 & N101;
  assign N98 = N97 & shamt_i[0];
  assign N529 = N98 & shamt_i[1];
  assign N99 = ~shamt_i[5];
  assign N100 = ~shamt_i[4];
  assign N101 = ~shamt_i[2];
  assign N102 = N106 & N107;
  assign N103 = N102 & shamt_i[3];
  assign N104 = N103 & shamt_i[2];
  assign N105 = N104 & N108;
  assign N530 = N105 & N109;
  assign N106 = ~shamt_i[5];
  assign N107 = ~shamt_i[4];
  assign N108 = ~shamt_i[0];
  assign N109 = ~shamt_i[1];
  assign N110 = N114 & N115;
  assign N111 = N110 & shamt_i[3];
  assign N112 = N111 & shamt_i[2];
  assign N113 = N112 & shamt_i[0];
  assign N531 = N113 & N116;
  assign N114 = ~shamt_i[5];
  assign N115 = ~shamt_i[4];
  assign N116 = ~shamt_i[1];
  assign N117 = N121 & N122;
  assign N118 = N117 & shamt_i[3];
  assign N119 = N118 & shamt_i[2];
  assign N120 = N119 & N123;
  assign N532 = N120 & shamt_i[1];
  assign N121 = ~shamt_i[5];
  assign N122 = ~shamt_i[4];
  assign N123 = ~shamt_i[0];
  assign N124 = N128 & N129;
  assign N125 = N124 & shamt_i[3];
  assign N126 = N125 & shamt_i[2];
  assign N127 = N126 & shamt_i[0];
  assign N533 = N127 & shamt_i[1];
  assign N128 = ~shamt_i[5];
  assign N129 = ~shamt_i[4];
  assign N130 = N134 & shamt_i[4];
  assign N131 = N130 & N135;
  assign N132 = N131 & N136;
  assign N133 = N132 & N137;
  assign N534 = N133 & N138;
  assign N134 = ~shamt_i[5];
  assign N135 = ~shamt_i[3];
  assign N136 = ~shamt_i[2];
  assign N137 = ~shamt_i[0];
  assign N138 = ~shamt_i[1];
  assign N139 = N143 & shamt_i[4];
  assign N140 = N139 & N144;
  assign N141 = N140 & N145;
  assign N142 = N141 & shamt_i[0];
  assign N535 = N142 & N146;
  assign N143 = ~shamt_i[5];
  assign N144 = ~shamt_i[3];
  assign N145 = ~shamt_i[2];
  assign N146 = ~shamt_i[1];
  assign N147 = N151 & shamt_i[4];
  assign N148 = N147 & N152;
  assign N149 = N148 & N153;
  assign N150 = N149 & N154;
  assign N536 = N150 & shamt_i[1];
  assign N151 = ~shamt_i[5];
  assign N152 = ~shamt_i[3];
  assign N153 = ~shamt_i[2];
  assign N154 = ~shamt_i[0];
  assign N155 = N159 & shamt_i[4];
  assign N156 = N155 & N160;
  assign N157 = N156 & N161;
  assign N158 = N157 & shamt_i[0];
  assign N537 = N158 & shamt_i[1];
  assign N159 = ~shamt_i[5];
  assign N160 = ~shamt_i[3];
  assign N161 = ~shamt_i[2];
  assign N162 = N166 & shamt_i[4];
  assign N163 = N162 & N167;
  assign N164 = N163 & shamt_i[2];
  assign N165 = N164 & N168;
  assign N538 = N165 & N169;
  assign N166 = ~shamt_i[5];
  assign N167 = ~shamt_i[3];
  assign N168 = ~shamt_i[0];
  assign N169 = ~shamt_i[1];
  assign N170 = N174 & shamt_i[4];
  assign N171 = N170 & N175;
  assign N172 = N171 & shamt_i[2];
  assign N173 = N172 & shamt_i[0];
  assign N539 = N173 & N176;
  assign N174 = ~shamt_i[5];
  assign N175 = ~shamt_i[3];
  assign N176 = ~shamt_i[1];
  assign N177 = N181 & shamt_i[4];
  assign N178 = N177 & N182;
  assign N179 = N178 & shamt_i[2];
  assign N180 = N179 & N183;
  assign N540 = N180 & shamt_i[1];
  assign N181 = ~shamt_i[5];
  assign N182 = ~shamt_i[3];
  assign N183 = ~shamt_i[0];
  assign N184 = N188 & shamt_i[4];
  assign N185 = N184 & N189;
  assign N186 = N185 & shamt_i[2];
  assign N187 = N186 & shamt_i[0];
  assign N541 = N187 & shamt_i[1];
  assign N188 = ~shamt_i[5];
  assign N189 = ~shamt_i[3];
  assign N190 = N194 & shamt_i[4];
  assign N191 = N190 & shamt_i[3];
  assign N192 = N191 & N195;
  assign N193 = N192 & N196;
  assign N542 = N193 & N197;
  assign N194 = ~shamt_i[5];
  assign N195 = ~shamt_i[2];
  assign N196 = ~shamt_i[0];
  assign N197 = ~shamt_i[1];
  assign N198 = N202 & shamt_i[4];
  assign N199 = N198 & shamt_i[3];
  assign N200 = N199 & N203;
  assign N201 = N200 & shamt_i[0];
  assign N543 = N201 & N204;
  assign N202 = ~shamt_i[5];
  assign N203 = ~shamt_i[2];
  assign N204 = ~shamt_i[1];
  assign N205 = N209 & shamt_i[4];
  assign N206 = N205 & shamt_i[3];
  assign N207 = N206 & N210;
  assign N208 = N207 & N211;
  assign N544 = N208 & shamt_i[1];
  assign N209 = ~shamt_i[5];
  assign N210 = ~shamt_i[2];
  assign N211 = ~shamt_i[0];
  assign N212 = N216 & shamt_i[4];
  assign N213 = N212 & shamt_i[3];
  assign N214 = N213 & N217;
  assign N215 = N214 & shamt_i[0];
  assign N545 = N215 & shamt_i[1];
  assign N216 = ~shamt_i[5];
  assign N217 = ~shamt_i[2];
  assign N218 = N222 & shamt_i[4];
  assign N219 = N218 & shamt_i[3];
  assign N220 = N219 & shamt_i[2];
  assign N221 = N220 & N223;
  assign N546 = N221 & N224;
  assign N222 = ~shamt_i[5];
  assign N223 = ~shamt_i[0];
  assign N224 = ~shamt_i[1];
  assign N225 = N229 & shamt_i[4];
  assign N226 = N225 & shamt_i[3];
  assign N227 = N226 & shamt_i[2];
  assign N228 = N227 & shamt_i[0];
  assign N547 = N228 & N230;
  assign N229 = ~shamt_i[5];
  assign N230 = ~shamt_i[1];
  assign N231 = N235 & shamt_i[4];
  assign N232 = N231 & shamt_i[3];
  assign N233 = N232 & shamt_i[2];
  assign N234 = N233 & N236;
  assign N548 = N234 & shamt_i[1];
  assign N235 = ~shamt_i[5];
  assign N236 = ~shamt_i[0];
  assign N237 = N241 & shamt_i[4];
  assign N238 = N237 & shamt_i[3];
  assign N239 = N238 & shamt_i[2];
  assign N240 = N239 & shamt_i[0];
  assign N549 = N240 & shamt_i[1];
  assign N241 = ~shamt_i[5];
  assign N242 = shamt_i[5] & N246;
  assign N243 = N242 & N247;
  assign N244 = N243 & N248;
  assign N245 = N244 & N249;
  assign N550 = N245 & N250;
  assign N246 = ~shamt_i[4];
  assign N247 = ~shamt_i[3];
  assign N248 = ~shamt_i[2];
  assign N249 = ~shamt_i[0];
  assign N250 = ~shamt_i[1];
  assign N251 = shamt_i[5] & N255;
  assign N252 = N251 & N256;
  assign N253 = N252 & N257;
  assign N254 = N253 & shamt_i[0];
  assign N551 = N254 & N258;
  assign N255 = ~shamt_i[4];
  assign N256 = ~shamt_i[3];
  assign N257 = ~shamt_i[2];
  assign N258 = ~shamt_i[1];
  assign N259 = shamt_i[5] & N263;
  assign N260 = N259 & N264;
  assign N261 = N260 & N265;
  assign N262 = N261 & N266;
  assign N552 = N262 & shamt_i[1];
  assign N263 = ~shamt_i[4];
  assign N264 = ~shamt_i[3];
  assign N265 = ~shamt_i[2];
  assign N266 = ~shamt_i[0];
  assign N267 = shamt_i[5] & N271;
  assign N268 = N267 & N272;
  assign N269 = N268 & N273;
  assign N270 = N269 & shamt_i[0];
  assign N553 = N270 & shamt_i[1];
  assign N271 = ~shamt_i[4];
  assign N272 = ~shamt_i[3];
  assign N273 = ~shamt_i[2];
  assign N274 = shamt_i[5] & N278;
  assign N275 = N274 & N279;
  assign N276 = N275 & shamt_i[2];
  assign N277 = N276 & N280;
  assign N554 = N277 & N281;
  assign N278 = ~shamt_i[4];
  assign N279 = ~shamt_i[3];
  assign N280 = ~shamt_i[0];
  assign N281 = ~shamt_i[1];
  assign N282 = shamt_i[5] & N286;
  assign N283 = N282 & N287;
  assign N284 = N283 & shamt_i[2];
  assign N285 = N284 & shamt_i[0];
  assign N555 = N285 & N288;
  assign N286 = ~shamt_i[4];
  assign N287 = ~shamt_i[3];
  assign N288 = ~shamt_i[1];
  assign N289 = shamt_i[5] & N293;
  assign N290 = N289 & N294;
  assign N291 = N290 & shamt_i[2];
  assign N292 = N291 & N295;
  assign N556 = N292 & shamt_i[1];
  assign N293 = ~shamt_i[4];
  assign N294 = ~shamt_i[3];
  assign N295 = ~shamt_i[0];
  assign N296 = shamt_i[5] & N300;
  assign N297 = N296 & N301;
  assign N298 = N297 & shamt_i[2];
  assign N299 = N298 & shamt_i[0];
  assign N557 = N299 & shamt_i[1];
  assign N300 = ~shamt_i[4];
  assign N301 = ~shamt_i[3];
  assign N302 = shamt_i[5] & N306;
  assign N303 = N302 & shamt_i[3];
  assign N304 = N303 & N307;
  assign N305 = N304 & N308;
  assign N558 = N305 & N309;
  assign N306 = ~shamt_i[4];
  assign N307 = ~shamt_i[2];
  assign N308 = ~shamt_i[0];
  assign N309 = ~shamt_i[1];
  assign N310 = shamt_i[5] & N314;
  assign N311 = N310 & shamt_i[3];
  assign N312 = N311 & N315;
  assign N313 = N312 & shamt_i[0];
  assign N559 = N313 & N316;
  assign N314 = ~shamt_i[4];
  assign N315 = ~shamt_i[2];
  assign N316 = ~shamt_i[1];
  assign N317 = shamt_i[5] & N321;
  assign N318 = N317 & shamt_i[3];
  assign N319 = N318 & N322;
  assign N320 = N319 & N323;
  assign N560 = N320 & shamt_i[1];
  assign N321 = ~shamt_i[4];
  assign N322 = ~shamt_i[2];
  assign N323 = ~shamt_i[0];
  assign N324 = shamt_i[5] & N328;
  assign N325 = N324 & shamt_i[3];
  assign N326 = N325 & N329;
  assign N327 = N326 & shamt_i[0];
  assign N561 = N327 & shamt_i[1];
  assign N328 = ~shamt_i[4];
  assign N329 = ~shamt_i[2];
  assign N330 = shamt_i[5] & N334;
  assign N331 = N330 & shamt_i[3];
  assign N332 = N331 & shamt_i[2];
  assign N333 = N332 & N335;
  assign N562 = N333 & N336;
  assign N334 = ~shamt_i[4];
  assign N335 = ~shamt_i[0];
  assign N336 = ~shamt_i[1];
  assign N337 = shamt_i[5] & N341;
  assign N338 = N337 & shamt_i[3];
  assign N339 = N338 & shamt_i[2];
  assign N340 = N339 & shamt_i[0];
  assign N563 = N340 & N342;
  assign N341 = ~shamt_i[4];
  assign N342 = ~shamt_i[1];
  assign N343 = shamt_i[5] & N347;
  assign N344 = N343 & shamt_i[3];
  assign N345 = N344 & shamt_i[2];
  assign N346 = N345 & N348;
  assign N564 = N346 & shamt_i[1];
  assign N347 = ~shamt_i[4];
  assign N348 = ~shamt_i[0];
  assign N349 = shamt_i[5] & N353;
  assign N350 = N349 & shamt_i[3];
  assign N351 = N350 & shamt_i[2];
  assign N352 = N351 & shamt_i[0];
  assign N565 = N352 & shamt_i[1];
  assign N353 = ~shamt_i[4];
  assign N354 = shamt_i[5] & shamt_i[4];
  assign N355 = N354 & N358;
  assign N356 = N355 & N359;
  assign N357 = N356 & N360;
  assign N566 = N357 & N361;
  assign N358 = ~shamt_i[3];
  assign N359 = ~shamt_i[2];
  assign N360 = ~shamt_i[0];
  assign N361 = ~shamt_i[1];
  assign N362 = shamt_i[5] & shamt_i[4];
  assign N363 = N362 & N366;
  assign N364 = N363 & N367;
  assign N365 = N364 & shamt_i[0];
  assign N567 = N365 & N368;
  assign N366 = ~shamt_i[3];
  assign N367 = ~shamt_i[2];
  assign N368 = ~shamt_i[1];
  assign N369 = shamt_i[5] & shamt_i[4];
  assign N370 = N369 & N373;
  assign N371 = N370 & N374;
  assign N372 = N371 & N375;
  assign N568 = N372 & shamt_i[1];
  assign N373 = ~shamt_i[3];
  assign N374 = ~shamt_i[2];
  assign N375 = ~shamt_i[0];
  assign N376 = shamt_i[5] & shamt_i[4];
  assign N377 = N376 & N380;
  assign N378 = N377 & N381;
  assign N379 = N378 & shamt_i[0];
  assign N569 = N379 & shamt_i[1];
  assign N380 = ~shamt_i[3];
  assign N381 = ~shamt_i[2];
  assign N382 = shamt_i[5] & shamt_i[4];
  assign N383 = N382 & N386;
  assign N384 = N383 & shamt_i[2];
  assign N385 = N384 & N387;
  assign N570 = N385 & N388;
  assign N386 = ~shamt_i[3];
  assign N387 = ~shamt_i[0];
  assign N388 = ~shamt_i[1];
  assign N389 = shamt_i[5] & shamt_i[4];
  assign N390 = N389 & N393;
  assign N391 = N390 & shamt_i[2];
  assign N392 = N391 & shamt_i[0];
  assign N571 = N392 & N394;
  assign N393 = ~shamt_i[3];
  assign N394 = ~shamt_i[1];
  assign N395 = shamt_i[5] & shamt_i[4];
  assign N396 = N395 & N399;
  assign N397 = N396 & shamt_i[2];
  assign N398 = N397 & N400;
  assign N572 = N398 & shamt_i[1];
  assign N399 = ~shamt_i[3];
  assign N400 = ~shamt_i[0];
  assign N401 = shamt_i[5] & shamt_i[4];
  assign N402 = N401 & N405;
  assign N403 = N402 & shamt_i[2];
  assign N404 = N403 & shamt_i[0];
  assign N573 = N404 & shamt_i[1];
  assign N405 = ~shamt_i[3];
  assign N406 = shamt_i[5] & shamt_i[4];
  assign N407 = N406 & shamt_i[3];
  assign N408 = N407 & N410;
  assign N409 = N408 & N411;
  assign N574 = N409 & N412;
  assign N410 = ~shamt_i[2];
  assign N411 = ~shamt_i[0];
  assign N412 = ~shamt_i[1];
  assign N413 = shamt_i[5] & shamt_i[4];
  assign N414 = N413 & shamt_i[3];
  assign N415 = N414 & N417;
  assign N416 = N415 & shamt_i[0];
  assign N575 = N416 & N418;
  assign N417 = ~shamt_i[2];
  assign N418 = ~shamt_i[1];
  assign N419 = shamt_i[5] & shamt_i[4];
  assign N420 = N419 & shamt_i[3];
  assign N421 = N420 & N423;
  assign N422 = N421 & N424;
  assign N576 = N422 & shamt_i[1];
  assign N423 = ~shamt_i[2];
  assign N424 = ~shamt_i[0];
  assign N425 = shamt_i[5] & shamt_i[4];
  assign N426 = N425 & shamt_i[3];
  assign N427 = N426 & N429;
  assign N428 = N427 & shamt_i[0];
  assign N577 = N428 & shamt_i[1];
  assign N429 = ~shamt_i[2];
  assign N430 = shamt_i[5] & shamt_i[4];
  assign N431 = N430 & shamt_i[3];
  assign N432 = N431 & shamt_i[2];
  assign N433 = N432 & N434;
  assign N578 = N433 & N435;
  assign N434 = ~shamt_i[0];
  assign N435 = ~shamt_i[1];
  assign N436 = shamt_i[5] & shamt_i[4];
  assign N437 = N436 & shamt_i[3];
  assign N438 = N437 & shamt_i[2];
  assign N439 = N438 & shamt_i[0];
  assign N579 = N439 & N440;
  assign N440 = ~shamt_i[1];
  assign N441 = shamt_i[5] & shamt_i[4];
  assign N442 = N441 & shamt_i[3];
  assign N443 = N442 & shamt_i[2];
  assign N444 = N443 & N445;
  assign N580 = N444 & shamt_i[1];
  assign N445 = ~shamt_i[0];
  assign N446 = shamt_i[5] & shamt_i[4];
  assign N447 = N446 & shamt_i[3];
  assign N448 = N447 & shamt_i[2];
  assign N449 = N448 & shamt_i[0];
  assign N581 = N449 & shamt_i[1];
  assign sticky_o = (N450)? scan_out[63] : 
                    (N517)? N582 : 1'b0;
  assign N450 = N516;
  assign N582 = (N451)? 1'b0 : 
                (N452)? scan_out[0] : 
                (N453)? scan_out[1] : 
                (N454)? scan_out[2] : 
                (N455)? scan_out[3] : 
                (N456)? scan_out[4] : 
                (N457)? scan_out[5] : 
                (N458)? scan_out[6] : 
                (N459)? scan_out[7] : 
                (N460)? scan_out[8] : 
                (N461)? scan_out[9] : 
                (N462)? scan_out[10] : 
                (N463)? scan_out[11] : 
                (N464)? scan_out[12] : 
                (N465)? scan_out[13] : 
                (N466)? scan_out[14] : 
                (N467)? scan_out[15] : 
                (N468)? scan_out[16] : 
                (N469)? scan_out[17] : 
                (N470)? scan_out[18] : 
                (N471)? scan_out[19] : 
                (N472)? scan_out[20] : 
                (N473)? scan_out[21] : 
                (N474)? scan_out[22] : 
                (N475)? scan_out[23] : 
                (N476)? scan_out[24] : 
                (N477)? scan_out[25] : 
                (N478)? scan_out[26] : 
                (N479)? scan_out[27] : 
                (N480)? scan_out[28] : 
                (N481)? scan_out[29] : 
                (N482)? scan_out[30] : 
                (N483)? scan_out[31] : 
                (N484)? scan_out[32] : 
                (N485)? scan_out[33] : 
                (N486)? scan_out[34] : 
                (N487)? scan_out[35] : 
                (N488)? scan_out[36] : 
                (N489)? scan_out[37] : 
                (N490)? scan_out[38] : 
                (N491)? scan_out[39] : 
                (N492)? scan_out[40] : 
                (N493)? scan_out[41] : 
                (N494)? scan_out[42] : 
                (N495)? scan_out[43] : 
                (N496)? scan_out[44] : 
                (N497)? scan_out[45] : 
                (N498)? scan_out[46] : 
                (N499)? scan_out[47] : 
                (N500)? scan_out[48] : 
                (N501)? scan_out[49] : 
                (N502)? scan_out[50] : 
                (N503)? scan_out[51] : 
                (N504)? scan_out[52] : 
                (N505)? scan_out[53] : 
                (N506)? scan_out[54] : 
                (N507)? scan_out[55] : 
                (N508)? scan_out[56] : 
                (N509)? scan_out[57] : 
                (N510)? scan_out[58] : 
                (N511)? scan_out[59] : 
                (N512)? scan_out[60] : 
                (N513)? scan_out[61] : 
                (N514)? scan_out[62] : 
                (N515)? scan_out[63] : 1'b0;
  assign N451 = N518;
  assign N452 = N519;
  assign N453 = N520;
  assign N454 = N521;
  assign N455 = N522;
  assign N456 = N523;
  assign N457 = N524;
  assign N458 = N525;
  assign N459 = N526;
  assign N460 = N527;
  assign N461 = N528;
  assign N462 = N529;
  assign N463 = N530;
  assign N464 = N531;
  assign N465 = N532;
  assign N466 = N533;
  assign N467 = N534;
  assign N468 = N535;
  assign N469 = N536;
  assign N470 = N537;
  assign N471 = N538;
  assign N472 = N539;
  assign N473 = N540;
  assign N474 = N541;
  assign N475 = N542;
  assign N476 = N543;
  assign N477 = N544;
  assign N478 = N545;
  assign N479 = N546;
  assign N480 = N547;
  assign N481 = N548;
  assign N482 = N549;
  assign N483 = N550;
  assign N484 = N551;
  assign N485 = N552;
  assign N486 = N553;
  assign N487 = N554;
  assign N488 = N555;
  assign N489 = N556;
  assign N490 = N557;
  assign N491 = N558;
  assign N492 = N559;
  assign N493 = N560;
  assign N494 = N561;
  assign N495 = N562;
  assign N496 = N563;
  assign N497 = N564;
  assign N498 = N565;
  assign N499 = N566;
  assign N500 = N567;
  assign N501 = N568;
  assign N502 = N569;
  assign N503 = N570;
  assign N504 = N571;
  assign N505 = N572;
  assign N506 = N573;
  assign N507 = N574;
  assign N508 = N575;
  assign N509 = N576;
  assign N510 = N577;
  assign N511 = N578;
  assign N512 = N579;
  assign N513 = N580;
  assign N514 = N581;
  assign N515 = shamt_i[6];
  assign N517 = ~N516;

endmodule

