

module top
(
  vec_i,
  fwd_o,
  fwd_datapath_o,
  bk_o,
  bk_datapath_o
);

  input [7:0] vec_i;
  output [23:0] fwd_o;
  output [23:0] fwd_datapath_o;
  output [23:0] bk_o;
  output [23:0] bk_datapath_o;

  bsg_scatter_gather
  wrapper
  (
    .vec_i(vec_i),
    .fwd_o(fwd_o),
    .fwd_datapath_o(fwd_datapath_o),
    .bk_o(bk_o),
    .bk_datapath_o(bk_datapath_o)
  );


endmodule



module bsg_scatter_gather
(
  vec_i,
  fwd_o,
  fwd_datapath_o,
  bk_o,
  bk_datapath_o
);

  input [7:0] vec_i;
  output [23:0] fwd_o;
  output [23:0] fwd_datapath_o;
  output [23:0] bk_o;
  output [23:0] bk_datapath_o;
  wire [23:0] fwd_o,fwd_datapath_o,bk_o,bk_datapath_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491;
  assign bk_datapath_o[0] = 1'b0;
  assign bk_datapath_o[1] = 1'b0;
  assign bk_datapath_o[2] = 1'b0;
  assign bk_datapath_o[4] = 1'b0;
  assign bk_datapath_o[5] = 1'b0;
  assign bk_datapath_o[8] = 1'b0;
  assign bk_datapath_o[11] = 1'b0;
  assign fwd_datapath_o[14] = 1'b0;
  assign fwd_datapath_o[17] = 1'b0;
  assign fwd_datapath_o[19] = 1'b0;
  assign fwd_datapath_o[20] = 1'b0;
  assign fwd_datapath_o[21] = 1'b0;
  assign fwd_datapath_o[22] = 1'b0;
  assign fwd_datapath_o[23] = 1'b0;
  assign N1028 = N1020 & N1021;
  assign N1029 = N1022 & N1023;
  assign N1030 = N1024 & N1025;
  assign N1031 = N1026 & N1027;
  assign N1032 = N1028 & N1029;
  assign N1033 = N1030 & N1031;
  assign N1034 = N1032 & N1033;
  assign N1035 = vec_i[7] | vec_i[6];
  assign N1036 = vec_i[5] | vec_i[4];
  assign N1037 = vec_i[3] | vec_i[2];
  assign N1038 = vec_i[1] | N1027;
  assign N1039 = N1035 | N1036;
  assign N1040 = N1037 | N1038;
  assign N1041 = N1039 | N1040;
  assign N1043 = vec_i[7] | vec_i[6];
  assign N1044 = vec_i[5] | vec_i[4];
  assign N1045 = vec_i[3] | vec_i[2];
  assign N1046 = N1026 | vec_i[0];
  assign N1047 = N1043 | N1044;
  assign N1048 = N1045 | N1046;
  assign N1049 = N1047 | N1048;
  assign N1051 = vec_i[7] | vec_i[6];
  assign N1052 = vec_i[5] | vec_i[4];
  assign N1053 = vec_i[3] | vec_i[2];
  assign N1054 = N1026 | N1027;
  assign N1055 = N1051 | N1052;
  assign N1056 = N1053 | N1054;
  assign N1057 = N1055 | N1056;
  assign N1059 = vec_i[3] | N1025;
  assign N1060 = vec_i[1] | vec_i[0];
  assign N1061 = N1059 | N1060;
  assign N1062 = N1055 | N1061;
  assign N1064 = vec_i[3] | N1025;
  assign N1065 = vec_i[1] | N1027;
  assign N1066 = N1064 | N1065;
  assign N1067 = N1055 | N1066;
  assign N1069 = vec_i[3] | N1025;
  assign N1070 = N1026 | vec_i[0];
  assign N1071 = N1069 | N1070;
  assign N1072 = N1055 | N1071;
  assign N1074 = vec_i[3] | N1025;
  assign N1075 = N1026 | N1027;
  assign N1076 = N1074 | N1075;
  assign N1077 = N1055 | N1076;
  assign N1079 = N1024 | vec_i[2];
  assign N1080 = vec_i[1] | vec_i[0];
  assign N1081 = N1079 | N1080;
  assign N1082 = N1055 | N1081;
  assign N1084 = N1024 | vec_i[2];
  assign N1085 = vec_i[1] | N1027;
  assign N1086 = N1084 | N1085;
  assign N1087 = N1055 | N1086;
  assign N1089 = N1024 | vec_i[2];
  assign N1090 = N1026 | vec_i[0];
  assign N1091 = N1089 | N1090;
  assign N1092 = N1055 | N1091;
  assign N1094 = N1024 | vec_i[2];
  assign N1095 = N1026 | N1027;
  assign N1096 = N1094 | N1095;
  assign N1097 = N1055 | N1096;
  assign N1099 = N1024 | N1025;
  assign N1100 = vec_i[1] | vec_i[0];
  assign N1101 = N1099 | N1100;
  assign N1102 = N1055 | N1101;
  assign N1104 = N1099 | N1085;
  assign N1105 = N1055 | N1104;
  assign N1107 = N1099 | N1090;
  assign N1108 = N1055 | N1107;
  assign N1110 = N1099 | N1095;
  assign N1111 = N1055 | N1110;
  assign N1113 = vec_i[5] | N1023;
  assign N1114 = N1051 | N1113;
  assign N1115 = N1053 | N1100;
  assign N1116 = N1114 | N1115;
  assign N1118 = vec_i[5] | N1023;
  assign N1119 = N1051 | N1118;
  assign N1120 = N1053 | N1085;
  assign N1121 = N1119 | N1120;
  assign N1123 = vec_i[5] | N1023;
  assign N1124 = N1051 | N1123;
  assign N1125 = N1053 | N1090;
  assign N1126 = N1124 | N1125;
  assign N1128 = vec_i[5] | N1023;
  assign N1129 = N1051 | N1128;
  assign N1130 = N1053 | N1095;
  assign N1131 = N1129 | N1130;
  assign N1133 = vec_i[5] | N1023;
  assign N1134 = vec_i[3] | N1025;
  assign N1135 = N1051 | N1133;
  assign N1136 = N1134 | N1100;
  assign N1137 = N1135 | N1136;
  assign N1139 = N1134 | N1085;
  assign N1140 = N1135 | N1139;
  assign N1142 = N1134 | N1090;
  assign N1143 = N1135 | N1142;
  assign N1145 = N1134 | N1095;
  assign N1146 = N1135 | N1145;
  assign N1148 = N1024 | vec_i[2];
  assign N1149 = N1148 | N1100;
  assign N1150 = N1135 | N1149;
  assign N1152 = N1148 | N1085;
  assign N1153 = N1135 | N1152;
  assign N1155 = N1148 | N1090;
  assign N1156 = N1135 | N1155;
  assign N1158 = N1148 | N1095;
  assign N1159 = N1135 | N1158;
  assign N1161 = N1135 | N1101;
  assign N1163 = N1135 | N1104;
  assign N1165 = N1135 | N1107;
  assign N1167 = N1135 | N1110;
  assign N1169 = N1022 | vec_i[4];
  assign N1170 = N1051 | N1169;
  assign N1171 = N1170 | N1115;
  assign N1173 = N1022 | vec_i[4];
  assign N1174 = vec_i[1] | N1027;
  assign N1175 = N1051 | N1173;
  assign N1176 = N1053 | N1174;
  assign N1177 = N1175 | N1176;
  assign N1179 = N1022 | vec_i[4];
  assign N1180 = N1026 | vec_i[0];
  assign N1181 = N1051 | N1179;
  assign N1182 = N1053 | N1180;
  assign N1183 = N1181 | N1182;
  assign N1185 = N1022 | vec_i[4];
  assign N1186 = N1051 | N1185;
  assign N1187 = N1053 | N1075;
  assign N1188 = N1186 | N1187;
  assign N1190 = N1022 | vec_i[4];
  assign N1191 = N1051 | N1190;
  assign N1192 = N1074 | N1100;
  assign N1193 = N1191 | N1192;
  assign N1195 = N1074 | N1174;
  assign N1196 = N1191 | N1195;
  assign N1198 = N1074 | N1180;
  assign N1199 = N1191 | N1198;
  assign N1201 = N1191 | N1076;
  assign N1203 = N1094 | N1100;
  assign N1204 = N1191 | N1203;
  assign N1206 = N1094 | N1174;
  assign N1207 = N1191 | N1206;
  assign N1209 = N1094 | N1180;
  assign N1210 = N1191 | N1209;
  assign N1212 = N1094 | N1075;
  assign N1213 = N1191 | N1212;
  assign N1215 = N1024 | N1025;
  assign N1216 = N1215 | N1100;
  assign N1217 = N1191 | N1216;
  assign N1219 = N1215 | N1174;
  assign N1220 = N1191 | N1219;
  assign N1222 = N1215 | N1180;
  assign N1223 = N1191 | N1222;
  assign N1225 = N1215 | N1075;
  assign N1226 = N1191 | N1225;
  assign N1228 = N1022 | N1023;
  assign N1229 = N1051 | N1228;
  assign N1230 = N1229 | N1115;
  assign N1232 = N1229 | N1176;
  assign N1234 = N1229 | N1182;
  assign N1236 = N1229 | N1187;
  assign N1238 = N1229 | N1192;
  assign N1240 = N1229 | N1195;
  assign N1242 = N1229 | N1198;
  assign N1244 = N1043 | N1228;
  assign N1245 = N1244 | N1076;
  assign N1247 = N1244 | N1203;
  assign N1249 = N1244 | N1206;
  assign N1251 = N1244 | N1209;
  assign N1253 = N1244 | N1212;
  assign N1255 = N1244 | N1216;
  assign N1257 = N1244 | N1219;
  assign N1259 = N1244 | N1222;
  assign N1261 = N1244 | N1225;
  assign N1263 = vec_i[7] | N1021;
  assign N1264 = N1263 | N1052;
  assign N1265 = N1264 | N1115;
  assign N1267 = vec_i[7] | N1021;
  assign N1268 = N1267 | N1052;
  assign N1269 = N1268 | N1176;
  assign N1271 = vec_i[7] | N1021;
  assign N1272 = N1271 | N1052;
  assign N1273 = N1272 | N1182;
  assign N1275 = vec_i[7] | N1021;
  assign N1276 = N1275 | N1052;
  assign N1277 = N1276 | N1187;
  assign N1279 = vec_i[7] | N1021;
  assign N1280 = N1279 | N1052;
  assign N1281 = N1280 | N1192;
  assign N1283 = N1280 | N1195;
  assign N1285 = N1280 | N1198;
  assign N1287 = N1280 | N1076;
  assign N1289 = N1280 | N1203;
  assign N1291 = N1280 | N1206;
  assign N1293 = N1280 | N1209;
  assign N1295 = N1280 | N1212;
  assign N1297 = N1280 | N1216;
  assign N1299 = N1280 | N1219;
  assign N1301 = N1280 | N1222;
  assign N1303 = N1280 | N1225;
  assign N1305 = N1275 | N1128;
  assign N1306 = N1305 | N1115;
  assign N1308 = N1305 | N1176;
  assign N1310 = N1305 | N1182;
  assign N1312 = N1305 | N1187;
  assign N1314 = N1305 | N1192;
  assign N1316 = N1305 | N1195;
  assign N1318 = N1305 | N1198;
  assign N1320 = N1305 | N1076;
  assign N1322 = N1305 | N1203;
  assign N1324 = N1305 | N1206;
  assign N1326 = N1305 | N1209;
  assign N1328 = N1305 | N1212;
  assign N1330 = N1305 | N1216;
  assign N1332 = N1305 | N1219;
  assign N1334 = N1305 | N1222;
  assign N1336 = N1305 | N1225;
  assign N1338 = N1275 | N1185;
  assign N1339 = N1338 | N1115;
  assign N1341 = N1338 | N1176;
  assign N1343 = N1338 | N1182;
  assign N1345 = N1338 | N1187;
  assign N1347 = N1338 | N1192;
  assign N1349 = N1338 | N1195;
  assign N1351 = N1338 | N1198;
  assign N1353 = N1338 | N1076;
  assign N1355 = N1338 | N1203;
  assign N1357 = N1338 | N1206;
  assign N1359 = N1338 | N1209;
  assign N1361 = N1338 | N1212;
  assign N1363 = N1338 | N1216;
  assign N1365 = N1338 | N1219;
  assign N1367 = N1338 | N1222;
  assign N1369 = N1338 | N1225;
  assign N1371 = N1275 | N1228;
  assign N1372 = N1371 | N1115;
  assign N1374 = N1371 | N1176;
  assign N1376 = N1371 | N1182;
  assign N1378 = N1371 | N1187;
  assign N1380 = N1371 | N1192;
  assign N1382 = N1371 | N1195;
  assign N1384 = N1371 | N1198;
  assign N1386 = N1371 | N1076;
  assign N1388 = N1371 | N1203;
  assign N1390 = N1371 | N1206;
  assign N1392 = N1371 | N1209;
  assign N1394 = N1371 | N1212;
  assign N1396 = N1371 | N1216;
  assign N1398 = N1371 | N1219;
  assign N1400 = N1371 | N1222;
  assign N1402 = N1371 | N1225;
  assign N1404 = N1020 | vec_i[6];
  assign N1405 = N1404 | N1052;
  assign N1406 = N1405 | N1115;
  assign N1408 = N1020 | vec_i[6];
  assign N1409 = N1408 | N1052;
  assign N1410 = N1409 | N1176;
  assign N1412 = N1020 | vec_i[6];
  assign N1413 = N1412 | N1052;
  assign N1414 = N1413 | N1182;
  assign N1416 = N1020 | vec_i[6];
  assign N1417 = N1416 | N1052;
  assign N1418 = N1417 | N1187;
  assign N1420 = N1020 | vec_i[6];
  assign N1421 = N1420 | N1052;
  assign N1422 = N1421 | N1192;
  assign N1424 = N1421 | N1195;
  assign N1426 = N1421 | N1198;
  assign N1428 = N1421 | N1076;
  assign N1430 = N1421 | N1203;
  assign N1432 = N1421 | N1206;
  assign N1434 = N1421 | N1209;
  assign N1436 = N1421 | N1212;
  assign N1438 = N1421 | N1216;
  assign N1440 = N1421 | N1219;
  assign N1442 = N1421 | N1222;
  assign N1444 = N1421 | N1225;
  assign N1446 = N1416 | N1128;
  assign N1447 = N1446 | N1115;
  assign N1449 = N1446 | N1176;
  assign N1451 = N1446 | N1182;
  assign N1453 = N1446 | N1187;
  assign N1455 = N1446 | N1192;
  assign N1457 = N1446 | N1195;
  assign N1459 = N1446 | N1198;
  assign N1461 = N1446 | N1076;
  assign N1463 = N1446 | N1203;
  assign N1465 = N1446 | N1206;
  assign N1467 = N1446 | N1209;
  assign N1469 = N1446 | N1212;
  assign N1471 = N1446 | N1216;
  assign N1473 = N1446 | N1219;
  assign N1475 = N1446 | N1222;
  assign N1477 = N1446 | N1225;
  assign N1479 = N1416 | N1185;
  assign N1480 = N1479 | N1115;
  assign N1482 = N1479 | N1176;
  assign N1484 = N1479 | N1182;
  assign N1486 = N1479 | N1187;
  assign N1488 = N1479 | N1192;
  assign N1490 = N1479 | N1195;
  assign N1492 = N1479 | N1198;
  assign N1494 = N1479 | N1076;
  assign N1496 = N1479 | N1203;
  assign N1498 = N1479 | N1206;
  assign N1500 = N1479 | N1209;
  assign N1502 = N1479 | N1212;
  assign N1504 = N1479 | N1216;
  assign N1506 = N1479 | N1219;
  assign N1508 = N1479 | N1222;
  assign N1510 = N1479 | N1225;
  assign N1512 = N1416 | N1228;
  assign N1513 = N1512 | N1115;
  assign N1515 = N1512 | N1176;
  assign N1517 = N1512 | N1182;
  assign N1519 = N1512 | N1187;
  assign N1521 = N1512 | N1192;
  assign N1523 = N1512 | N1195;
  assign N1525 = N1512 | N1198;
  assign N1527 = N1512 | N1076;
  assign N1529 = N1512 | N1203;
  assign N1531 = N1512 | N1206;
  assign N1533 = N1512 | N1209;
  assign N1535 = N1512 | N1212;
  assign N1537 = N1512 | N1216;
  assign N1539 = N1512 | N1219;
  assign N1541 = N1512 | N1222;
  assign N1543 = N1512 | N1225;
  assign N1545 = N1020 | N1021;
  assign N1546 = N1545 | N1052;
  assign N1547 = N1546 | N1115;
  assign N1549 = N1546 | N1176;
  assign N1551 = N1546 | N1182;
  assign N1553 = N1546 | N1187;
  assign N1555 = N1546 | N1192;
  assign N1557 = N1546 | N1195;
  assign N1559 = N1546 | N1198;
  assign N1561 = N1545 | N1044;
  assign N1562 = N1561 | N1076;
  assign N1564 = N1561 | N1203;
  assign N1566 = N1561 | N1206;
  assign N1568 = N1561 | N1209;
  assign N1570 = N1561 | N1212;
  assign N1572 = N1561 | N1216;
  assign N1574 = N1561 | N1219;
  assign N1576 = N1561 | N1222;
  assign N1578 = N1561 | N1225;
  assign N1580 = N1545 | N1128;
  assign N1581 = N1580 | N1115;
  assign N1583 = N1580 | N1176;
  assign N1585 = N1580 | N1182;
  assign N1587 = N1045 | N1075;
  assign N1588 = N1580 | N1587;
  assign N1590 = N1580 | N1192;
  assign N1592 = N1580 | N1195;
  assign N1594 = N1580 | N1198;
  assign N1596 = N1580 | N1076;
  assign N1598 = N1580 | N1203;
  assign N1600 = N1580 | N1206;
  assign N1602 = N1580 | N1209;
  assign N1604 = N1580 | N1212;
  assign N1606 = N1215 | N1080;
  assign N1607 = N1580 | N1606;
  assign N1609 = N1580 | N1219;
  assign N1611 = N1580 | N1222;
  assign N1613 = N1580 | N1225;
  assign N1615 = N1545 | N1185;
  assign N1616 = N1045 | N1080;
  assign N1617 = N1615 | N1616;
  assign N1619 = N1045 | N1174;
  assign N1620 = N1615 | N1619;
  assign N1622 = N1045 | N1180;
  assign N1623 = N1615 | N1622;
  assign N1625 = N1615 | N1587;
  assign N1627 = N1074 | N1080;
  assign N1628 = N1615 | N1627;
  assign N1630 = N1615 | N1195;
  assign N1632 = N1615 | N1198;
  assign N1634 = N1026 | N1027;
  assign N1635 = N1069 | N1634;
  assign N1636 = N1615 | N1635;
  assign N1638 = N1094 | N1080;
  assign N1639 = N1615 | N1638;
  assign N1641 = N1094 | N1065;
  assign N1642 = N1615 | N1641;
  assign N1644 = N1094 | N1070;
  assign N1645 = N1615 | N1644;
  assign N1647 = N1089 | N1634;
  assign N1648 = N1615 | N1647;
  assign N1650 = N1024 | N1025;
  assign N1651 = N1650 | N1080;
  assign N1652 = N1615 | N1651;
  assign N1654 = N1650 | N1065;
  assign N1655 = N1615 | N1654;
  assign N1657 = N1650 | N1070;
  assign N1658 = N1615 | N1657;
  assign N1660 = N1650 | N1634;
  assign N1661 = N1615 | N1660;
  assign N1663 = N1545 | N1228;
  assign N1664 = N1663 | N1616;
  assign N1666 = N1045 | N1065;
  assign N1667 = N1663 | N1666;
  assign N1669 = N1045 | N1070;
  assign N1670 = N1663 | N1669;
  assign N1672 = N1020 | N1021;
  assign N1673 = N1022 | N1023;
  assign N1674 = N1672 | N1673;
  assign N1675 = N1045 | N1634;
  assign N1676 = N1674 | N1675;
  assign N1678 = N1069 | N1080;
  assign N1679 = N1674 | N1678;
  assign N1681 = N1069 | N1065;
  assign N1682 = N1674 | N1681;
  assign N1684 = N1674 | N1071;
  assign N1686 = N1674 | N1635;
  assign N1688 = N1089 | N1080;
  assign N1689 = N1674 | N1688;
  assign N1691 = N1089 | N1065;
  assign N1692 = N1674 | N1691;
  assign N1694 = N1089 | N1070;
  assign N1695 = N1674 | N1694;
  assign N1697 = N1674 | N1647;
  assign N1699 = N1674 | N1651;
  assign N1701 = N1674 | N1654;
  assign N1703 = N1674 | N1657;
  assign N1705 = vec_i[7] & vec_i[6];
  assign N1706 = vec_i[5] & vec_i[4];
  assign N1707 = vec_i[3] & vec_i[2];
  assign N1708 = vec_i[1] & vec_i[0];
  assign N1709 = N1705 & N1706;
  assign N1710 = N1707 & N1708;
  assign N1711 = N1709 & N1710;
  assign N1712 = N1020 & N1021;
  assign N1713 = N1022 & N1023;
  assign N1714 = N1024 & N1025;
  assign N1715 = N1026 & N1027;
  assign N1716 = N1712 & N1713;
  assign N1717 = N1714 & N1715;
  assign N1718 = N1716 & N1717;
  assign N1719 = N1047 | N1666;
  assign N1721 = N1047 | N1669;
  assign N1723 = N1047 | N1675;
  assign N1725 = N1047 | N1678;
  assign N1727 = N1047 | N1681;
  assign N1729 = N1047 | N1071;
  assign N1731 = N1047 | N1635;
  assign N1733 = N1047 | N1688;
  assign N1735 = N1047 | N1691;
  assign N1737 = N1047 | N1694;
  assign N1739 = N1047 | N1647;
  assign N1741 = N1047 | N1651;
  assign N1743 = N1047 | N1654;
  assign N1745 = N1047 | N1657;
  assign N1747 = N1047 | N1660;
  assign N1749 = N1779 | N1616;
  assign N1751 = N1779 | N1666;
  assign N1753 = N1779 | N1669;
  assign N1755 = N1779 | N1675;
  assign N1757 = N1779 | N1678;
  assign N1759 = N1779 | N1681;
  assign N1761 = N1779 | N1071;
  assign N1763 = N1779 | N1635;
  assign N1765 = N1779 | N1688;
  assign N1767 = N1779 | N1691;
  assign N1769 = N1779 | N1694;
  assign N1771 = N1779 | N1647;
  assign N1773 = N1779 | N1651;
  assign N1775 = N1779 | N1654;
  assign N1777 = N1779 | N1657;
  assign N1779 = N1043 | N1123;
  assign N1780 = N1779 | N1660;
  assign N1782 = N1796 | N1616;
  assign N1784 = N1796 | N1666;
  assign N1786 = N1796 | N1669;
  assign N1788 = N1796 | N1675;
  assign N1790 = N1796 | N1678;
  assign N1792 = N1796 | N1681;
  assign N1794 = N1796 | N1071;
  assign N1796 = N1043 | N1179;
  assign N1797 = N1796 | N1635;
  assign N1799 = N1796 | N1688;
  assign N1801 = N1796 | N1691;
  assign N1803 = N1796 | N1694;
  assign N1805 = N1796 | N1647;
  assign N1807 = N1796 | N1651;
  assign N1809 = N1796 | N1654;
  assign N1811 = N1796 | N1657;
  assign N1813 = N1796 | N1660;
  assign N1815 = N1845 | N1616;
  assign N1817 = N1845 | N1666;
  assign N1819 = N1845 | N1669;
  assign N1821 = N1845 | N1675;
  assign N1823 = N1845 | N1678;
  assign N1825 = N1845 | N1681;
  assign N1827 = N1845 | N1071;
  assign N1829 = N1845 | N1635;
  assign N1831 = N1845 | N1688;
  assign N1833 = N1845 | N1691;
  assign N1835 = N1845 | N1694;
  assign N1837 = N1845 | N1647;
  assign N1839 = N1845 | N1651;
  assign N1841 = N1845 | N1654;
  assign N1843 = N1845 | N1657;
  assign N1845 = N1043 | N1673;
  assign N1846 = N1845 | N1660;
  assign N1848 = N1862 | N1616;
  assign N1850 = N1862 | N1666;
  assign N1852 = N1862 | N1669;
  assign N1854 = N1862 | N1675;
  assign N1856 = N1862 | N1678;
  assign N1858 = N1862 | N1681;
  assign N1860 = N1862 | N1071;
  assign N1862 = N1271 | N1044;
  assign N1863 = N1862 | N1635;
  assign N1865 = N1862 | N1688;
  assign N1867 = N1862 | N1691;
  assign N1869 = N1862 | N1694;
  assign N1871 = N1862 | N1647;
  assign N1873 = N1862 | N1651;
  assign N1875 = N1862 | N1654;
  assign N1877 = N1862 | N1657;
  assign N1879 = N1862 | N1660;
  assign N1881 = N1911 | N1616;
  assign N1883 = N1911 | N1666;
  assign N1885 = N1911 | N1669;
  assign N1887 = N1911 | N1675;
  assign N1889 = N1911 | N1678;
  assign N1891 = N1911 | N1681;
  assign N1893 = N1911 | N1071;
  assign N1895 = N1911 | N1635;
  assign N1897 = N1911 | N1688;
  assign N1899 = N1911 | N1691;
  assign N1901 = N1911 | N1694;
  assign N1903 = N1911 | N1647;
  assign N1905 = N1911 | N1651;
  assign N1907 = N1911 | N1654;
  assign N1909 = N1911 | N1657;
  assign N1911 = N1271 | N1123;
  assign N1912 = N1911 | N1660;
  assign N1914 = N1928 | N1616;
  assign N1916 = N1928 | N1666;
  assign N1918 = N1928 | N1669;
  assign N1920 = N1928 | N1675;
  assign N1922 = N1928 | N1678;
  assign N1924 = N1928 | N1681;
  assign N1926 = N1928 | N1071;
  assign N1928 = N1271 | N1179;
  assign N1929 = N1928 | N1635;
  assign N1931 = N1928 | N1688;
  assign N1933 = N1928 | N1691;
  assign N1935 = N1928 | N1694;
  assign N1937 = N1928 | N1647;
  assign N1939 = N1928 | N1651;
  assign N1941 = N1928 | N1654;
  assign N1943 = N1928 | N1657;
  assign N1945 = N1928 | N1660;
  assign N1947 = N1977 | N1616;
  assign N1949 = N1977 | N1666;
  assign N1951 = N1977 | N1669;
  assign N1953 = N1977 | N1675;
  assign N1955 = N1977 | N1678;
  assign N1957 = N1977 | N1681;
  assign N1959 = N1977 | N1071;
  assign N1961 = N1977 | N1635;
  assign N1963 = N1977 | N1688;
  assign N1965 = N1977 | N1691;
  assign N1967 = N1977 | N1694;
  assign N1969 = N1977 | N1647;
  assign N1971 = N1977 | N1651;
  assign N1973 = N1977 | N1654;
  assign N1975 = N1977 | N1657;
  assign N1977 = N1271 | N1673;
  assign N1978 = N1977 | N1660;
  assign N1980 = N1994 | N1616;
  assign N1982 = N1994 | N1666;
  assign N1984 = N1994 | N1669;
  assign N1986 = N1994 | N1675;
  assign N1988 = N1994 | N1678;
  assign N1990 = N1994 | N1681;
  assign N1992 = N1994 | N1071;
  assign N1994 = N1412 | N1044;
  assign N1995 = N1994 | N1635;
  assign N1997 = N1994 | N1688;
  assign N1999 = N1994 | N1691;
  assign N2001 = N1994 | N1694;
  assign N2003 = N1994 | N1647;
  assign N2005 = N1994 | N1651;
  assign N2007 = N1994 | N1654;
  assign N2009 = N1994 | N1657;
  assign N2011 = N1994 | N1660;
  assign N2013 = N2043 | N1616;
  assign N2015 = N2043 | N1666;
  assign N2017 = N2043 | N1669;
  assign N2019 = N2043 | N1675;
  assign N2021 = N2043 | N1678;
  assign N2023 = N2043 | N1681;
  assign N2025 = N2043 | N1071;
  assign N2027 = N2043 | N1635;
  assign N2029 = N2043 | N1688;
  assign N2031 = N2043 | N1691;
  assign N2033 = N2043 | N1694;
  assign N2035 = N2043 | N1647;
  assign N2037 = N2043 | N1651;
  assign N2039 = N2043 | N1654;
  assign N2041 = N2043 | N1657;
  assign N2043 = N1412 | N1123;
  assign N2044 = N2043 | N1660;
  assign N2046 = N2060 | N1616;
  assign N2048 = N2060 | N1666;
  assign N2050 = N2060 | N1669;
  assign N2052 = N2060 | N1675;
  assign N2054 = N2060 | N1678;
  assign N2056 = N2060 | N1681;
  assign N2058 = N2060 | N1071;
  assign N2060 = N1412 | N1179;
  assign N2061 = N2060 | N1635;
  assign N2063 = N2060 | N1688;
  assign N2065 = N2060 | N1691;
  assign N2067 = N2060 | N1694;
  assign N2069 = N2060 | N1647;
  assign N2071 = N2060 | N1651;
  assign N2073 = N1650 | N2253;
  assign N2074 = N2060 | N2073;
  assign N2076 = N2060 | N2295;
  assign N2078 = N2060 | N2298;
  assign N2080 = N1412 | N1673;
  assign N2081 = N2080 | N1616;
  assign N2083 = N2080 | N2254;
  assign N2085 = N2080 | N2258;
  assign N2087 = N2080 | N2261;
  assign N2089 = N2080 | N2264;
  assign N2091 = N2080 | N2267;
  assign N2093 = N2111 | N2270;
  assign N2095 = N2111 | N2273;
  assign N2097 = N2111 | N2276;
  assign N2099 = N2111 | N2279;
  assign N2101 = N2111 | N2282;
  assign N2103 = N2111 | N2285;
  assign N2105 = N2111 | N2289;
  assign N2107 = N2111 | N2292;
  assign N2109 = N2111 | N2295;
  assign N2111 = N1412 | N2376;
  assign N2112 = N2111 | N2298;
  assign N2114 = N2128 | N1616;
  assign N2116 = N2128 | N2254;
  assign N2118 = N2128 | N2258;
  assign N2120 = N2128 | N2261;
  assign N2122 = N2128 | N2264;
  assign N2124 = N2128 | N2267;
  assign N2126 = N2128 | N2270;
  assign N2128 = N1672 | N1044;
  assign N2129 = N2128 | N2273;
  assign N2131 = N2128 | N2276;
  assign N2133 = N2128 | N2279;
  assign N2135 = N2128 | N2282;
  assign N2137 = N2128 | N2285;
  assign N2139 = N2128 | N2289;
  assign N2141 = N2128 | N2292;
  assign N2143 = N2128 | N2295;
  assign N2145 = N2128 | N2298;
  assign N2147 = N1672 | N1118;
  assign N2148 = N2147 | N1616;
  assign N2150 = N2147 | N2254;
  assign N2152 = N2147 | N2258;
  assign N2154 = N2147 | N2261;
  assign N2156 = N2147 | N2264;
  assign N2158 = N2147 | N2267;
  assign N2160 = N2179 | N2270;
  assign N2162 = N2179 | N2273;
  assign N2164 = N2179 | N2276;
  assign N2166 = N2179 | N2279;
  assign N2168 = N2179 | N2282;
  assign N2170 = N2179 | N2285;
  assign N2172 = N2179 | N2289;
  assign N2174 = N2179 | N2292;
  assign N2176 = N2179 | N2295;
  assign N2178 = N1020 | N1021;
  assign N2179 = N2178 | N1118;
  assign N2180 = N2179 | N2298;
  assign N2182 = N2196 | N1616;
  assign N2184 = N2196 | N2254;
  assign N2186 = N2196 | N2258;
  assign N2188 = N2196 | N2261;
  assign N2190 = N2196 | N2264;
  assign N2192 = N2196 | N2267;
  assign N2194 = N2196 | N2270;
  assign N2196 = N2178 | N1173;
  assign N2197 = N2196 | N2273;
  assign N2199 = N2196 | N2276;
  assign N2201 = N2196 | N2279;
  assign N2203 = N2196 | N2282;
  assign N2205 = N2196 | N2285;
  assign N2207 = N2196 | N2289;
  assign N2209 = N2196 | N2292;
  assign N2211 = N2196 | N2295;
  assign N2213 = N2196 | N2298;
  assign N2215 = N2229 | N1616;
  assign N2217 = N2229 | N2254;
  assign N2219 = N2229 | N2258;
  assign N2221 = N2229 | N2261;
  assign N2223 = N2229 | N2264;
  assign N2225 = N2229 | N2267;
  assign N2227 = N2229 | N2270;
  assign N2229 = N2178 | N2376;
  assign N2230 = N2229 | N2273;
  assign N2232 = N2229 | N2276;
  assign N2234 = N2229 | N2279;
  assign N2236 = N2229 | N2282;
  assign N2238 = N2229 | N2285;
  assign N2240 = N2229 | N2289;
  assign N2242 = N2229 | N2292;
  assign N2244 = N2229 | N2295;
  assign N2246 = N1020 & N1021;
  assign N2247 = N1022 & N1023;
  assign N2248 = N1024 & N1025;
  assign N2249 = N1026 & N1027;
  assign N2250 = N2246 & N2247;
  assign N2251 = N2248 & N2249;
  assign N2252 = N2250 & N2251;
  assign N2253 = vec_i[1] | N1027;
  assign N2254 = N1045 | N2253;
  assign N2255 = N1047 | N2254;
  assign N2257 = N1026 | vec_i[0];
  assign N2258 = N1045 | N2257;
  assign N2259 = N1047 | N2258;
  assign N2261 = N1045 | N1054;
  assign N2262 = N1047 | N2261;
  assign N2264 = N1064 | N1080;
  assign N2265 = N1047 | N2264;
  assign N2267 = N1064 | N2253;
  assign N2268 = N1047 | N2267;
  assign N2270 = N1064 | N2257;
  assign N2271 = N1047 | N2270;
  assign N2273 = N1064 | N1054;
  assign N2274 = N1047 | N2273;
  assign N2276 = N1084 | N1080;
  assign N2277 = N1047 | N2276;
  assign N2279 = N1084 | N2253;
  assign N2280 = N1047 | N2279;
  assign N2282 = N1084 | N2257;
  assign N2283 = N1047 | N2282;
  assign N2285 = N1084 | N1054;
  assign N2286 = N1047 | N2285;
  assign N2288 = N1024 | N1025;
  assign N2289 = N2288 | N1080;
  assign N2290 = N1047 | N2289;
  assign N2292 = N2288 | N2253;
  assign N2293 = N1047 | N2292;
  assign N2295 = N2288 | N2257;
  assign N2296 = N1047 | N2295;
  assign N2298 = N2288 | N1054;
  assign N2299 = N1047 | N2298;
  assign N2301 = N2309 | N1616;
  assign N2303 = N2309 | N2254;
  assign N2305 = N2309 | N2258;
  assign N2307 = N2309 | N2261;
  assign N2309 = N1043 | N1118;
  assign N2310 = N2309 | N2264;
  assign N2312 = N2309 | N2267;
  assign N2314 = N2309 | N2270;
  assign N2316 = N2309 | N2273;
  assign N2318 = N2309 | N2276;
  assign N2320 = N2309 | N2279;
  assign N2322 = N2309 | N2282;
  assign N2324 = N2309 | N2285;
  assign N2326 = N1035 | N1118;
  assign N2327 = N2326 | N2289;
  assign N2329 = N2326 | N2292;
  assign N2331 = N2326 | N2295;
  assign N2333 = N2326 | N2298;
  assign N2335 = N2343 | N1616;
  assign N2337 = N2343 | N2254;
  assign N2339 = N2343 | N2258;
  assign N2341 = N2343 | N2261;
  assign N2343 = N1035 | N1173;
  assign N2344 = N2343 | N2264;
  assign N2346 = N2343 | N2267;
  assign N2348 = N2343 | N2270;
  assign N2350 = N2343 | N2273;
  assign N2352 = N2343 | N2276;
  assign N2354 = N2343 | N2279;
  assign N2356 = N2343 | N2282;
  assign N2358 = N2343 | N2285;
  assign N2360 = N2343 | N2289;
  assign N2362 = N2343 | N2292;
  assign N2364 = N2343 | N2295;
  assign N2366 = N2343 | N2298;
  assign N2368 = N2377 | N1616;
  assign N2370 = N2377 | N2254;
  assign N2372 = N2377 | N2258;
  assign N2374 = N2377 | N2261;
  assign N2376 = N1022 | N1023;
  assign N2377 = N1035 | N2376;
  assign N2378 = N2377 | N2264;
  assign N2380 = N2377 | N2267;
  assign N2382 = N2377 | N2270;
  assign N2384 = N2377 | N2273;
  assign N2386 = N2377 | N2276;
  assign N2388 = N2377 | N2279;
  assign N2390 = N2377 | N2282;
  assign N2392 = N2377 | N2285;
  assign N2394 = N2377 | N2289;
  assign N2396 = N2377 | N2292;
  assign N2398 = N2377 | N2295;
  assign N2400 = N2377 | N2298;
  assign N2402 = N1267 | N1044;
  assign N2403 = N2402 | N1616;
  assign N2405 = N2402 | N2254;
  assign N2407 = N2402 | N2258;
  assign N2409 = N2402 | N2261;
  assign N2411 = N2402 | N2264;
  assign N2413 = N2402 | N2267;
  assign N2415 = N2402 | N2270;
  assign N2417 = N2402 | N2273;
  assign N2419 = N2402 | N2276;
  assign N2421 = N2402 | N2279;
  assign N2423 = N2402 | N2282;
  assign N2425 = N2402 | N2285;
  assign N2427 = N1267 | N1036;
  assign N2428 = N2427 | N2289;
  assign N2430 = N2427 | N2292;
  assign N2432 = N2427 | N2295;
  assign N2434 = N2427 | N2298;
  assign N2436 = N2444 | N1616;
  assign N2438 = N2444 | N2254;
  assign N2440 = N2444 | N2258;
  assign N2442 = N2444 | N2261;
  assign N2444 = N1267 | N1118;
  assign N2445 = N2444 | N2264;
  assign N2447 = N2444 | N2267;
  assign N2449 = N2444 | N2270;
  assign N2451 = N2444 | N2273;
  assign N2453 = N2444 | N2276;
  assign N2455 = N2444 | N2279;
  assign N2457 = N2444 | N2282;
  assign N2459 = N2444 | N2285;
  assign N2461 = N2444 | N2289;
  assign N2463 = N2444 | N2292;
  assign N2465 = N2444 | N2295;
  assign N2467 = N2444 | N2298;
  assign N2469 = N2477 | N1616;
  assign N2471 = N2477 | N2254;
  assign N2473 = N2477 | N2258;
  assign N2475 = N2477 | N2261;
  assign N2477 = N1267 | N1173;
  assign N2478 = N2477 | N2264;
  assign N2480 = N2477 | N2267;
  assign N2482 = N2477 | N2270;
  assign N2484 = N2477 | N2273;
  assign N2486 = N2477 | N2276;
  assign N2488 = N2477 | N2279;
  assign N2490 = N2477 | N2282;
  assign N2492 = N2477 | N2285;
  assign N2494 = N2477 | N2289;
  assign N2496 = N2477 | N2292;
  assign N2498 = N2477 | N2295;
  assign N2500 = N2477 | N2298;
  assign N2502 = N2513 | N2551;
  assign N2504 = N1037 | N2253;
  assign N2505 = N2513 | N2504;
  assign N2507 = N1037 | N2257;
  assign N2508 = N2513 | N2507;
  assign N2510 = N1037 | N2809;
  assign N2511 = N2513 | N2510;
  assign N2513 = N1267 | N2376;
  assign N2514 = N1064 | N1060;
  assign N2515 = N2513 | N2514;
  assign N2517 = N1059 | N1038;
  assign N2518 = N2513 | N2517;
  assign N2520 = N1059 | N1046;
  assign N2521 = N2513 | N2520;
  assign N2523 = N1059 | N2809;
  assign N2524 = N2513 | N2523;
  assign N2526 = N1084 | N1060;
  assign N2527 = N2513 | N2526;
  assign N2529 = N1079 | N1038;
  assign N2530 = N2539 | N2529;
  assign N2532 = N1079 | N1046;
  assign N2533 = N2539 | N2532;
  assign N2535 = N2539 | N2810;
  assign N2537 = N1022 | N1023;
  assign N2538 = N1024 | N1025;
  assign N2539 = N1263 | N2537;
  assign N2540 = N2538 | N1060;
  assign N2541 = N2539 | N2540;
  assign N2543 = N2539 | N2815;
  assign N2545 = N2539 | N2818;
  assign N2547 = N2538 | N2809;
  assign N2548 = N2539 | N2547;
  assign N2550 = N1408 | N1036;
  assign N2551 = N1037 | N1060;
  assign N2552 = N2550 | N2551;
  assign N2554 = N2550 | N1040;
  assign N2556 = N1037 | N1046;
  assign N2557 = N2550 | N2556;
  assign N2559 = N2550 | N2510;
  assign N2561 = N2550 | N1061;
  assign N2563 = N2550 | N2517;
  assign N2565 = N2550 | N2520;
  assign N2567 = N2550 | N2523;
  assign N2569 = N1079 | N1060;
  assign N2570 = N2550 | N2569;
  assign N2572 = N2550 | N2529;
  assign N2574 = N2550 | N2532;
  assign N2576 = N2550 | N2810;
  assign N2578 = N2550 | N2540;
  assign N2580 = N2550 | N2815;
  assign N2582 = N2550 | N2818;
  assign N2584 = N2550 | N2547;
  assign N2586 = N2594 | N2551;
  assign N2588 = N2594 | N1040;
  assign N2590 = N2594 | N2556;
  assign N2592 = N2594 | N2510;
  assign N2594 = N1408 | N1113;
  assign N2595 = N2594 | N1061;
  assign N2597 = N2594 | N2517;
  assign N2599 = N2594 | N2520;
  assign N2601 = N2594 | N2523;
  assign N2603 = N2594 | N2569;
  assign N2605 = N2594 | N2529;
  assign N2607 = N2594 | N2532;
  assign N2609 = N2594 | N2810;
  assign N2611 = N2594 | N2540;
  assign N2613 = N2594 | N2815;
  assign N2615 = N2594 | N2818;
  assign N2617 = N2594 | N2547;
  assign N2619 = N2627 | N2551;
  assign N2621 = N2627 | N1040;
  assign N2623 = N2627 | N2556;
  assign N2625 = N2627 | N2510;
  assign N2627 = N1408 | N1169;
  assign N2628 = N2627 | N1061;
  assign N2630 = N2627 | N2517;
  assign N2632 = N2627 | N2520;
  assign N2634 = N2627 | N2523;
  assign N2636 = N2627 | N2569;
  assign N2638 = N2627 | N2529;
  assign N2640 = N2627 | N2532;
  assign N2642 = N2627 | N2810;
  assign N2644 = N2627 | N2540;
  assign N2646 = N2627 | N2815;
  assign N2648 = N2627 | N2818;
  assign N2650 = N2627 | N2547;
  assign N2652 = N2660 | N2551;
  assign N2654 = N2660 | N1040;
  assign N2656 = N2660 | N2556;
  assign N2658 = N2660 | N2510;
  assign N2660 = N1408 | N2537;
  assign N2661 = N2660 | N1061;
  assign N2663 = N2660 | N2517;
  assign N2665 = N2660 | N2520;
  assign N2667 = N2660 | N2523;
  assign N2669 = N2660 | N2569;
  assign N2671 = N2677 | N2529;
  assign N2673 = N2677 | N2532;
  assign N2675 = N2677 | N2810;
  assign N2677 = N1404 | N2537;
  assign N2678 = N2677 | N2540;
  assign N2680 = N2677 | N2815;
  assign N2682 = N2677 | N2818;
  assign N2684 = N2677 | N2547;
  assign N2686 = N1020 | N1021;
  assign N2687 = N2686 | N1036;
  assign N2688 = N2687 | N2551;
  assign N2690 = N2687 | N1040;
  assign N2692 = N2687 | N2556;
  assign N2694 = N2687 | N2510;
  assign N2696 = N2687 | N1061;
  assign N2698 = N2687 | N2517;
  assign N2700 = N2687 | N2520;
  assign N2702 = N2687 | N2523;
  assign N2704 = N2687 | N2569;
  assign N2706 = N2687 | N2529;
  assign N2708 = N2687 | N2532;
  assign N2710 = N2687 | N2810;
  assign N2712 = N2687 | N2540;
  assign N2714 = N2687 | N2815;
  assign N2716 = N2687 | N2818;
  assign N2718 = N2687 | N2547;
  assign N2720 = N2728 | N2551;
  assign N2722 = N2728 | N1040;
  assign N2724 = N2728 | N2556;
  assign N2726 = N2728 | N2510;
  assign N2728 = N2686 | N1113;
  assign N2729 = N2728 | N1061;
  assign N2731 = N2728 | N2517;
  assign N2733 = N2728 | N2520;
  assign N2735 = N2728 | N2523;
  assign N2737 = N2728 | N2569;
  assign N2739 = N2728 | N2529;
  assign N2741 = N2728 | N2532;
  assign N2743 = N2728 | N2810;
  assign N2745 = N2728 | N2540;
  assign N2747 = N2728 | N2815;
  assign N2749 = N2728 | N2818;
  assign N2751 = N2728 | N2547;
  assign N2753 = N2761 | N2551;
  assign N2755 = N2761 | N1040;
  assign N2757 = N2761 | N2556;
  assign N2759 = N2761 | N2510;
  assign N2761 = N2686 | N1169;
  assign N2762 = N2761 | N1061;
  assign N2764 = N2761 | N2517;
  assign N2766 = N2761 | N2520;
  assign N2768 = N2761 | N2523;
  assign N2770 = N2761 | N2569;
  assign N2772 = N2761 | N2529;
  assign N2774 = N2761 | N2532;
  assign N2776 = N2761 | N2810;
  assign N2778 = N2761 | N2540;
  assign N2780 = N2761 | N2815;
  assign N2782 = N2761 | N2818;
  assign N2784 = N2761 | N2547;
  assign N2786 = N2794 | N2551;
  assign N2788 = N2794 | N1040;
  assign N2790 = N2794 | N2556;
  assign N2792 = N2794 | N2510;
  assign N2794 = N2686 | N2537;
  assign N2795 = N2794 | N1061;
  assign N2797 = N2794 | N2517;
  assign N2799 = N2794 | N2520;
  assign N2801 = N2794 | N2523;
  assign N2803 = N2794 | N2569;
  assign N2805 = N2794 | N2529;
  assign N2807 = N2794 | N2532;
  assign N2809 = N1026 | N1027;
  assign N2810 = N1079 | N2809;
  assign N2811 = N2794 | N2810;
  assign N2813 = N2794 | N2540;
  assign N2815 = N2538 | N1038;
  assign N2816 = N2794 | N2815;
  assign N2818 = N2538 | N1046;
  assign N2819 = N2794 | N2818;
  assign N2821 = N1020 & N1021;
  assign N2822 = N1022 & N1023;
  assign N2823 = N1024 & N1025;
  assign N2824 = N1026 & N1027;
  assign N2825 = N2821 & N2822;
  assign N2826 = N2823 & N2824;
  assign N2827 = N2825 & N2826;
  assign N2828 = N1039 | N2556;
  assign N2830 = N1039 | N2510;
  assign N2832 = N1039 | N1061;
  assign N2834 = N1039 | N2517;
  assign N2836 = N1039 | N2520;
  assign N2838 = N1039 | N2523;
  assign N2840 = N1039 | N2569;
  assign N2842 = N1039 | N2529;
  assign N2844 = N1039 | N2532;
  assign N2846 = N1039 | N2810;
  assign N2848 = N1039 | N2540;
  assign N2850 = N1039 | N2815;
  assign N2852 = N1039 | N2818;
  assign N2854 = N1039 | N2547;
  assign N2856 = N2864 | N2551;
  assign N2858 = N2864 | N1040;
  assign N2860 = N2864 | N2556;
  assign N2862 = N2864 | N2510;
  assign N2864 = N1035 | N1113;
  assign N2865 = N2864 | N1061;
  assign N2867 = N2864 | N2517;
  assign N2869 = N2864 | N2520;
  assign N2871 = N2864 | N2523;
  assign N2873 = N2864 | N2569;
  assign N2875 = N2864 | N2529;
  assign N2877 = N2864 | N2532;
  assign N2879 = N2864 | N2810;
  assign N2881 = N2864 | N2540;
  assign N2883 = N2864 | N2815;
  assign N2885 = N2864 | N2818;
  assign N2887 = N2864 | N2547;
  assign N2889 = N2897 | N2551;
  assign N2891 = N2897 | N1040;
  assign N2893 = N2897 | N2556;
  assign N2895 = N2897 | N2510;
  assign N2897 = N1035 | N1169;
  assign N2898 = N2897 | N1061;
  assign N2900 = N2897 | N2517;
  assign N2902 = N2897 | N2520;
  assign N2904 = N2897 | N2523;
  assign N2906 = N2897 | N2569;
  assign N2908 = N2897 | N2529;
  assign N2910 = N2897 | N2532;
  assign N2912 = N2897 | N2810;
  assign N2914 = N2897 | N2540;
  assign N2916 = N2897 | N2815;
  assign N2918 = N2897 | N2818;
  assign N2920 = N2897 | N2547;
  assign N2922 = N2930 | N2551;
  assign N2924 = N2930 | N1040;
  assign N2926 = N2930 | N2556;
  assign N2928 = N2930 | N2510;
  assign N2930 = N1035 | N2537;
  assign N2931 = N2930 | N1061;
  assign N2933 = N2930 | N2517;
  assign N2935 = N2930 | N2520;
  assign N2937 = N2930 | N2523;
  assign N2939 = N2930 | N2569;
  assign N2941 = N1079 | N3375;
  assign N2942 = N2930 | N2941;
  assign N2944 = N1079 | N3365;
  assign N2945 = N2930 | N2944;
  assign N2947 = N1079 | N3369;
  assign N2948 = N2930 | N2947;
  assign N2950 = N1022 | N1023;
  assign N2951 = N1024 | N1025;
  assign N2952 = N1035 | N2950;
  assign N2953 = N2951 | N1060;
  assign N2954 = N2952 | N2953;
  assign N2956 = N2952 | N3376;
  assign N2958 = N2952 | N3379;
  assign N2960 = N2951 | N3369;
  assign N2961 = N2952 | N2960;
  assign N2963 = N1263 | N1036;
  assign N2964 = N2963 | N2551;
  assign N2966 = N1037 | N3375;
  assign N2967 = N2963 | N2966;
  assign N2969 = N1037 | N3365;
  assign N2970 = N2963 | N2969;
  assign N2972 = N1037 | N3369;
  assign N2973 = N2963 | N2972;
  assign N2975 = vec_i[3] | N1025;
  assign N2976 = N2975 | N1060;
  assign N2977 = N2963 | N2976;
  assign N2979 = N2975 | N3375;
  assign N2980 = N2963 | N2979;
  assign N2982 = N2975 | N3365;
  assign N2983 = N2963 | N2982;
  assign N2985 = N2975 | N3369;
  assign N2986 = N2963 | N2985;
  assign N2988 = N1024 | vec_i[2];
  assign N2989 = N2988 | N1060;
  assign N2990 = N2963 | N2989;
  assign N2992 = N2988 | N3375;
  assign N2993 = N2963 | N2992;
  assign N2995 = N2963 | N3366;
  assign N2997 = N2963 | N3370;
  assign N2999 = N2963 | N2953;
  assign N3001 = N2963 | N3376;
  assign N3003 = N2963 | N3379;
  assign N3005 = N2963 | N2960;
  assign N3007 = N3016 | N2551;
  assign N3009 = N3016 | N2966;
  assign N3011 = N3016 | N2969;
  assign N3013 = N3016 | N2972;
  assign N3015 = vec_i[5] | N1023;
  assign N3016 = N1263 | N3015;
  assign N3017 = N3016 | N2976;
  assign N3019 = N3016 | N2979;
  assign N3021 = N3016 | N2982;
  assign N3023 = N3016 | N2985;
  assign N3025 = N3016 | N2989;
  assign N3027 = N3016 | N2992;
  assign N3029 = N3016 | N3366;
  assign N3031 = N3016 | N3370;
  assign N3033 = vec_i[7] | N1021;
  assign N3034 = N3033 | N3015;
  assign N3035 = N3034 | N2953;
  assign N3037 = N3034 | N3376;
  assign N3039 = N3034 | N3379;
  assign N3041 = N3034 | N2960;
  assign N3043 = N3052 | N2551;
  assign N3045 = N3052 | N2966;
  assign N3047 = N3052 | N2969;
  assign N3049 = N3052 | N2972;
  assign N3051 = N1022 | vec_i[4];
  assign N3052 = N3033 | N3051;
  assign N3053 = N3052 | N2976;
  assign N3055 = N3052 | N2979;
  assign N3057 = N3052 | N2982;
  assign N3059 = N3052 | N2985;
  assign N3061 = N3052 | N2989;
  assign N3063 = N3052 | N2992;
  assign N3065 = N3052 | N3366;
  assign N3067 = N3052 | N3370;
  assign N3069 = N3052 | N2953;
  assign N3071 = N3052 | N3376;
  assign N3073 = N3052 | N3379;
  assign N3075 = N3052 | N2960;
  assign N3077 = N3085 | N2551;
  assign N3079 = N3085 | N2966;
  assign N3081 = N3085 | N2969;
  assign N3083 = N3085 | N2972;
  assign N3085 = N3033 | N2950;
  assign N3086 = N3085 | N2976;
  assign N3088 = N3085 | N2979;
  assign N3090 = N3085 | N2982;
  assign N3092 = N3085 | N2985;
  assign N3094 = N3085 | N2989;
  assign N3096 = N3085 | N2992;
  assign N3098 = N3085 | N3366;
  assign N3100 = N3085 | N3370;
  assign N3102 = N3085 | N2953;
  assign N3104 = N3085 | N3376;
  assign N3106 = N3085 | N3379;
  assign N3108 = N3085 | N2960;
  assign N3110 = N1404 | N1036;
  assign N3111 = N3110 | N2551;
  assign N3113 = N3110 | N2966;
  assign N3115 = N3110 | N2969;
  assign N3117 = N3110 | N2972;
  assign N3119 = N3110 | N2976;
  assign N3121 = N3110 | N2979;
  assign N3123 = N3110 | N2982;
  assign N3125 = N3110 | N2985;
  assign N3127 = N3110 | N2989;
  assign N3129 = N3110 | N2992;
  assign N3131 = N3110 | N3366;
  assign N3133 = N3110 | N3370;
  assign N3135 = N3110 | N2953;
  assign N3137 = N3110 | N3376;
  assign N3139 = N3110 | N3379;
  assign N3141 = N3110 | N2960;
  assign N3143 = N3151 | N2551;
  assign N3145 = N3151 | N2966;
  assign N3147 = N3151 | N2969;
  assign N3149 = N3151 | N2972;
  assign N3151 = N1404 | N3015;
  assign N3152 = N3151 | N2976;
  assign N3154 = N3151 | N2979;
  assign N3156 = N3151 | N2982;
  assign N3158 = N3151 | N2985;
  assign N3160 = N3151 | N2989;
  assign N3162 = N3151 | N2992;
  assign N3164 = N3151 | N3366;
  assign N3166 = N3151 | N3370;
  assign N3168 = N1020 | vec_i[6];
  assign N3169 = N3168 | N3015;
  assign N3170 = N3169 | N2953;
  assign N3172 = N3169 | N3376;
  assign N3174 = N3169 | N3379;
  assign N3176 = N3169 | N2960;
  assign N3178 = N3186 | N2551;
  assign N3180 = N3186 | N2966;
  assign N3182 = N3186 | N2969;
  assign N3184 = N3186 | N2972;
  assign N3186 = N3168 | N3051;
  assign N3187 = N3186 | N2976;
  assign N3189 = N3186 | N2979;
  assign N3191 = N3186 | N2982;
  assign N3193 = N3186 | N2985;
  assign N3195 = N3186 | N2989;
  assign N3197 = N3186 | N2992;
  assign N3199 = N3186 | N3366;
  assign N3201 = N3186 | N3370;
  assign N3203 = N3186 | N2953;
  assign N3205 = N3186 | N3376;
  assign N3207 = N3186 | N3379;
  assign N3209 = N3186 | N2960;
  assign N3211 = N3219 | N2551;
  assign N3213 = N3219 | N2966;
  assign N3215 = N3219 | N2969;
  assign N3217 = N3219 | N2972;
  assign N3219 = N3168 | N2950;
  assign N3220 = N3219 | N2976;
  assign N3222 = N3219 | N2979;
  assign N3224 = N3219 | N2982;
  assign N3226 = N3219 | N2985;
  assign N3228 = N3219 | N2989;
  assign N3230 = N3219 | N2992;
  assign N3232 = N3219 | N3366;
  assign N3234 = N3219 | N3370;
  assign N3236 = N3219 | N2953;
  assign N3238 = N3219 | N3376;
  assign N3240 = N3219 | N3379;
  assign N3242 = N3219 | N2960;
  assign N3244 = N1020 | N1021;
  assign N3245 = N3244 | N1036;
  assign N3246 = N3245 | N2551;
  assign N3248 = N3245 | N2966;
  assign N3250 = N3245 | N2969;
  assign N3252 = N3245 | N2972;
  assign N3254 = N3245 | N2976;
  assign N3256 = N3245 | N2979;
  assign N3258 = N3245 | N2982;
  assign N3260 = N3245 | N2985;
  assign N3262 = N3245 | N2989;
  assign N3264 = N3245 | N2992;
  assign N3266 = N3245 | N3366;
  assign N3268 = N3245 | N3370;
  assign N3270 = N3245 | N2953;
  assign N3272 = N3245 | N3376;
  assign N3274 = N3245 | N3379;
  assign N3276 = N3245 | N2960;
  assign N3278 = N3286 | N2551;
  assign N3280 = N3286 | N2966;
  assign N3282 = N3286 | N2969;
  assign N3284 = N3286 | N2972;
  assign N3286 = N3244 | N3015;
  assign N3287 = N3286 | N2976;
  assign N3289 = N3286 | N2979;
  assign N3291 = N3286 | N2982;
  assign N3293 = N3286 | N2985;
  assign N3295 = N3286 | N2989;
  assign N3297 = N3286 | N2992;
  assign N3299 = N3286 | N3366;
  assign N3301 = N3286 | N3370;
  assign N3303 = N3286 | N2953;
  assign N3305 = N3286 | N3376;
  assign N3307 = N3286 | N3379;
  assign N3309 = N3286 | N2960;
  assign N3311 = N3319 | N2551;
  assign N3313 = N3319 | N2966;
  assign N3315 = N3319 | N2969;
  assign N3317 = N3319 | N2972;
  assign N3319 = N3244 | N3051;
  assign N3320 = N3319 | N2976;
  assign N3322 = N3319 | N2979;
  assign N3324 = N3319 | N2982;
  assign N3326 = N3319 | N2985;
  assign N3328 = N3319 | N2989;
  assign N3330 = N3319 | N2992;
  assign N3332 = N3319 | N3366;
  assign N3334 = N3319 | N3370;
  assign N3336 = N3319 | N2953;
  assign N3338 = N3319 | N3376;
  assign N3340 = N3319 | N3379;
  assign N3342 = N3319 | N2960;
  assign N3344 = N3352 | N2551;
  assign N3346 = N3352 | N2966;
  assign N3348 = N3352 | N2969;
  assign N3350 = N3352 | N2972;
  assign N3352 = N3244 | N2950;
  assign N3353 = N3352 | N2976;
  assign N3355 = N3352 | N2979;
  assign N3357 = N3352 | N2982;
  assign N3359 = N3352 | N2985;
  assign N3361 = N3352 | N2989;
  assign N3363 = N3352 | N2992;
  assign N3365 = N1026 | vec_i[0];
  assign N3366 = N2988 | N3365;
  assign N3367 = N3352 | N3366;
  assign N3369 = N1026 | N1027;
  assign N3370 = N2988 | N3369;
  assign N3371 = N3352 | N3370;
  assign N3373 = N3352 | N2953;
  assign N3375 = vec_i[1] | N1027;
  assign N3376 = N2951 | N3375;
  assign N3377 = N3352 | N3376;
  assign N3379 = N2951 | N3365;
  assign N3380 = N3352 | N3379;
  assign N3382 = N2252 | N2266 | (N2278 | N2291) | N2311;
  assign N3383 = N2319 | N2328 | (N2345 | N2353) | N2361;
  assign N3384 = N2379 | N2387 | (N2395 | N2404) | N2412;
  assign N3385 = N2420 | N2429 | (N2446 | N2454) | N2462;
  assign N3386 = N2479 | N2487 | (N2495 | N2516) | N2528;
  assign N3387 = N2542 | N2553 | (N2562 | N2571) | N2579;
  assign N3388 = N2596 | N2604 | (N2612 | N2629) | N2637;
  assign N3389 = N2645 | N2662 | (N2670 | N2679) | N2689;
  assign N3390 = N2697 | N2705 | (N2713 | N2730) | N2738;
  assign N3391 = N2746 | N2763 | (N2771 | N2779) | N2796;
  assign N3392 = N2804 | N2814;
  assign N3393 = N3382 | N3383 | (N3384 | N3385) | N3386;
  assign N3394 = N3387 | N3388 | (N3389 | N3390) | N3391;
  assign fwd_o[1] = N3393 | N3394 | N3392;
  assign N3395 = N2252 | N2302 | (N2336 | N2369) | N2404;
  assign N3396 = N2437 | N2470 | (N2503 | N2553) | N2587;
  assign N3397 = N2620 | N2653 | (N2689 | N2721) | N2754;
  assign fwd_o[2] = N3395 | N3396 | (N3397 | N2787);
  assign N3398 = N2833 | N2841 | (N2849 | N2866) | N2874;
  assign N3399 = N2882 | N2899 | (N2907 | N2915) | N2932;
  assign N3400 = N2940 | N2955 | (N2965 | N2978) | N2991;
  assign N3401 = N3000 | N3018 | (N3026 | N3036) | N3054;
  assign N3402 = N3062 | N3070 | (N3087 | N3095) | N3103;
  assign N3403 = N3112 | N3120 | (N3128 | N3136) | N3153;
  assign N3404 = N3161 | N3171 | (N3188 | N3196) | N3204;
  assign N3405 = N3221 | N3229 | (N3237 | N3247) | N3255;
  assign N3406 = N3263 | N3271 | (N3288 | N3296) | N3304;
  assign N3407 = N3321 | N3329 | (N3337 | N3354) | N3362;
  assign N3408 = N3398 | N3399 | (N3400 | N3401) | N3402;
  assign N3409 = N3403 | N3404 | (N3405 | N3406) | N3407;
  assign fwd_datapath_o[1] = N3408 | N3409 | N3374;
  assign N3410 = N3233 | N3235 | (N3237 | N3239) | N3241;
  assign N3411 = N2857 | N2890 | (N2923 | N2965) | N3008;
  assign N3412 = N3044 | N3078 | (N3112 | N3144) | N3179;
  assign N3413 = N3212 | N3247 | (N3279 | N3312) | N3345;
  assign fwd_datapath_o[2] = N3411 | N3412 | N3413;
  assign N3414 = N2892 | N2894 | (N2899 | N2907) | N2923;
  assign N3415 = N2968 | N2971 | (N2978 | N2991) | N3008;
  assign N3416 = N3044 | N3046 | (N3048 | N3054) | N3062;
  assign N3417 = N3078 | N3114 | (N3116 | N3120) | N3128;
  assign N3418 = N3144 | N3179 | (N3181 | N3183) | N3188;
  assign N3419 = N3196 | N3212 | (N3247 | N3249) | N3251;
  assign N3420 = N3255 | N3263 | (N3279 | N3312) | N3314;
  assign N3421 = N3316 | N3321 | (N3329 | N3345);
  assign N3422 = N3414 | N3415 | (N3416 | N3417) | N3418;
  assign N3423 = N3419 | N3420 | N3421;
  assign fwd_datapath_o[5] = N3422 | N3423;
  assign N3424 = N2974 | N2981 | (N2984 | N2994) | N2996;
  assign N3425 = N3000 | N3010 | (N3012 | N3018) | N3026;
  assign N3426 = N3046 | N3048 | (N3054 | N3062) | N3078;
  assign N3427 = N3118 | N3122 | (N3124 | N3130) | N3132;
  assign N3428 = N3136 | N3146 | (N3148 | N3153) | N3161;
  assign N3429 = N3181 | N3183 | (N3188 | N3196) | N3212;
  assign N3430 = N3249 | N3251 | (N3253 | N3255) | N3257;
  assign N3431 = N3259 | N3263 | (N3265 | N3267) | N3271;
  assign N3432 = N3279 | N3281 | (N3283 | N3288) | N3296;
  assign N3433 = N3312 | N3314 | (N3316 | N3321) | N3329;
  assign N3434 = N3424 | N3425 | (N3426 | N3427) | N3428;
  assign N3435 = N3429 | N3430 | (N3431 | N3432) | N3433;
  assign fwd_datapath_o[8] = N3434 | N3435 | N3345;
  assign N3436 = N3126 | N3134 | (N3138 | N3140) | N3150;
  assign N3437 = N3155 | N3157 | (N3163 | N3165) | N3171;
  assign N3438 = N3185 | N3190 | (N3192 | N3198) | N3200;
  assign N3439 = N3204 | N3214 | (N3216 | N3221) | N3229;
  assign N3440 = N3253 | N3257 | (N3259 | N3265) | N3267;
  assign N3441 = N3271 | N3281 | (N3283 | N3288) | N3296;
  assign N3442 = N3314 | N3316 | (N3321 | N3329) | N3345;
  assign N3443 = N3436 | N3437 | (N3438 | N3439) | N3440;
  assign N3444 = N3441 | N3442;
  assign fwd_datapath_o[11] = N3443 | N3444;
  assign N3445 = N2921 | N2938 | (N2949 | N2957) | N2959;
  assign N3446 = N3076 | N3093 | (N3101 | N3105) | N3107;
  assign N3447 = N3142 | N3159 | (N3167 | N3173) | N3175;
  assign N3448 = N3194 | N3202 | (N3206 | N3208) | N3210;
  assign N3449 = N3218 | N3223 | (N3225 | N3227) | N3231;
  assign N3450 = N3261 | N3269 | (N3273 | N3275) | N3285;
  assign N3451 = N3290 | N3292 | (N3298 | N3300) | N3304;
  assign N3452 = N3318 | N3323 | (N3325 | N3331) | N3333;
  assign N3453 = N3337 | N3343 | (N3347 | N3349) | N3354;
  assign N3454 = N3360 | N3362 | (N3372 | N3378) | N3381;
  assign N3455 = N3445 | N3446 | (N3447 | N3448) | N3449;
  assign N3456 = N3410 | N3450 | (N3451 | N3452) | N3453;
  assign fwd_datapath_o[12] = N3455 | N3456 | N3454;
  assign N3457 = N3042 | N3076 | (N3093 | N3101) | N3105;
  assign N3458 = N3107 | N3310 | (N3343 | N3360) | N3372;
  assign N3459 = N3378 | N3381;
  assign fwd_datapath_o[15] = N3457 | N3458 | N3459;
  assign N3460 = N3177 | N3210 | (N3227 | N3235) | N3239;
  assign N3461 = N3241 | N3277 | (N3294 | N3302) | N3306;
  assign N3462 = N3308 | N3327 | (N3335 | N3339) | N3341;
  assign N3463 = N3351 | N3356 | (N3358 | N3364) | N3368;
  assign fwd_datapath_o[16] = N3460 | N3461 | (N3462 | N3463) | N3374;
  assign N3464 = N3243 | N3310 | (N3343 | N3360) | N3372;
  assign fwd_datapath_o[18] = N3464 | N3459;
  assign N3465 = N1732 | N1748 | (N1764 | N1781) | N1798;
  assign N3466 = N1814 | N1830 | (N1847 | N1864) | N1880;
  assign N3467 = N1896 | N1913 | (N1930 | N1946) | N1962;
  assign N3468 = N1979 | N1996 | (N2012 | N2028) | N2045;
  assign N3469 = N2062 | N2079 | (N2096 | N2113) | N2130;
  assign N3470 = N2146 | N2163 | (N2181 | N2198) | N2214;
  assign N3471 = N2231 | N1711;
  assign N3472 = N3465 | N3466 | (N3467 | N3468) | N3469;
  assign N3473 = N3470 | N3471;
  assign bk_datapath_o[7] = N3472 | N3473;
  assign N3474 = N1781 | N1847 | (N1913 | N1979) | N2045;
  assign N3475 = N2113 | N2181 | N1711;
  assign bk_datapath_o[14] = N3474 | N3475;
  assign N3476 = N1814 | N1830 | (N1838 | N1842) | N1844;
  assign N3477 = N1847 | N1946 | (N1962 | N1970) | N1974;
  assign N3478 = N1976 | N1979 | (N2079 | N2096) | N2104;
  assign N3479 = N2108 | N2110 | (N2113 | N2214) | N2231;
  assign N3480 = N2239 | N2243 | (N2245 | N1711);
  assign bk_datapath_o[17] = N3476 | N3477 | (N3478 | N3479) | N3480;
  assign N3481 = N1880 | N1896 | (N1904 | N1908) | N1910;
  assign N3482 = N1913 | N1930 | (N1938 | N1942) | N1944;
  assign N3483 = N1946 | N1954 | (N1958 | N1960) | N1962;
  assign N3484 = N1966 | N1968 | (N1970 | N1972) | N1974;
  assign N3485 = N1976 | N1979 | (N2146 | N2163) | N2171;
  assign N3486 = N2175 | N2177 | (N2181 | N2198) | N2206;
  assign N3487 = N2210 | N2212 | (N2214 | N2222) | N2226;
  assign N3488 = N2228 | N2231 | (N2235 | N2237) | N2239;
  assign N3489 = N2241 | N2243 | (N2245 | N1711);
  assign N3490 = N3481 | N3482 | (N3483 | N3484) | N3485;
  assign N3491 = N3486 | N3487 | (N3488 | N3489);
  assign bk_datapath_o[20] = N3490 | N3491;
  assign bk_o[23] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b0 : 
                    (N129)? 1'b0 : 
                    (N130)? 1'b0 : 
                    (N131)? 1'b0 : 
                    (N132)? 1'b0 : 
                    (N133)? 1'b0 : 
                    (N134)? 1'b0 : 
                    (N135)? 1'b0 : 
                    (N136)? 1'b0 : 
                    (N137)? 1'b0 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b0 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b0 : 
                    (N142)? 1'b0 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b0 : 
                    (N145)? 1'b0 : 
                    (N146)? 1'b0 : 
                    (N147)? 1'b0 : 
                    (N148)? 1'b0 : 
                    (N149)? 1'b0 : 
                    (N150)? 1'b0 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b0 : 
                    (N161)? 1'b0 : 
                    (N162)? 1'b0 : 
                    (N163)? 1'b0 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b0 : 
                    (N166)? 1'b0 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b0 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b0 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b0 : 
                    (N196)? 1'b0 : 
                    (N197)? 1'b0 : 
                    (N198)? 1'b0 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b0 : 
                    (N201)? 1'b0 : 
                    (N202)? 1'b0 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b0 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b0 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b1 : 1'b0;
  assign N0 = N1034;
  assign N1 = N1042;
  assign N2 = N1050;
  assign N3 = N1058;
  assign N4 = N1063;
  assign N5 = N1068;
  assign N6 = N1073;
  assign N7 = N1078;
  assign N8 = N1083;
  assign N9 = N1088;
  assign N10 = N1093;
  assign N11 = N1098;
  assign N12 = N1103;
  assign N13 = N1106;
  assign N14 = N1109;
  assign N15 = N1112;
  assign N16 = N1117;
  assign N17 = N1122;
  assign N18 = N1127;
  assign N19 = N1132;
  assign N20 = N1138;
  assign N21 = N1141;
  assign N22 = N1144;
  assign N23 = N1147;
  assign N24 = N1151;
  assign N25 = N1154;
  assign N26 = N1157;
  assign N27 = N1160;
  assign N28 = N1162;
  assign N29 = N1164;
  assign N30 = N1166;
  assign N31 = N1168;
  assign N32 = N1172;
  assign N33 = N1178;
  assign N34 = N1184;
  assign N35 = N1189;
  assign N36 = N1194;
  assign N37 = N1197;
  assign N38 = N1200;
  assign N39 = N1202;
  assign N40 = N1205;
  assign N41 = N1208;
  assign N42 = N1211;
  assign N43 = N1214;
  assign N44 = N1218;
  assign N45 = N1221;
  assign N46 = N1224;
  assign N47 = N1227;
  assign N48 = N1231;
  assign N49 = N1233;
  assign N50 = N1235;
  assign N51 = N1237;
  assign N52 = N1239;
  assign N53 = N1241;
  assign N54 = N1243;
  assign N55 = N1246;
  assign N56 = N1248;
  assign N57 = N1250;
  assign N58 = N1252;
  assign N59 = N1254;
  assign N60 = N1256;
  assign N61 = N1258;
  assign N62 = N1260;
  assign N63 = N1262;
  assign N64 = N1266;
  assign N65 = N1270;
  assign N66 = N1274;
  assign N67 = N1278;
  assign N68 = N1282;
  assign N69 = N1284;
  assign N70 = N1286;
  assign N71 = N1288;
  assign N72 = N1290;
  assign N73 = N1292;
  assign N74 = N1294;
  assign N75 = N1296;
  assign N76 = N1298;
  assign N77 = N1300;
  assign N78 = N1302;
  assign N79 = N1304;
  assign N80 = N1307;
  assign N81 = N1309;
  assign N82 = N1311;
  assign N83 = N1313;
  assign N84 = N1315;
  assign N85 = N1317;
  assign N86 = N1319;
  assign N87 = N1321;
  assign N88 = N1323;
  assign N89 = N1325;
  assign N90 = N1327;
  assign N91 = N1329;
  assign N92 = N1331;
  assign N93 = N1333;
  assign N94 = N1335;
  assign N95 = N1337;
  assign N96 = N1340;
  assign N97 = N1342;
  assign N98 = N1344;
  assign N99 = N1346;
  assign N100 = N1348;
  assign N101 = N1350;
  assign N102 = N1352;
  assign N103 = N1354;
  assign N104 = N1356;
  assign N105 = N1358;
  assign N106 = N1360;
  assign N107 = N1362;
  assign N108 = N1364;
  assign N109 = N1366;
  assign N110 = N1368;
  assign N111 = N1370;
  assign N112 = N1373;
  assign N113 = N1375;
  assign N114 = N1377;
  assign N115 = N1379;
  assign N116 = N1381;
  assign N117 = N1383;
  assign N118 = N1385;
  assign N119 = N1387;
  assign N120 = N1389;
  assign N121 = N1391;
  assign N122 = N1393;
  assign N123 = N1395;
  assign N124 = N1397;
  assign N125 = N1399;
  assign N126 = N1401;
  assign N127 = N1403;
  assign N128 = N1407;
  assign N129 = N1411;
  assign N130 = N1415;
  assign N131 = N1419;
  assign N132 = N1423;
  assign N133 = N1425;
  assign N134 = N1427;
  assign N135 = N1429;
  assign N136 = N1431;
  assign N137 = N1433;
  assign N138 = N1435;
  assign N139 = N1437;
  assign N140 = N1439;
  assign N141 = N1441;
  assign N142 = N1443;
  assign N143 = N1445;
  assign N144 = N1448;
  assign N145 = N1450;
  assign N146 = N1452;
  assign N147 = N1454;
  assign N148 = N1456;
  assign N149 = N1458;
  assign N150 = N1460;
  assign N151 = N1462;
  assign N152 = N1464;
  assign N153 = N1466;
  assign N154 = N1468;
  assign N155 = N1470;
  assign N156 = N1472;
  assign N157 = N1474;
  assign N158 = N1476;
  assign N159 = N1478;
  assign N160 = N1481;
  assign N161 = N1483;
  assign N162 = N1485;
  assign N163 = N1487;
  assign N164 = N1489;
  assign N165 = N1491;
  assign N166 = N1493;
  assign N167 = N1495;
  assign N168 = N1497;
  assign N169 = N1499;
  assign N170 = N1501;
  assign N171 = N1503;
  assign N172 = N1505;
  assign N173 = N1507;
  assign N174 = N1509;
  assign N175 = N1511;
  assign N176 = N1514;
  assign N177 = N1516;
  assign N178 = N1518;
  assign N179 = N1520;
  assign N180 = N1522;
  assign N181 = N1524;
  assign N182 = N1526;
  assign N183 = N1528;
  assign N184 = N1530;
  assign N185 = N1532;
  assign N186 = N1534;
  assign N187 = N1536;
  assign N188 = N1538;
  assign N189 = N1540;
  assign N190 = N1542;
  assign N191 = N1544;
  assign N192 = N1548;
  assign N193 = N1550;
  assign N194 = N1552;
  assign N195 = N1554;
  assign N196 = N1556;
  assign N197 = N1558;
  assign N198 = N1560;
  assign N199 = N1563;
  assign N200 = N1565;
  assign N201 = N1567;
  assign N202 = N1569;
  assign N203 = N1571;
  assign N204 = N1573;
  assign N205 = N1575;
  assign N206 = N1577;
  assign N207 = N1579;
  assign N208 = N1582;
  assign N209 = N1584;
  assign N210 = N1586;
  assign N211 = N1589;
  assign N212 = N1591;
  assign N213 = N1593;
  assign N214 = N1595;
  assign N215 = N1597;
  assign N216 = N1599;
  assign N217 = N1601;
  assign N218 = N1603;
  assign N219 = N1605;
  assign N220 = N1608;
  assign N221 = N1610;
  assign N222 = N1612;
  assign N223 = N1614;
  assign N224 = N1618;
  assign N225 = N1621;
  assign N226 = N1624;
  assign N227 = N1626;
  assign N228 = N1629;
  assign N229 = N1631;
  assign N230 = N1633;
  assign N231 = N1637;
  assign N232 = N1640;
  assign N233 = N1643;
  assign N234 = N1646;
  assign N235 = N1649;
  assign N236 = N1653;
  assign N237 = N1656;
  assign N238 = N1659;
  assign N239 = N1662;
  assign N240 = N1665;
  assign N241 = N1668;
  assign N242 = N1671;
  assign N243 = N1677;
  assign N244 = N1680;
  assign N245 = N1683;
  assign N246 = N1685;
  assign N247 = N1687;
  assign N248 = N1690;
  assign N249 = N1693;
  assign N250 = N1696;
  assign N251 = N1698;
  assign N252 = N1700;
  assign N253 = N1702;
  assign N254 = N1704;
  assign N255 = N1711;
  assign bk_o[22] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b0 : 
                    (N129)? 1'b0 : 
                    (N130)? 1'b0 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b0 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b0 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b0 : 
                    (N144)? 1'b0 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b0 : 
                    (N158)? 1'b0 : 
                    (N159)? 1'b0 : 
                    (N160)? 1'b0 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b0 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b0 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b0 : 
                    (N174)? 1'b0 : 
                    (N175)? 1'b0 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b0 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b0 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b0 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b0 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b0 : 
                    (N215)? 1'b0 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b0 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[21] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b0 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b0 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b0 : 
                    (N134)? 1'b0 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b0 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b0 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b0 : 
                    (N146)? 1'b0 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b0 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b0 : 
                    (N158)? 1'b0 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b0 : 
                    (N162)? 1'b0 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b0 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b0 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b0 : 
                    (N174)? 1'b0 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b0 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b0 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b0 : 
                    (N200)? 1'b0 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b0 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b0 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b0 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b0 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[20] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b0 : 
                    (N65)? 1'b0 : 
                    (N66)? 1'b0 : 
                    (N67)? 1'b0 : 
                    (N68)? 1'b0 : 
                    (N69)? 1'b0 : 
                    (N70)? 1'b0 : 
                    (N71)? 1'b0 : 
                    (N72)? 1'b0 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N75)? 1'b0 : 
                    (N76)? 1'b0 : 
                    (N77)? 1'b0 : 
                    (N78)? 1'b0 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b0 : 
                    (N82)? 1'b0 : 
                    (N83)? 1'b0 : 
                    (N84)? 1'b0 : 
                    (N85)? 1'b0 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b0 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b0 : 
                    (N98)? 1'b0 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b0 : 
                    (N102)? 1'b0 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b0 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b0 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b0 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b0 : 
                    (N196)? 1'b0 : 
                    (N197)? 1'b0 : 
                    (N198)? 1'b0 : 
                    (N199)? 1'b0 : 
                    (N200)? 1'b0 : 
                    (N201)? 1'b0 : 
                    (N202)? 1'b0 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b0 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b0 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b0 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b0 : 
                    (N228)? 1'b0 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[19] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b0 : 
                    (N65)? 1'b0 : 
                    (N66)? 1'b0 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b0 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b0 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b0 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b0 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b0 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b0 : 
                    (N94)? 1'b0 : 
                    (N95)? 1'b0 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b0 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b0 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b0 : 
                    (N110)? 1'b0 : 
                    (N111)? 1'b0 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b0 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b0 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b0 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b0 : 
                    (N194)? 1'b0 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b0 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b0 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b0 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b0 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[18] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b0 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b0 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b0 : 
                    (N70)? 1'b0 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b0 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b0 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b0 : 
                    (N82)? 1'b0 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b0 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b0 : 
                    (N88)? 1'b0 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b0 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b0 : 
                    (N94)? 1'b0 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b0 : 
                    (N98)? 1'b0 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b0 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b0 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b0 : 
                    (N110)? 1'b0 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b0 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b0 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b0 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b0 : 
                    (N198)? 1'b0 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b0 : 
                    (N202)? 1'b0 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b0 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b0 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b0 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b0 : 1'b0;
  assign bk_o[17] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b0 : 
                    (N33)? 1'b0 : 
                    (N34)? 1'b0 : 
                    (N35)? 1'b0 : 
                    (N36)? 1'b0 : 
                    (N37)? 1'b0 : 
                    (N38)? 1'b0 : 
                    (N39)? 1'b0 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b0 : 
                    (N42)? 1'b0 : 
                    (N43)? 1'b0 : 
                    (N44)? 1'b0 : 
                    (N45)? 1'b0 : 
                    (N46)? 1'b0 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b0 : 
                    (N51)? 1'b0 : 
                    (N52)? 1'b0 : 
                    (N53)? 1'b0 : 
                    (N54)? 1'b0 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b0 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b0 : 
                    (N98)? 1'b0 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b0 : 
                    (N102)? 1'b0 : 
                    (N103)? 1'b0 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b0 : 
                    (N108)? 1'b0 : 
                    (N109)? 1'b0 : 
                    (N110)? 1'b0 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b0 : 
                    (N117)? 1'b0 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b0 : 
                    (N161)? 1'b0 : 
                    (N162)? 1'b0 : 
                    (N163)? 1'b0 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b0 : 
                    (N166)? 1'b0 : 
                    (N167)? 1'b0 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b0 : 
                    (N172)? 1'b0 : 
                    (N173)? 1'b0 : 
                    (N174)? 1'b0 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b0 : 
                    (N228)? 1'b0 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b0 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[16] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b0 : 
                    (N33)? 1'b0 : 
                    (N34)? 1'b0 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b0 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b0 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b0 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b0 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b0 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b0 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b0 : 
                    (N98)? 1'b0 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b0 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b0 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b0 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b0 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b0 : 
                    (N161)? 1'b0 : 
                    (N162)? 1'b0 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b0 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b0 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b0 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b0 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b0 : 
                    (N226)? 1'b0 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b0 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b0 : 1'b0;
  assign bk_o[15] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b0 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b0 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b0 : 
                    (N38)? 1'b0 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b0 : 
                    (N42)? 1'b0 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b0 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b0 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b0 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b0 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b0 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b0 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b0 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b0 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b0 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b0 : 
                    (N102)? 1'b0 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b0 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b0 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b0 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b0 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b0 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b0 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b0 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b0 : 
                    (N166)? 1'b0 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b0 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b0 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b0 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b0 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b0 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b0 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b0 : 
                    (N230)? 1'b0 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[14] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b0 : 
                    (N17)? 1'b0 : 
                    (N18)? 1'b0 : 
                    (N19)? 1'b0 : 
                    (N20)? 1'b0 : 
                    (N21)? 1'b0 : 
                    (N22)? 1'b0 : 
                    (N23)? 1'b0 : 
                    (N24)? 1'b0 : 
                    (N25)? 1'b0 : 
                    (N26)? 1'b0 : 
                    (N27)? 1'b0 : 
                    (N28)? 1'b0 : 
                    (N29)? 1'b0 : 
                    (N30)? 1'b0 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b0 : 
                    (N51)? 1'b0 : 
                    (N52)? 1'b0 : 
                    (N53)? 1'b0 : 
                    (N54)? 1'b0 : 
                    (N55)? 1'b0 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b0 : 
                    (N59)? 1'b0 : 
                    (N60)? 1'b0 : 
                    (N61)? 1'b0 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b0 : 
                    (N82)? 1'b0 : 
                    (N83)? 1'b0 : 
                    (N84)? 1'b0 : 
                    (N85)? 1'b0 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b0 : 
                    (N88)? 1'b0 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b0 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b0 : 
                    (N94)? 1'b0 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b0 : 
                    (N117)? 1'b0 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b0 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b0 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b0 : 
                    (N145)? 1'b0 : 
                    (N146)? 1'b0 : 
                    (N147)? 1'b0 : 
                    (N148)? 1'b0 : 
                    (N149)? 1'b0 : 
                    (N150)? 1'b0 : 
                    (N151)? 1'b0 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b0 : 
                    (N158)? 1'b0 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b0 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b0 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b0 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b0 : 
                    (N215)? 1'b0 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b0 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[13] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b0 : 
                    (N17)? 1'b0 : 
                    (N18)? 1'b0 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b0 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b0 : 
                    (N25)? 1'b1 : 
                    (N26)? 1'b1 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b1 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b0 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b0 : 
                    (N50)? 1'b0 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b0 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b1 : 
                    (N58)? 1'b1 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b1 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b0 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b0 : 
                    (N82)? 1'b0 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b0 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b0 : 
                    (N89)? 1'b1 : 
                    (N90)? 1'b1 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b1 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b0 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b0 : 
                    (N114)? 1'b0 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b0 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b1 : 
                    (N122)? 1'b1 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b1 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b0 : 
                    (N145)? 1'b0 : 
                    (N146)? 1'b0 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b0 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b1 : 
                    (N154)? 1'b1 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b1 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b0 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b0 : 
                    (N178)? 1'b0 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b0 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b1 : 
                    (N186)? 1'b1 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b1 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b0 : 
                    (N210)? 1'b0 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b0 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b1 : 
                    (N218)? 1'b1 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b1 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b0 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b0 : 
                    (N242)? 1'b0 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b0 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b1 : 
                    (N250)? 1'b1 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b1 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b0 : 1'b0;
  assign bk_o[12] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b1 : 
                    (N9)? 1'b1 : 
                    (N10)? 1'b1 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b1 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b0 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b0 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b0 : 
                    (N22)? 1'b0 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b1 : 
                    (N25)? 1'b0 : 
                    (N26)? 1'b0 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b0 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b0 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b1 : 
                    (N41)? 1'b1 : 
                    (N42)? 1'b1 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b1 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b0 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b0 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b0 : 
                    (N54)? 1'b0 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b1 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b0 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b0 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b1 : 
                    (N73)? 1'b1 : 
                    (N74)? 1'b1 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b1 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b0 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b0 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b0 : 
                    (N86)? 1'b0 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b1 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b0 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b1 : 
                    (N105)? 1'b1 : 
                    (N106)? 1'b1 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b1 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b0 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b0 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b0 : 
                    (N118)? 1'b0 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b1 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b1 : 
                    (N137)? 1'b1 : 
                    (N138)? 1'b1 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b1 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b0 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b0 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b0 : 
                    (N150)? 1'b0 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b1 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b0 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b1 : 
                    (N169)? 1'b1 : 
                    (N170)? 1'b1 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b1 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b0 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b0 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b0 : 
                    (N182)? 1'b0 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b1 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b1 : 
                    (N201)? 1'b1 : 
                    (N202)? 1'b1 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b1 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b0 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b0 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b0 : 
                    (N214)? 1'b0 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b1 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b0 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b1 : 
                    (N233)? 1'b1 : 
                    (N234)? 1'b1 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b1 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b0 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b0 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b0 : 
                    (N246)? 1'b0 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b1 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b0 : 1'b0;
  assign bk_o[11] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b0 : 
                    (N9)? 1'b0 : 
                    (N10)? 1'b0 : 
                    (N11)? 1'b0 : 
                    (N12)? 1'b0 : 
                    (N13)? 1'b0 : 
                    (N14)? 1'b0 : 
                    (N15)? 1'b0 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b0 : 
                    (N25)? 1'b0 : 
                    (N26)? 1'b0 : 
                    (N27)? 1'b0 : 
                    (N28)? 1'b0 : 
                    (N29)? 1'b0 : 
                    (N30)? 1'b0 : 
                    (N31)? 1'b0 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b0 : 
                    (N42)? 1'b0 : 
                    (N43)? 1'b0 : 
                    (N44)? 1'b0 : 
                    (N45)? 1'b0 : 
                    (N46)? 1'b0 : 
                    (N47)? 1'b0 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b0 : 
                    (N59)? 1'b0 : 
                    (N60)? 1'b0 : 
                    (N61)? 1'b0 : 
                    (N62)? 1'b0 : 
                    (N63)? 1'b0 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b0 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N75)? 1'b0 : 
                    (N76)? 1'b0 : 
                    (N77)? 1'b0 : 
                    (N78)? 1'b0 : 
                    (N79)? 1'b0 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b0 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b0 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b0 : 
                    (N94)? 1'b0 : 
                    (N95)? 1'b0 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b0 : 
                    (N108)? 1'b0 : 
                    (N109)? 1'b0 : 
                    (N110)? 1'b0 : 
                    (N111)? 1'b0 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b0 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b0 : 
                    (N126)? 1'b0 : 
                    (N127)? 1'b0 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b0 : 
                    (N137)? 1'b0 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b0 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b0 : 
                    (N142)? 1'b0 : 
                    (N143)? 1'b0 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b0 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b0 : 
                    (N158)? 1'b0 : 
                    (N159)? 1'b0 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b0 : 
                    (N172)? 1'b0 : 
                    (N173)? 1'b0 : 
                    (N174)? 1'b0 : 
                    (N175)? 1'b0 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b0 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b0 : 
                    (N190)? 1'b0 : 
                    (N191)? 1'b0 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b0 : 
                    (N201)? 1'b0 : 
                    (N202)? 1'b0 : 
                    (N203)? 1'b0 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b0 : 
                    (N206)? 1'b0 : 
                    (N207)? 1'b0 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b0 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b0 : 
                    (N222)? 1'b0 : 
                    (N223)? 1'b0 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b0 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b0 : 
                    (N238)? 1'b0 : 
                    (N239)? 1'b0 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b0 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b0 : 
                    (N254)? 1'b0 : 
                    (N255)? 1'b0 : 1'b0;
  assign bk_o[10] = (N0)? 1'b1 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b1 : 
                    (N4)? 1'b1 : 
                    (N5)? 1'b1 : 
                    (N6)? 1'b1 : 
                    (N7)? 1'b1 : 
                    (N8)? 1'b0 : 
                    (N9)? 1'b0 : 
                    (N10)? 1'b0 : 
                    (N11)? 1'b1 : 
                    (N12)? 1'b0 : 
                    (N13)? 1'b1 : 
                    (N14)? 1'b1 : 
                    (N15)? 1'b1 : 
                    (N16)? 1'b1 : 
                    (N17)? 1'b1 : 
                    (N18)? 1'b1 : 
                    (N19)? 1'b1 : 
                    (N20)? 1'b1 : 
                    (N21)? 1'b1 : 
                    (N22)? 1'b1 : 
                    (N23)? 1'b1 : 
                    (N24)? 1'b0 : 
                    (N25)? 1'b0 : 
                    (N26)? 1'b0 : 
                    (N27)? 1'b1 : 
                    (N28)? 1'b0 : 
                    (N29)? 1'b1 : 
                    (N30)? 1'b1 : 
                    (N31)? 1'b1 : 
                    (N32)? 1'b1 : 
                    (N33)? 1'b1 : 
                    (N34)? 1'b1 : 
                    (N35)? 1'b1 : 
                    (N36)? 1'b1 : 
                    (N37)? 1'b1 : 
                    (N38)? 1'b1 : 
                    (N39)? 1'b1 : 
                    (N40)? 1'b0 : 
                    (N41)? 1'b0 : 
                    (N42)? 1'b0 : 
                    (N43)? 1'b1 : 
                    (N44)? 1'b0 : 
                    (N45)? 1'b1 : 
                    (N46)? 1'b1 : 
                    (N47)? 1'b1 : 
                    (N48)? 1'b1 : 
                    (N49)? 1'b1 : 
                    (N50)? 1'b1 : 
                    (N51)? 1'b1 : 
                    (N52)? 1'b1 : 
                    (N53)? 1'b1 : 
                    (N54)? 1'b1 : 
                    (N55)? 1'b1 : 
                    (N56)? 1'b0 : 
                    (N57)? 1'b0 : 
                    (N58)? 1'b0 : 
                    (N59)? 1'b1 : 
                    (N60)? 1'b0 : 
                    (N61)? 1'b1 : 
                    (N62)? 1'b1 : 
                    (N63)? 1'b1 : 
                    (N64)? 1'b1 : 
                    (N65)? 1'b1 : 
                    (N66)? 1'b1 : 
                    (N67)? 1'b1 : 
                    (N68)? 1'b1 : 
                    (N69)? 1'b1 : 
                    (N70)? 1'b1 : 
                    (N71)? 1'b1 : 
                    (N72)? 1'b0 : 
                    (N73)? 1'b0 : 
                    (N74)? 1'b0 : 
                    (N75)? 1'b1 : 
                    (N76)? 1'b0 : 
                    (N77)? 1'b1 : 
                    (N78)? 1'b1 : 
                    (N79)? 1'b1 : 
                    (N80)? 1'b1 : 
                    (N81)? 1'b1 : 
                    (N82)? 1'b1 : 
                    (N83)? 1'b1 : 
                    (N84)? 1'b1 : 
                    (N85)? 1'b1 : 
                    (N86)? 1'b1 : 
                    (N87)? 1'b1 : 
                    (N88)? 1'b0 : 
                    (N89)? 1'b0 : 
                    (N90)? 1'b0 : 
                    (N91)? 1'b1 : 
                    (N92)? 1'b0 : 
                    (N93)? 1'b1 : 
                    (N94)? 1'b1 : 
                    (N95)? 1'b1 : 
                    (N96)? 1'b1 : 
                    (N97)? 1'b1 : 
                    (N98)? 1'b1 : 
                    (N99)? 1'b1 : 
                    (N100)? 1'b1 : 
                    (N101)? 1'b1 : 
                    (N102)? 1'b1 : 
                    (N103)? 1'b1 : 
                    (N104)? 1'b0 : 
                    (N105)? 1'b0 : 
                    (N106)? 1'b0 : 
                    (N107)? 1'b1 : 
                    (N108)? 1'b0 : 
                    (N109)? 1'b1 : 
                    (N110)? 1'b1 : 
                    (N111)? 1'b1 : 
                    (N112)? 1'b1 : 
                    (N113)? 1'b1 : 
                    (N114)? 1'b1 : 
                    (N115)? 1'b1 : 
                    (N116)? 1'b1 : 
                    (N117)? 1'b1 : 
                    (N118)? 1'b1 : 
                    (N119)? 1'b1 : 
                    (N120)? 1'b0 : 
                    (N121)? 1'b0 : 
                    (N122)? 1'b0 : 
                    (N123)? 1'b1 : 
                    (N124)? 1'b0 : 
                    (N125)? 1'b1 : 
                    (N126)? 1'b1 : 
                    (N127)? 1'b1 : 
                    (N128)? 1'b1 : 
                    (N129)? 1'b1 : 
                    (N130)? 1'b1 : 
                    (N131)? 1'b1 : 
                    (N132)? 1'b1 : 
                    (N133)? 1'b1 : 
                    (N134)? 1'b1 : 
                    (N135)? 1'b1 : 
                    (N136)? 1'b0 : 
                    (N137)? 1'b0 : 
                    (N138)? 1'b0 : 
                    (N139)? 1'b1 : 
                    (N140)? 1'b0 : 
                    (N141)? 1'b1 : 
                    (N142)? 1'b1 : 
                    (N143)? 1'b1 : 
                    (N144)? 1'b1 : 
                    (N145)? 1'b1 : 
                    (N146)? 1'b1 : 
                    (N147)? 1'b1 : 
                    (N148)? 1'b1 : 
                    (N149)? 1'b1 : 
                    (N150)? 1'b1 : 
                    (N151)? 1'b1 : 
                    (N152)? 1'b0 : 
                    (N153)? 1'b0 : 
                    (N154)? 1'b0 : 
                    (N155)? 1'b1 : 
                    (N156)? 1'b0 : 
                    (N157)? 1'b1 : 
                    (N158)? 1'b1 : 
                    (N159)? 1'b1 : 
                    (N160)? 1'b1 : 
                    (N161)? 1'b1 : 
                    (N162)? 1'b1 : 
                    (N163)? 1'b1 : 
                    (N164)? 1'b1 : 
                    (N165)? 1'b1 : 
                    (N166)? 1'b1 : 
                    (N167)? 1'b1 : 
                    (N168)? 1'b0 : 
                    (N169)? 1'b0 : 
                    (N170)? 1'b0 : 
                    (N171)? 1'b1 : 
                    (N172)? 1'b0 : 
                    (N173)? 1'b1 : 
                    (N174)? 1'b1 : 
                    (N175)? 1'b1 : 
                    (N176)? 1'b1 : 
                    (N177)? 1'b1 : 
                    (N178)? 1'b1 : 
                    (N179)? 1'b1 : 
                    (N180)? 1'b1 : 
                    (N181)? 1'b1 : 
                    (N182)? 1'b1 : 
                    (N183)? 1'b1 : 
                    (N184)? 1'b0 : 
                    (N185)? 1'b0 : 
                    (N186)? 1'b0 : 
                    (N187)? 1'b1 : 
                    (N188)? 1'b0 : 
                    (N189)? 1'b1 : 
                    (N190)? 1'b1 : 
                    (N191)? 1'b1 : 
                    (N192)? 1'b1 : 
                    (N193)? 1'b1 : 
                    (N194)? 1'b1 : 
                    (N195)? 1'b1 : 
                    (N196)? 1'b1 : 
                    (N197)? 1'b1 : 
                    (N198)? 1'b1 : 
                    (N199)? 1'b1 : 
                    (N200)? 1'b0 : 
                    (N201)? 1'b0 : 
                    (N202)? 1'b0 : 
                    (N203)? 1'b1 : 
                    (N204)? 1'b0 : 
                    (N205)? 1'b1 : 
                    (N206)? 1'b1 : 
                    (N207)? 1'b1 : 
                    (N208)? 1'b1 : 
                    (N209)? 1'b1 : 
                    (N210)? 1'b1 : 
                    (N211)? 1'b1 : 
                    (N212)? 1'b1 : 
                    (N213)? 1'b1 : 
                    (N214)? 1'b1 : 
                    (N215)? 1'b1 : 
                    (N216)? 1'b0 : 
                    (N217)? 1'b0 : 
                    (N218)? 1'b0 : 
                    (N219)? 1'b1 : 
                    (N220)? 1'b0 : 
                    (N221)? 1'b1 : 
                    (N222)? 1'b1 : 
                    (N223)? 1'b1 : 
                    (N224)? 1'b1 : 
                    (N225)? 1'b1 : 
                    (N226)? 1'b1 : 
                    (N227)? 1'b1 : 
                    (N228)? 1'b1 : 
                    (N229)? 1'b1 : 
                    (N230)? 1'b1 : 
                    (N231)? 1'b1 : 
                    (N232)? 1'b0 : 
                    (N233)? 1'b0 : 
                    (N234)? 1'b0 : 
                    (N235)? 1'b1 : 
                    (N236)? 1'b0 : 
                    (N237)? 1'b1 : 
                    (N238)? 1'b1 : 
                    (N239)? 1'b1 : 
                    (N240)? 1'b1 : 
                    (N241)? 1'b1 : 
                    (N242)? 1'b1 : 
                    (N243)? 1'b1 : 
                    (N244)? 1'b1 : 
                    (N245)? 1'b1 : 
                    (N246)? 1'b1 : 
                    (N247)? 1'b1 : 
                    (N248)? 1'b0 : 
                    (N249)? 1'b0 : 
                    (N250)? 1'b0 : 
                    (N251)? 1'b1 : 
                    (N252)? 1'b0 : 
                    (N253)? 1'b1 : 
                    (N254)? 1'b1 : 
                    (N255)? 1'b1 : 1'b0;
  assign bk_o[9] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b1 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b1 : 
                   (N6)? 1'b1 : 
                   (N7)? 1'b1 : 
                   (N8)? 1'b0 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b0 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b0 : 
                   (N14)? 1'b0 : 
                   (N15)? 1'b1 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b1 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b1 : 
                   (N22)? 1'b1 : 
                   (N23)? 1'b1 : 
                   (N24)? 1'b0 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b0 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b0 : 
                   (N30)? 1'b0 : 
                   (N31)? 1'b1 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b1 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b1 : 
                   (N38)? 1'b1 : 
                   (N39)? 1'b1 : 
                   (N40)? 1'b0 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b0 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b0 : 
                   (N46)? 1'b0 : 
                   (N47)? 1'b1 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b1 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b1 : 
                   (N54)? 1'b1 : 
                   (N55)? 1'b1 : 
                   (N56)? 1'b0 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b0 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b0 : 
                   (N62)? 1'b0 : 
                   (N63)? 1'b1 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b1 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b1 : 
                   (N70)? 1'b1 : 
                   (N71)? 1'b1 : 
                   (N72)? 1'b0 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b0 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b0 : 
                   (N78)? 1'b0 : 
                   (N79)? 1'b1 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b1 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b1 : 
                   (N86)? 1'b1 : 
                   (N87)? 1'b1 : 
                   (N88)? 1'b0 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b0 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b0 : 
                   (N94)? 1'b0 : 
                   (N95)? 1'b1 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b1 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b1 : 
                   (N102)? 1'b1 : 
                   (N103)? 1'b1 : 
                   (N104)? 1'b0 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b0 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b0 : 
                   (N110)? 1'b0 : 
                   (N111)? 1'b1 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b1 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b1 : 
                   (N118)? 1'b1 : 
                   (N119)? 1'b1 : 
                   (N120)? 1'b0 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b0 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b0 : 
                   (N126)? 1'b0 : 
                   (N127)? 1'b1 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b1 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b1 : 
                   (N134)? 1'b1 : 
                   (N135)? 1'b1 : 
                   (N136)? 1'b0 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b0 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b0 : 
                   (N142)? 1'b0 : 
                   (N143)? 1'b1 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b1 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b1 : 
                   (N150)? 1'b1 : 
                   (N151)? 1'b1 : 
                   (N152)? 1'b0 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b0 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b0 : 
                   (N158)? 1'b0 : 
                   (N159)? 1'b1 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b1 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b1 : 
                   (N166)? 1'b1 : 
                   (N167)? 1'b1 : 
                   (N168)? 1'b0 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b0 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b0 : 
                   (N174)? 1'b0 : 
                   (N175)? 1'b1 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b1 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b1 : 
                   (N182)? 1'b1 : 
                   (N183)? 1'b1 : 
                   (N184)? 1'b0 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b0 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b0 : 
                   (N190)? 1'b0 : 
                   (N191)? 1'b1 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b1 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b1 : 
                   (N198)? 1'b1 : 
                   (N199)? 1'b1 : 
                   (N200)? 1'b0 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b0 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b0 : 
                   (N206)? 1'b0 : 
                   (N207)? 1'b1 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b1 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b1 : 
                   (N214)? 1'b1 : 
                   (N215)? 1'b1 : 
                   (N216)? 1'b0 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b0 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b0 : 
                   (N222)? 1'b0 : 
                   (N223)? 1'b1 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b1 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b1 : 
                   (N230)? 1'b1 : 
                   (N231)? 1'b1 : 
                   (N232)? 1'b0 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b0 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b0 : 
                   (N238)? 1'b0 : 
                   (N239)? 1'b1 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b1 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b1 : 
                   (N246)? 1'b1 : 
                   (N247)? 1'b1 : 
                   (N248)? 1'b0 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b0 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b0 : 
                   (N254)? 1'b0 : 
                   (N255)? 1'b1 : 1'b0;
  assign bk_o[8] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b1 : 
                   (N4)? 1'b0 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b0 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b1 : 
                   (N12)? 1'b0 : 
                   (N13)? 1'b0 : 
                   (N14)? 1'b0 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b1 : 
                   (N20)? 1'b0 : 
                   (N21)? 1'b0 : 
                   (N22)? 1'b0 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b1 : 
                   (N28)? 1'b0 : 
                   (N29)? 1'b0 : 
                   (N30)? 1'b0 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b1 : 
                   (N36)? 1'b0 : 
                   (N37)? 1'b0 : 
                   (N38)? 1'b0 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b1 : 
                   (N44)? 1'b0 : 
                   (N45)? 1'b0 : 
                   (N46)? 1'b0 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b1 : 
                   (N52)? 1'b0 : 
                   (N53)? 1'b0 : 
                   (N54)? 1'b0 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b1 : 
                   (N60)? 1'b0 : 
                   (N61)? 1'b0 : 
                   (N62)? 1'b0 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b1 : 
                   (N68)? 1'b0 : 
                   (N69)? 1'b0 : 
                   (N70)? 1'b0 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b1 : 
                   (N76)? 1'b0 : 
                   (N77)? 1'b0 : 
                   (N78)? 1'b0 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b1 : 
                   (N84)? 1'b0 : 
                   (N85)? 1'b0 : 
                   (N86)? 1'b0 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b1 : 
                   (N92)? 1'b0 : 
                   (N93)? 1'b0 : 
                   (N94)? 1'b0 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b1 : 
                   (N100)? 1'b0 : 
                   (N101)? 1'b0 : 
                   (N102)? 1'b0 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b1 : 
                   (N108)? 1'b0 : 
                   (N109)? 1'b0 : 
                   (N110)? 1'b0 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b1 : 
                   (N116)? 1'b0 : 
                   (N117)? 1'b0 : 
                   (N118)? 1'b0 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b1 : 
                   (N124)? 1'b0 : 
                   (N125)? 1'b0 : 
                   (N126)? 1'b0 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b1 : 
                   (N132)? 1'b0 : 
                   (N133)? 1'b0 : 
                   (N134)? 1'b0 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b1 : 
                   (N140)? 1'b0 : 
                   (N141)? 1'b0 : 
                   (N142)? 1'b0 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b1 : 
                   (N148)? 1'b0 : 
                   (N149)? 1'b0 : 
                   (N150)? 1'b0 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b1 : 
                   (N156)? 1'b0 : 
                   (N157)? 1'b0 : 
                   (N158)? 1'b0 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b1 : 
                   (N164)? 1'b0 : 
                   (N165)? 1'b0 : 
                   (N166)? 1'b0 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b1 : 
                   (N172)? 1'b0 : 
                   (N173)? 1'b0 : 
                   (N174)? 1'b0 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b1 : 
                   (N180)? 1'b0 : 
                   (N181)? 1'b0 : 
                   (N182)? 1'b0 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b1 : 
                   (N188)? 1'b0 : 
                   (N189)? 1'b0 : 
                   (N190)? 1'b0 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b1 : 
                   (N196)? 1'b0 : 
                   (N197)? 1'b0 : 
                   (N198)? 1'b0 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b1 : 
                   (N204)? 1'b0 : 
                   (N205)? 1'b0 : 
                   (N206)? 1'b0 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b1 : 
                   (N212)? 1'b0 : 
                   (N213)? 1'b0 : 
                   (N214)? 1'b0 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b1 : 
                   (N220)? 1'b0 : 
                   (N221)? 1'b0 : 
                   (N222)? 1'b0 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b1 : 
                   (N228)? 1'b0 : 
                   (N229)? 1'b0 : 
                   (N230)? 1'b0 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b1 : 
                   (N236)? 1'b0 : 
                   (N237)? 1'b0 : 
                   (N238)? 1'b0 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b1 : 
                   (N244)? 1'b0 : 
                   (N245)? 1'b0 : 
                   (N246)? 1'b0 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b1 : 
                   (N252)? 1'b0 : 
                   (N253)? 1'b0 : 
                   (N254)? 1'b0 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_o[7] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b1 : 
                   (N4)? 1'b0 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b0 : 
                   (N7)? 1'b1 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b1 : 
                   (N12)? 1'b0 : 
                   (N13)? 1'b0 : 
                   (N14)? 1'b0 : 
                   (N15)? 1'b1 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b1 : 
                   (N20)? 1'b0 : 
                   (N21)? 1'b0 : 
                   (N22)? 1'b0 : 
                   (N23)? 1'b1 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b1 : 
                   (N28)? 1'b0 : 
                   (N29)? 1'b0 : 
                   (N30)? 1'b0 : 
                   (N31)? 1'b1 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b1 : 
                   (N36)? 1'b0 : 
                   (N37)? 1'b0 : 
                   (N38)? 1'b0 : 
                   (N39)? 1'b1 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b1 : 
                   (N44)? 1'b0 : 
                   (N45)? 1'b0 : 
                   (N46)? 1'b0 : 
                   (N47)? 1'b1 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b1 : 
                   (N52)? 1'b0 : 
                   (N53)? 1'b0 : 
                   (N54)? 1'b0 : 
                   (N55)? 1'b1 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b1 : 
                   (N60)? 1'b0 : 
                   (N61)? 1'b0 : 
                   (N62)? 1'b0 : 
                   (N63)? 1'b1 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b1 : 
                   (N68)? 1'b0 : 
                   (N69)? 1'b0 : 
                   (N70)? 1'b0 : 
                   (N71)? 1'b1 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b1 : 
                   (N76)? 1'b0 : 
                   (N77)? 1'b0 : 
                   (N78)? 1'b0 : 
                   (N79)? 1'b1 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b1 : 
                   (N84)? 1'b0 : 
                   (N85)? 1'b0 : 
                   (N86)? 1'b0 : 
                   (N87)? 1'b1 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b1 : 
                   (N92)? 1'b0 : 
                   (N93)? 1'b0 : 
                   (N94)? 1'b0 : 
                   (N95)? 1'b1 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b1 : 
                   (N100)? 1'b0 : 
                   (N101)? 1'b0 : 
                   (N102)? 1'b0 : 
                   (N103)? 1'b1 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b1 : 
                   (N108)? 1'b0 : 
                   (N109)? 1'b0 : 
                   (N110)? 1'b0 : 
                   (N111)? 1'b1 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b1 : 
                   (N116)? 1'b0 : 
                   (N117)? 1'b0 : 
                   (N118)? 1'b0 : 
                   (N119)? 1'b1 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b1 : 
                   (N124)? 1'b0 : 
                   (N125)? 1'b0 : 
                   (N126)? 1'b0 : 
                   (N127)? 1'b1 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b1 : 
                   (N132)? 1'b0 : 
                   (N133)? 1'b0 : 
                   (N134)? 1'b0 : 
                   (N135)? 1'b1 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b1 : 
                   (N140)? 1'b0 : 
                   (N141)? 1'b0 : 
                   (N142)? 1'b0 : 
                   (N143)? 1'b1 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b1 : 
                   (N148)? 1'b0 : 
                   (N149)? 1'b0 : 
                   (N150)? 1'b0 : 
                   (N151)? 1'b1 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b1 : 
                   (N156)? 1'b0 : 
                   (N157)? 1'b0 : 
                   (N158)? 1'b0 : 
                   (N159)? 1'b1 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b1 : 
                   (N164)? 1'b0 : 
                   (N165)? 1'b0 : 
                   (N166)? 1'b0 : 
                   (N167)? 1'b1 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b1 : 
                   (N172)? 1'b0 : 
                   (N173)? 1'b0 : 
                   (N174)? 1'b0 : 
                   (N175)? 1'b1 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b1 : 
                   (N180)? 1'b0 : 
                   (N181)? 1'b0 : 
                   (N182)? 1'b0 : 
                   (N183)? 1'b1 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b1 : 
                   (N188)? 1'b0 : 
                   (N189)? 1'b0 : 
                   (N190)? 1'b0 : 
                   (N191)? 1'b1 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b1 : 
                   (N196)? 1'b0 : 
                   (N197)? 1'b0 : 
                   (N198)? 1'b0 : 
                   (N199)? 1'b1 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b1 : 
                   (N204)? 1'b0 : 
                   (N205)? 1'b0 : 
                   (N206)? 1'b0 : 
                   (N207)? 1'b1 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b1 : 
                   (N212)? 1'b0 : 
                   (N213)? 1'b0 : 
                   (N214)? 1'b0 : 
                   (N215)? 1'b1 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b1 : 
                   (N220)? 1'b0 : 
                   (N221)? 1'b0 : 
                   (N222)? 1'b0 : 
                   (N223)? 1'b1 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b1 : 
                   (N228)? 1'b0 : 
                   (N229)? 1'b0 : 
                   (N230)? 1'b0 : 
                   (N231)? 1'b1 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b1 : 
                   (N236)? 1'b0 : 
                   (N237)? 1'b0 : 
                   (N238)? 1'b0 : 
                   (N239)? 1'b1 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b1 : 
                   (N244)? 1'b0 : 
                   (N245)? 1'b0 : 
                   (N246)? 1'b0 : 
                   (N247)? 1'b1 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b1 : 
                   (N252)? 1'b0 : 
                   (N253)? 1'b0 : 
                   (N254)? 1'b0 : 
                   (N255)? 1'b1 : 1'b0;
  assign bk_o[6] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b1 : 
                   (N4)? 1'b0 : 
                   (N5)? 1'b1 : 
                   (N6)? 1'b1 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b1 : 
                   (N12)? 1'b0 : 
                   (N13)? 1'b1 : 
                   (N14)? 1'b1 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b1 : 
                   (N20)? 1'b0 : 
                   (N21)? 1'b1 : 
                   (N22)? 1'b1 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b1 : 
                   (N28)? 1'b0 : 
                   (N29)? 1'b1 : 
                   (N30)? 1'b1 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b1 : 
                   (N36)? 1'b0 : 
                   (N37)? 1'b1 : 
                   (N38)? 1'b1 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b1 : 
                   (N44)? 1'b0 : 
                   (N45)? 1'b1 : 
                   (N46)? 1'b1 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b1 : 
                   (N52)? 1'b0 : 
                   (N53)? 1'b1 : 
                   (N54)? 1'b1 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b1 : 
                   (N60)? 1'b0 : 
                   (N61)? 1'b1 : 
                   (N62)? 1'b1 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b1 : 
                   (N68)? 1'b0 : 
                   (N69)? 1'b1 : 
                   (N70)? 1'b1 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b1 : 
                   (N76)? 1'b0 : 
                   (N77)? 1'b1 : 
                   (N78)? 1'b1 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b1 : 
                   (N84)? 1'b0 : 
                   (N85)? 1'b1 : 
                   (N86)? 1'b1 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b1 : 
                   (N92)? 1'b0 : 
                   (N93)? 1'b1 : 
                   (N94)? 1'b1 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b1 : 
                   (N100)? 1'b0 : 
                   (N101)? 1'b1 : 
                   (N102)? 1'b1 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b1 : 
                   (N108)? 1'b0 : 
                   (N109)? 1'b1 : 
                   (N110)? 1'b1 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b1 : 
                   (N116)? 1'b0 : 
                   (N117)? 1'b1 : 
                   (N118)? 1'b1 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b1 : 
                   (N124)? 1'b0 : 
                   (N125)? 1'b1 : 
                   (N126)? 1'b1 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b1 : 
                   (N132)? 1'b0 : 
                   (N133)? 1'b1 : 
                   (N134)? 1'b1 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b1 : 
                   (N140)? 1'b0 : 
                   (N141)? 1'b1 : 
                   (N142)? 1'b1 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b1 : 
                   (N148)? 1'b0 : 
                   (N149)? 1'b1 : 
                   (N150)? 1'b1 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b1 : 
                   (N156)? 1'b0 : 
                   (N157)? 1'b1 : 
                   (N158)? 1'b1 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b1 : 
                   (N164)? 1'b0 : 
                   (N165)? 1'b1 : 
                   (N166)? 1'b1 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b1 : 
                   (N172)? 1'b0 : 
                   (N173)? 1'b1 : 
                   (N174)? 1'b1 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b1 : 
                   (N180)? 1'b0 : 
                   (N181)? 1'b1 : 
                   (N182)? 1'b1 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b1 : 
                   (N188)? 1'b0 : 
                   (N189)? 1'b1 : 
                   (N190)? 1'b1 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b1 : 
                   (N196)? 1'b0 : 
                   (N197)? 1'b1 : 
                   (N198)? 1'b1 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b1 : 
                   (N204)? 1'b0 : 
                   (N205)? 1'b1 : 
                   (N206)? 1'b1 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b1 : 
                   (N212)? 1'b0 : 
                   (N213)? 1'b1 : 
                   (N214)? 1'b1 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b1 : 
                   (N220)? 1'b0 : 
                   (N221)? 1'b1 : 
                   (N222)? 1'b1 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b1 : 
                   (N228)? 1'b0 : 
                   (N229)? 1'b1 : 
                   (N230)? 1'b1 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b1 : 
                   (N236)? 1'b0 : 
                   (N237)? 1'b1 : 
                   (N238)? 1'b1 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b1 : 
                   (N244)? 1'b0 : 
                   (N245)? 1'b1 : 
                   (N246)? 1'b1 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b1 : 
                   (N252)? 1'b0 : 
                   (N253)? 1'b1 : 
                   (N254)? 1'b1 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_o[5] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b1 : 
                   (N6)? 1'b0 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b0 : 
                   (N11)? 1'b0 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b1 : 
                   (N14)? 1'b0 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b0 : 
                   (N19)? 1'b0 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b1 : 
                   (N22)? 1'b0 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b0 : 
                   (N27)? 1'b0 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b1 : 
                   (N30)? 1'b0 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b0 : 
                   (N35)? 1'b0 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b1 : 
                   (N38)? 1'b0 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b0 : 
                   (N43)? 1'b0 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b1 : 
                   (N46)? 1'b0 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b0 : 
                   (N51)? 1'b0 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b1 : 
                   (N54)? 1'b0 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b0 : 
                   (N59)? 1'b0 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b1 : 
                   (N62)? 1'b0 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b0 : 
                   (N67)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b1 : 
                   (N70)? 1'b0 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b0 : 
                   (N75)? 1'b0 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b1 : 
                   (N78)? 1'b0 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b0 : 
                   (N83)? 1'b0 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b1 : 
                   (N86)? 1'b0 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b0 : 
                   (N91)? 1'b0 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b1 : 
                   (N94)? 1'b0 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b0 : 
                   (N99)? 1'b0 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b1 : 
                   (N102)? 1'b0 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b0 : 
                   (N107)? 1'b0 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b1 : 
                   (N110)? 1'b0 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b0 : 
                   (N115)? 1'b0 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b1 : 
                   (N118)? 1'b0 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b0 : 
                   (N123)? 1'b0 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b1 : 
                   (N126)? 1'b0 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b0 : 
                   (N131)? 1'b0 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b1 : 
                   (N134)? 1'b0 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b0 : 
                   (N139)? 1'b0 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b1 : 
                   (N142)? 1'b0 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b0 : 
                   (N147)? 1'b0 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b1 : 
                   (N150)? 1'b0 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b0 : 
                   (N155)? 1'b0 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b1 : 
                   (N158)? 1'b0 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b0 : 
                   (N163)? 1'b0 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b1 : 
                   (N166)? 1'b0 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b0 : 
                   (N171)? 1'b0 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b1 : 
                   (N174)? 1'b0 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b0 : 
                   (N179)? 1'b0 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b1 : 
                   (N182)? 1'b0 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b0 : 
                   (N187)? 1'b0 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b1 : 
                   (N190)? 1'b0 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b0 : 
                   (N195)? 1'b0 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b1 : 
                   (N198)? 1'b0 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b0 : 
                   (N203)? 1'b0 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b1 : 
                   (N206)? 1'b0 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b0 : 
                   (N211)? 1'b0 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b1 : 
                   (N214)? 1'b0 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b0 : 
                   (N219)? 1'b0 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b1 : 
                   (N222)? 1'b0 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b0 : 
                   (N227)? 1'b0 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b1 : 
                   (N230)? 1'b0 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b0 : 
                   (N235)? 1'b0 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b1 : 
                   (N238)? 1'b0 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b0 : 
                   (N243)? 1'b0 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b1 : 
                   (N246)? 1'b0 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b0 : 
                   (N251)? 1'b0 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b1 : 
                   (N254)? 1'b0 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_o[4] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b1 : 
                   (N6)? 1'b0 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b0 : 
                   (N11)? 1'b0 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b1 : 
                   (N14)? 1'b0 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b0 : 
                   (N19)? 1'b0 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b1 : 
                   (N22)? 1'b0 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b0 : 
                   (N27)? 1'b0 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b1 : 
                   (N30)? 1'b0 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b0 : 
                   (N35)? 1'b0 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b1 : 
                   (N38)? 1'b0 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b0 : 
                   (N43)? 1'b0 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b1 : 
                   (N46)? 1'b0 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b0 : 
                   (N51)? 1'b0 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b1 : 
                   (N54)? 1'b0 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b0 : 
                   (N59)? 1'b0 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b1 : 
                   (N62)? 1'b0 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b0 : 
                   (N67)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b1 : 
                   (N70)? 1'b0 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b0 : 
                   (N75)? 1'b0 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b1 : 
                   (N78)? 1'b0 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b0 : 
                   (N83)? 1'b0 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b1 : 
                   (N86)? 1'b0 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b0 : 
                   (N91)? 1'b0 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b1 : 
                   (N94)? 1'b0 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b0 : 
                   (N99)? 1'b0 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b1 : 
                   (N102)? 1'b0 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b0 : 
                   (N107)? 1'b0 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b1 : 
                   (N110)? 1'b0 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b0 : 
                   (N115)? 1'b0 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b1 : 
                   (N118)? 1'b0 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b0 : 
                   (N123)? 1'b0 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b1 : 
                   (N126)? 1'b0 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b0 : 
                   (N131)? 1'b0 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b1 : 
                   (N134)? 1'b0 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b0 : 
                   (N139)? 1'b0 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b1 : 
                   (N142)? 1'b0 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b0 : 
                   (N147)? 1'b0 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b1 : 
                   (N150)? 1'b0 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b0 : 
                   (N155)? 1'b0 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b1 : 
                   (N158)? 1'b0 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b0 : 
                   (N163)? 1'b0 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b1 : 
                   (N166)? 1'b0 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b0 : 
                   (N171)? 1'b0 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b1 : 
                   (N174)? 1'b0 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b0 : 
                   (N179)? 1'b0 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b1 : 
                   (N182)? 1'b0 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b0 : 
                   (N187)? 1'b0 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b1 : 
                   (N190)? 1'b0 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b0 : 
                   (N195)? 1'b0 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b1 : 
                   (N198)? 1'b0 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b0 : 
                   (N203)? 1'b0 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b1 : 
                   (N206)? 1'b0 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b0 : 
                   (N211)? 1'b0 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b1 : 
                   (N214)? 1'b0 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b0 : 
                   (N219)? 1'b0 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b1 : 
                   (N222)? 1'b0 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b0 : 
                   (N227)? 1'b0 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b1 : 
                   (N230)? 1'b0 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b0 : 
                   (N235)? 1'b0 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b1 : 
                   (N238)? 1'b0 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b0 : 
                   (N243)? 1'b0 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b1 : 
                   (N246)? 1'b0 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b0 : 
                   (N251)? 1'b0 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b1 : 
                   (N254)? 1'b0 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_o[3] = (N0)? 1'b1 : 
                   (N1)? 1'b1 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b1 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b1 : 
                   (N6)? 1'b0 : 
                   (N7)? 1'b1 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b1 : 
                   (N10)? 1'b0 : 
                   (N11)? 1'b1 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b1 : 
                   (N14)? 1'b0 : 
                   (N15)? 1'b1 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b1 : 
                   (N18)? 1'b0 : 
                   (N19)? 1'b1 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b1 : 
                   (N22)? 1'b0 : 
                   (N23)? 1'b1 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b1 : 
                   (N26)? 1'b0 : 
                   (N27)? 1'b1 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b1 : 
                   (N30)? 1'b0 : 
                   (N31)? 1'b1 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b1 : 
                   (N34)? 1'b0 : 
                   (N35)? 1'b1 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b1 : 
                   (N38)? 1'b0 : 
                   (N39)? 1'b1 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b1 : 
                   (N42)? 1'b0 : 
                   (N43)? 1'b1 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b1 : 
                   (N46)? 1'b0 : 
                   (N47)? 1'b1 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b1 : 
                   (N50)? 1'b0 : 
                   (N51)? 1'b1 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b1 : 
                   (N54)? 1'b0 : 
                   (N55)? 1'b1 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b1 : 
                   (N58)? 1'b0 : 
                   (N59)? 1'b1 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b1 : 
                   (N62)? 1'b0 : 
                   (N63)? 1'b1 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b1 : 
                   (N66)? 1'b0 : 
                   (N67)? 1'b1 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b1 : 
                   (N70)? 1'b0 : 
                   (N71)? 1'b1 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b1 : 
                   (N74)? 1'b0 : 
                   (N75)? 1'b1 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b1 : 
                   (N78)? 1'b0 : 
                   (N79)? 1'b1 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b1 : 
                   (N82)? 1'b0 : 
                   (N83)? 1'b1 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b1 : 
                   (N86)? 1'b0 : 
                   (N87)? 1'b1 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b1 : 
                   (N90)? 1'b0 : 
                   (N91)? 1'b1 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b1 : 
                   (N94)? 1'b0 : 
                   (N95)? 1'b1 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b1 : 
                   (N98)? 1'b0 : 
                   (N99)? 1'b1 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b1 : 
                   (N102)? 1'b0 : 
                   (N103)? 1'b1 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b1 : 
                   (N106)? 1'b0 : 
                   (N107)? 1'b1 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b1 : 
                   (N110)? 1'b0 : 
                   (N111)? 1'b1 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b1 : 
                   (N114)? 1'b0 : 
                   (N115)? 1'b1 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b1 : 
                   (N118)? 1'b0 : 
                   (N119)? 1'b1 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b1 : 
                   (N122)? 1'b0 : 
                   (N123)? 1'b1 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b1 : 
                   (N126)? 1'b0 : 
                   (N127)? 1'b1 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b1 : 
                   (N130)? 1'b0 : 
                   (N131)? 1'b1 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b1 : 
                   (N134)? 1'b0 : 
                   (N135)? 1'b1 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b1 : 
                   (N138)? 1'b0 : 
                   (N139)? 1'b1 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b1 : 
                   (N142)? 1'b0 : 
                   (N143)? 1'b1 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b1 : 
                   (N146)? 1'b0 : 
                   (N147)? 1'b1 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b1 : 
                   (N150)? 1'b0 : 
                   (N151)? 1'b1 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b1 : 
                   (N154)? 1'b0 : 
                   (N155)? 1'b1 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b1 : 
                   (N158)? 1'b0 : 
                   (N159)? 1'b1 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b1 : 
                   (N162)? 1'b0 : 
                   (N163)? 1'b1 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b1 : 
                   (N166)? 1'b0 : 
                   (N167)? 1'b1 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b1 : 
                   (N170)? 1'b0 : 
                   (N171)? 1'b1 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b1 : 
                   (N174)? 1'b0 : 
                   (N175)? 1'b1 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b1 : 
                   (N178)? 1'b0 : 
                   (N179)? 1'b1 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b1 : 
                   (N182)? 1'b0 : 
                   (N183)? 1'b1 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b1 : 
                   (N186)? 1'b0 : 
                   (N187)? 1'b1 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b1 : 
                   (N190)? 1'b0 : 
                   (N191)? 1'b1 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b1 : 
                   (N194)? 1'b0 : 
                   (N195)? 1'b1 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b1 : 
                   (N198)? 1'b0 : 
                   (N199)? 1'b1 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b1 : 
                   (N202)? 1'b0 : 
                   (N203)? 1'b1 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b1 : 
                   (N206)? 1'b0 : 
                   (N207)? 1'b1 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b1 : 
                   (N210)? 1'b0 : 
                   (N211)? 1'b1 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b1 : 
                   (N214)? 1'b0 : 
                   (N215)? 1'b1 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b1 : 
                   (N218)? 1'b0 : 
                   (N219)? 1'b1 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b1 : 
                   (N222)? 1'b0 : 
                   (N223)? 1'b1 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b1 : 
                   (N226)? 1'b0 : 
                   (N227)? 1'b1 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b1 : 
                   (N230)? 1'b0 : 
                   (N231)? 1'b1 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b1 : 
                   (N234)? 1'b0 : 
                   (N235)? 1'b1 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b1 : 
                   (N238)? 1'b0 : 
                   (N239)? 1'b1 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b1 : 
                   (N242)? 1'b0 : 
                   (N243)? 1'b1 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b1 : 
                   (N246)? 1'b0 : 
                   (N247)? 1'b1 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b1 : 
                   (N250)? 1'b0 : 
                   (N251)? 1'b1 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b1 : 
                   (N254)? 1'b0 : 
                   (N255)? 1'b1 : 1'b0;
  assign bk_o[2] = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b0 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b1 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b0 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b0 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b0 : 
                   (N14)? 1'b1 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b0 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b0 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b0 : 
                   (N22)? 1'b1 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b0 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b0 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b0 : 
                   (N30)? 1'b1 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b0 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b0 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b0 : 
                   (N38)? 1'b1 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b0 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b0 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b0 : 
                   (N46)? 1'b1 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b0 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b0 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b0 : 
                   (N54)? 1'b1 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b0 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b0 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b0 : 
                   (N62)? 1'b1 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b0 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b0 : 
                   (N70)? 1'b1 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b0 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b0 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b0 : 
                   (N78)? 1'b1 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b0 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b0 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b0 : 
                   (N86)? 1'b1 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b0 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b0 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b0 : 
                   (N94)? 1'b1 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b0 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b0 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b0 : 
                   (N102)? 1'b1 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b0 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b0 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b0 : 
                   (N110)? 1'b1 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b0 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b0 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b0 : 
                   (N118)? 1'b1 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b0 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b0 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b0 : 
                   (N126)? 1'b1 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b0 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b0 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b0 : 
                   (N134)? 1'b1 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b0 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b0 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b0 : 
                   (N142)? 1'b1 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b0 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b0 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b0 : 
                   (N150)? 1'b1 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b0 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b0 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b0 : 
                   (N158)? 1'b1 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b0 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b0 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b0 : 
                   (N166)? 1'b1 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b0 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b0 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b0 : 
                   (N174)? 1'b1 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b0 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b0 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b0 : 
                   (N182)? 1'b1 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b0 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b0 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b0 : 
                   (N190)? 1'b1 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b0 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b0 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b0 : 
                   (N198)? 1'b1 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b0 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b0 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b0 : 
                   (N206)? 1'b1 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b0 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b0 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b0 : 
                   (N214)? 1'b1 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b0 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b0 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b0 : 
                   (N222)? 1'b1 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b0 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b0 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b0 : 
                   (N230)? 1'b1 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b0 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b0 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b0 : 
                   (N238)? 1'b1 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b0 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b0 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b0 : 
                   (N246)? 1'b1 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b0 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b0 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b0 : 
                   (N254)? 1'b1 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_o[1] = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b0 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b1 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b0 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b0 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b0 : 
                   (N14)? 1'b1 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b0 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b0 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b0 : 
                   (N22)? 1'b1 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b0 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b0 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b0 : 
                   (N30)? 1'b1 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b0 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b0 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b0 : 
                   (N38)? 1'b1 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b0 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b0 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b0 : 
                   (N46)? 1'b1 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b0 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b0 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b0 : 
                   (N54)? 1'b1 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b0 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b0 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b0 : 
                   (N62)? 1'b1 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b0 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b0 : 
                   (N70)? 1'b1 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b0 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b0 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b0 : 
                   (N78)? 1'b1 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b0 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b0 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b0 : 
                   (N86)? 1'b1 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b0 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b0 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b0 : 
                   (N94)? 1'b1 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b0 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b0 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b0 : 
                   (N102)? 1'b1 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b0 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b0 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b0 : 
                   (N110)? 1'b1 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b0 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b0 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b0 : 
                   (N118)? 1'b1 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b0 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b0 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b0 : 
                   (N126)? 1'b1 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b0 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b0 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b0 : 
                   (N134)? 1'b1 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b0 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b0 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b0 : 
                   (N142)? 1'b1 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b0 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b0 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b0 : 
                   (N150)? 1'b1 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b0 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b0 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b0 : 
                   (N158)? 1'b1 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b0 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b0 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b0 : 
                   (N166)? 1'b1 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b0 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b0 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b0 : 
                   (N174)? 1'b1 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b0 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b0 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b0 : 
                   (N182)? 1'b1 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b0 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b0 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b0 : 
                   (N190)? 1'b1 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b0 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b0 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b0 : 
                   (N198)? 1'b1 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b0 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b0 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b0 : 
                   (N206)? 1'b1 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b0 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b0 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b0 : 
                   (N214)? 1'b1 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b0 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b0 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b0 : 
                   (N222)? 1'b1 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b0 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b0 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b0 : 
                   (N230)? 1'b1 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b0 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b0 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b0 : 
                   (N238)? 1'b1 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b0 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b0 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b0 : 
                   (N246)? 1'b1 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b0 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b0 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b0 : 
                   (N254)? 1'b1 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_o[0] = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b1 : 
                   (N3)? 1'b0 : 
                   (N4)? 1'b1 : 
                   (N5)? 1'b0 : 
                   (N6)? 1'b1 : 
                   (N7)? 1'b0 : 
                   (N8)? 1'b1 : 
                   (N9)? 1'b0 : 
                   (N10)? 1'b1 : 
                   (N11)? 1'b0 : 
                   (N12)? 1'b1 : 
                   (N13)? 1'b0 : 
                   (N14)? 1'b1 : 
                   (N15)? 1'b0 : 
                   (N16)? 1'b1 : 
                   (N17)? 1'b0 : 
                   (N18)? 1'b1 : 
                   (N19)? 1'b0 : 
                   (N20)? 1'b1 : 
                   (N21)? 1'b0 : 
                   (N22)? 1'b1 : 
                   (N23)? 1'b0 : 
                   (N24)? 1'b1 : 
                   (N25)? 1'b0 : 
                   (N26)? 1'b1 : 
                   (N27)? 1'b0 : 
                   (N28)? 1'b1 : 
                   (N29)? 1'b0 : 
                   (N30)? 1'b1 : 
                   (N31)? 1'b0 : 
                   (N32)? 1'b1 : 
                   (N33)? 1'b0 : 
                   (N34)? 1'b1 : 
                   (N35)? 1'b0 : 
                   (N36)? 1'b1 : 
                   (N37)? 1'b0 : 
                   (N38)? 1'b1 : 
                   (N39)? 1'b0 : 
                   (N40)? 1'b1 : 
                   (N41)? 1'b0 : 
                   (N42)? 1'b1 : 
                   (N43)? 1'b0 : 
                   (N44)? 1'b1 : 
                   (N45)? 1'b0 : 
                   (N46)? 1'b1 : 
                   (N47)? 1'b0 : 
                   (N48)? 1'b1 : 
                   (N49)? 1'b0 : 
                   (N50)? 1'b1 : 
                   (N51)? 1'b0 : 
                   (N52)? 1'b1 : 
                   (N53)? 1'b0 : 
                   (N54)? 1'b1 : 
                   (N55)? 1'b0 : 
                   (N56)? 1'b1 : 
                   (N57)? 1'b0 : 
                   (N58)? 1'b1 : 
                   (N59)? 1'b0 : 
                   (N60)? 1'b1 : 
                   (N61)? 1'b0 : 
                   (N62)? 1'b1 : 
                   (N63)? 1'b0 : 
                   (N64)? 1'b1 : 
                   (N65)? 1'b0 : 
                   (N66)? 1'b1 : 
                   (N67)? 1'b0 : 
                   (N68)? 1'b1 : 
                   (N69)? 1'b0 : 
                   (N70)? 1'b1 : 
                   (N71)? 1'b0 : 
                   (N72)? 1'b1 : 
                   (N73)? 1'b0 : 
                   (N74)? 1'b1 : 
                   (N75)? 1'b0 : 
                   (N76)? 1'b1 : 
                   (N77)? 1'b0 : 
                   (N78)? 1'b1 : 
                   (N79)? 1'b0 : 
                   (N80)? 1'b1 : 
                   (N81)? 1'b0 : 
                   (N82)? 1'b1 : 
                   (N83)? 1'b0 : 
                   (N84)? 1'b1 : 
                   (N85)? 1'b0 : 
                   (N86)? 1'b1 : 
                   (N87)? 1'b0 : 
                   (N88)? 1'b1 : 
                   (N89)? 1'b0 : 
                   (N90)? 1'b1 : 
                   (N91)? 1'b0 : 
                   (N92)? 1'b1 : 
                   (N93)? 1'b0 : 
                   (N94)? 1'b1 : 
                   (N95)? 1'b0 : 
                   (N96)? 1'b1 : 
                   (N97)? 1'b0 : 
                   (N98)? 1'b1 : 
                   (N99)? 1'b0 : 
                   (N100)? 1'b1 : 
                   (N101)? 1'b0 : 
                   (N102)? 1'b1 : 
                   (N103)? 1'b0 : 
                   (N104)? 1'b1 : 
                   (N105)? 1'b0 : 
                   (N106)? 1'b1 : 
                   (N107)? 1'b0 : 
                   (N108)? 1'b1 : 
                   (N109)? 1'b0 : 
                   (N110)? 1'b1 : 
                   (N111)? 1'b0 : 
                   (N112)? 1'b1 : 
                   (N113)? 1'b0 : 
                   (N114)? 1'b1 : 
                   (N115)? 1'b0 : 
                   (N116)? 1'b1 : 
                   (N117)? 1'b0 : 
                   (N118)? 1'b1 : 
                   (N119)? 1'b0 : 
                   (N120)? 1'b1 : 
                   (N121)? 1'b0 : 
                   (N122)? 1'b1 : 
                   (N123)? 1'b0 : 
                   (N124)? 1'b1 : 
                   (N125)? 1'b0 : 
                   (N126)? 1'b1 : 
                   (N127)? 1'b0 : 
                   (N128)? 1'b1 : 
                   (N129)? 1'b0 : 
                   (N130)? 1'b1 : 
                   (N131)? 1'b0 : 
                   (N132)? 1'b1 : 
                   (N133)? 1'b0 : 
                   (N134)? 1'b1 : 
                   (N135)? 1'b0 : 
                   (N136)? 1'b1 : 
                   (N137)? 1'b0 : 
                   (N138)? 1'b1 : 
                   (N139)? 1'b0 : 
                   (N140)? 1'b1 : 
                   (N141)? 1'b0 : 
                   (N142)? 1'b1 : 
                   (N143)? 1'b0 : 
                   (N144)? 1'b1 : 
                   (N145)? 1'b0 : 
                   (N146)? 1'b1 : 
                   (N147)? 1'b0 : 
                   (N148)? 1'b1 : 
                   (N149)? 1'b0 : 
                   (N150)? 1'b1 : 
                   (N151)? 1'b0 : 
                   (N152)? 1'b1 : 
                   (N153)? 1'b0 : 
                   (N154)? 1'b1 : 
                   (N155)? 1'b0 : 
                   (N156)? 1'b1 : 
                   (N157)? 1'b0 : 
                   (N158)? 1'b1 : 
                   (N159)? 1'b0 : 
                   (N160)? 1'b1 : 
                   (N161)? 1'b0 : 
                   (N162)? 1'b1 : 
                   (N163)? 1'b0 : 
                   (N164)? 1'b1 : 
                   (N165)? 1'b0 : 
                   (N166)? 1'b1 : 
                   (N167)? 1'b0 : 
                   (N168)? 1'b1 : 
                   (N169)? 1'b0 : 
                   (N170)? 1'b1 : 
                   (N171)? 1'b0 : 
                   (N172)? 1'b1 : 
                   (N173)? 1'b0 : 
                   (N174)? 1'b1 : 
                   (N175)? 1'b0 : 
                   (N176)? 1'b1 : 
                   (N177)? 1'b0 : 
                   (N178)? 1'b1 : 
                   (N179)? 1'b0 : 
                   (N180)? 1'b1 : 
                   (N181)? 1'b0 : 
                   (N182)? 1'b1 : 
                   (N183)? 1'b0 : 
                   (N184)? 1'b1 : 
                   (N185)? 1'b0 : 
                   (N186)? 1'b1 : 
                   (N187)? 1'b0 : 
                   (N188)? 1'b1 : 
                   (N189)? 1'b0 : 
                   (N190)? 1'b1 : 
                   (N191)? 1'b0 : 
                   (N192)? 1'b1 : 
                   (N193)? 1'b0 : 
                   (N194)? 1'b1 : 
                   (N195)? 1'b0 : 
                   (N196)? 1'b1 : 
                   (N197)? 1'b0 : 
                   (N198)? 1'b1 : 
                   (N199)? 1'b0 : 
                   (N200)? 1'b1 : 
                   (N201)? 1'b0 : 
                   (N202)? 1'b1 : 
                   (N203)? 1'b0 : 
                   (N204)? 1'b1 : 
                   (N205)? 1'b0 : 
                   (N206)? 1'b1 : 
                   (N207)? 1'b0 : 
                   (N208)? 1'b1 : 
                   (N209)? 1'b0 : 
                   (N210)? 1'b1 : 
                   (N211)? 1'b0 : 
                   (N212)? 1'b1 : 
                   (N213)? 1'b0 : 
                   (N214)? 1'b1 : 
                   (N215)? 1'b0 : 
                   (N216)? 1'b1 : 
                   (N217)? 1'b0 : 
                   (N218)? 1'b1 : 
                   (N219)? 1'b0 : 
                   (N220)? 1'b1 : 
                   (N221)? 1'b0 : 
                   (N222)? 1'b1 : 
                   (N223)? 1'b0 : 
                   (N224)? 1'b1 : 
                   (N225)? 1'b0 : 
                   (N226)? 1'b1 : 
                   (N227)? 1'b0 : 
                   (N228)? 1'b1 : 
                   (N229)? 1'b0 : 
                   (N230)? 1'b1 : 
                   (N231)? 1'b0 : 
                   (N232)? 1'b1 : 
                   (N233)? 1'b0 : 
                   (N234)? 1'b1 : 
                   (N235)? 1'b0 : 
                   (N236)? 1'b1 : 
                   (N237)? 1'b0 : 
                   (N238)? 1'b1 : 
                   (N239)? 1'b0 : 
                   (N240)? 1'b1 : 
                   (N241)? 1'b0 : 
                   (N242)? 1'b1 : 
                   (N243)? 1'b0 : 
                   (N244)? 1'b1 : 
                   (N245)? 1'b0 : 
                   (N246)? 1'b1 : 
                   (N247)? 1'b0 : 
                   (N248)? 1'b1 : 
                   (N249)? 1'b0 : 
                   (N250)? 1'b1 : 
                   (N251)? 1'b0 : 
                   (N252)? 1'b1 : 
                   (N253)? 1'b0 : 
                   (N254)? 1'b1 : 
                   (N255)? 1'b0 : 1'b0;
  assign bk_datapath_o[23] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b0 : 
                             (N370)? 1'b0 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b0 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b0 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b0 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b0 : 
                             (N382)? 1'b0 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b1 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b1 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b1 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b1 : 
                             (N414)? 1'b1 : 
                             (N415)? 1'b1 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b1 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b1 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b1 : 
                             (N430)? 1'b1 : 
                             (N431)? 1'b1 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b0 : 
                             (N434)? 1'b0 : 
                             (N435)? 1'b1 : 
                             (N436)? 1'b0 : 
                             (N437)? 1'b1 : 
                             (N438)? 1'b1 : 
                             (N439)? 1'b1 : 
                             (N440)? 1'b0 : 
                             (N441)? 1'b1 : 
                             (N442)? 1'b1 : 
                             (N443)? 1'b1 : 
                             (N444)? 1'b1 : 
                             (N445)? 1'b1 : 
                             (N446)? 1'b1 : 
                             (N447)? 1'b1 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b1 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b1 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b1 : 
                             (N462)? 1'b1 : 
                             (N463)? 1'b1 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b0 : 
                             (N466)? 1'b0 : 
                             (N467)? 1'b1 : 
                             (N468)? 1'b0 : 
                             (N469)? 1'b1 : 
                             (N470)? 1'b1 : 
                             (N471)? 1'b1 : 
                             (N472)? 1'b0 : 
                             (N473)? 1'b1 : 
                             (N474)? 1'b1 : 
                             (N475)? 1'b1 : 
                             (N476)? 1'b1 : 
                             (N477)? 1'b1 : 
                             (N478)? 1'b1 : 
                             (N479)? 1'b1 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b0 : 
                             (N482)? 1'b0 : 
                             (N483)? 1'b1 : 
                             (N484)? 1'b0 : 
                             (N485)? 1'b1 : 
                             (N486)? 1'b1 : 
                             (N487)? 1'b1 : 
                             (N488)? 1'b0 : 
                             (N489)? 1'b1 : 
                             (N490)? 1'b1 : 
                             (N491)? 1'b1 : 
                             (N492)? 1'b1 : 
                             (N493)? 1'b1 : 
                             (N494)? 1'b1 : 
                             (N495)? 1'b1 : 
                             (N496)? 1'b0 : 
                             (N497)? 1'b1 : 
                             (N498)? 1'b1 : 
                             (N499)? 1'b1 : 
                             (N500)? 1'b1 : 
                             (N501)? 1'b1 : 
                             (N502)? 1'b1 : 
                             (N503)? 1'b1 : 
                             (N504)? 1'b1 : 
                             (N505)? 1'b1 : 
                             (N506)? 1'b1 : 
                             (N507)? 1'b1 : 
                             (N508)? 1'b1 : 
                             (N509)? 1'b1 : 
                             (N510)? 1'b1 : 
                             (N255)? 1'b1 : 1'b0;
  assign N256 = N1718;
  assign N257 = N1720;
  assign N258 = N1722;
  assign N259 = N1724;
  assign N260 = N1726;
  assign N261 = N1728;
  assign N262 = N1730;
  assign N263 = N1732;
  assign N264 = N1734;
  assign N265 = N1736;
  assign N266 = N1738;
  assign N267 = N1740;
  assign N268 = N1742;
  assign N269 = N1744;
  assign N270 = N1746;
  assign N271 = N1748;
  assign N272 = N1750;
  assign N273 = N1752;
  assign N274 = N1754;
  assign N275 = N1756;
  assign N276 = N1758;
  assign N277 = N1760;
  assign N278 = N1762;
  assign N279 = N1764;
  assign N280 = N1766;
  assign N281 = N1768;
  assign N282 = N1770;
  assign N283 = N1772;
  assign N284 = N1774;
  assign N285 = N1776;
  assign N286 = N1778;
  assign N287 = N1781;
  assign N288 = N1783;
  assign N289 = N1785;
  assign N290 = N1787;
  assign N291 = N1789;
  assign N292 = N1791;
  assign N293 = N1793;
  assign N294 = N1795;
  assign N295 = N1798;
  assign N296 = N1800;
  assign N297 = N1802;
  assign N298 = N1804;
  assign N299 = N1806;
  assign N300 = N1808;
  assign N301 = N1810;
  assign N302 = N1812;
  assign N303 = N1814;
  assign N304 = N1816;
  assign N305 = N1818;
  assign N306 = N1820;
  assign N307 = N1822;
  assign N308 = N1824;
  assign N309 = N1826;
  assign N310 = N1828;
  assign N311 = N1830;
  assign N312 = N1832;
  assign N313 = N1834;
  assign N314 = N1836;
  assign N315 = N1838;
  assign N316 = N1840;
  assign N317 = N1842;
  assign N318 = N1844;
  assign N319 = N1847;
  assign N320 = N1849;
  assign N321 = N1851;
  assign N322 = N1853;
  assign N323 = N1855;
  assign N324 = N1857;
  assign N325 = N1859;
  assign N326 = N1861;
  assign N327 = N1864;
  assign N328 = N1866;
  assign N329 = N1868;
  assign N330 = N1870;
  assign N331 = N1872;
  assign N332 = N1874;
  assign N333 = N1876;
  assign N334 = N1878;
  assign N335 = N1880;
  assign N336 = N1882;
  assign N337 = N1884;
  assign N338 = N1886;
  assign N339 = N1888;
  assign N340 = N1890;
  assign N341 = N1892;
  assign N342 = N1894;
  assign N343 = N1896;
  assign N344 = N1898;
  assign N345 = N1900;
  assign N346 = N1902;
  assign N347 = N1904;
  assign N348 = N1906;
  assign N349 = N1908;
  assign N350 = N1910;
  assign N351 = N1913;
  assign N352 = N1915;
  assign N353 = N1917;
  assign N354 = N1919;
  assign N355 = N1921;
  assign N356 = N1923;
  assign N357 = N1925;
  assign N358 = N1927;
  assign N359 = N1930;
  assign N360 = N1932;
  assign N361 = N1934;
  assign N362 = N1936;
  assign N363 = N1938;
  assign N364 = N1940;
  assign N365 = N1942;
  assign N366 = N1944;
  assign N367 = N1946;
  assign N368 = N1948;
  assign N369 = N1950;
  assign N370 = N1952;
  assign N371 = N1954;
  assign N372 = N1956;
  assign N373 = N1958;
  assign N374 = N1960;
  assign N375 = N1962;
  assign N376 = N1964;
  assign N377 = N1966;
  assign N378 = N1968;
  assign N379 = N1970;
  assign N380 = N1972;
  assign N381 = N1974;
  assign N382 = N1976;
  assign N383 = N1979;
  assign N384 = N1981;
  assign N385 = N1983;
  assign N386 = N1985;
  assign N387 = N1987;
  assign N388 = N1989;
  assign N389 = N1991;
  assign N390 = N1993;
  assign N391 = N1996;
  assign N392 = N1998;
  assign N393 = N2000;
  assign N394 = N2002;
  assign N395 = N2004;
  assign N396 = N2006;
  assign N397 = N2008;
  assign N398 = N2010;
  assign N399 = N2012;
  assign N400 = N2014;
  assign N401 = N2016;
  assign N402 = N2018;
  assign N403 = N2020;
  assign N404 = N2022;
  assign N405 = N2024;
  assign N406 = N2026;
  assign N407 = N2028;
  assign N408 = N2030;
  assign N409 = N2032;
  assign N410 = N2034;
  assign N411 = N2036;
  assign N412 = N2038;
  assign N413 = N2040;
  assign N414 = N2042;
  assign N415 = N2045;
  assign N416 = N2047;
  assign N417 = N2049;
  assign N418 = N2051;
  assign N419 = N2053;
  assign N420 = N2055;
  assign N421 = N2057;
  assign N422 = N2059;
  assign N423 = N2062;
  assign N424 = N2064;
  assign N425 = N2066;
  assign N426 = N2068;
  assign N427 = N2070;
  assign N428 = N2072;
  assign N429 = N2075;
  assign N430 = N2077;
  assign N431 = N2079;
  assign N432 = N2082;
  assign N433 = N2084;
  assign N434 = N2086;
  assign N435 = N2088;
  assign N436 = N2090;
  assign N437 = N2092;
  assign N438 = N2094;
  assign N439 = N2096;
  assign N440 = N2098;
  assign N441 = N2100;
  assign N442 = N2102;
  assign N443 = N2104;
  assign N444 = N2106;
  assign N445 = N2108;
  assign N446 = N2110;
  assign N447 = N2113;
  assign N448 = N2115;
  assign N449 = N2117;
  assign N450 = N2119;
  assign N451 = N2121;
  assign N452 = N2123;
  assign N453 = N2125;
  assign N454 = N2127;
  assign N455 = N2130;
  assign N456 = N2132;
  assign N457 = N2134;
  assign N458 = N2136;
  assign N459 = N2138;
  assign N460 = N2140;
  assign N461 = N2142;
  assign N462 = N2144;
  assign N463 = N2146;
  assign N464 = N2149;
  assign N465 = N2151;
  assign N466 = N2153;
  assign N467 = N2155;
  assign N468 = N2157;
  assign N469 = N2159;
  assign N470 = N2161;
  assign N471 = N2163;
  assign N472 = N2165;
  assign N473 = N2167;
  assign N474 = N2169;
  assign N475 = N2171;
  assign N476 = N2173;
  assign N477 = N2175;
  assign N478 = N2177;
  assign N479 = N2181;
  assign N480 = N2183;
  assign N481 = N2185;
  assign N482 = N2187;
  assign N483 = N2189;
  assign N484 = N2191;
  assign N485 = N2193;
  assign N486 = N2195;
  assign N487 = N2198;
  assign N488 = N2200;
  assign N489 = N2202;
  assign N490 = N2204;
  assign N491 = N2206;
  assign N492 = N2208;
  assign N493 = N2210;
  assign N494 = N2212;
  assign N495 = N2214;
  assign N496 = N2216;
  assign N497 = N2218;
  assign N498 = N2220;
  assign N499 = N2222;
  assign N500 = N2224;
  assign N501 = N2226;
  assign N502 = N2228;
  assign N503 = N2231;
  assign N504 = N2233;
  assign N505 = N2235;
  assign N506 = N2237;
  assign N507 = N2239;
  assign N508 = N2241;
  assign N509 = N2243;
  assign N510 = N2245;
  assign bk_datapath_o[22] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b0 : 
                             (N370)? 1'b0 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b0 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b0 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b0 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b0 : 
                             (N382)? 1'b0 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b1 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b1 : 
                             (N390)? 1'b1 : 
                             (N391)? 1'b1 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b1 : 
                             (N394)? 1'b1 : 
                             (N395)? 1'b1 : 
                             (N396)? 1'b1 : 
                             (N397)? 1'b1 : 
                             (N398)? 1'b1 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b1 : 
                             (N402)? 1'b1 : 
                             (N403)? 1'b1 : 
                             (N404)? 1'b1 : 
                             (N405)? 1'b1 : 
                             (N406)? 1'b1 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b1 : 
                             (N409)? 1'b1 : 
                             (N410)? 1'b1 : 
                             (N411)? 1'b0 : 
                             (N412)? 1'b1 : 
                             (N413)? 1'b0 : 
                             (N414)? 1'b0 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b1 : 
                             (N418)? 1'b1 : 
                             (N419)? 1'b1 : 
                             (N420)? 1'b1 : 
                             (N421)? 1'b1 : 
                             (N422)? 1'b1 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b1 : 
                             (N425)? 1'b1 : 
                             (N426)? 1'b1 : 
                             (N427)? 1'b0 : 
                             (N428)? 1'b1 : 
                             (N429)? 1'b0 : 
                             (N430)? 1'b0 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b1 : 
                             (N433)? 1'b1 : 
                             (N434)? 1'b1 : 
                             (N435)? 1'b0 : 
                             (N436)? 1'b1 : 
                             (N437)? 1'b0 : 
                             (N438)? 1'b0 : 
                             (N439)? 1'b0 : 
                             (N440)? 1'b1 : 
                             (N441)? 1'b0 : 
                             (N442)? 1'b0 : 
                             (N443)? 1'b0 : 
                             (N444)? 1'b0 : 
                             (N445)? 1'b0 : 
                             (N446)? 1'b0 : 
                             (N447)? 1'b1 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b1 : 
                             (N450)? 1'b1 : 
                             (N451)? 1'b1 : 
                             (N452)? 1'b1 : 
                             (N453)? 1'b1 : 
                             (N454)? 1'b1 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b1 : 
                             (N457)? 1'b1 : 
                             (N458)? 1'b1 : 
                             (N459)? 1'b0 : 
                             (N460)? 1'b1 : 
                             (N461)? 1'b0 : 
                             (N462)? 1'b0 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b1 : 
                             (N465)? 1'b1 : 
                             (N466)? 1'b1 : 
                             (N467)? 1'b0 : 
                             (N468)? 1'b1 : 
                             (N469)? 1'b0 : 
                             (N470)? 1'b0 : 
                             (N471)? 1'b0 : 
                             (N472)? 1'b1 : 
                             (N473)? 1'b0 : 
                             (N474)? 1'b0 : 
                             (N475)? 1'b0 : 
                             (N476)? 1'b0 : 
                             (N477)? 1'b0 : 
                             (N478)? 1'b0 : 
                             (N479)? 1'b1 : 
                             (N480)? 1'b1 : 
                             (N481)? 1'b1 : 
                             (N482)? 1'b1 : 
                             (N483)? 1'b0 : 
                             (N484)? 1'b1 : 
                             (N485)? 1'b0 : 
                             (N486)? 1'b0 : 
                             (N487)? 1'b0 : 
                             (N488)? 1'b1 : 
                             (N489)? 1'b0 : 
                             (N490)? 1'b0 : 
                             (N491)? 1'b0 : 
                             (N492)? 1'b0 : 
                             (N493)? 1'b0 : 
                             (N494)? 1'b0 : 
                             (N495)? 1'b1 : 
                             (N496)? 1'b1 : 
                             (N497)? 1'b0 : 
                             (N498)? 1'b0 : 
                             (N499)? 1'b0 : 
                             (N500)? 1'b0 : 
                             (N501)? 1'b0 : 
                             (N502)? 1'b0 : 
                             (N503)? 1'b1 : 
                             (N504)? 1'b0 : 
                             (N505)? 1'b0 : 
                             (N506)? 1'b0 : 
                             (N507)? 1'b1 : 
                             (N508)? 1'b0 : 
                             (N509)? 1'b1 : 
                             (N510)? 1'b1 : 
                             (N255)? 1'b1 : 1'b0;
  assign bk_datapath_o[21] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b0 : 
                             (N370)? 1'b0 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b0 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b0 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b0 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b0 : 
                             (N382)? 1'b0 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b1 : 
                             (N386)? 1'b1 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b1 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b1 : 
                             (N392)? 1'b1 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b1 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b1 : 
                             (N398)? 1'b1 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b1 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b1 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b1 : 
                             (N406)? 1'b1 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b1 : 
                             (N410)? 1'b1 : 
                             (N411)? 1'b0 : 
                             (N412)? 1'b1 : 
                             (N413)? 1'b0 : 
                             (N414)? 1'b0 : 
                             (N415)? 1'b1 : 
                             (N416)? 1'b1 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b1 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b1 : 
                             (N422)? 1'b1 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b1 : 
                             (N426)? 1'b1 : 
                             (N427)? 1'b0 : 
                             (N428)? 1'b1 : 
                             (N429)? 1'b0 : 
                             (N430)? 1'b0 : 
                             (N431)? 1'b1 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b1 : 
                             (N434)? 1'b1 : 
                             (N435)? 1'b0 : 
                             (N436)? 1'b1 : 
                             (N437)? 1'b0 : 
                             (N438)? 1'b0 : 
                             (N439)? 1'b1 : 
                             (N440)? 1'b1 : 
                             (N441)? 1'b0 : 
                             (N442)? 1'b0 : 
                             (N443)? 1'b1 : 
                             (N444)? 1'b0 : 
                             (N445)? 1'b1 : 
                             (N446)? 1'b1 : 
                             (N447)? 1'b0 : 
                             (N448)? 1'b1 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b1 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b1 : 
                             (N454)? 1'b1 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b1 : 
                             (N458)? 1'b1 : 
                             (N459)? 1'b0 : 
                             (N460)? 1'b1 : 
                             (N461)? 1'b0 : 
                             (N462)? 1'b0 : 
                             (N463)? 1'b1 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b1 : 
                             (N466)? 1'b1 : 
                             (N467)? 1'b0 : 
                             (N468)? 1'b1 : 
                             (N469)? 1'b0 : 
                             (N470)? 1'b0 : 
                             (N471)? 1'b1 : 
                             (N472)? 1'b1 : 
                             (N473)? 1'b0 : 
                             (N474)? 1'b0 : 
                             (N475)? 1'b1 : 
                             (N476)? 1'b0 : 
                             (N477)? 1'b1 : 
                             (N478)? 1'b1 : 
                             (N479)? 1'b0 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b1 : 
                             (N482)? 1'b1 : 
                             (N483)? 1'b0 : 
                             (N484)? 1'b1 : 
                             (N485)? 1'b0 : 
                             (N486)? 1'b0 : 
                             (N487)? 1'b1 : 
                             (N488)? 1'b1 : 
                             (N489)? 1'b0 : 
                             (N490)? 1'b0 : 
                             (N491)? 1'b1 : 
                             (N492)? 1'b0 : 
                             (N493)? 1'b1 : 
                             (N494)? 1'b1 : 
                             (N495)? 1'b0 : 
                             (N496)? 1'b1 : 
                             (N497)? 1'b0 : 
                             (N498)? 1'b0 : 
                             (N499)? 1'b1 : 
                             (N500)? 1'b0 : 
                             (N501)? 1'b1 : 
                             (N502)? 1'b1 : 
                             (N503)? 1'b0 : 
                             (N504)? 1'b0 : 
                             (N505)? 1'b1 : 
                             (N506)? 1'b1 : 
                             (N507)? 1'b0 : 
                             (N508)? 1'b1 : 
                             (N509)? 1'b0 : 
                             (N510)? 1'b0 : 
                             (N255)? 1'b1 : 1'b0;
  assign bk_datapath_o[19] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b1 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b1 : 
                             (N326)? 1'b1 : 
                             (N327)? 1'b1 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b1 : 
                             (N330)? 1'b1 : 
                             (N331)? 1'b1 : 
                             (N332)? 1'b1 : 
                             (N333)? 1'b1 : 
                             (N334)? 1'b1 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b1 : 
                             (N338)? 1'b1 : 
                             (N339)? 1'b1 : 
                             (N340)? 1'b1 : 
                             (N341)? 1'b1 : 
                             (N342)? 1'b1 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b1 : 
                             (N345)? 1'b1 : 
                             (N346)? 1'b1 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b1 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b1 : 
                             (N354)? 1'b1 : 
                             (N355)? 1'b1 : 
                             (N356)? 1'b1 : 
                             (N357)? 1'b1 : 
                             (N358)? 1'b1 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b1 : 
                             (N361)? 1'b1 : 
                             (N362)? 1'b1 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b1 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b1 : 
                             (N369)? 1'b1 : 
                             (N370)? 1'b1 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b1 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b1 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b0 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b0 : 
                             (N382)? 1'b0 : 
                             (N383)? 1'b1 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b0 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b0 : 
                             (N414)? 1'b0 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b0 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b0 : 
                             (N430)? 1'b0 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b0 : 
                             (N434)? 1'b0 : 
                             (N435)? 1'b0 : 
                             (N436)? 1'b0 : 
                             (N437)? 1'b0 : 
                             (N438)? 1'b0 : 
                             (N439)? 1'b0 : 
                             (N440)? 1'b0 : 
                             (N441)? 1'b0 : 
                             (N442)? 1'b0 : 
                             (N443)? 1'b0 : 
                             (N444)? 1'b0 : 
                             (N445)? 1'b0 : 
                             (N446)? 1'b0 : 
                             (N447)? 1'b0 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b1 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b1 : 
                             (N454)? 1'b1 : 
                             (N455)? 1'b1 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b1 : 
                             (N458)? 1'b1 : 
                             (N459)? 1'b1 : 
                             (N460)? 1'b1 : 
                             (N461)? 1'b1 : 
                             (N462)? 1'b1 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b1 : 
                             (N466)? 1'b1 : 
                             (N467)? 1'b1 : 
                             (N468)? 1'b1 : 
                             (N469)? 1'b1 : 
                             (N470)? 1'b1 : 
                             (N471)? 1'b0 : 
                             (N472)? 1'b1 : 
                             (N473)? 1'b1 : 
                             (N474)? 1'b1 : 
                             (N475)? 1'b0 : 
                             (N476)? 1'b1 : 
                             (N477)? 1'b0 : 
                             (N478)? 1'b0 : 
                             (N479)? 1'b0 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b1 : 
                             (N482)? 1'b1 : 
                             (N483)? 1'b1 : 
                             (N484)? 1'b1 : 
                             (N485)? 1'b1 : 
                             (N486)? 1'b1 : 
                             (N487)? 1'b0 : 
                             (N488)? 1'b1 : 
                             (N489)? 1'b1 : 
                             (N490)? 1'b1 : 
                             (N491)? 1'b0 : 
                             (N492)? 1'b1 : 
                             (N493)? 1'b0 : 
                             (N494)? 1'b0 : 
                             (N495)? 1'b0 : 
                             (N496)? 1'b1 : 
                             (N497)? 1'b1 : 
                             (N498)? 1'b1 : 
                             (N499)? 1'b0 : 
                             (N500)? 1'b1 : 
                             (N501)? 1'b0 : 
                             (N502)? 1'b0 : 
                             (N503)? 1'b0 : 
                             (N504)? 1'b1 : 
                             (N505)? 1'b0 : 
                             (N506)? 1'b0 : 
                             (N507)? 1'b0 : 
                             (N508)? 1'b0 : 
                             (N509)? 1'b0 : 
                             (N510)? 1'b0 : 
                             (N255)? 1'b1 : 1'b0;
  assign bk_datapath_o[18] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b1 : 
                             (N322)? 1'b1 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b1 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b1 : 
                             (N328)? 1'b1 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b1 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b1 : 
                             (N334)? 1'b1 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b1 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b1 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b1 : 
                             (N342)? 1'b1 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b1 : 
                             (N346)? 1'b1 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b1 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b1 : 
                             (N352)? 1'b1 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b1 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b1 : 
                             (N358)? 1'b1 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b1 : 
                             (N362)? 1'b1 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b1 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b1 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b1 : 
                             (N370)? 1'b1 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b1 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b1 : 
                             (N376)? 1'b1 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b1 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b1 : 
                             (N382)? 1'b1 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b0 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b0 : 
                             (N414)? 1'b0 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b0 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b0 : 
                             (N430)? 1'b0 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b0 : 
                             (N434)? 1'b0 : 
                             (N435)? 1'b0 : 
                             (N436)? 1'b0 : 
                             (N437)? 1'b0 : 
                             (N438)? 1'b0 : 
                             (N439)? 1'b0 : 
                             (N440)? 1'b0 : 
                             (N441)? 1'b0 : 
                             (N442)? 1'b0 : 
                             (N443)? 1'b0 : 
                             (N444)? 1'b0 : 
                             (N445)? 1'b0 : 
                             (N446)? 1'b0 : 
                             (N447)? 1'b0 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b1 : 
                             (N450)? 1'b1 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b1 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b1 : 
                             (N456)? 1'b1 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b1 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b1 : 
                             (N462)? 1'b1 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b1 : 
                             (N465)? 1'b0 : 
                             (N466)? 1'b0 : 
                             (N467)? 1'b1 : 
                             (N468)? 1'b0 : 
                             (N469)? 1'b1 : 
                             (N470)? 1'b1 : 
                             (N471)? 1'b0 : 
                             (N472)? 1'b0 : 
                             (N473)? 1'b1 : 
                             (N474)? 1'b1 : 
                             (N475)? 1'b0 : 
                             (N476)? 1'b1 : 
                             (N477)? 1'b0 : 
                             (N478)? 1'b0 : 
                             (N479)? 1'b1 : 
                             (N480)? 1'b1 : 
                             (N481)? 1'b0 : 
                             (N482)? 1'b0 : 
                             (N483)? 1'b1 : 
                             (N484)? 1'b0 : 
                             (N485)? 1'b1 : 
                             (N486)? 1'b1 : 
                             (N487)? 1'b0 : 
                             (N488)? 1'b0 : 
                             (N489)? 1'b1 : 
                             (N490)? 1'b1 : 
                             (N491)? 1'b0 : 
                             (N492)? 1'b1 : 
                             (N493)? 1'b0 : 
                             (N494)? 1'b0 : 
                             (N495)? 1'b1 : 
                             (N496)? 1'b0 : 
                             (N497)? 1'b1 : 
                             (N498)? 1'b1 : 
                             (N499)? 1'b0 : 
                             (N500)? 1'b1 : 
                             (N501)? 1'b0 : 
                             (N502)? 1'b0 : 
                             (N503)? 1'b1 : 
                             (N504)? 1'b1 : 
                             (N505)? 1'b0 : 
                             (N506)? 1'b0 : 
                             (N507)? 1'b1 : 
                             (N508)? 1'b0 : 
                             (N509)? 1'b1 : 
                             (N510)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign bk_datapath_o[16] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b1 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b1 : 
                             (N294)? 1'b1 : 
                             (N295)? 1'b1 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b1 : 
                             (N298)? 1'b1 : 
                             (N299)? 1'b1 : 
                             (N300)? 1'b1 : 
                             (N301)? 1'b1 : 
                             (N302)? 1'b1 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b1 : 
                             (N306)? 1'b1 : 
                             (N307)? 1'b1 : 
                             (N308)? 1'b1 : 
                             (N309)? 1'b1 : 
                             (N310)? 1'b1 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b1 : 
                             (N313)? 1'b1 : 
                             (N314)? 1'b1 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b1 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b1 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b1 : 
                             (N358)? 1'b1 : 
                             (N359)? 1'b1 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b1 : 
                             (N362)? 1'b1 : 
                             (N363)? 1'b1 : 
                             (N364)? 1'b1 : 
                             (N365)? 1'b1 : 
                             (N366)? 1'b1 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b1 : 
                             (N370)? 1'b1 : 
                             (N371)? 1'b1 : 
                             (N372)? 1'b1 : 
                             (N373)? 1'b1 : 
                             (N374)? 1'b1 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b1 : 
                             (N377)? 1'b1 : 
                             (N378)? 1'b1 : 
                             (N379)? 1'b0 : 
                             (N380)? 1'b1 : 
                             (N381)? 1'b0 : 
                             (N382)? 1'b0 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b0 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b0 : 
                             (N414)? 1'b0 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b1 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b1 : 
                             (N422)? 1'b1 : 
                             (N423)? 1'b1 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b1 : 
                             (N426)? 1'b1 : 
                             (N427)? 1'b1 : 
                             (N428)? 1'b1 : 
                             (N429)? 1'b1 : 
                             (N430)? 1'b1 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b1 : 
                             (N434)? 1'b1 : 
                             (N435)? 1'b1 : 
                             (N436)? 1'b1 : 
                             (N437)? 1'b1 : 
                             (N438)? 1'b1 : 
                             (N439)? 1'b0 : 
                             (N440)? 1'b1 : 
                             (N441)? 1'b1 : 
                             (N442)? 1'b1 : 
                             (N443)? 1'b0 : 
                             (N444)? 1'b1 : 
                             (N445)? 1'b0 : 
                             (N446)? 1'b0 : 
                             (N447)? 1'b0 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b0 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b0 : 
                             (N462)? 1'b0 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b0 : 
                             (N466)? 1'b0 : 
                             (N467)? 1'b0 : 
                             (N468)? 1'b0 : 
                             (N469)? 1'b0 : 
                             (N470)? 1'b0 : 
                             (N471)? 1'b0 : 
                             (N472)? 1'b0 : 
                             (N473)? 1'b0 : 
                             (N474)? 1'b0 : 
                             (N475)? 1'b0 : 
                             (N476)? 1'b0 : 
                             (N477)? 1'b0 : 
                             (N478)? 1'b0 : 
                             (N479)? 1'b0 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b0 : 
                             (N482)? 1'b0 : 
                             (N483)? 1'b1 : 
                             (N484)? 1'b0 : 
                             (N485)? 1'b1 : 
                             (N486)? 1'b1 : 
                             (N487)? 1'b1 : 
                             (N488)? 1'b0 : 
                             (N489)? 1'b1 : 
                             (N490)? 1'b1 : 
                             (N491)? 1'b1 : 
                             (N492)? 1'b1 : 
                             (N493)? 1'b1 : 
                             (N494)? 1'b1 : 
                             (N495)? 1'b0 : 
                             (N496)? 1'b0 : 
                             (N497)? 1'b1 : 
                             (N498)? 1'b1 : 
                             (N499)? 1'b1 : 
                             (N500)? 1'b1 : 
                             (N501)? 1'b1 : 
                             (N502)? 1'b1 : 
                             (N503)? 1'b0 : 
                             (N504)? 1'b1 : 
                             (N505)? 1'b1 : 
                             (N506)? 1'b1 : 
                             (N507)? 1'b0 : 
                             (N508)? 1'b1 : 
                             (N509)? 1'b0 : 
                             (N510)? 1'b0 : 
                             (N255)? 1'b0 : 1'b0;
  assign bk_datapath_o[15] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b0 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b0 : 
                             (N286)? 1'b0 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b1 : 
                             (N290)? 1'b1 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b1 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b1 : 
                             (N296)? 1'b1 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b1 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b1 : 
                             (N302)? 1'b1 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b1 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b1 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b1 : 
                             (N310)? 1'b1 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b1 : 
                             (N314)? 1'b1 : 
                             (N315)? 1'b0 : 
                             (N316)? 1'b1 : 
                             (N317)? 1'b0 : 
                             (N318)? 1'b0 : 
                             (N319)? 1'b1 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b0 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b0 : 
                             (N350)? 1'b0 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b1 : 
                             (N354)? 1'b1 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b1 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b1 : 
                             (N360)? 1'b1 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b1 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b1 : 
                             (N366)? 1'b1 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b1 : 
                             (N369)? 1'b0 : 
                             (N370)? 1'b0 : 
                             (N371)? 1'b1 : 
                             (N372)? 1'b0 : 
                             (N373)? 1'b1 : 
                             (N374)? 1'b1 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b0 : 
                             (N377)? 1'b1 : 
                             (N378)? 1'b1 : 
                             (N379)? 1'b0 : 
                             (N380)? 1'b1 : 
                             (N381)? 1'b0 : 
                             (N382)? 1'b0 : 
                             (N383)? 1'b1 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b0 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b0 : 
                             (N414)? 1'b0 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b1 : 
                             (N418)? 1'b1 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b1 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b1 : 
                             (N424)? 1'b1 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b1 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b1 : 
                             (N430)? 1'b1 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b1 : 
                             (N433)? 1'b0 : 
                             (N434)? 1'b0 : 
                             (N435)? 1'b1 : 
                             (N436)? 1'b0 : 
                             (N437)? 1'b1 : 
                             (N438)? 1'b1 : 
                             (N439)? 1'b0 : 
                             (N440)? 1'b0 : 
                             (N441)? 1'b1 : 
                             (N442)? 1'b1 : 
                             (N443)? 1'b0 : 
                             (N444)? 1'b1 : 
                             (N445)? 1'b0 : 
                             (N446)? 1'b0 : 
                             (N447)? 1'b1 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b0 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b0 : 
                             (N462)? 1'b0 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b0 : 
                             (N466)? 1'b0 : 
                             (N467)? 1'b0 : 
                             (N468)? 1'b0 : 
                             (N469)? 1'b0 : 
                             (N470)? 1'b0 : 
                             (N471)? 1'b0 : 
                             (N472)? 1'b0 : 
                             (N473)? 1'b0 : 
                             (N474)? 1'b0 : 
                             (N475)? 1'b0 : 
                             (N476)? 1'b0 : 
                             (N477)? 1'b0 : 
                             (N478)? 1'b0 : 
                             (N479)? 1'b0 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b1 : 
                             (N482)? 1'b1 : 
                             (N483)? 1'b0 : 
                             (N484)? 1'b1 : 
                             (N485)? 1'b0 : 
                             (N486)? 1'b0 : 
                             (N487)? 1'b1 : 
                             (N488)? 1'b1 : 
                             (N489)? 1'b0 : 
                             (N490)? 1'b0 : 
                             (N491)? 1'b1 : 
                             (N492)? 1'b0 : 
                             (N493)? 1'b1 : 
                             (N494)? 1'b1 : 
                             (N495)? 1'b0 : 
                             (N496)? 1'b1 : 
                             (N497)? 1'b0 : 
                             (N498)? 1'b0 : 
                             (N499)? 1'b1 : 
                             (N500)? 1'b0 : 
                             (N501)? 1'b1 : 
                             (N502)? 1'b1 : 
                             (N503)? 1'b0 : 
                             (N504)? 1'b0 : 
                             (N505)? 1'b1 : 
                             (N506)? 1'b1 : 
                             (N507)? 1'b0 : 
                             (N508)? 1'b1 : 
                             (N509)? 1'b0 : 
                             (N510)? 1'b0 : 
                             (N255)? 1'b1 : 1'b0;
  assign bk_datapath_o[13] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b1 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b1 : 
                             (N278)? 1'b1 : 
                             (N279)? 1'b1 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b1 : 
                             (N282)? 1'b1 : 
                             (N283)? 1'b1 : 
                             (N284)? 1'b1 : 
                             (N285)? 1'b1 : 
                             (N286)? 1'b1 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b1 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b1 : 
                             (N310)? 1'b1 : 
                             (N311)? 1'b1 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b1 : 
                             (N314)? 1'b1 : 
                             (N315)? 1'b1 : 
                             (N316)? 1'b1 : 
                             (N317)? 1'b1 : 
                             (N318)? 1'b1 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b1 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b1 : 
                             (N342)? 1'b1 : 
                             (N343)? 1'b1 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b1 : 
                             (N346)? 1'b1 : 
                             (N347)? 1'b1 : 
                             (N348)? 1'b1 : 
                             (N349)? 1'b1 : 
                             (N350)? 1'b1 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b0 : 
                             (N370)? 1'b0 : 
                             (N371)? 1'b1 : 
                             (N372)? 1'b0 : 
                             (N373)? 1'b1 : 
                             (N374)? 1'b1 : 
                             (N375)? 1'b1 : 
                             (N376)? 1'b0 : 
                             (N377)? 1'b1 : 
                             (N378)? 1'b1 : 
                             (N379)? 1'b1 : 
                             (N380)? 1'b1 : 
                             (N381)? 1'b1 : 
                             (N382)? 1'b1 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b1 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b1 : 
                             (N406)? 1'b1 : 
                             (N407)? 1'b1 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b1 : 
                             (N410)? 1'b1 : 
                             (N411)? 1'b1 : 
                             (N412)? 1'b1 : 
                             (N413)? 1'b1 : 
                             (N414)? 1'b1 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b0 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b0 : 
                             (N430)? 1'b0 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b0 : 
                             (N434)? 1'b0 : 
                             (N435)? 1'b1 : 
                             (N436)? 1'b0 : 
                             (N437)? 1'b1 : 
                             (N438)? 1'b1 : 
                             (N439)? 1'b1 : 
                             (N440)? 1'b0 : 
                             (N441)? 1'b1 : 
                             (N442)? 1'b1 : 
                             (N443)? 1'b1 : 
                             (N444)? 1'b1 : 
                             (N445)? 1'b1 : 
                             (N446)? 1'b1 : 
                             (N447)? 1'b0 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b0 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b0 : 
                             (N462)? 1'b0 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b0 : 
                             (N466)? 1'b0 : 
                             (N467)? 1'b1 : 
                             (N468)? 1'b0 : 
                             (N469)? 1'b1 : 
                             (N470)? 1'b1 : 
                             (N471)? 1'b1 : 
                             (N472)? 1'b0 : 
                             (N473)? 1'b1 : 
                             (N474)? 1'b1 : 
                             (N475)? 1'b1 : 
                             (N476)? 1'b1 : 
                             (N477)? 1'b1 : 
                             (N478)? 1'b1 : 
                             (N479)? 1'b0 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b0 : 
                             (N482)? 1'b0 : 
                             (N483)? 1'b0 : 
                             (N484)? 1'b0 : 
                             (N485)? 1'b0 : 
                             (N486)? 1'b0 : 
                             (N487)? 1'b0 : 
                             (N488)? 1'b0 : 
                             (N489)? 1'b0 : 
                             (N490)? 1'b0 : 
                             (N491)? 1'b0 : 
                             (N492)? 1'b0 : 
                             (N493)? 1'b0 : 
                             (N494)? 1'b0 : 
                             (N495)? 1'b0 : 
                             (N496)? 1'b0 : 
                             (N497)? 1'b0 : 
                             (N498)? 1'b0 : 
                             (N499)? 1'b1 : 
                             (N500)? 1'b0 : 
                             (N501)? 1'b1 : 
                             (N502)? 1'b1 : 
                             (N503)? 1'b1 : 
                             (N504)? 1'b0 : 
                             (N505)? 1'b1 : 
                             (N506)? 1'b1 : 
                             (N507)? 1'b1 : 
                             (N508)? 1'b1 : 
                             (N509)? 1'b1 : 
                             (N510)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign bk_datapath_o[12] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b0 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b0 : 
                             (N270)? 1'b0 : 
                             (N271)? 1'b0 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b1 : 
                             (N274)? 1'b1 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b1 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b1 : 
                             (N280)? 1'b1 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b1 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b1 : 
                             (N286)? 1'b1 : 
                             (N287)? 1'b0 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b0 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b0 : 
                             (N302)? 1'b0 : 
                             (N303)? 1'b0 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b1 : 
                             (N306)? 1'b1 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b1 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b1 : 
                             (N312)? 1'b1 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b1 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b1 : 
                             (N318)? 1'b1 : 
                             (N319)? 1'b0 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b0 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b0 : 
                             (N334)? 1'b0 : 
                             (N335)? 1'b0 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b1 : 
                             (N338)? 1'b1 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b1 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b1 : 
                             (N344)? 1'b1 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b1 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b1 : 
                             (N350)? 1'b1 : 
                             (N351)? 1'b0 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b0 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b0 : 
                             (N366)? 1'b0 : 
                             (N367)? 1'b0 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b1 : 
                             (N370)? 1'b1 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b1 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b1 : 
                             (N376)? 1'b1 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b1 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b1 : 
                             (N382)? 1'b1 : 
                             (N383)? 1'b0 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b0 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b0 : 
                             (N398)? 1'b0 : 
                             (N399)? 1'b0 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b1 : 
                             (N402)? 1'b1 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b1 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b1 : 
                             (N408)? 1'b1 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b1 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b1 : 
                             (N414)? 1'b1 : 
                             (N415)? 1'b0 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b0 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b0 : 
                             (N430)? 1'b0 : 
                             (N431)? 1'b0 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b1 : 
                             (N434)? 1'b1 : 
                             (N435)? 1'b0 : 
                             (N436)? 1'b1 : 
                             (N437)? 1'b0 : 
                             (N438)? 1'b0 : 
                             (N439)? 1'b1 : 
                             (N440)? 1'b1 : 
                             (N441)? 1'b0 : 
                             (N442)? 1'b0 : 
                             (N443)? 1'b1 : 
                             (N444)? 1'b0 : 
                             (N445)? 1'b1 : 
                             (N446)? 1'b1 : 
                             (N447)? 1'b0 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b0 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b0 : 
                             (N462)? 1'b0 : 
                             (N463)? 1'b0 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b1 : 
                             (N466)? 1'b1 : 
                             (N467)? 1'b0 : 
                             (N468)? 1'b1 : 
                             (N469)? 1'b0 : 
                             (N470)? 1'b0 : 
                             (N471)? 1'b1 : 
                             (N472)? 1'b1 : 
                             (N473)? 1'b0 : 
                             (N474)? 1'b0 : 
                             (N475)? 1'b1 : 
                             (N476)? 1'b0 : 
                             (N477)? 1'b1 : 
                             (N478)? 1'b1 : 
                             (N479)? 1'b0 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b0 : 
                             (N482)? 1'b0 : 
                             (N483)? 1'b0 : 
                             (N484)? 1'b0 : 
                             (N485)? 1'b0 : 
                             (N486)? 1'b0 : 
                             (N487)? 1'b0 : 
                             (N488)? 1'b0 : 
                             (N489)? 1'b0 : 
                             (N490)? 1'b0 : 
                             (N491)? 1'b0 : 
                             (N492)? 1'b0 : 
                             (N493)? 1'b0 : 
                             (N494)? 1'b0 : 
                             (N495)? 1'b0 : 
                             (N496)? 1'b0 : 
                             (N497)? 1'b1 : 
                             (N498)? 1'b1 : 
                             (N499)? 1'b0 : 
                             (N500)? 1'b1 : 
                             (N501)? 1'b0 : 
                             (N502)? 1'b0 : 
                             (N503)? 1'b1 : 
                             (N504)? 1'b1 : 
                             (N505)? 1'b0 : 
                             (N506)? 1'b0 : 
                             (N507)? 1'b1 : 
                             (N508)? 1'b0 : 
                             (N509)? 1'b1 : 
                             (N510)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign bk_datapath_o[10] = (N256)? 1'b0 : 
                             (N257)? 1'b0 : 
                             (N258)? 1'b0 : 
                             (N259)? 1'b0 : 
                             (N260)? 1'b0 : 
                             (N261)? 1'b0 : 
                             (N262)? 1'b0 : 
                             (N263)? 1'b0 : 
                             (N264)? 1'b0 : 
                             (N265)? 1'b0 : 
                             (N266)? 1'b0 : 
                             (N267)? 1'b1 : 
                             (N268)? 1'b0 : 
                             (N269)? 1'b1 : 
                             (N270)? 1'b1 : 
                             (N271)? 1'b1 : 
                             (N272)? 1'b0 : 
                             (N273)? 1'b0 : 
                             (N274)? 1'b0 : 
                             (N275)? 1'b0 : 
                             (N276)? 1'b0 : 
                             (N277)? 1'b0 : 
                             (N278)? 1'b0 : 
                             (N279)? 1'b0 : 
                             (N280)? 1'b0 : 
                             (N281)? 1'b0 : 
                             (N282)? 1'b0 : 
                             (N283)? 1'b1 : 
                             (N284)? 1'b0 : 
                             (N285)? 1'b1 : 
                             (N286)? 1'b1 : 
                             (N287)? 1'b1 : 
                             (N288)? 1'b0 : 
                             (N289)? 1'b0 : 
                             (N290)? 1'b0 : 
                             (N291)? 1'b0 : 
                             (N292)? 1'b0 : 
                             (N293)? 1'b0 : 
                             (N294)? 1'b0 : 
                             (N295)? 1'b0 : 
                             (N296)? 1'b0 : 
                             (N297)? 1'b0 : 
                             (N298)? 1'b0 : 
                             (N299)? 1'b1 : 
                             (N300)? 1'b0 : 
                             (N301)? 1'b1 : 
                             (N302)? 1'b1 : 
                             (N303)? 1'b1 : 
                             (N304)? 1'b0 : 
                             (N305)? 1'b0 : 
                             (N306)? 1'b0 : 
                             (N307)? 1'b0 : 
                             (N308)? 1'b0 : 
                             (N309)? 1'b0 : 
                             (N310)? 1'b0 : 
                             (N311)? 1'b0 : 
                             (N312)? 1'b0 : 
                             (N313)? 1'b0 : 
                             (N314)? 1'b0 : 
                             (N315)? 1'b1 : 
                             (N316)? 1'b0 : 
                             (N317)? 1'b1 : 
                             (N318)? 1'b1 : 
                             (N319)? 1'b1 : 
                             (N320)? 1'b0 : 
                             (N321)? 1'b0 : 
                             (N322)? 1'b0 : 
                             (N323)? 1'b0 : 
                             (N324)? 1'b0 : 
                             (N325)? 1'b0 : 
                             (N326)? 1'b0 : 
                             (N327)? 1'b0 : 
                             (N328)? 1'b0 : 
                             (N329)? 1'b0 : 
                             (N330)? 1'b0 : 
                             (N331)? 1'b1 : 
                             (N332)? 1'b0 : 
                             (N333)? 1'b1 : 
                             (N334)? 1'b1 : 
                             (N335)? 1'b1 : 
                             (N336)? 1'b0 : 
                             (N337)? 1'b0 : 
                             (N338)? 1'b0 : 
                             (N339)? 1'b0 : 
                             (N340)? 1'b0 : 
                             (N341)? 1'b0 : 
                             (N342)? 1'b0 : 
                             (N343)? 1'b0 : 
                             (N344)? 1'b0 : 
                             (N345)? 1'b0 : 
                             (N346)? 1'b0 : 
                             (N347)? 1'b1 : 
                             (N348)? 1'b0 : 
                             (N349)? 1'b1 : 
                             (N350)? 1'b1 : 
                             (N351)? 1'b1 : 
                             (N352)? 1'b0 : 
                             (N353)? 1'b0 : 
                             (N354)? 1'b0 : 
                             (N355)? 1'b0 : 
                             (N356)? 1'b0 : 
                             (N357)? 1'b0 : 
                             (N358)? 1'b0 : 
                             (N359)? 1'b0 : 
                             (N360)? 1'b0 : 
                             (N361)? 1'b0 : 
                             (N362)? 1'b0 : 
                             (N363)? 1'b1 : 
                             (N364)? 1'b0 : 
                             (N365)? 1'b1 : 
                             (N366)? 1'b1 : 
                             (N367)? 1'b1 : 
                             (N368)? 1'b0 : 
                             (N369)? 1'b0 : 
                             (N370)? 1'b0 : 
                             (N371)? 1'b0 : 
                             (N372)? 1'b0 : 
                             (N373)? 1'b0 : 
                             (N374)? 1'b0 : 
                             (N375)? 1'b0 : 
                             (N376)? 1'b0 : 
                             (N377)? 1'b0 : 
                             (N378)? 1'b0 : 
                             (N379)? 1'b1 : 
                             (N380)? 1'b0 : 
                             (N381)? 1'b1 : 
                             (N382)? 1'b1 : 
                             (N383)? 1'b1 : 
                             (N384)? 1'b0 : 
                             (N385)? 1'b0 : 
                             (N386)? 1'b0 : 
                             (N387)? 1'b0 : 
                             (N388)? 1'b0 : 
                             (N389)? 1'b0 : 
                             (N390)? 1'b0 : 
                             (N391)? 1'b0 : 
                             (N392)? 1'b0 : 
                             (N393)? 1'b0 : 
                             (N394)? 1'b0 : 
                             (N395)? 1'b1 : 
                             (N396)? 1'b0 : 
                             (N397)? 1'b1 : 
                             (N398)? 1'b1 : 
                             (N399)? 1'b1 : 
                             (N400)? 1'b0 : 
                             (N401)? 1'b0 : 
                             (N402)? 1'b0 : 
                             (N403)? 1'b0 : 
                             (N404)? 1'b0 : 
                             (N405)? 1'b0 : 
                             (N406)? 1'b0 : 
                             (N407)? 1'b0 : 
                             (N408)? 1'b0 : 
                             (N409)? 1'b0 : 
                             (N410)? 1'b0 : 
                             (N411)? 1'b1 : 
                             (N412)? 1'b0 : 
                             (N413)? 1'b1 : 
                             (N414)? 1'b1 : 
                             (N415)? 1'b1 : 
                             (N416)? 1'b0 : 
                             (N417)? 1'b0 : 
                             (N418)? 1'b0 : 
                             (N419)? 1'b0 : 
                             (N420)? 1'b0 : 
                             (N421)? 1'b0 : 
                             (N422)? 1'b0 : 
                             (N423)? 1'b0 : 
                             (N424)? 1'b0 : 
                             (N425)? 1'b0 : 
                             (N426)? 1'b0 : 
                             (N427)? 1'b1 : 
                             (N428)? 1'b0 : 
                             (N429)? 1'b1 : 
                             (N430)? 1'b1 : 
                             (N431)? 1'b1 : 
                             (N432)? 1'b0 : 
                             (N433)? 1'b0 : 
                             (N434)? 1'b0 : 
                             (N435)? 1'b0 : 
                             (N436)? 1'b0 : 
                             (N437)? 1'b0 : 
                             (N438)? 1'b0 : 
                             (N439)? 1'b0 : 
                             (N440)? 1'b0 : 
                             (N441)? 1'b0 : 
                             (N442)? 1'b0 : 
                             (N443)? 1'b1 : 
                             (N444)? 1'b0 : 
                             (N445)? 1'b1 : 
                             (N446)? 1'b1 : 
                             (N447)? 1'b1 : 
                             (N448)? 1'b0 : 
                             (N449)? 1'b0 : 
                             (N450)? 1'b0 : 
                             (N451)? 1'b0 : 
                             (N452)? 1'b0 : 
                             (N453)? 1'b0 : 
                             (N454)? 1'b0 : 
                             (N455)? 1'b0 : 
                             (N456)? 1'b0 : 
                             (N457)? 1'b0 : 
                             (N458)? 1'b0 : 
                             (N459)? 1'b1 : 
                             (N460)? 1'b0 : 
                             (N461)? 1'b1 : 
                             (N462)? 1'b1 : 
                             (N463)? 1'b1 : 
                             (N464)? 1'b0 : 
                             (N465)? 1'b0 : 
                             (N466)? 1'b0 : 
                             (N467)? 1'b0 : 
                             (N468)? 1'b0 : 
                             (N469)? 1'b0 : 
                             (N470)? 1'b0 : 
                             (N471)? 1'b0 : 
                             (N472)? 1'b0 : 
                             (N473)? 1'b0 : 
                             (N474)? 1'b0 : 
                             (N475)? 1'b1 : 
                             (N476)? 1'b0 : 
                             (N477)? 1'b1 : 
                             (N478)? 1'b1 : 
                             (N479)? 1'b1 : 
                             (N480)? 1'b0 : 
                             (N481)? 1'b0 : 
                             (N482)? 1'b0 : 
                             (N483)? 1'b0 : 
                             (N484)? 1'b0 : 
                             (N485)? 1'b0 : 
                             (N486)? 1'b0 : 
                             (N487)? 1'b0 : 
                             (N488)? 1'b0 : 
                             (N489)? 1'b0 : 
                             (N490)? 1'b0 : 
                             (N491)? 1'b1 : 
                             (N492)? 1'b0 : 
                             (N493)? 1'b1 : 
                             (N494)? 1'b1 : 
                             (N495)? 1'b1 : 
                             (N496)? 1'b0 : 
                             (N497)? 1'b0 : 
                             (N498)? 1'b0 : 
                             (N499)? 1'b0 : 
                             (N500)? 1'b0 : 
                             (N501)? 1'b0 : 
                             (N502)? 1'b0 : 
                             (N503)? 1'b0 : 
                             (N504)? 1'b0 : 
                             (N505)? 1'b0 : 
                             (N506)? 1'b0 : 
                             (N507)? 1'b1 : 
                             (N508)? 1'b0 : 
                             (N509)? 1'b1 : 
                             (N510)? 1'b1 : 
                             (N255)? 1'b1 : 1'b0;
  assign bk_datapath_o[9] = (N256)? 1'b0 : 
                            (N257)? 1'b0 : 
                            (N258)? 1'b0 : 
                            (N259)? 1'b0 : 
                            (N260)? 1'b0 : 
                            (N261)? 1'b0 : 
                            (N262)? 1'b0 : 
                            (N263)? 1'b0 : 
                            (N264)? 1'b0 : 
                            (N265)? 1'b1 : 
                            (N266)? 1'b1 : 
                            (N267)? 1'b0 : 
                            (N268)? 1'b1 : 
                            (N269)? 1'b0 : 
                            (N270)? 1'b0 : 
                            (N271)? 1'b1 : 
                            (N272)? 1'b0 : 
                            (N273)? 1'b0 : 
                            (N274)? 1'b0 : 
                            (N275)? 1'b0 : 
                            (N276)? 1'b0 : 
                            (N277)? 1'b0 : 
                            (N278)? 1'b0 : 
                            (N279)? 1'b0 : 
                            (N280)? 1'b0 : 
                            (N281)? 1'b1 : 
                            (N282)? 1'b1 : 
                            (N283)? 1'b0 : 
                            (N284)? 1'b1 : 
                            (N285)? 1'b0 : 
                            (N286)? 1'b0 : 
                            (N287)? 1'b1 : 
                            (N288)? 1'b0 : 
                            (N289)? 1'b0 : 
                            (N290)? 1'b0 : 
                            (N291)? 1'b0 : 
                            (N292)? 1'b0 : 
                            (N293)? 1'b0 : 
                            (N294)? 1'b0 : 
                            (N295)? 1'b0 : 
                            (N296)? 1'b0 : 
                            (N297)? 1'b1 : 
                            (N298)? 1'b1 : 
                            (N299)? 1'b0 : 
                            (N300)? 1'b1 : 
                            (N301)? 1'b0 : 
                            (N302)? 1'b0 : 
                            (N303)? 1'b1 : 
                            (N304)? 1'b0 : 
                            (N305)? 1'b0 : 
                            (N306)? 1'b0 : 
                            (N307)? 1'b0 : 
                            (N308)? 1'b0 : 
                            (N309)? 1'b0 : 
                            (N310)? 1'b0 : 
                            (N311)? 1'b0 : 
                            (N312)? 1'b0 : 
                            (N313)? 1'b1 : 
                            (N314)? 1'b1 : 
                            (N315)? 1'b0 : 
                            (N316)? 1'b1 : 
                            (N317)? 1'b0 : 
                            (N318)? 1'b0 : 
                            (N319)? 1'b1 : 
                            (N320)? 1'b0 : 
                            (N321)? 1'b0 : 
                            (N322)? 1'b0 : 
                            (N323)? 1'b0 : 
                            (N324)? 1'b0 : 
                            (N325)? 1'b0 : 
                            (N326)? 1'b0 : 
                            (N327)? 1'b0 : 
                            (N328)? 1'b0 : 
                            (N329)? 1'b1 : 
                            (N330)? 1'b1 : 
                            (N331)? 1'b0 : 
                            (N332)? 1'b1 : 
                            (N333)? 1'b0 : 
                            (N334)? 1'b0 : 
                            (N335)? 1'b1 : 
                            (N336)? 1'b0 : 
                            (N337)? 1'b0 : 
                            (N338)? 1'b0 : 
                            (N339)? 1'b0 : 
                            (N340)? 1'b0 : 
                            (N341)? 1'b0 : 
                            (N342)? 1'b0 : 
                            (N343)? 1'b0 : 
                            (N344)? 1'b0 : 
                            (N345)? 1'b1 : 
                            (N346)? 1'b1 : 
                            (N347)? 1'b0 : 
                            (N348)? 1'b1 : 
                            (N349)? 1'b0 : 
                            (N350)? 1'b0 : 
                            (N351)? 1'b1 : 
                            (N352)? 1'b0 : 
                            (N353)? 1'b0 : 
                            (N354)? 1'b0 : 
                            (N355)? 1'b0 : 
                            (N356)? 1'b0 : 
                            (N357)? 1'b0 : 
                            (N358)? 1'b0 : 
                            (N359)? 1'b0 : 
                            (N360)? 1'b0 : 
                            (N361)? 1'b1 : 
                            (N362)? 1'b1 : 
                            (N363)? 1'b0 : 
                            (N364)? 1'b1 : 
                            (N365)? 1'b0 : 
                            (N366)? 1'b0 : 
                            (N367)? 1'b1 : 
                            (N368)? 1'b0 : 
                            (N369)? 1'b0 : 
                            (N370)? 1'b0 : 
                            (N371)? 1'b0 : 
                            (N372)? 1'b0 : 
                            (N373)? 1'b0 : 
                            (N374)? 1'b0 : 
                            (N375)? 1'b0 : 
                            (N376)? 1'b0 : 
                            (N377)? 1'b1 : 
                            (N378)? 1'b1 : 
                            (N379)? 1'b0 : 
                            (N380)? 1'b1 : 
                            (N381)? 1'b0 : 
                            (N382)? 1'b0 : 
                            (N383)? 1'b1 : 
                            (N384)? 1'b0 : 
                            (N385)? 1'b0 : 
                            (N386)? 1'b0 : 
                            (N387)? 1'b0 : 
                            (N388)? 1'b0 : 
                            (N389)? 1'b0 : 
                            (N390)? 1'b0 : 
                            (N391)? 1'b0 : 
                            (N392)? 1'b0 : 
                            (N393)? 1'b1 : 
                            (N394)? 1'b1 : 
                            (N395)? 1'b0 : 
                            (N396)? 1'b1 : 
                            (N397)? 1'b0 : 
                            (N398)? 1'b0 : 
                            (N399)? 1'b1 : 
                            (N400)? 1'b0 : 
                            (N401)? 1'b0 : 
                            (N402)? 1'b0 : 
                            (N403)? 1'b0 : 
                            (N404)? 1'b0 : 
                            (N405)? 1'b0 : 
                            (N406)? 1'b0 : 
                            (N407)? 1'b0 : 
                            (N408)? 1'b0 : 
                            (N409)? 1'b1 : 
                            (N410)? 1'b1 : 
                            (N411)? 1'b0 : 
                            (N412)? 1'b1 : 
                            (N413)? 1'b0 : 
                            (N414)? 1'b0 : 
                            (N415)? 1'b1 : 
                            (N416)? 1'b0 : 
                            (N417)? 1'b0 : 
                            (N418)? 1'b0 : 
                            (N419)? 1'b0 : 
                            (N420)? 1'b0 : 
                            (N421)? 1'b0 : 
                            (N422)? 1'b0 : 
                            (N423)? 1'b0 : 
                            (N424)? 1'b0 : 
                            (N425)? 1'b1 : 
                            (N426)? 1'b1 : 
                            (N427)? 1'b0 : 
                            (N428)? 1'b1 : 
                            (N429)? 1'b0 : 
                            (N430)? 1'b0 : 
                            (N431)? 1'b1 : 
                            (N432)? 1'b0 : 
                            (N433)? 1'b0 : 
                            (N434)? 1'b0 : 
                            (N435)? 1'b0 : 
                            (N436)? 1'b0 : 
                            (N437)? 1'b0 : 
                            (N438)? 1'b0 : 
                            (N439)? 1'b0 : 
                            (N440)? 1'b0 : 
                            (N441)? 1'b1 : 
                            (N442)? 1'b1 : 
                            (N443)? 1'b0 : 
                            (N444)? 1'b1 : 
                            (N445)? 1'b0 : 
                            (N446)? 1'b0 : 
                            (N447)? 1'b1 : 
                            (N448)? 1'b0 : 
                            (N449)? 1'b0 : 
                            (N450)? 1'b0 : 
                            (N451)? 1'b0 : 
                            (N452)? 1'b0 : 
                            (N453)? 1'b0 : 
                            (N454)? 1'b0 : 
                            (N455)? 1'b0 : 
                            (N456)? 1'b0 : 
                            (N457)? 1'b1 : 
                            (N458)? 1'b1 : 
                            (N459)? 1'b0 : 
                            (N460)? 1'b1 : 
                            (N461)? 1'b0 : 
                            (N462)? 1'b0 : 
                            (N463)? 1'b1 : 
                            (N464)? 1'b0 : 
                            (N465)? 1'b0 : 
                            (N466)? 1'b0 : 
                            (N467)? 1'b0 : 
                            (N468)? 1'b0 : 
                            (N469)? 1'b0 : 
                            (N470)? 1'b0 : 
                            (N471)? 1'b0 : 
                            (N472)? 1'b0 : 
                            (N473)? 1'b1 : 
                            (N474)? 1'b1 : 
                            (N475)? 1'b0 : 
                            (N476)? 1'b1 : 
                            (N477)? 1'b0 : 
                            (N478)? 1'b0 : 
                            (N479)? 1'b1 : 
                            (N480)? 1'b0 : 
                            (N481)? 1'b0 : 
                            (N482)? 1'b0 : 
                            (N483)? 1'b0 : 
                            (N484)? 1'b0 : 
                            (N485)? 1'b0 : 
                            (N486)? 1'b0 : 
                            (N487)? 1'b0 : 
                            (N488)? 1'b0 : 
                            (N489)? 1'b1 : 
                            (N490)? 1'b1 : 
                            (N491)? 1'b0 : 
                            (N492)? 1'b1 : 
                            (N493)? 1'b0 : 
                            (N494)? 1'b0 : 
                            (N495)? 1'b1 : 
                            (N496)? 1'b0 : 
                            (N497)? 1'b0 : 
                            (N498)? 1'b0 : 
                            (N499)? 1'b0 : 
                            (N500)? 1'b0 : 
                            (N501)? 1'b0 : 
                            (N502)? 1'b0 : 
                            (N503)? 1'b0 : 
                            (N504)? 1'b0 : 
                            (N505)? 1'b1 : 
                            (N506)? 1'b1 : 
                            (N507)? 1'b0 : 
                            (N508)? 1'b1 : 
                            (N509)? 1'b0 : 
                            (N510)? 1'b0 : 
                            (N255)? 1'b1 : 1'b0;
  assign bk_datapath_o[6] = (N256)? 1'b0 : 
                            (N257)? 1'b0 : 
                            (N258)? 1'b0 : 
                            (N259)? 1'b0 : 
                            (N260)? 1'b0 : 
                            (N261)? 1'b1 : 
                            (N262)? 1'b1 : 
                            (N263)? 1'b0 : 
                            (N264)? 1'b0 : 
                            (N265)? 1'b0 : 
                            (N266)? 1'b0 : 
                            (N267)? 1'b0 : 
                            (N268)? 1'b0 : 
                            (N269)? 1'b1 : 
                            (N270)? 1'b1 : 
                            (N271)? 1'b0 : 
                            (N272)? 1'b0 : 
                            (N273)? 1'b0 : 
                            (N274)? 1'b0 : 
                            (N275)? 1'b0 : 
                            (N276)? 1'b0 : 
                            (N277)? 1'b1 : 
                            (N278)? 1'b1 : 
                            (N279)? 1'b0 : 
                            (N280)? 1'b0 : 
                            (N281)? 1'b0 : 
                            (N282)? 1'b0 : 
                            (N283)? 1'b0 : 
                            (N284)? 1'b0 : 
                            (N285)? 1'b1 : 
                            (N286)? 1'b1 : 
                            (N287)? 1'b0 : 
                            (N288)? 1'b0 : 
                            (N289)? 1'b0 : 
                            (N290)? 1'b0 : 
                            (N291)? 1'b0 : 
                            (N292)? 1'b0 : 
                            (N293)? 1'b1 : 
                            (N294)? 1'b1 : 
                            (N295)? 1'b0 : 
                            (N296)? 1'b0 : 
                            (N297)? 1'b0 : 
                            (N298)? 1'b0 : 
                            (N299)? 1'b0 : 
                            (N300)? 1'b0 : 
                            (N301)? 1'b1 : 
                            (N302)? 1'b1 : 
                            (N303)? 1'b0 : 
                            (N304)? 1'b0 : 
                            (N305)? 1'b0 : 
                            (N306)? 1'b0 : 
                            (N307)? 1'b0 : 
                            (N308)? 1'b0 : 
                            (N309)? 1'b1 : 
                            (N310)? 1'b1 : 
                            (N311)? 1'b0 : 
                            (N312)? 1'b0 : 
                            (N313)? 1'b0 : 
                            (N314)? 1'b0 : 
                            (N315)? 1'b0 : 
                            (N316)? 1'b0 : 
                            (N317)? 1'b1 : 
                            (N318)? 1'b1 : 
                            (N319)? 1'b0 : 
                            (N320)? 1'b0 : 
                            (N321)? 1'b0 : 
                            (N322)? 1'b0 : 
                            (N323)? 1'b0 : 
                            (N324)? 1'b0 : 
                            (N325)? 1'b1 : 
                            (N326)? 1'b1 : 
                            (N327)? 1'b0 : 
                            (N328)? 1'b0 : 
                            (N329)? 1'b0 : 
                            (N330)? 1'b0 : 
                            (N331)? 1'b0 : 
                            (N332)? 1'b0 : 
                            (N333)? 1'b1 : 
                            (N334)? 1'b1 : 
                            (N335)? 1'b0 : 
                            (N336)? 1'b0 : 
                            (N337)? 1'b0 : 
                            (N338)? 1'b0 : 
                            (N339)? 1'b0 : 
                            (N340)? 1'b0 : 
                            (N341)? 1'b1 : 
                            (N342)? 1'b1 : 
                            (N343)? 1'b0 : 
                            (N344)? 1'b0 : 
                            (N345)? 1'b0 : 
                            (N346)? 1'b0 : 
                            (N347)? 1'b0 : 
                            (N348)? 1'b0 : 
                            (N349)? 1'b1 : 
                            (N350)? 1'b1 : 
                            (N351)? 1'b0 : 
                            (N352)? 1'b0 : 
                            (N353)? 1'b0 : 
                            (N354)? 1'b0 : 
                            (N355)? 1'b0 : 
                            (N356)? 1'b0 : 
                            (N357)? 1'b1 : 
                            (N358)? 1'b1 : 
                            (N359)? 1'b0 : 
                            (N360)? 1'b0 : 
                            (N361)? 1'b0 : 
                            (N362)? 1'b0 : 
                            (N363)? 1'b0 : 
                            (N364)? 1'b0 : 
                            (N365)? 1'b1 : 
                            (N366)? 1'b1 : 
                            (N367)? 1'b0 : 
                            (N368)? 1'b0 : 
                            (N369)? 1'b0 : 
                            (N370)? 1'b0 : 
                            (N371)? 1'b0 : 
                            (N372)? 1'b0 : 
                            (N373)? 1'b1 : 
                            (N374)? 1'b1 : 
                            (N375)? 1'b0 : 
                            (N376)? 1'b0 : 
                            (N377)? 1'b0 : 
                            (N378)? 1'b0 : 
                            (N379)? 1'b0 : 
                            (N380)? 1'b0 : 
                            (N381)? 1'b1 : 
                            (N382)? 1'b1 : 
                            (N383)? 1'b0 : 
                            (N384)? 1'b0 : 
                            (N385)? 1'b0 : 
                            (N386)? 1'b0 : 
                            (N387)? 1'b0 : 
                            (N388)? 1'b0 : 
                            (N389)? 1'b1 : 
                            (N390)? 1'b1 : 
                            (N391)? 1'b0 : 
                            (N392)? 1'b0 : 
                            (N393)? 1'b0 : 
                            (N394)? 1'b0 : 
                            (N395)? 1'b0 : 
                            (N396)? 1'b0 : 
                            (N397)? 1'b1 : 
                            (N398)? 1'b1 : 
                            (N399)? 1'b0 : 
                            (N400)? 1'b0 : 
                            (N401)? 1'b0 : 
                            (N402)? 1'b0 : 
                            (N403)? 1'b0 : 
                            (N404)? 1'b0 : 
                            (N405)? 1'b1 : 
                            (N406)? 1'b1 : 
                            (N407)? 1'b0 : 
                            (N408)? 1'b0 : 
                            (N409)? 1'b0 : 
                            (N410)? 1'b0 : 
                            (N411)? 1'b0 : 
                            (N412)? 1'b0 : 
                            (N413)? 1'b1 : 
                            (N414)? 1'b1 : 
                            (N415)? 1'b0 : 
                            (N416)? 1'b0 : 
                            (N417)? 1'b0 : 
                            (N418)? 1'b0 : 
                            (N419)? 1'b0 : 
                            (N420)? 1'b0 : 
                            (N421)? 1'b1 : 
                            (N422)? 1'b1 : 
                            (N423)? 1'b0 : 
                            (N424)? 1'b0 : 
                            (N425)? 1'b0 : 
                            (N426)? 1'b0 : 
                            (N427)? 1'b0 : 
                            (N428)? 1'b0 : 
                            (N429)? 1'b1 : 
                            (N430)? 1'b1 : 
                            (N431)? 1'b0 : 
                            (N432)? 1'b0 : 
                            (N433)? 1'b0 : 
                            (N434)? 1'b0 : 
                            (N435)? 1'b0 : 
                            (N436)? 1'b0 : 
                            (N437)? 1'b1 : 
                            (N438)? 1'b1 : 
                            (N439)? 1'b0 : 
                            (N440)? 1'b0 : 
                            (N441)? 1'b0 : 
                            (N442)? 1'b0 : 
                            (N443)? 1'b0 : 
                            (N444)? 1'b0 : 
                            (N445)? 1'b1 : 
                            (N446)? 1'b1 : 
                            (N447)? 1'b0 : 
                            (N448)? 1'b0 : 
                            (N449)? 1'b0 : 
                            (N450)? 1'b0 : 
                            (N451)? 1'b0 : 
                            (N452)? 1'b0 : 
                            (N453)? 1'b1 : 
                            (N454)? 1'b1 : 
                            (N455)? 1'b0 : 
                            (N456)? 1'b0 : 
                            (N457)? 1'b0 : 
                            (N458)? 1'b0 : 
                            (N459)? 1'b0 : 
                            (N460)? 1'b0 : 
                            (N461)? 1'b1 : 
                            (N462)? 1'b1 : 
                            (N463)? 1'b0 : 
                            (N464)? 1'b0 : 
                            (N465)? 1'b0 : 
                            (N466)? 1'b0 : 
                            (N467)? 1'b0 : 
                            (N468)? 1'b0 : 
                            (N469)? 1'b1 : 
                            (N470)? 1'b1 : 
                            (N471)? 1'b0 : 
                            (N472)? 1'b0 : 
                            (N473)? 1'b0 : 
                            (N474)? 1'b0 : 
                            (N475)? 1'b0 : 
                            (N476)? 1'b0 : 
                            (N477)? 1'b1 : 
                            (N478)? 1'b1 : 
                            (N479)? 1'b0 : 
                            (N480)? 1'b0 : 
                            (N481)? 1'b0 : 
                            (N482)? 1'b0 : 
                            (N483)? 1'b0 : 
                            (N484)? 1'b0 : 
                            (N485)? 1'b1 : 
                            (N486)? 1'b1 : 
                            (N487)? 1'b0 : 
                            (N488)? 1'b0 : 
                            (N489)? 1'b0 : 
                            (N490)? 1'b0 : 
                            (N491)? 1'b0 : 
                            (N492)? 1'b0 : 
                            (N493)? 1'b1 : 
                            (N494)? 1'b1 : 
                            (N495)? 1'b0 : 
                            (N496)? 1'b0 : 
                            (N497)? 1'b0 : 
                            (N498)? 1'b0 : 
                            (N499)? 1'b0 : 
                            (N500)? 1'b0 : 
                            (N501)? 1'b1 : 
                            (N502)? 1'b1 : 
                            (N503)? 1'b0 : 
                            (N504)? 1'b0 : 
                            (N505)? 1'b0 : 
                            (N506)? 1'b0 : 
                            (N507)? 1'b0 : 
                            (N508)? 1'b0 : 
                            (N509)? 1'b1 : 
                            (N510)? 1'b1 : 
                            (N255)? 1'b0 : 1'b0;
  assign bk_datapath_o[3] = (N256)? 1'b0 : 
                            (N257)? 1'b0 : 
                            (N258)? 1'b0 : 
                            (N259)? 1'b1 : 
                            (N260)? 1'b0 : 
                            (N261)? 1'b0 : 
                            (N262)? 1'b0 : 
                            (N263)? 1'b1 : 
                            (N264)? 1'b0 : 
                            (N265)? 1'b0 : 
                            (N266)? 1'b0 : 
                            (N267)? 1'b1 : 
                            (N268)? 1'b0 : 
                            (N269)? 1'b0 : 
                            (N270)? 1'b0 : 
                            (N271)? 1'b1 : 
                            (N272)? 1'b0 : 
                            (N273)? 1'b0 : 
                            (N274)? 1'b0 : 
                            (N275)? 1'b1 : 
                            (N276)? 1'b0 : 
                            (N277)? 1'b0 : 
                            (N278)? 1'b0 : 
                            (N279)? 1'b1 : 
                            (N280)? 1'b0 : 
                            (N281)? 1'b0 : 
                            (N282)? 1'b0 : 
                            (N283)? 1'b1 : 
                            (N284)? 1'b0 : 
                            (N285)? 1'b0 : 
                            (N286)? 1'b0 : 
                            (N287)? 1'b1 : 
                            (N288)? 1'b0 : 
                            (N289)? 1'b0 : 
                            (N290)? 1'b0 : 
                            (N291)? 1'b1 : 
                            (N292)? 1'b0 : 
                            (N293)? 1'b0 : 
                            (N294)? 1'b0 : 
                            (N295)? 1'b1 : 
                            (N296)? 1'b0 : 
                            (N297)? 1'b0 : 
                            (N298)? 1'b0 : 
                            (N299)? 1'b1 : 
                            (N300)? 1'b0 : 
                            (N301)? 1'b0 : 
                            (N302)? 1'b0 : 
                            (N303)? 1'b1 : 
                            (N304)? 1'b0 : 
                            (N305)? 1'b0 : 
                            (N306)? 1'b0 : 
                            (N307)? 1'b1 : 
                            (N308)? 1'b0 : 
                            (N309)? 1'b0 : 
                            (N310)? 1'b0 : 
                            (N311)? 1'b1 : 
                            (N312)? 1'b0 : 
                            (N313)? 1'b0 : 
                            (N314)? 1'b0 : 
                            (N315)? 1'b1 : 
                            (N316)? 1'b0 : 
                            (N317)? 1'b0 : 
                            (N318)? 1'b0 : 
                            (N319)? 1'b1 : 
                            (N320)? 1'b0 : 
                            (N321)? 1'b0 : 
                            (N322)? 1'b0 : 
                            (N323)? 1'b1 : 
                            (N324)? 1'b0 : 
                            (N325)? 1'b0 : 
                            (N326)? 1'b0 : 
                            (N327)? 1'b1 : 
                            (N328)? 1'b0 : 
                            (N329)? 1'b0 : 
                            (N330)? 1'b0 : 
                            (N331)? 1'b1 : 
                            (N332)? 1'b0 : 
                            (N333)? 1'b0 : 
                            (N334)? 1'b0 : 
                            (N335)? 1'b1 : 
                            (N336)? 1'b0 : 
                            (N337)? 1'b0 : 
                            (N338)? 1'b0 : 
                            (N339)? 1'b1 : 
                            (N340)? 1'b0 : 
                            (N341)? 1'b0 : 
                            (N342)? 1'b0 : 
                            (N343)? 1'b1 : 
                            (N344)? 1'b0 : 
                            (N345)? 1'b0 : 
                            (N346)? 1'b0 : 
                            (N347)? 1'b1 : 
                            (N348)? 1'b0 : 
                            (N349)? 1'b0 : 
                            (N350)? 1'b0 : 
                            (N351)? 1'b1 : 
                            (N352)? 1'b0 : 
                            (N353)? 1'b0 : 
                            (N354)? 1'b0 : 
                            (N355)? 1'b1 : 
                            (N356)? 1'b0 : 
                            (N357)? 1'b0 : 
                            (N358)? 1'b0 : 
                            (N359)? 1'b1 : 
                            (N360)? 1'b0 : 
                            (N361)? 1'b0 : 
                            (N362)? 1'b0 : 
                            (N363)? 1'b1 : 
                            (N364)? 1'b0 : 
                            (N365)? 1'b0 : 
                            (N366)? 1'b0 : 
                            (N367)? 1'b1 : 
                            (N368)? 1'b0 : 
                            (N369)? 1'b0 : 
                            (N370)? 1'b0 : 
                            (N371)? 1'b1 : 
                            (N372)? 1'b0 : 
                            (N373)? 1'b0 : 
                            (N374)? 1'b0 : 
                            (N375)? 1'b1 : 
                            (N376)? 1'b0 : 
                            (N377)? 1'b0 : 
                            (N378)? 1'b0 : 
                            (N379)? 1'b1 : 
                            (N380)? 1'b0 : 
                            (N381)? 1'b0 : 
                            (N382)? 1'b0 : 
                            (N383)? 1'b1 : 
                            (N384)? 1'b0 : 
                            (N385)? 1'b0 : 
                            (N386)? 1'b0 : 
                            (N387)? 1'b1 : 
                            (N388)? 1'b0 : 
                            (N389)? 1'b0 : 
                            (N390)? 1'b0 : 
                            (N391)? 1'b1 : 
                            (N392)? 1'b0 : 
                            (N393)? 1'b0 : 
                            (N394)? 1'b0 : 
                            (N395)? 1'b1 : 
                            (N396)? 1'b0 : 
                            (N397)? 1'b0 : 
                            (N398)? 1'b0 : 
                            (N399)? 1'b1 : 
                            (N400)? 1'b0 : 
                            (N401)? 1'b0 : 
                            (N402)? 1'b0 : 
                            (N403)? 1'b1 : 
                            (N404)? 1'b0 : 
                            (N405)? 1'b0 : 
                            (N406)? 1'b0 : 
                            (N407)? 1'b1 : 
                            (N408)? 1'b0 : 
                            (N409)? 1'b0 : 
                            (N410)? 1'b0 : 
                            (N411)? 1'b1 : 
                            (N412)? 1'b0 : 
                            (N413)? 1'b0 : 
                            (N414)? 1'b0 : 
                            (N415)? 1'b1 : 
                            (N416)? 1'b0 : 
                            (N417)? 1'b0 : 
                            (N418)? 1'b0 : 
                            (N419)? 1'b1 : 
                            (N420)? 1'b0 : 
                            (N421)? 1'b0 : 
                            (N422)? 1'b0 : 
                            (N423)? 1'b1 : 
                            (N424)? 1'b0 : 
                            (N425)? 1'b0 : 
                            (N426)? 1'b0 : 
                            (N427)? 1'b1 : 
                            (N428)? 1'b0 : 
                            (N429)? 1'b0 : 
                            (N430)? 1'b0 : 
                            (N431)? 1'b1 : 
                            (N432)? 1'b0 : 
                            (N433)? 1'b0 : 
                            (N434)? 1'b0 : 
                            (N435)? 1'b1 : 
                            (N436)? 1'b0 : 
                            (N437)? 1'b0 : 
                            (N438)? 1'b0 : 
                            (N439)? 1'b1 : 
                            (N440)? 1'b0 : 
                            (N441)? 1'b0 : 
                            (N442)? 1'b0 : 
                            (N443)? 1'b1 : 
                            (N444)? 1'b0 : 
                            (N445)? 1'b0 : 
                            (N446)? 1'b0 : 
                            (N447)? 1'b1 : 
                            (N448)? 1'b0 : 
                            (N449)? 1'b0 : 
                            (N450)? 1'b0 : 
                            (N451)? 1'b1 : 
                            (N452)? 1'b0 : 
                            (N453)? 1'b0 : 
                            (N454)? 1'b0 : 
                            (N455)? 1'b1 : 
                            (N456)? 1'b0 : 
                            (N457)? 1'b0 : 
                            (N458)? 1'b0 : 
                            (N459)? 1'b1 : 
                            (N460)? 1'b0 : 
                            (N461)? 1'b0 : 
                            (N462)? 1'b0 : 
                            (N463)? 1'b1 : 
                            (N464)? 1'b0 : 
                            (N465)? 1'b0 : 
                            (N466)? 1'b0 : 
                            (N467)? 1'b1 : 
                            (N468)? 1'b0 : 
                            (N469)? 1'b0 : 
                            (N470)? 1'b0 : 
                            (N471)? 1'b1 : 
                            (N472)? 1'b0 : 
                            (N473)? 1'b0 : 
                            (N474)? 1'b0 : 
                            (N475)? 1'b1 : 
                            (N476)? 1'b0 : 
                            (N477)? 1'b0 : 
                            (N478)? 1'b0 : 
                            (N479)? 1'b1 : 
                            (N480)? 1'b0 : 
                            (N481)? 1'b0 : 
                            (N482)? 1'b0 : 
                            (N483)? 1'b1 : 
                            (N484)? 1'b0 : 
                            (N485)? 1'b0 : 
                            (N486)? 1'b0 : 
                            (N487)? 1'b1 : 
                            (N488)? 1'b0 : 
                            (N489)? 1'b0 : 
                            (N490)? 1'b0 : 
                            (N491)? 1'b1 : 
                            (N492)? 1'b0 : 
                            (N493)? 1'b0 : 
                            (N494)? 1'b0 : 
                            (N495)? 1'b1 : 
                            (N496)? 1'b0 : 
                            (N497)? 1'b0 : 
                            (N498)? 1'b0 : 
                            (N499)? 1'b1 : 
                            (N500)? 1'b0 : 
                            (N501)? 1'b0 : 
                            (N502)? 1'b0 : 
                            (N503)? 1'b1 : 
                            (N504)? 1'b0 : 
                            (N505)? 1'b0 : 
                            (N506)? 1'b0 : 
                            (N507)? 1'b1 : 
                            (N508)? 1'b0 : 
                            (N509)? 1'b0 : 
                            (N510)? 1'b0 : 
                            (N255)? 1'b1 : 1'b0;
  assign fwd_o[23] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b1 : 
                     (N736)? 1'b1 : 
                     (N737)? 1'b1 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b1 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b1 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b0 : 
                     (N752)? 1'b0 : 
                     (N753)? 1'b0 : 
                     (N754)? 1'b0 : 
                     (N755)? 1'b0 : 
                     (N756)? 1'b0 : 
                     (N757)? 1'b0 : 
                     (N758)? 1'b0 : 
                     (N759)? 1'b0 : 
                     (N760)? 1'b0 : 
                     (N761)? 1'b0 : 
                     (N762)? 1'b0 : 
                     (N763)? 1'b0 : 
                     (N764)? 1'b0 : 
                     (N765)? 1'b0 : 
                     (N255)? 1'b1 : 1'b0;
  assign N511 = N2252;
  assign N512 = N2256;
  assign N513 = N2260;
  assign N514 = N2263;
  assign N515 = N2266;
  assign N516 = N2269;
  assign N517 = N2272;
  assign N518 = N2275;
  assign N519 = N2278;
  assign N520 = N2281;
  assign N521 = N2284;
  assign N522 = N2287;
  assign N523 = N2291;
  assign N524 = N2294;
  assign N525 = N2297;
  assign N526 = N2300;
  assign N527 = N2302;
  assign N528 = N2304;
  assign N529 = N2306;
  assign N530 = N2308;
  assign N531 = N2311;
  assign N532 = N2313;
  assign N533 = N2315;
  assign N534 = N2317;
  assign N535 = N2319;
  assign N536 = N2321;
  assign N537 = N2323;
  assign N538 = N2325;
  assign N539 = N2328;
  assign N540 = N2330;
  assign N541 = N2332;
  assign N542 = N2334;
  assign N543 = N2336;
  assign N544 = N2338;
  assign N545 = N2340;
  assign N546 = N2342;
  assign N547 = N2345;
  assign N548 = N2347;
  assign N549 = N2349;
  assign N550 = N2351;
  assign N551 = N2353;
  assign N552 = N2355;
  assign N553 = N2357;
  assign N554 = N2359;
  assign N555 = N2361;
  assign N556 = N2363;
  assign N557 = N2365;
  assign N558 = N2367;
  assign N559 = N2369;
  assign N560 = N2371;
  assign N561 = N2373;
  assign N562 = N2375;
  assign N563 = N2379;
  assign N564 = N2381;
  assign N565 = N2383;
  assign N566 = N2385;
  assign N567 = N2387;
  assign N568 = N2389;
  assign N569 = N2391;
  assign N570 = N2393;
  assign N571 = N2395;
  assign N572 = N2397;
  assign N573 = N2399;
  assign N574 = N2401;
  assign N575 = N2404;
  assign N576 = N2406;
  assign N577 = N2408;
  assign N578 = N2410;
  assign N579 = N2412;
  assign N580 = N2414;
  assign N581 = N2416;
  assign N582 = N2418;
  assign N583 = N2420;
  assign N584 = N2422;
  assign N585 = N2424;
  assign N586 = N2426;
  assign N587 = N2429;
  assign N588 = N2431;
  assign N589 = N2433;
  assign N590 = N2435;
  assign N591 = N2437;
  assign N592 = N2439;
  assign N593 = N2441;
  assign N594 = N2443;
  assign N595 = N2446;
  assign N596 = N2448;
  assign N597 = N2450;
  assign N598 = N2452;
  assign N599 = N2454;
  assign N600 = N2456;
  assign N601 = N2458;
  assign N602 = N2460;
  assign N603 = N2462;
  assign N604 = N2464;
  assign N605 = N2466;
  assign N606 = N2468;
  assign N607 = N2470;
  assign N608 = N2472;
  assign N609 = N2474;
  assign N610 = N2476;
  assign N611 = N2479;
  assign N612 = N2481;
  assign N613 = N2483;
  assign N614 = N2485;
  assign N615 = N2487;
  assign N616 = N2489;
  assign N617 = N2491;
  assign N618 = N2493;
  assign N619 = N2495;
  assign N620 = N2497;
  assign N621 = N2499;
  assign N622 = N2501;
  assign N623 = N2503;
  assign N624 = N2506;
  assign N625 = N2509;
  assign N626 = N2512;
  assign N627 = N2516;
  assign N628 = N2519;
  assign N629 = N2522;
  assign N630 = N2525;
  assign N631 = N2528;
  assign N632 = N2531;
  assign N633 = N2534;
  assign N634 = N2536;
  assign N635 = N2542;
  assign N636 = N2544;
  assign N637 = N2546;
  assign N638 = N2549;
  assign N639 = N2553;
  assign N640 = N2555;
  assign N641 = N2558;
  assign N642 = N2560;
  assign N643 = N2562;
  assign N644 = N2564;
  assign N645 = N2566;
  assign N646 = N2568;
  assign N647 = N2571;
  assign N648 = N2573;
  assign N649 = N2575;
  assign N650 = N2577;
  assign N651 = N2579;
  assign N652 = N2581;
  assign N653 = N2583;
  assign N654 = N2585;
  assign N655 = N2587;
  assign N656 = N2589;
  assign N657 = N2591;
  assign N658 = N2593;
  assign N659 = N2596;
  assign N660 = N2598;
  assign N661 = N2600;
  assign N662 = N2602;
  assign N663 = N2604;
  assign N664 = N2606;
  assign N665 = N2608;
  assign N666 = N2610;
  assign N667 = N2612;
  assign N668 = N2614;
  assign N669 = N2616;
  assign N670 = N2618;
  assign N671 = N2620;
  assign N672 = N2622;
  assign N673 = N2624;
  assign N674 = N2626;
  assign N675 = N2629;
  assign N676 = N2631;
  assign N677 = N2633;
  assign N678 = N2635;
  assign N679 = N2637;
  assign N680 = N2639;
  assign N681 = N2641;
  assign N682 = N2643;
  assign N683 = N2645;
  assign N684 = N2647;
  assign N685 = N2649;
  assign N686 = N2651;
  assign N687 = N2653;
  assign N688 = N2655;
  assign N689 = N2657;
  assign N690 = N2659;
  assign N691 = N2662;
  assign N692 = N2664;
  assign N693 = N2666;
  assign N694 = N2668;
  assign N695 = N2670;
  assign N696 = N2672;
  assign N697 = N2674;
  assign N698 = N2676;
  assign N699 = N2679;
  assign N700 = N2681;
  assign N701 = N2683;
  assign N702 = N2685;
  assign N703 = N2689;
  assign N704 = N2691;
  assign N705 = N2693;
  assign N706 = N2695;
  assign N707 = N2697;
  assign N708 = N2699;
  assign N709 = N2701;
  assign N710 = N2703;
  assign N711 = N2705;
  assign N712 = N2707;
  assign N713 = N2709;
  assign N714 = N2711;
  assign N715 = N2713;
  assign N716 = N2715;
  assign N717 = N2717;
  assign N718 = N2719;
  assign N719 = N2721;
  assign N720 = N2723;
  assign N721 = N2725;
  assign N722 = N2727;
  assign N723 = N2730;
  assign N724 = N2732;
  assign N725 = N2734;
  assign N726 = N2736;
  assign N727 = N2738;
  assign N728 = N2740;
  assign N729 = N2742;
  assign N730 = N2744;
  assign N731 = N2746;
  assign N732 = N2748;
  assign N733 = N2750;
  assign N734 = N2752;
  assign N735 = N2754;
  assign N736 = N2756;
  assign N737 = N2758;
  assign N738 = N2760;
  assign N739 = N2763;
  assign N740 = N2765;
  assign N741 = N2767;
  assign N742 = N2769;
  assign N743 = N2771;
  assign N744 = N2773;
  assign N745 = N2775;
  assign N746 = N2777;
  assign N747 = N2779;
  assign N748 = N2781;
  assign N749 = N2783;
  assign N750 = N2785;
  assign N751 = N2787;
  assign N752 = N2789;
  assign N753 = N2791;
  assign N754 = N2793;
  assign N755 = N2796;
  assign N756 = N2798;
  assign N757 = N2800;
  assign N758 = N2802;
  assign N759 = N2804;
  assign N760 = N2806;
  assign N761 = N2808;
  assign N762 = N2812;
  assign N763 = N2814;
  assign N764 = N2817;
  assign N765 = N2820;
  assign fwd_o[22] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b0 : 
                     (N704)? 1'b0 : 
                     (N705)? 1'b0 : 
                     (N706)? 1'b0 : 
                     (N707)? 1'b0 : 
                     (N708)? 1'b0 : 
                     (N709)? 1'b0 : 
                     (N710)? 1'b0 : 
                     (N711)? 1'b0 : 
                     (N712)? 1'b0 : 
                     (N713)? 1'b0 : 
                     (N714)? 1'b0 : 
                     (N715)? 1'b0 : 
                     (N716)? 1'b0 : 
                     (N717)? 1'b0 : 
                     (N718)? 1'b0 : 
                     (N719)? 1'b0 : 
                     (N720)? 1'b0 : 
                     (N721)? 1'b0 : 
                     (N722)? 1'b0 : 
                     (N723)? 1'b0 : 
                     (N724)? 1'b0 : 
                     (N725)? 1'b0 : 
                     (N726)? 1'b0 : 
                     (N727)? 1'b0 : 
                     (N728)? 1'b0 : 
                     (N729)? 1'b0 : 
                     (N730)? 1'b0 : 
                     (N731)? 1'b0 : 
                     (N732)? 1'b0 : 
                     (N733)? 1'b0 : 
                     (N734)? 1'b0 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b0 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b0 : 
                     (N741)? 1'b0 : 
                     (N742)? 1'b0 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b0 : 
                     (N745)? 1'b0 : 
                     (N746)? 1'b0 : 
                     (N747)? 1'b0 : 
                     (N748)? 1'b0 : 
                     (N749)? 1'b0 : 
                     (N750)? 1'b0 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b0 : 
                     (N764)? 1'b0 : 
                     (N765)? 1'b0 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[21] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b0 : 
                     (N640)? 1'b0 : 
                     (N641)? 1'b0 : 
                     (N642)? 1'b0 : 
                     (N643)? 1'b0 : 
                     (N644)? 1'b0 : 
                     (N645)? 1'b0 : 
                     (N646)? 1'b0 : 
                     (N647)? 1'b0 : 
                     (N648)? 1'b0 : 
                     (N649)? 1'b0 : 
                     (N650)? 1'b0 : 
                     (N651)? 1'b0 : 
                     (N652)? 1'b0 : 
                     (N653)? 1'b0 : 
                     (N654)? 1'b0 : 
                     (N655)? 1'b0 : 
                     (N656)? 1'b0 : 
                     (N657)? 1'b0 : 
                     (N658)? 1'b0 : 
                     (N659)? 1'b0 : 
                     (N660)? 1'b0 : 
                     (N661)? 1'b0 : 
                     (N662)? 1'b0 : 
                     (N663)? 1'b0 : 
                     (N664)? 1'b0 : 
                     (N665)? 1'b0 : 
                     (N666)? 1'b0 : 
                     (N667)? 1'b0 : 
                     (N668)? 1'b0 : 
                     (N669)? 1'b0 : 
                     (N670)? 1'b0 : 
                     (N671)? 1'b0 : 
                     (N672)? 1'b0 : 
                     (N673)? 1'b0 : 
                     (N674)? 1'b0 : 
                     (N675)? 1'b0 : 
                     (N676)? 1'b0 : 
                     (N677)? 1'b0 : 
                     (N678)? 1'b0 : 
                     (N679)? 1'b0 : 
                     (N680)? 1'b0 : 
                     (N681)? 1'b0 : 
                     (N682)? 1'b0 : 
                     (N683)? 1'b0 : 
                     (N684)? 1'b0 : 
                     (N685)? 1'b0 : 
                     (N686)? 1'b0 : 
                     (N687)? 1'b0 : 
                     (N688)? 1'b0 : 
                     (N689)? 1'b0 : 
                     (N690)? 1'b0 : 
                     (N691)? 1'b0 : 
                     (N692)? 1'b0 : 
                     (N693)? 1'b0 : 
                     (N694)? 1'b0 : 
                     (N695)? 1'b0 : 
                     (N696)? 1'b0 : 
                     (N697)? 1'b0 : 
                     (N698)? 1'b0 : 
                     (N699)? 1'b0 : 
                     (N700)? 1'b0 : 
                     (N701)? 1'b0 : 
                     (N702)? 1'b0 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b0 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b0 : 
                     (N741)? 1'b0 : 
                     (N742)? 1'b0 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b0 : 
                     (N745)? 1'b0 : 
                     (N746)? 1'b0 : 
                     (N747)? 1'b0 : 
                     (N748)? 1'b0 : 
                     (N749)? 1'b0 : 
                     (N750)? 1'b0 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b0 : 
                     (N760)? 1'b0 : 
                     (N761)? 1'b0 : 
                     (N762)? 1'b0 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b0 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[20] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b1 : 
                     (N736)? 1'b1 : 
                     (N737)? 1'b1 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b1 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b1 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b0 : 
                     (N752)? 1'b0 : 
                     (N753)? 1'b0 : 
                     (N754)? 1'b0 : 
                     (N755)? 1'b0 : 
                     (N756)? 1'b0 : 
                     (N757)? 1'b0 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b0 : 
                     (N760)? 1'b0 : 
                     (N761)? 1'b0 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b0 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[19] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b0 : 
                     (N704)? 1'b0 : 
                     (N705)? 1'b0 : 
                     (N706)? 1'b0 : 
                     (N707)? 1'b0 : 
                     (N708)? 1'b0 : 
                     (N709)? 1'b0 : 
                     (N710)? 1'b0 : 
                     (N711)? 1'b0 : 
                     (N712)? 1'b0 : 
                     (N713)? 1'b0 : 
                     (N714)? 1'b0 : 
                     (N715)? 1'b0 : 
                     (N716)? 1'b0 : 
                     (N717)? 1'b0 : 
                     (N718)? 1'b0 : 
                     (N719)? 1'b0 : 
                     (N720)? 1'b0 : 
                     (N721)? 1'b0 : 
                     (N722)? 1'b0 : 
                     (N723)? 1'b0 : 
                     (N724)? 1'b0 : 
                     (N725)? 1'b0 : 
                     (N726)? 1'b0 : 
                     (N727)? 1'b0 : 
                     (N728)? 1'b0 : 
                     (N729)? 1'b0 : 
                     (N730)? 1'b0 : 
                     (N731)? 1'b0 : 
                     (N732)? 1'b0 : 
                     (N733)? 1'b0 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b0 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b0 : 
                     (N741)? 1'b0 : 
                     (N742)? 1'b0 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b0 : 
                     (N745)? 1'b0 : 
                     (N746)? 1'b0 : 
                     (N747)? 1'b0 : 
                     (N748)? 1'b0 : 
                     (N749)? 1'b0 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b0 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[18] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b0 : 
                     (N639)? 1'b0 : 
                     (N640)? 1'b0 : 
                     (N641)? 1'b0 : 
                     (N642)? 1'b0 : 
                     (N643)? 1'b0 : 
                     (N644)? 1'b0 : 
                     (N645)? 1'b0 : 
                     (N646)? 1'b0 : 
                     (N647)? 1'b0 : 
                     (N648)? 1'b0 : 
                     (N649)? 1'b0 : 
                     (N650)? 1'b0 : 
                     (N651)? 1'b0 : 
                     (N652)? 1'b0 : 
                     (N653)? 1'b0 : 
                     (N654)? 1'b0 : 
                     (N655)? 1'b0 : 
                     (N656)? 1'b0 : 
                     (N657)? 1'b0 : 
                     (N658)? 1'b0 : 
                     (N659)? 1'b0 : 
                     (N660)? 1'b0 : 
                     (N661)? 1'b0 : 
                     (N662)? 1'b0 : 
                     (N663)? 1'b0 : 
                     (N664)? 1'b0 : 
                     (N665)? 1'b0 : 
                     (N666)? 1'b0 : 
                     (N667)? 1'b0 : 
                     (N668)? 1'b0 : 
                     (N669)? 1'b0 : 
                     (N670)? 1'b0 : 
                     (N671)? 1'b0 : 
                     (N672)? 1'b0 : 
                     (N673)? 1'b0 : 
                     (N674)? 1'b0 : 
                     (N675)? 1'b0 : 
                     (N676)? 1'b0 : 
                     (N677)? 1'b0 : 
                     (N678)? 1'b0 : 
                     (N679)? 1'b0 : 
                     (N680)? 1'b0 : 
                     (N681)? 1'b0 : 
                     (N682)? 1'b0 : 
                     (N683)? 1'b0 : 
                     (N684)? 1'b0 : 
                     (N685)? 1'b0 : 
                     (N686)? 1'b0 : 
                     (N687)? 1'b0 : 
                     (N688)? 1'b0 : 
                     (N689)? 1'b0 : 
                     (N690)? 1'b0 : 
                     (N691)? 1'b0 : 
                     (N692)? 1'b0 : 
                     (N693)? 1'b0 : 
                     (N694)? 1'b0 : 
                     (N695)? 1'b0 : 
                     (N696)? 1'b0 : 
                     (N697)? 1'b0 : 
                     (N698)? 1'b0 : 
                     (N699)? 1'b0 : 
                     (N700)? 1'b0 : 
                     (N701)? 1'b0 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b0 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b0 : 
                     (N741)? 1'b0 : 
                     (N742)? 1'b0 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b0 : 
                     (N745)? 1'b0 : 
                     (N746)? 1'b0 : 
                     (N747)? 1'b0 : 
                     (N748)? 1'b0 : 
                     (N749)? 1'b0 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b0 : 
                     (N760)? 1'b0 : 
                     (N761)? 1'b0 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b0 : 1'b0;
  assign fwd_o[17] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b1 : 
                     (N736)? 1'b1 : 
                     (N737)? 1'b1 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b1 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b1 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b0 : 
                     (N752)? 1'b0 : 
                     (N753)? 1'b0 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b0 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b0 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[16] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b0 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b0 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b0 : 
                     (N703)? 1'b0 : 
                     (N704)? 1'b0 : 
                     (N705)? 1'b0 : 
                     (N706)? 1'b0 : 
                     (N707)? 1'b0 : 
                     (N708)? 1'b0 : 
                     (N709)? 1'b0 : 
                     (N710)? 1'b0 : 
                     (N711)? 1'b0 : 
                     (N712)? 1'b0 : 
                     (N713)? 1'b0 : 
                     (N714)? 1'b0 : 
                     (N715)? 1'b0 : 
                     (N716)? 1'b0 : 
                     (N717)? 1'b0 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b0 : 
                     (N720)? 1'b0 : 
                     (N721)? 1'b0 : 
                     (N722)? 1'b0 : 
                     (N723)? 1'b0 : 
                     (N724)? 1'b0 : 
                     (N725)? 1'b0 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b0 : 
                     (N728)? 1'b0 : 
                     (N729)? 1'b0 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b0 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b0 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b0 : 
                     (N741)? 1'b0 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b0 : 
                     (N745)? 1'b0 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b0 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b0 : 1'b0;
  assign fwd_o[15] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b0 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b0 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b0 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b0 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b0 : 
                     (N637)? 1'b0 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b0 : 
                     (N640)? 1'b0 : 
                     (N641)? 1'b0 : 
                     (N642)? 1'b0 : 
                     (N643)? 1'b0 : 
                     (N644)? 1'b0 : 
                     (N645)? 1'b0 : 
                     (N646)? 1'b0 : 
                     (N647)? 1'b0 : 
                     (N648)? 1'b0 : 
                     (N649)? 1'b0 : 
                     (N650)? 1'b0 : 
                     (N651)? 1'b0 : 
                     (N652)? 1'b0 : 
                     (N653)? 1'b0 : 
                     (N654)? 1'b0 : 
                     (N655)? 1'b0 : 
                     (N656)? 1'b0 : 
                     (N657)? 1'b0 : 
                     (N658)? 1'b0 : 
                     (N659)? 1'b0 : 
                     (N660)? 1'b0 : 
                     (N661)? 1'b0 : 
                     (N662)? 1'b0 : 
                     (N663)? 1'b0 : 
                     (N664)? 1'b0 : 
                     (N665)? 1'b0 : 
                     (N666)? 1'b0 : 
                     (N667)? 1'b0 : 
                     (N668)? 1'b0 : 
                     (N669)? 1'b0 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b0 : 
                     (N672)? 1'b0 : 
                     (N673)? 1'b0 : 
                     (N674)? 1'b0 : 
                     (N675)? 1'b0 : 
                     (N676)? 1'b0 : 
                     (N677)? 1'b0 : 
                     (N678)? 1'b0 : 
                     (N679)? 1'b0 : 
                     (N680)? 1'b0 : 
                     (N681)? 1'b0 : 
                     (N682)? 1'b0 : 
                     (N683)? 1'b0 : 
                     (N684)? 1'b0 : 
                     (N685)? 1'b0 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b0 : 
                     (N688)? 1'b0 : 
                     (N689)? 1'b0 : 
                     (N690)? 1'b0 : 
                     (N691)? 1'b0 : 
                     (N692)? 1'b0 : 
                     (N693)? 1'b0 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b0 : 
                     (N696)? 1'b0 : 
                     (N697)? 1'b0 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b0 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b0 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b0 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b0 : 
                     (N741)? 1'b0 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b0 : 
                     (N745)? 1'b0 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b0 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b0 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b0 : 
                     (N759)? 1'b0 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b0 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b0 : 
                     (N765)? 1'b0 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[14] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b1 : 
                     (N736)? 1'b1 : 
                     (N737)? 1'b1 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b1 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b1 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b0 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[13] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b0 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b0 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b0 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b0 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b0 : 
                     (N573)? 1'b0 : 
                     (N574)? 1'b0 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b0 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b0 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b0 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b0 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b0 : 
                     (N637)? 1'b0 : 
                     (N638)? 1'b0 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b0 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b0 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b0 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b0 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b0 : 
                     (N701)? 1'b0 : 
                     (N702)? 1'b0 : 
                     (N703)? 1'b0 : 
                     (N704)? 1'b0 : 
                     (N705)? 1'b0 : 
                     (N706)? 1'b0 : 
                     (N707)? 1'b0 : 
                     (N708)? 1'b0 : 
                     (N709)? 1'b0 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b0 : 
                     (N712)? 1'b0 : 
                     (N713)? 1'b0 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b0 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b0 : 
                     (N720)? 1'b0 : 
                     (N721)? 1'b0 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b0 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b0 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b0 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b0 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b0 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b0 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b0 : 
                     (N765)? 1'b0 : 
                     (N255)? 1'b0 : 1'b0;
  assign fwd_o[12] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b0 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b0 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b0 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b0 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b0 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b0 : 
                     (N605)? 1'b0 : 
                     (N606)? 1'b0 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b0 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b0 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b0 : 
                     (N621)? 1'b0 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b0 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b0 : 
                     (N629)? 1'b0 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b0 : 
                     (N633)? 1'b0 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b0 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b0 : 
                     (N639)? 1'b0 : 
                     (N640)? 1'b0 : 
                     (N641)? 1'b0 : 
                     (N642)? 1'b0 : 
                     (N643)? 1'b0 : 
                     (N644)? 1'b0 : 
                     (N645)? 1'b0 : 
                     (N646)? 1'b0 : 
                     (N647)? 1'b0 : 
                     (N648)? 1'b0 : 
                     (N649)? 1'b0 : 
                     (N650)? 1'b0 : 
                     (N651)? 1'b0 : 
                     (N652)? 1'b0 : 
                     (N653)? 1'b0 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b0 : 
                     (N656)? 1'b0 : 
                     (N657)? 1'b0 : 
                     (N658)? 1'b0 : 
                     (N659)? 1'b0 : 
                     (N660)? 1'b0 : 
                     (N661)? 1'b0 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b0 : 
                     (N664)? 1'b0 : 
                     (N665)? 1'b0 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b0 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b0 : 
                     (N671)? 1'b0 : 
                     (N672)? 1'b0 : 
                     (N673)? 1'b0 : 
                     (N674)? 1'b0 : 
                     (N675)? 1'b0 : 
                     (N676)? 1'b0 : 
                     (N677)? 1'b0 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b0 : 
                     (N680)? 1'b0 : 
                     (N681)? 1'b0 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b0 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b0 : 
                     (N688)? 1'b0 : 
                     (N689)? 1'b0 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b0 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b0 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b0 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b0 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b0 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b0 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b0 : 
                     (N733)? 1'b0 : 
                     (N734)? 1'b0 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b0 : 
                     (N737)? 1'b0 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b0 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b0 : 
                     (N743)? 1'b0 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b0 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b0 : 
                     (N749)? 1'b0 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b0 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b0 : 
                     (N757)? 1'b0 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b0 : 
                     (N761)? 1'b0 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b0 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b0 : 1'b0;
  assign fwd_o[11] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b0 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b1 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b1 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b1 : 
                     (N541)? 1'b1 : 
                     (N542)? 1'b0 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b1 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b1 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b1 : 
                     (N557)? 1'b1 : 
                     (N558)? 1'b0 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b1 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b1 : 
                     (N565)? 1'b1 : 
                     (N566)? 1'b1 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b1 : 
                     (N569)? 1'b1 : 
                     (N570)? 1'b1 : 
                     (N571)? 1'b1 : 
                     (N572)? 1'b1 : 
                     (N573)? 1'b1 : 
                     (N574)? 1'b0 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b0 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b1 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b1 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b1 : 
                     (N605)? 1'b1 : 
                     (N606)? 1'b0 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b1 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b1 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b1 : 
                     (N621)? 1'b1 : 
                     (N622)? 1'b0 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b1 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b1 : 
                     (N629)? 1'b1 : 
                     (N630)? 1'b1 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b1 : 
                     (N633)? 1'b1 : 
                     (N634)? 1'b1 : 
                     (N635)? 1'b1 : 
                     (N636)? 1'b1 : 
                     (N637)? 1'b1 : 
                     (N638)? 1'b0 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b0 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b1 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b1 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b1 : 
                     (N669)? 1'b1 : 
                     (N670)? 1'b0 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b1 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b1 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b1 : 
                     (N685)? 1'b1 : 
                     (N686)? 1'b0 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b1 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b1 : 
                     (N693)? 1'b1 : 
                     (N694)? 1'b1 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b1 : 
                     (N697)? 1'b1 : 
                     (N698)? 1'b1 : 
                     (N699)? 1'b1 : 
                     (N700)? 1'b1 : 
                     (N701)? 1'b1 : 
                     (N702)? 1'b0 : 
                     (N703)? 1'b1 : 
                     (N704)? 1'b1 : 
                     (N705)? 1'b1 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b1 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b1 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b0 : 
                     (N719)? 1'b1 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b1 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b1 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b1 : 
                     (N733)? 1'b1 : 
                     (N734)? 1'b0 : 
                     (N735)? 1'b1 : 
                     (N736)? 1'b1 : 
                     (N737)? 1'b1 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b1 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b1 : 
                     (N743)? 1'b1 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b1 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b1 : 
                     (N749)? 1'b1 : 
                     (N750)? 1'b0 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b1 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b1 : 
                     (N757)? 1'b1 : 
                     (N758)? 1'b1 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b1 : 
                     (N761)? 1'b1 : 
                     (N762)? 1'b1 : 
                     (N763)? 1'b1 : 
                     (N764)? 1'b1 : 
                     (N765)? 1'b1 : 
                     (N255)? 1'b0 : 1'b0;
  assign fwd_o[10] = (N511)? 1'b1 : 
                     (N512)? 1'b1 : 
                     (N513)? 1'b1 : 
                     (N514)? 1'b1 : 
                     (N515)? 1'b1 : 
                     (N516)? 1'b1 : 
                     (N517)? 1'b1 : 
                     (N518)? 1'b1 : 
                     (N519)? 1'b1 : 
                     (N520)? 1'b1 : 
                     (N521)? 1'b1 : 
                     (N522)? 1'b1 : 
                     (N523)? 1'b1 : 
                     (N524)? 1'b1 : 
                     (N525)? 1'b1 : 
                     (N526)? 1'b1 : 
                     (N527)? 1'b1 : 
                     (N528)? 1'b1 : 
                     (N529)? 1'b1 : 
                     (N530)? 1'b1 : 
                     (N531)? 1'b1 : 
                     (N532)? 1'b1 : 
                     (N533)? 1'b1 : 
                     (N534)? 1'b0 : 
                     (N535)? 1'b1 : 
                     (N536)? 1'b1 : 
                     (N537)? 1'b1 : 
                     (N538)? 1'b0 : 
                     (N539)? 1'b1 : 
                     (N540)? 1'b0 : 
                     (N541)? 1'b0 : 
                     (N542)? 1'b1 : 
                     (N543)? 1'b1 : 
                     (N544)? 1'b1 : 
                     (N545)? 1'b1 : 
                     (N546)? 1'b1 : 
                     (N547)? 1'b1 : 
                     (N548)? 1'b1 : 
                     (N549)? 1'b1 : 
                     (N550)? 1'b0 : 
                     (N551)? 1'b1 : 
                     (N552)? 1'b1 : 
                     (N553)? 1'b1 : 
                     (N554)? 1'b0 : 
                     (N555)? 1'b1 : 
                     (N556)? 1'b0 : 
                     (N557)? 1'b0 : 
                     (N558)? 1'b1 : 
                     (N559)? 1'b1 : 
                     (N560)? 1'b1 : 
                     (N561)? 1'b1 : 
                     (N562)? 1'b0 : 
                     (N563)? 1'b1 : 
                     (N564)? 1'b0 : 
                     (N565)? 1'b0 : 
                     (N566)? 1'b0 : 
                     (N567)? 1'b1 : 
                     (N568)? 1'b0 : 
                     (N569)? 1'b0 : 
                     (N570)? 1'b0 : 
                     (N571)? 1'b0 : 
                     (N572)? 1'b0 : 
                     (N573)? 1'b0 : 
                     (N574)? 1'b1 : 
                     (N575)? 1'b1 : 
                     (N576)? 1'b1 : 
                     (N577)? 1'b1 : 
                     (N578)? 1'b1 : 
                     (N579)? 1'b1 : 
                     (N580)? 1'b1 : 
                     (N581)? 1'b1 : 
                     (N582)? 1'b1 : 
                     (N583)? 1'b1 : 
                     (N584)? 1'b1 : 
                     (N585)? 1'b1 : 
                     (N586)? 1'b1 : 
                     (N587)? 1'b1 : 
                     (N588)? 1'b1 : 
                     (N589)? 1'b1 : 
                     (N590)? 1'b1 : 
                     (N591)? 1'b1 : 
                     (N592)? 1'b1 : 
                     (N593)? 1'b1 : 
                     (N594)? 1'b1 : 
                     (N595)? 1'b1 : 
                     (N596)? 1'b1 : 
                     (N597)? 1'b1 : 
                     (N598)? 1'b0 : 
                     (N599)? 1'b1 : 
                     (N600)? 1'b1 : 
                     (N601)? 1'b1 : 
                     (N602)? 1'b0 : 
                     (N603)? 1'b1 : 
                     (N604)? 1'b0 : 
                     (N605)? 1'b0 : 
                     (N606)? 1'b1 : 
                     (N607)? 1'b1 : 
                     (N608)? 1'b1 : 
                     (N609)? 1'b1 : 
                     (N610)? 1'b1 : 
                     (N611)? 1'b1 : 
                     (N612)? 1'b1 : 
                     (N613)? 1'b1 : 
                     (N614)? 1'b0 : 
                     (N615)? 1'b1 : 
                     (N616)? 1'b1 : 
                     (N617)? 1'b1 : 
                     (N618)? 1'b0 : 
                     (N619)? 1'b1 : 
                     (N620)? 1'b0 : 
                     (N621)? 1'b0 : 
                     (N622)? 1'b1 : 
                     (N623)? 1'b1 : 
                     (N624)? 1'b1 : 
                     (N625)? 1'b1 : 
                     (N626)? 1'b0 : 
                     (N627)? 1'b1 : 
                     (N628)? 1'b0 : 
                     (N629)? 1'b0 : 
                     (N630)? 1'b0 : 
                     (N631)? 1'b1 : 
                     (N632)? 1'b0 : 
                     (N633)? 1'b0 : 
                     (N634)? 1'b0 : 
                     (N635)? 1'b0 : 
                     (N636)? 1'b0 : 
                     (N637)? 1'b0 : 
                     (N638)? 1'b1 : 
                     (N639)? 1'b1 : 
                     (N640)? 1'b1 : 
                     (N641)? 1'b1 : 
                     (N642)? 1'b1 : 
                     (N643)? 1'b1 : 
                     (N644)? 1'b1 : 
                     (N645)? 1'b1 : 
                     (N646)? 1'b1 : 
                     (N647)? 1'b1 : 
                     (N648)? 1'b1 : 
                     (N649)? 1'b1 : 
                     (N650)? 1'b1 : 
                     (N651)? 1'b1 : 
                     (N652)? 1'b1 : 
                     (N653)? 1'b1 : 
                     (N654)? 1'b1 : 
                     (N655)? 1'b1 : 
                     (N656)? 1'b1 : 
                     (N657)? 1'b1 : 
                     (N658)? 1'b1 : 
                     (N659)? 1'b1 : 
                     (N660)? 1'b1 : 
                     (N661)? 1'b1 : 
                     (N662)? 1'b0 : 
                     (N663)? 1'b1 : 
                     (N664)? 1'b1 : 
                     (N665)? 1'b1 : 
                     (N666)? 1'b0 : 
                     (N667)? 1'b1 : 
                     (N668)? 1'b0 : 
                     (N669)? 1'b0 : 
                     (N670)? 1'b1 : 
                     (N671)? 1'b1 : 
                     (N672)? 1'b1 : 
                     (N673)? 1'b1 : 
                     (N674)? 1'b1 : 
                     (N675)? 1'b1 : 
                     (N676)? 1'b1 : 
                     (N677)? 1'b1 : 
                     (N678)? 1'b0 : 
                     (N679)? 1'b1 : 
                     (N680)? 1'b1 : 
                     (N681)? 1'b1 : 
                     (N682)? 1'b0 : 
                     (N683)? 1'b1 : 
                     (N684)? 1'b0 : 
                     (N685)? 1'b0 : 
                     (N686)? 1'b1 : 
                     (N687)? 1'b1 : 
                     (N688)? 1'b1 : 
                     (N689)? 1'b1 : 
                     (N690)? 1'b0 : 
                     (N691)? 1'b1 : 
                     (N692)? 1'b0 : 
                     (N693)? 1'b0 : 
                     (N694)? 1'b0 : 
                     (N695)? 1'b1 : 
                     (N696)? 1'b0 : 
                     (N697)? 1'b0 : 
                     (N698)? 1'b0 : 
                     (N699)? 1'b0 : 
                     (N700)? 1'b0 : 
                     (N701)? 1'b0 : 
                     (N702)? 1'b1 : 
                     (N703)? 1'b0 : 
                     (N704)? 1'b0 : 
                     (N705)? 1'b0 : 
                     (N706)? 1'b1 : 
                     (N707)? 1'b0 : 
                     (N708)? 1'b1 : 
                     (N709)? 1'b1 : 
                     (N710)? 1'b1 : 
                     (N711)? 1'b0 : 
                     (N712)? 1'b1 : 
                     (N713)? 1'b1 : 
                     (N714)? 1'b1 : 
                     (N715)? 1'b1 : 
                     (N716)? 1'b1 : 
                     (N717)? 1'b1 : 
                     (N718)? 1'b1 : 
                     (N719)? 1'b0 : 
                     (N720)? 1'b1 : 
                     (N721)? 1'b1 : 
                     (N722)? 1'b1 : 
                     (N723)? 1'b1 : 
                     (N724)? 1'b1 : 
                     (N725)? 1'b1 : 
                     (N726)? 1'b0 : 
                     (N727)? 1'b1 : 
                     (N728)? 1'b1 : 
                     (N729)? 1'b1 : 
                     (N730)? 1'b0 : 
                     (N731)? 1'b1 : 
                     (N732)? 1'b0 : 
                     (N733)? 1'b0 : 
                     (N734)? 1'b1 : 
                     (N735)? 1'b0 : 
                     (N736)? 1'b1 : 
                     (N737)? 1'b1 : 
                     (N738)? 1'b1 : 
                     (N739)? 1'b1 : 
                     (N740)? 1'b1 : 
                     (N741)? 1'b1 : 
                     (N742)? 1'b0 : 
                     (N743)? 1'b1 : 
                     (N744)? 1'b1 : 
                     (N745)? 1'b1 : 
                     (N746)? 1'b0 : 
                     (N747)? 1'b1 : 
                     (N748)? 1'b0 : 
                     (N749)? 1'b0 : 
                     (N750)? 1'b1 : 
                     (N751)? 1'b1 : 
                     (N752)? 1'b1 : 
                     (N753)? 1'b1 : 
                     (N754)? 1'b0 : 
                     (N755)? 1'b1 : 
                     (N756)? 1'b0 : 
                     (N757)? 1'b0 : 
                     (N758)? 1'b0 : 
                     (N759)? 1'b1 : 
                     (N760)? 1'b0 : 
                     (N761)? 1'b0 : 
                     (N762)? 1'b0 : 
                     (N763)? 1'b0 : 
                     (N764)? 1'b0 : 
                     (N765)? 1'b0 : 
                     (N255)? 1'b1 : 1'b0;
  assign fwd_o[9] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b1 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b1 : 
                    (N517)? 1'b1 : 
                    (N518)? 1'b1 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b1 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b1 : 
                    (N523)? 1'b1 : 
                    (N524)? 1'b1 : 
                    (N525)? 1'b1 : 
                    (N526)? 1'b1 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b1 : 
                    (N529)? 1'b1 : 
                    (N530)? 1'b1 : 
                    (N531)? 1'b1 : 
                    (N532)? 1'b1 : 
                    (N533)? 1'b1 : 
                    (N534)? 1'b0 : 
                    (N535)? 1'b1 : 
                    (N536)? 1'b1 : 
                    (N537)? 1'b1 : 
                    (N538)? 1'b0 : 
                    (N539)? 1'b1 : 
                    (N540)? 1'b0 : 
                    (N541)? 1'b0 : 
                    (N542)? 1'b1 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b1 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b1 : 
                    (N547)? 1'b1 : 
                    (N548)? 1'b1 : 
                    (N549)? 1'b1 : 
                    (N550)? 1'b1 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N553)? 1'b1 : 
                    (N554)? 1'b1 : 
                    (N555)? 1'b1 : 
                    (N556)? 1'b1 : 
                    (N557)? 1'b1 : 
                    (N558)? 1'b1 : 
                    (N559)? 1'b1 : 
                    (N560)? 1'b1 : 
                    (N561)? 1'b1 : 
                    (N562)? 1'b1 : 
                    (N563)? 1'b1 : 
                    (N564)? 1'b1 : 
                    (N565)? 1'b1 : 
                    (N566)? 1'b0 : 
                    (N567)? 1'b1 : 
                    (N568)? 1'b1 : 
                    (N569)? 1'b1 : 
                    (N570)? 1'b0 : 
                    (N571)? 1'b1 : 
                    (N572)? 1'b0 : 
                    (N573)? 1'b0 : 
                    (N574)? 1'b1 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b1 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b1 : 
                    (N579)? 1'b1 : 
                    (N580)? 1'b1 : 
                    (N581)? 1'b1 : 
                    (N582)? 1'b0 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b1 : 
                    (N585)? 1'b1 : 
                    (N586)? 1'b0 : 
                    (N587)? 1'b1 : 
                    (N588)? 1'b0 : 
                    (N589)? 1'b0 : 
                    (N590)? 1'b1 : 
                    (N591)? 1'b1 : 
                    (N592)? 1'b1 : 
                    (N593)? 1'b1 : 
                    (N594)? 1'b0 : 
                    (N595)? 1'b1 : 
                    (N596)? 1'b0 : 
                    (N597)? 1'b0 : 
                    (N598)? 1'b0 : 
                    (N599)? 1'b1 : 
                    (N600)? 1'b0 : 
                    (N601)? 1'b0 : 
                    (N602)? 1'b0 : 
                    (N603)? 1'b0 : 
                    (N604)? 1'b0 : 
                    (N605)? 1'b0 : 
                    (N606)? 1'b1 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b1 : 
                    (N609)? 1'b1 : 
                    (N610)? 1'b0 : 
                    (N611)? 1'b1 : 
                    (N612)? 1'b0 : 
                    (N613)? 1'b0 : 
                    (N614)? 1'b1 : 
                    (N615)? 1'b1 : 
                    (N616)? 1'b0 : 
                    (N617)? 1'b0 : 
                    (N618)? 1'b1 : 
                    (N619)? 1'b0 : 
                    (N620)? 1'b1 : 
                    (N621)? 1'b1 : 
                    (N622)? 1'b1 : 
                    (N623)? 1'b1 : 
                    (N624)? 1'b0 : 
                    (N625)? 1'b0 : 
                    (N626)? 1'b1 : 
                    (N627)? 1'b0 : 
                    (N628)? 1'b1 : 
                    (N629)? 1'b1 : 
                    (N630)? 1'b0 : 
                    (N631)? 1'b0 : 
                    (N632)? 1'b1 : 
                    (N633)? 1'b1 : 
                    (N634)? 1'b0 : 
                    (N635)? 1'b1 : 
                    (N636)? 1'b0 : 
                    (N637)? 1'b0 : 
                    (N638)? 1'b1 : 
                    (N639)? 1'b0 : 
                    (N640)? 1'b0 : 
                    (N641)? 1'b0 : 
                    (N642)? 1'b0 : 
                    (N643)? 1'b0 : 
                    (N644)? 1'b0 : 
                    (N645)? 1'b0 : 
                    (N646)? 1'b1 : 
                    (N647)? 1'b0 : 
                    (N648)? 1'b0 : 
                    (N649)? 1'b0 : 
                    (N650)? 1'b1 : 
                    (N651)? 1'b0 : 
                    (N652)? 1'b1 : 
                    (N653)? 1'b1 : 
                    (N654)? 1'b1 : 
                    (N655)? 1'b0 : 
                    (N656)? 1'b0 : 
                    (N657)? 1'b0 : 
                    (N658)? 1'b1 : 
                    (N659)? 1'b0 : 
                    (N660)? 1'b1 : 
                    (N661)? 1'b1 : 
                    (N662)? 1'b0 : 
                    (N663)? 1'b0 : 
                    (N664)? 1'b1 : 
                    (N665)? 1'b1 : 
                    (N666)? 1'b0 : 
                    (N667)? 1'b1 : 
                    (N668)? 1'b0 : 
                    (N669)? 1'b0 : 
                    (N670)? 1'b1 : 
                    (N671)? 1'b0 : 
                    (N672)? 1'b0 : 
                    (N673)? 1'b0 : 
                    (N674)? 1'b1 : 
                    (N675)? 1'b0 : 
                    (N676)? 1'b1 : 
                    (N677)? 1'b1 : 
                    (N678)? 1'b1 : 
                    (N679)? 1'b0 : 
                    (N680)? 1'b1 : 
                    (N681)? 1'b1 : 
                    (N682)? 1'b1 : 
                    (N683)? 1'b1 : 
                    (N684)? 1'b1 : 
                    (N685)? 1'b1 : 
                    (N686)? 1'b1 : 
                    (N687)? 1'b0 : 
                    (N688)? 1'b1 : 
                    (N689)? 1'b1 : 
                    (N690)? 1'b1 : 
                    (N691)? 1'b1 : 
                    (N692)? 1'b1 : 
                    (N693)? 1'b1 : 
                    (N694)? 1'b0 : 
                    (N695)? 1'b1 : 
                    (N696)? 1'b1 : 
                    (N697)? 1'b1 : 
                    (N698)? 1'b0 : 
                    (N699)? 1'b1 : 
                    (N700)? 1'b0 : 
                    (N701)? 1'b0 : 
                    (N702)? 1'b1 : 
                    (N703)? 1'b1 : 
                    (N704)? 1'b1 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b1 : 
                    (N707)? 1'b1 : 
                    (N708)? 1'b1 : 
                    (N709)? 1'b1 : 
                    (N710)? 1'b0 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b1 : 
                    (N713)? 1'b1 : 
                    (N714)? 1'b0 : 
                    (N715)? 1'b1 : 
                    (N716)? 1'b0 : 
                    (N717)? 1'b0 : 
                    (N718)? 1'b1 : 
                    (N719)? 1'b1 : 
                    (N720)? 1'b1 : 
                    (N721)? 1'b1 : 
                    (N722)? 1'b0 : 
                    (N723)? 1'b1 : 
                    (N724)? 1'b0 : 
                    (N725)? 1'b0 : 
                    (N726)? 1'b0 : 
                    (N727)? 1'b1 : 
                    (N728)? 1'b0 : 
                    (N729)? 1'b0 : 
                    (N730)? 1'b0 : 
                    (N731)? 1'b0 : 
                    (N732)? 1'b0 : 
                    (N733)? 1'b0 : 
                    (N734)? 1'b1 : 
                    (N735)? 1'b0 : 
                    (N736)? 1'b1 : 
                    (N737)? 1'b1 : 
                    (N738)? 1'b0 : 
                    (N739)? 1'b1 : 
                    (N740)? 1'b0 : 
                    (N741)? 1'b0 : 
                    (N742)? 1'b1 : 
                    (N743)? 1'b1 : 
                    (N744)? 1'b0 : 
                    (N745)? 1'b0 : 
                    (N746)? 1'b1 : 
                    (N747)? 1'b0 : 
                    (N748)? 1'b1 : 
                    (N749)? 1'b1 : 
                    (N750)? 1'b1 : 
                    (N751)? 1'b1 : 
                    (N752)? 1'b0 : 
                    (N753)? 1'b0 : 
                    (N754)? 1'b1 : 
                    (N755)? 1'b0 : 
                    (N756)? 1'b1 : 
                    (N757)? 1'b1 : 
                    (N758)? 1'b0 : 
                    (N759)? 1'b0 : 
                    (N760)? 1'b1 : 
                    (N761)? 1'b1 : 
                    (N762)? 1'b0 : 
                    (N763)? 1'b1 : 
                    (N764)? 1'b0 : 
                    (N765)? 1'b0 : 
                    (N255)? 1'b1 : 1'b0;
  assign fwd_o[8] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b1 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b1 : 
                    (N517)? 1'b1 : 
                    (N518)? 1'b0 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b1 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b0 : 
                    (N523)? 1'b1 : 
                    (N524)? 1'b0 : 
                    (N525)? 1'b0 : 
                    (N526)? 1'b0 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b1 : 
                    (N529)? 1'b1 : 
                    (N530)? 1'b1 : 
                    (N531)? 1'b1 : 
                    (N532)? 1'b1 : 
                    (N533)? 1'b1 : 
                    (N534)? 1'b0 : 
                    (N535)? 1'b1 : 
                    (N536)? 1'b1 : 
                    (N537)? 1'b1 : 
                    (N538)? 1'b0 : 
                    (N539)? 1'b1 : 
                    (N540)? 1'b0 : 
                    (N541)? 1'b0 : 
                    (N542)? 1'b0 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b1 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b1 : 
                    (N547)? 1'b1 : 
                    (N548)? 1'b1 : 
                    (N549)? 1'b1 : 
                    (N550)? 1'b0 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N553)? 1'b1 : 
                    (N554)? 1'b0 : 
                    (N555)? 1'b1 : 
                    (N556)? 1'b0 : 
                    (N557)? 1'b0 : 
                    (N558)? 1'b0 : 
                    (N559)? 1'b1 : 
                    (N560)? 1'b1 : 
                    (N561)? 1'b1 : 
                    (N562)? 1'b1 : 
                    (N563)? 1'b1 : 
                    (N564)? 1'b1 : 
                    (N565)? 1'b1 : 
                    (N566)? 1'b0 : 
                    (N567)? 1'b1 : 
                    (N568)? 1'b1 : 
                    (N569)? 1'b1 : 
                    (N570)? 1'b0 : 
                    (N571)? 1'b1 : 
                    (N572)? 1'b0 : 
                    (N573)? 1'b0 : 
                    (N574)? 1'b0 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b1 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b1 : 
                    (N579)? 1'b1 : 
                    (N580)? 1'b1 : 
                    (N581)? 1'b1 : 
                    (N582)? 1'b0 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b1 : 
                    (N585)? 1'b1 : 
                    (N586)? 1'b0 : 
                    (N587)? 1'b1 : 
                    (N588)? 1'b0 : 
                    (N589)? 1'b0 : 
                    (N590)? 1'b0 : 
                    (N591)? 1'b1 : 
                    (N592)? 1'b1 : 
                    (N593)? 1'b1 : 
                    (N594)? 1'b1 : 
                    (N595)? 1'b1 : 
                    (N596)? 1'b1 : 
                    (N597)? 1'b1 : 
                    (N598)? 1'b0 : 
                    (N599)? 1'b1 : 
                    (N600)? 1'b1 : 
                    (N601)? 1'b1 : 
                    (N602)? 1'b0 : 
                    (N603)? 1'b1 : 
                    (N604)? 1'b0 : 
                    (N605)? 1'b0 : 
                    (N606)? 1'b0 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b1 : 
                    (N609)? 1'b1 : 
                    (N610)? 1'b1 : 
                    (N611)? 1'b1 : 
                    (N612)? 1'b1 : 
                    (N613)? 1'b1 : 
                    (N614)? 1'b0 : 
                    (N615)? 1'b1 : 
                    (N616)? 1'b1 : 
                    (N617)? 1'b1 : 
                    (N618)? 1'b0 : 
                    (N619)? 1'b1 : 
                    (N620)? 1'b0 : 
                    (N621)? 1'b0 : 
                    (N622)? 1'b0 : 
                    (N623)? 1'b1 : 
                    (N624)? 1'b1 : 
                    (N625)? 1'b1 : 
                    (N626)? 1'b1 : 
                    (N627)? 1'b1 : 
                    (N628)? 1'b1 : 
                    (N629)? 1'b1 : 
                    (N630)? 1'b0 : 
                    (N631)? 1'b1 : 
                    (N632)? 1'b1 : 
                    (N633)? 1'b1 : 
                    (N634)? 1'b0 : 
                    (N635)? 1'b1 : 
                    (N636)? 1'b0 : 
                    (N637)? 1'b0 : 
                    (N638)? 1'b0 : 
                    (N639)? 1'b1 : 
                    (N640)? 1'b1 : 
                    (N641)? 1'b1 : 
                    (N642)? 1'b1 : 
                    (N643)? 1'b1 : 
                    (N644)? 1'b1 : 
                    (N645)? 1'b1 : 
                    (N646)? 1'b0 : 
                    (N647)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N649)? 1'b1 : 
                    (N650)? 1'b0 : 
                    (N651)? 1'b1 : 
                    (N652)? 1'b0 : 
                    (N653)? 1'b0 : 
                    (N654)? 1'b0 : 
                    (N655)? 1'b1 : 
                    (N656)? 1'b1 : 
                    (N657)? 1'b1 : 
                    (N658)? 1'b1 : 
                    (N659)? 1'b1 : 
                    (N660)? 1'b1 : 
                    (N661)? 1'b1 : 
                    (N662)? 1'b0 : 
                    (N663)? 1'b1 : 
                    (N664)? 1'b1 : 
                    (N665)? 1'b1 : 
                    (N666)? 1'b0 : 
                    (N667)? 1'b1 : 
                    (N668)? 1'b0 : 
                    (N669)? 1'b0 : 
                    (N670)? 1'b0 : 
                    (N671)? 1'b1 : 
                    (N672)? 1'b1 : 
                    (N673)? 1'b1 : 
                    (N674)? 1'b1 : 
                    (N675)? 1'b1 : 
                    (N676)? 1'b1 : 
                    (N677)? 1'b1 : 
                    (N678)? 1'b0 : 
                    (N679)? 1'b1 : 
                    (N680)? 1'b1 : 
                    (N681)? 1'b1 : 
                    (N682)? 1'b0 : 
                    (N683)? 1'b1 : 
                    (N684)? 1'b0 : 
                    (N685)? 1'b0 : 
                    (N686)? 1'b0 : 
                    (N687)? 1'b1 : 
                    (N688)? 1'b1 : 
                    (N689)? 1'b1 : 
                    (N690)? 1'b1 : 
                    (N691)? 1'b1 : 
                    (N692)? 1'b1 : 
                    (N693)? 1'b1 : 
                    (N694)? 1'b0 : 
                    (N695)? 1'b1 : 
                    (N696)? 1'b1 : 
                    (N697)? 1'b1 : 
                    (N698)? 1'b0 : 
                    (N699)? 1'b1 : 
                    (N700)? 1'b0 : 
                    (N701)? 1'b0 : 
                    (N702)? 1'b0 : 
                    (N703)? 1'b1 : 
                    (N704)? 1'b1 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b1 : 
                    (N707)? 1'b1 : 
                    (N708)? 1'b1 : 
                    (N709)? 1'b1 : 
                    (N710)? 1'b0 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b1 : 
                    (N713)? 1'b1 : 
                    (N714)? 1'b0 : 
                    (N715)? 1'b1 : 
                    (N716)? 1'b0 : 
                    (N717)? 1'b0 : 
                    (N718)? 1'b0 : 
                    (N719)? 1'b1 : 
                    (N720)? 1'b1 : 
                    (N721)? 1'b1 : 
                    (N722)? 1'b1 : 
                    (N723)? 1'b1 : 
                    (N724)? 1'b1 : 
                    (N725)? 1'b1 : 
                    (N726)? 1'b0 : 
                    (N727)? 1'b1 : 
                    (N728)? 1'b1 : 
                    (N729)? 1'b1 : 
                    (N730)? 1'b0 : 
                    (N731)? 1'b1 : 
                    (N732)? 1'b0 : 
                    (N733)? 1'b0 : 
                    (N734)? 1'b0 : 
                    (N735)? 1'b1 : 
                    (N736)? 1'b1 : 
                    (N737)? 1'b1 : 
                    (N738)? 1'b1 : 
                    (N739)? 1'b1 : 
                    (N740)? 1'b1 : 
                    (N741)? 1'b1 : 
                    (N742)? 1'b0 : 
                    (N743)? 1'b1 : 
                    (N744)? 1'b1 : 
                    (N745)? 1'b1 : 
                    (N746)? 1'b0 : 
                    (N747)? 1'b1 : 
                    (N748)? 1'b0 : 
                    (N749)? 1'b0 : 
                    (N750)? 1'b0 : 
                    (N751)? 1'b1 : 
                    (N752)? 1'b1 : 
                    (N753)? 1'b1 : 
                    (N754)? 1'b1 : 
                    (N755)? 1'b1 : 
                    (N756)? 1'b1 : 
                    (N757)? 1'b1 : 
                    (N758)? 1'b0 : 
                    (N759)? 1'b1 : 
                    (N760)? 1'b1 : 
                    (N761)? 1'b1 : 
                    (N762)? 1'b0 : 
                    (N763)? 1'b1 : 
                    (N764)? 1'b0 : 
                    (N765)? 1'b0 : 
                    (N255)? 1'b0 : 1'b0;
  assign fwd_o[7] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b1 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b1 : 
                    (N517)? 1'b1 : 
                    (N518)? 1'b1 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b1 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b1 : 
                    (N523)? 1'b1 : 
                    (N524)? 1'b1 : 
                    (N525)? 1'b1 : 
                    (N526)? 1'b1 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b1 : 
                    (N529)? 1'b1 : 
                    (N530)? 1'b0 : 
                    (N531)? 1'b1 : 
                    (N532)? 1'b0 : 
                    (N533)? 1'b0 : 
                    (N534)? 1'b1 : 
                    (N535)? 1'b1 : 
                    (N536)? 1'b0 : 
                    (N537)? 1'b0 : 
                    (N538)? 1'b1 : 
                    (N539)? 1'b0 : 
                    (N540)? 1'b1 : 
                    (N541)? 1'b1 : 
                    (N542)? 1'b1 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b1 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b0 : 
                    (N547)? 1'b1 : 
                    (N548)? 1'b0 : 
                    (N549)? 1'b0 : 
                    (N550)? 1'b1 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b0 : 
                    (N553)? 1'b0 : 
                    (N554)? 1'b1 : 
                    (N555)? 1'b0 : 
                    (N556)? 1'b1 : 
                    (N557)? 1'b1 : 
                    (N558)? 1'b1 : 
                    (N559)? 1'b1 : 
                    (N560)? 1'b0 : 
                    (N561)? 1'b0 : 
                    (N562)? 1'b0 : 
                    (N563)? 1'b0 : 
                    (N564)? 1'b0 : 
                    (N565)? 1'b0 : 
                    (N566)? 1'b1 : 
                    (N567)? 1'b0 : 
                    (N568)? 1'b0 : 
                    (N569)? 1'b0 : 
                    (N570)? 1'b1 : 
                    (N571)? 1'b0 : 
                    (N572)? 1'b1 : 
                    (N573)? 1'b1 : 
                    (N574)? 1'b1 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b1 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b1 : 
                    (N579)? 1'b1 : 
                    (N580)? 1'b1 : 
                    (N581)? 1'b1 : 
                    (N582)? 1'b1 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b1 : 
                    (N585)? 1'b1 : 
                    (N586)? 1'b1 : 
                    (N587)? 1'b1 : 
                    (N588)? 1'b1 : 
                    (N589)? 1'b1 : 
                    (N590)? 1'b1 : 
                    (N591)? 1'b1 : 
                    (N592)? 1'b1 : 
                    (N593)? 1'b1 : 
                    (N594)? 1'b0 : 
                    (N595)? 1'b1 : 
                    (N596)? 1'b0 : 
                    (N597)? 1'b0 : 
                    (N598)? 1'b1 : 
                    (N599)? 1'b1 : 
                    (N600)? 1'b0 : 
                    (N601)? 1'b0 : 
                    (N602)? 1'b1 : 
                    (N603)? 1'b0 : 
                    (N604)? 1'b1 : 
                    (N605)? 1'b1 : 
                    (N606)? 1'b1 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b1 : 
                    (N609)? 1'b1 : 
                    (N610)? 1'b0 : 
                    (N611)? 1'b1 : 
                    (N612)? 1'b0 : 
                    (N613)? 1'b0 : 
                    (N614)? 1'b1 : 
                    (N615)? 1'b1 : 
                    (N616)? 1'b0 : 
                    (N617)? 1'b0 : 
                    (N618)? 1'b1 : 
                    (N619)? 1'b0 : 
                    (N620)? 1'b1 : 
                    (N621)? 1'b1 : 
                    (N622)? 1'b1 : 
                    (N623)? 1'b1 : 
                    (N624)? 1'b0 : 
                    (N625)? 1'b0 : 
                    (N626)? 1'b0 : 
                    (N627)? 1'b0 : 
                    (N628)? 1'b0 : 
                    (N629)? 1'b0 : 
                    (N630)? 1'b1 : 
                    (N631)? 1'b0 : 
                    (N632)? 1'b0 : 
                    (N633)? 1'b0 : 
                    (N634)? 1'b1 : 
                    (N635)? 1'b0 : 
                    (N636)? 1'b1 : 
                    (N637)? 1'b1 : 
                    (N638)? 1'b1 : 
                    (N639)? 1'b1 : 
                    (N640)? 1'b1 : 
                    (N641)? 1'b1 : 
                    (N642)? 1'b1 : 
                    (N643)? 1'b1 : 
                    (N644)? 1'b1 : 
                    (N645)? 1'b1 : 
                    (N646)? 1'b1 : 
                    (N647)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N649)? 1'b1 : 
                    (N650)? 1'b1 : 
                    (N651)? 1'b1 : 
                    (N652)? 1'b1 : 
                    (N653)? 1'b1 : 
                    (N654)? 1'b1 : 
                    (N655)? 1'b1 : 
                    (N656)? 1'b1 : 
                    (N657)? 1'b1 : 
                    (N658)? 1'b0 : 
                    (N659)? 1'b1 : 
                    (N660)? 1'b0 : 
                    (N661)? 1'b0 : 
                    (N662)? 1'b1 : 
                    (N663)? 1'b1 : 
                    (N664)? 1'b0 : 
                    (N665)? 1'b0 : 
                    (N666)? 1'b1 : 
                    (N667)? 1'b0 : 
                    (N668)? 1'b1 : 
                    (N669)? 1'b1 : 
                    (N670)? 1'b1 : 
                    (N671)? 1'b1 : 
                    (N672)? 1'b1 : 
                    (N673)? 1'b1 : 
                    (N674)? 1'b0 : 
                    (N675)? 1'b1 : 
                    (N676)? 1'b0 : 
                    (N677)? 1'b0 : 
                    (N678)? 1'b1 : 
                    (N679)? 1'b1 : 
                    (N680)? 1'b0 : 
                    (N681)? 1'b0 : 
                    (N682)? 1'b1 : 
                    (N683)? 1'b0 : 
                    (N684)? 1'b1 : 
                    (N685)? 1'b1 : 
                    (N686)? 1'b1 : 
                    (N687)? 1'b1 : 
                    (N688)? 1'b0 : 
                    (N689)? 1'b0 : 
                    (N690)? 1'b0 : 
                    (N691)? 1'b0 : 
                    (N692)? 1'b0 : 
                    (N693)? 1'b0 : 
                    (N694)? 1'b1 : 
                    (N695)? 1'b0 : 
                    (N696)? 1'b0 : 
                    (N697)? 1'b0 : 
                    (N698)? 1'b1 : 
                    (N699)? 1'b0 : 
                    (N700)? 1'b1 : 
                    (N701)? 1'b1 : 
                    (N702)? 1'b1 : 
                    (N703)? 1'b0 : 
                    (N704)? 1'b1 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b1 : 
                    (N707)? 1'b1 : 
                    (N708)? 1'b1 : 
                    (N709)? 1'b1 : 
                    (N710)? 1'b1 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b1 : 
                    (N713)? 1'b1 : 
                    (N714)? 1'b1 : 
                    (N715)? 1'b1 : 
                    (N716)? 1'b1 : 
                    (N717)? 1'b1 : 
                    (N718)? 1'b1 : 
                    (N719)? 1'b1 : 
                    (N720)? 1'b1 : 
                    (N721)? 1'b1 : 
                    (N722)? 1'b0 : 
                    (N723)? 1'b1 : 
                    (N724)? 1'b0 : 
                    (N725)? 1'b0 : 
                    (N726)? 1'b1 : 
                    (N727)? 1'b1 : 
                    (N728)? 1'b0 : 
                    (N729)? 1'b0 : 
                    (N730)? 1'b1 : 
                    (N731)? 1'b0 : 
                    (N732)? 1'b1 : 
                    (N733)? 1'b1 : 
                    (N734)? 1'b1 : 
                    (N735)? 1'b1 : 
                    (N736)? 1'b1 : 
                    (N737)? 1'b1 : 
                    (N738)? 1'b0 : 
                    (N739)? 1'b1 : 
                    (N740)? 1'b0 : 
                    (N741)? 1'b0 : 
                    (N742)? 1'b1 : 
                    (N743)? 1'b1 : 
                    (N744)? 1'b0 : 
                    (N745)? 1'b0 : 
                    (N746)? 1'b1 : 
                    (N747)? 1'b0 : 
                    (N748)? 1'b1 : 
                    (N749)? 1'b1 : 
                    (N750)? 1'b1 : 
                    (N751)? 1'b1 : 
                    (N752)? 1'b0 : 
                    (N753)? 1'b0 : 
                    (N754)? 1'b0 : 
                    (N755)? 1'b0 : 
                    (N756)? 1'b0 : 
                    (N757)? 1'b0 : 
                    (N758)? 1'b1 : 
                    (N759)? 1'b0 : 
                    (N760)? 1'b0 : 
                    (N761)? 1'b0 : 
                    (N762)? 1'b1 : 
                    (N763)? 1'b0 : 
                    (N764)? 1'b1 : 
                    (N765)? 1'b1 : 
                    (N255)? 1'b1 : 1'b0;
  assign fwd_o[6] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b1 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b1 : 
                    (N517)? 1'b1 : 
                    (N518)? 1'b0 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b1 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b1 : 
                    (N523)? 1'b1 : 
                    (N524)? 1'b1 : 
                    (N525)? 1'b1 : 
                    (N526)? 1'b0 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b1 : 
                    (N529)? 1'b1 : 
                    (N530)? 1'b0 : 
                    (N531)? 1'b1 : 
                    (N532)? 1'b0 : 
                    (N533)? 1'b0 : 
                    (N534)? 1'b0 : 
                    (N535)? 1'b1 : 
                    (N536)? 1'b0 : 
                    (N537)? 1'b0 : 
                    (N538)? 1'b1 : 
                    (N539)? 1'b0 : 
                    (N540)? 1'b1 : 
                    (N541)? 1'b1 : 
                    (N542)? 1'b0 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b1 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b1 : 
                    (N547)? 1'b1 : 
                    (N548)? 1'b1 : 
                    (N549)? 1'b1 : 
                    (N550)? 1'b0 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N553)? 1'b1 : 
                    (N554)? 1'b1 : 
                    (N555)? 1'b1 : 
                    (N556)? 1'b1 : 
                    (N557)? 1'b1 : 
                    (N558)? 1'b0 : 
                    (N559)? 1'b1 : 
                    (N560)? 1'b1 : 
                    (N561)? 1'b1 : 
                    (N562)? 1'b0 : 
                    (N563)? 1'b1 : 
                    (N564)? 1'b0 : 
                    (N565)? 1'b0 : 
                    (N566)? 1'b0 : 
                    (N567)? 1'b1 : 
                    (N568)? 1'b0 : 
                    (N569)? 1'b0 : 
                    (N570)? 1'b1 : 
                    (N571)? 1'b0 : 
                    (N572)? 1'b1 : 
                    (N573)? 1'b1 : 
                    (N574)? 1'b0 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b1 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b0 : 
                    (N579)? 1'b1 : 
                    (N580)? 1'b0 : 
                    (N581)? 1'b0 : 
                    (N582)? 1'b0 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b0 : 
                    (N585)? 1'b0 : 
                    (N586)? 1'b1 : 
                    (N587)? 1'b0 : 
                    (N588)? 1'b1 : 
                    (N589)? 1'b1 : 
                    (N590)? 1'b0 : 
                    (N591)? 1'b1 : 
                    (N592)? 1'b0 : 
                    (N593)? 1'b0 : 
                    (N594)? 1'b0 : 
                    (N595)? 1'b0 : 
                    (N596)? 1'b0 : 
                    (N597)? 1'b0 : 
                    (N598)? 1'b0 : 
                    (N599)? 1'b0 : 
                    (N600)? 1'b0 : 
                    (N601)? 1'b0 : 
                    (N602)? 1'b1 : 
                    (N603)? 1'b0 : 
                    (N604)? 1'b1 : 
                    (N605)? 1'b1 : 
                    (N606)? 1'b0 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b0 : 
                    (N609)? 1'b0 : 
                    (N610)? 1'b1 : 
                    (N611)? 1'b0 : 
                    (N612)? 1'b1 : 
                    (N613)? 1'b1 : 
                    (N614)? 1'b0 : 
                    (N615)? 1'b0 : 
                    (N616)? 1'b1 : 
                    (N617)? 1'b1 : 
                    (N618)? 1'b1 : 
                    (N619)? 1'b1 : 
                    (N620)? 1'b1 : 
                    (N621)? 1'b1 : 
                    (N622)? 1'b0 : 
                    (N623)? 1'b0 : 
                    (N624)? 1'b1 : 
                    (N625)? 1'b1 : 
                    (N626)? 1'b0 : 
                    (N627)? 1'b1 : 
                    (N628)? 1'b0 : 
                    (N629)? 1'b0 : 
                    (N630)? 1'b0 : 
                    (N631)? 1'b1 : 
                    (N632)? 1'b0 : 
                    (N633)? 1'b0 : 
                    (N634)? 1'b1 : 
                    (N635)? 1'b0 : 
                    (N636)? 1'b1 : 
                    (N637)? 1'b1 : 
                    (N638)? 1'b0 : 
                    (N639)? 1'b0 : 
                    (N640)? 1'b0 : 
                    (N641)? 1'b0 : 
                    (N642)? 1'b1 : 
                    (N643)? 1'b0 : 
                    (N644)? 1'b1 : 
                    (N645)? 1'b1 : 
                    (N646)? 1'b0 : 
                    (N647)? 1'b0 : 
                    (N648)? 1'b1 : 
                    (N649)? 1'b1 : 
                    (N650)? 1'b1 : 
                    (N651)? 1'b1 : 
                    (N652)? 1'b1 : 
                    (N653)? 1'b1 : 
                    (N654)? 1'b0 : 
                    (N655)? 1'b0 : 
                    (N656)? 1'b1 : 
                    (N657)? 1'b1 : 
                    (N658)? 1'b0 : 
                    (N659)? 1'b1 : 
                    (N660)? 1'b0 : 
                    (N661)? 1'b0 : 
                    (N662)? 1'b0 : 
                    (N663)? 1'b1 : 
                    (N664)? 1'b0 : 
                    (N665)? 1'b0 : 
                    (N666)? 1'b1 : 
                    (N667)? 1'b0 : 
                    (N668)? 1'b1 : 
                    (N669)? 1'b1 : 
                    (N670)? 1'b0 : 
                    (N671)? 1'b0 : 
                    (N672)? 1'b1 : 
                    (N673)? 1'b1 : 
                    (N674)? 1'b1 : 
                    (N675)? 1'b1 : 
                    (N676)? 1'b1 : 
                    (N677)? 1'b1 : 
                    (N678)? 1'b0 : 
                    (N679)? 1'b1 : 
                    (N680)? 1'b1 : 
                    (N681)? 1'b1 : 
                    (N682)? 1'b1 : 
                    (N683)? 1'b1 : 
                    (N684)? 1'b1 : 
                    (N685)? 1'b1 : 
                    (N686)? 1'b0 : 
                    (N687)? 1'b1 : 
                    (N688)? 1'b1 : 
                    (N689)? 1'b1 : 
                    (N690)? 1'b0 : 
                    (N691)? 1'b1 : 
                    (N692)? 1'b0 : 
                    (N693)? 1'b0 : 
                    (N694)? 1'b0 : 
                    (N695)? 1'b1 : 
                    (N696)? 1'b0 : 
                    (N697)? 1'b0 : 
                    (N698)? 1'b1 : 
                    (N699)? 1'b0 : 
                    (N700)? 1'b1 : 
                    (N701)? 1'b1 : 
                    (N702)? 1'b0 : 
                    (N703)? 1'b1 : 
                    (N704)? 1'b1 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b0 : 
                    (N707)? 1'b1 : 
                    (N708)? 1'b0 : 
                    (N709)? 1'b0 : 
                    (N710)? 1'b0 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b0 : 
                    (N713)? 1'b0 : 
                    (N714)? 1'b1 : 
                    (N715)? 1'b0 : 
                    (N716)? 1'b1 : 
                    (N717)? 1'b1 : 
                    (N718)? 1'b0 : 
                    (N719)? 1'b1 : 
                    (N720)? 1'b0 : 
                    (N721)? 1'b0 : 
                    (N722)? 1'b0 : 
                    (N723)? 1'b0 : 
                    (N724)? 1'b0 : 
                    (N725)? 1'b0 : 
                    (N726)? 1'b0 : 
                    (N727)? 1'b0 : 
                    (N728)? 1'b0 : 
                    (N729)? 1'b0 : 
                    (N730)? 1'b1 : 
                    (N731)? 1'b0 : 
                    (N732)? 1'b1 : 
                    (N733)? 1'b1 : 
                    (N734)? 1'b0 : 
                    (N735)? 1'b1 : 
                    (N736)? 1'b0 : 
                    (N737)? 1'b0 : 
                    (N738)? 1'b1 : 
                    (N739)? 1'b0 : 
                    (N740)? 1'b1 : 
                    (N741)? 1'b1 : 
                    (N742)? 1'b0 : 
                    (N743)? 1'b0 : 
                    (N744)? 1'b1 : 
                    (N745)? 1'b1 : 
                    (N746)? 1'b1 : 
                    (N747)? 1'b1 : 
                    (N748)? 1'b1 : 
                    (N749)? 1'b1 : 
                    (N750)? 1'b0 : 
                    (N751)? 1'b0 : 
                    (N752)? 1'b1 : 
                    (N753)? 1'b1 : 
                    (N754)? 1'b0 : 
                    (N755)? 1'b1 : 
                    (N756)? 1'b0 : 
                    (N757)? 1'b0 : 
                    (N758)? 1'b0 : 
                    (N759)? 1'b1 : 
                    (N760)? 1'b0 : 
                    (N761)? 1'b0 : 
                    (N762)? 1'b1 : 
                    (N763)? 1'b0 : 
                    (N764)? 1'b1 : 
                    (N765)? 1'b1 : 
                    (N255)? 1'b0 : 1'b0;
  assign fwd_o[5] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b0 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b0 : 
                    (N517)? 1'b0 : 
                    (N518)? 1'b0 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b0 : 
                    (N521)? 1'b0 : 
                    (N522)? 1'b0 : 
                    (N523)? 1'b0 : 
                    (N524)? 1'b0 : 
                    (N525)? 1'b0 : 
                    (N526)? 1'b0 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b1 : 
                    (N529)? 1'b1 : 
                    (N530)? 1'b0 : 
                    (N531)? 1'b1 : 
                    (N532)? 1'b0 : 
                    (N533)? 1'b0 : 
                    (N534)? 1'b0 : 
                    (N535)? 1'b1 : 
                    (N536)? 1'b0 : 
                    (N537)? 1'b0 : 
                    (N538)? 1'b0 : 
                    (N539)? 1'b0 : 
                    (N540)? 1'b0 : 
                    (N541)? 1'b0 : 
                    (N542)? 1'b0 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b1 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b0 : 
                    (N547)? 1'b1 : 
                    (N548)? 1'b0 : 
                    (N549)? 1'b0 : 
                    (N550)? 1'b0 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b0 : 
                    (N553)? 1'b0 : 
                    (N554)? 1'b0 : 
                    (N555)? 1'b0 : 
                    (N556)? 1'b0 : 
                    (N557)? 1'b0 : 
                    (N558)? 1'b0 : 
                    (N559)? 1'b1 : 
                    (N560)? 1'b1 : 
                    (N561)? 1'b1 : 
                    (N562)? 1'b0 : 
                    (N563)? 1'b1 : 
                    (N564)? 1'b0 : 
                    (N565)? 1'b0 : 
                    (N566)? 1'b0 : 
                    (N567)? 1'b1 : 
                    (N568)? 1'b0 : 
                    (N569)? 1'b0 : 
                    (N570)? 1'b0 : 
                    (N571)? 1'b0 : 
                    (N572)? 1'b0 : 
                    (N573)? 1'b0 : 
                    (N574)? 1'b0 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b1 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b0 : 
                    (N579)? 1'b1 : 
                    (N580)? 1'b0 : 
                    (N581)? 1'b0 : 
                    (N582)? 1'b0 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b0 : 
                    (N585)? 1'b0 : 
                    (N586)? 1'b0 : 
                    (N587)? 1'b0 : 
                    (N588)? 1'b0 : 
                    (N589)? 1'b0 : 
                    (N590)? 1'b0 : 
                    (N591)? 1'b1 : 
                    (N592)? 1'b1 : 
                    (N593)? 1'b1 : 
                    (N594)? 1'b0 : 
                    (N595)? 1'b1 : 
                    (N596)? 1'b0 : 
                    (N597)? 1'b0 : 
                    (N598)? 1'b0 : 
                    (N599)? 1'b1 : 
                    (N600)? 1'b0 : 
                    (N601)? 1'b0 : 
                    (N602)? 1'b0 : 
                    (N603)? 1'b0 : 
                    (N604)? 1'b0 : 
                    (N605)? 1'b0 : 
                    (N606)? 1'b0 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b1 : 
                    (N609)? 1'b1 : 
                    (N610)? 1'b0 : 
                    (N611)? 1'b1 : 
                    (N612)? 1'b0 : 
                    (N613)? 1'b0 : 
                    (N614)? 1'b0 : 
                    (N615)? 1'b1 : 
                    (N616)? 1'b0 : 
                    (N617)? 1'b0 : 
                    (N618)? 1'b0 : 
                    (N619)? 1'b0 : 
                    (N620)? 1'b0 : 
                    (N621)? 1'b0 : 
                    (N622)? 1'b0 : 
                    (N623)? 1'b1 : 
                    (N624)? 1'b1 : 
                    (N625)? 1'b1 : 
                    (N626)? 1'b0 : 
                    (N627)? 1'b1 : 
                    (N628)? 1'b0 : 
                    (N629)? 1'b0 : 
                    (N630)? 1'b0 : 
                    (N631)? 1'b1 : 
                    (N632)? 1'b0 : 
                    (N633)? 1'b0 : 
                    (N634)? 1'b0 : 
                    (N635)? 1'b0 : 
                    (N636)? 1'b0 : 
                    (N637)? 1'b0 : 
                    (N638)? 1'b0 : 
                    (N639)? 1'b1 : 
                    (N640)? 1'b1 : 
                    (N641)? 1'b1 : 
                    (N642)? 1'b0 : 
                    (N643)? 1'b1 : 
                    (N644)? 1'b0 : 
                    (N645)? 1'b0 : 
                    (N646)? 1'b0 : 
                    (N647)? 1'b1 : 
                    (N648)? 1'b0 : 
                    (N649)? 1'b0 : 
                    (N650)? 1'b0 : 
                    (N651)? 1'b0 : 
                    (N652)? 1'b0 : 
                    (N653)? 1'b0 : 
                    (N654)? 1'b0 : 
                    (N655)? 1'b1 : 
                    (N656)? 1'b1 : 
                    (N657)? 1'b1 : 
                    (N658)? 1'b0 : 
                    (N659)? 1'b1 : 
                    (N660)? 1'b0 : 
                    (N661)? 1'b0 : 
                    (N662)? 1'b0 : 
                    (N663)? 1'b1 : 
                    (N664)? 1'b0 : 
                    (N665)? 1'b0 : 
                    (N666)? 1'b0 : 
                    (N667)? 1'b0 : 
                    (N668)? 1'b0 : 
                    (N669)? 1'b0 : 
                    (N670)? 1'b0 : 
                    (N671)? 1'b1 : 
                    (N672)? 1'b1 : 
                    (N673)? 1'b1 : 
                    (N674)? 1'b0 : 
                    (N675)? 1'b1 : 
                    (N676)? 1'b0 : 
                    (N677)? 1'b0 : 
                    (N678)? 1'b0 : 
                    (N679)? 1'b1 : 
                    (N680)? 1'b0 : 
                    (N681)? 1'b0 : 
                    (N682)? 1'b0 : 
                    (N683)? 1'b0 : 
                    (N684)? 1'b0 : 
                    (N685)? 1'b0 : 
                    (N686)? 1'b0 : 
                    (N687)? 1'b1 : 
                    (N688)? 1'b1 : 
                    (N689)? 1'b1 : 
                    (N690)? 1'b0 : 
                    (N691)? 1'b1 : 
                    (N692)? 1'b0 : 
                    (N693)? 1'b0 : 
                    (N694)? 1'b0 : 
                    (N695)? 1'b1 : 
                    (N696)? 1'b0 : 
                    (N697)? 1'b0 : 
                    (N698)? 1'b0 : 
                    (N699)? 1'b0 : 
                    (N700)? 1'b0 : 
                    (N701)? 1'b0 : 
                    (N702)? 1'b0 : 
                    (N703)? 1'b1 : 
                    (N704)? 1'b1 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b0 : 
                    (N707)? 1'b1 : 
                    (N708)? 1'b0 : 
                    (N709)? 1'b0 : 
                    (N710)? 1'b0 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b0 : 
                    (N713)? 1'b0 : 
                    (N714)? 1'b0 : 
                    (N715)? 1'b0 : 
                    (N716)? 1'b0 : 
                    (N717)? 1'b0 : 
                    (N718)? 1'b0 : 
                    (N719)? 1'b1 : 
                    (N720)? 1'b1 : 
                    (N721)? 1'b1 : 
                    (N722)? 1'b0 : 
                    (N723)? 1'b1 : 
                    (N724)? 1'b0 : 
                    (N725)? 1'b0 : 
                    (N726)? 1'b0 : 
                    (N727)? 1'b1 : 
                    (N728)? 1'b0 : 
                    (N729)? 1'b0 : 
                    (N730)? 1'b0 : 
                    (N731)? 1'b0 : 
                    (N732)? 1'b0 : 
                    (N733)? 1'b0 : 
                    (N734)? 1'b0 : 
                    (N735)? 1'b1 : 
                    (N736)? 1'b1 : 
                    (N737)? 1'b1 : 
                    (N738)? 1'b0 : 
                    (N739)? 1'b1 : 
                    (N740)? 1'b0 : 
                    (N741)? 1'b0 : 
                    (N742)? 1'b0 : 
                    (N743)? 1'b1 : 
                    (N744)? 1'b0 : 
                    (N745)? 1'b0 : 
                    (N746)? 1'b0 : 
                    (N747)? 1'b0 : 
                    (N748)? 1'b0 : 
                    (N749)? 1'b0 : 
                    (N750)? 1'b0 : 
                    (N751)? 1'b1 : 
                    (N752)? 1'b1 : 
                    (N753)? 1'b1 : 
                    (N754)? 1'b0 : 
                    (N755)? 1'b1 : 
                    (N756)? 1'b0 : 
                    (N757)? 1'b0 : 
                    (N758)? 1'b0 : 
                    (N759)? 1'b1 : 
                    (N760)? 1'b0 : 
                    (N761)? 1'b0 : 
                    (N762)? 1'b0 : 
                    (N763)? 1'b0 : 
                    (N764)? 1'b0 : 
                    (N765)? 1'b0 : 
                    (N255)? 1'b0 : 1'b0;
  assign fwd_o[4] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b0 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b1 : 
                    (N517)? 1'b1 : 
                    (N518)? 1'b0 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b1 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b0 : 
                    (N523)? 1'b1 : 
                    (N524)? 1'b1 : 
                    (N525)? 1'b1 : 
                    (N526)? 1'b0 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b0 : 
                    (N529)? 1'b0 : 
                    (N530)? 1'b0 : 
                    (N531)? 1'b0 : 
                    (N532)? 1'b1 : 
                    (N533)? 1'b1 : 
                    (N534)? 1'b0 : 
                    (N535)? 1'b0 : 
                    (N536)? 1'b1 : 
                    (N537)? 1'b1 : 
                    (N538)? 1'b0 : 
                    (N539)? 1'b1 : 
                    (N540)? 1'b1 : 
                    (N541)? 1'b1 : 
                    (N542)? 1'b0 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b0 : 
                    (N545)? 1'b0 : 
                    (N546)? 1'b0 : 
                    (N547)? 1'b0 : 
                    (N548)? 1'b1 : 
                    (N549)? 1'b1 : 
                    (N550)? 1'b0 : 
                    (N551)? 1'b0 : 
                    (N552)? 1'b1 : 
                    (N553)? 1'b1 : 
                    (N554)? 1'b0 : 
                    (N555)? 1'b1 : 
                    (N556)? 1'b1 : 
                    (N557)? 1'b1 : 
                    (N558)? 1'b0 : 
                    (N559)? 1'b0 : 
                    (N560)? 1'b0 : 
                    (N561)? 1'b0 : 
                    (N562)? 1'b0 : 
                    (N563)? 1'b0 : 
                    (N564)? 1'b1 : 
                    (N565)? 1'b1 : 
                    (N566)? 1'b0 : 
                    (N567)? 1'b0 : 
                    (N568)? 1'b1 : 
                    (N569)? 1'b1 : 
                    (N570)? 1'b0 : 
                    (N571)? 1'b1 : 
                    (N572)? 1'b1 : 
                    (N573)? 1'b1 : 
                    (N574)? 1'b0 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b1 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b0 : 
                    (N579)? 1'b1 : 
                    (N580)? 1'b1 : 
                    (N581)? 1'b1 : 
                    (N582)? 1'b0 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b1 : 
                    (N585)? 1'b1 : 
                    (N586)? 1'b0 : 
                    (N587)? 1'b1 : 
                    (N588)? 1'b1 : 
                    (N589)? 1'b1 : 
                    (N590)? 1'b0 : 
                    (N591)? 1'b1 : 
                    (N592)? 1'b0 : 
                    (N593)? 1'b0 : 
                    (N594)? 1'b0 : 
                    (N595)? 1'b0 : 
                    (N596)? 1'b1 : 
                    (N597)? 1'b1 : 
                    (N598)? 1'b0 : 
                    (N599)? 1'b0 : 
                    (N600)? 1'b1 : 
                    (N601)? 1'b1 : 
                    (N602)? 1'b0 : 
                    (N603)? 1'b1 : 
                    (N604)? 1'b1 : 
                    (N605)? 1'b1 : 
                    (N606)? 1'b0 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b0 : 
                    (N609)? 1'b0 : 
                    (N610)? 1'b0 : 
                    (N611)? 1'b0 : 
                    (N612)? 1'b1 : 
                    (N613)? 1'b1 : 
                    (N614)? 1'b0 : 
                    (N615)? 1'b0 : 
                    (N616)? 1'b1 : 
                    (N617)? 1'b1 : 
                    (N618)? 1'b0 : 
                    (N619)? 1'b1 : 
                    (N620)? 1'b1 : 
                    (N621)? 1'b1 : 
                    (N622)? 1'b0 : 
                    (N623)? 1'b0 : 
                    (N624)? 1'b0 : 
                    (N625)? 1'b0 : 
                    (N626)? 1'b0 : 
                    (N627)? 1'b0 : 
                    (N628)? 1'b1 : 
                    (N629)? 1'b1 : 
                    (N630)? 1'b0 : 
                    (N631)? 1'b0 : 
                    (N632)? 1'b1 : 
                    (N633)? 1'b1 : 
                    (N634)? 1'b0 : 
                    (N635)? 1'b1 : 
                    (N636)? 1'b1 : 
                    (N637)? 1'b1 : 
                    (N638)? 1'b0 : 
                    (N639)? 1'b1 : 
                    (N640)? 1'b1 : 
                    (N641)? 1'b1 : 
                    (N642)? 1'b0 : 
                    (N643)? 1'b1 : 
                    (N644)? 1'b1 : 
                    (N645)? 1'b1 : 
                    (N646)? 1'b0 : 
                    (N647)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N649)? 1'b1 : 
                    (N650)? 1'b0 : 
                    (N651)? 1'b1 : 
                    (N652)? 1'b1 : 
                    (N653)? 1'b1 : 
                    (N654)? 1'b0 : 
                    (N655)? 1'b1 : 
                    (N656)? 1'b0 : 
                    (N657)? 1'b0 : 
                    (N658)? 1'b0 : 
                    (N659)? 1'b0 : 
                    (N660)? 1'b1 : 
                    (N661)? 1'b1 : 
                    (N662)? 1'b0 : 
                    (N663)? 1'b0 : 
                    (N664)? 1'b1 : 
                    (N665)? 1'b1 : 
                    (N666)? 1'b0 : 
                    (N667)? 1'b1 : 
                    (N668)? 1'b1 : 
                    (N669)? 1'b1 : 
                    (N670)? 1'b0 : 
                    (N671)? 1'b1 : 
                    (N672)? 1'b0 : 
                    (N673)? 1'b0 : 
                    (N674)? 1'b0 : 
                    (N675)? 1'b0 : 
                    (N676)? 1'b1 : 
                    (N677)? 1'b1 : 
                    (N678)? 1'b0 : 
                    (N679)? 1'b0 : 
                    (N680)? 1'b1 : 
                    (N681)? 1'b1 : 
                    (N682)? 1'b0 : 
                    (N683)? 1'b1 : 
                    (N684)? 1'b1 : 
                    (N685)? 1'b1 : 
                    (N686)? 1'b0 : 
                    (N687)? 1'b0 : 
                    (N688)? 1'b0 : 
                    (N689)? 1'b0 : 
                    (N690)? 1'b0 : 
                    (N691)? 1'b0 : 
                    (N692)? 1'b1 : 
                    (N693)? 1'b1 : 
                    (N694)? 1'b0 : 
                    (N695)? 1'b0 : 
                    (N696)? 1'b1 : 
                    (N697)? 1'b1 : 
                    (N698)? 1'b0 : 
                    (N699)? 1'b1 : 
                    (N700)? 1'b1 : 
                    (N701)? 1'b1 : 
                    (N702)? 1'b0 : 
                    (N703)? 1'b1 : 
                    (N704)? 1'b1 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b0 : 
                    (N707)? 1'b1 : 
                    (N708)? 1'b1 : 
                    (N709)? 1'b1 : 
                    (N710)? 1'b0 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b1 : 
                    (N713)? 1'b1 : 
                    (N714)? 1'b0 : 
                    (N715)? 1'b1 : 
                    (N716)? 1'b1 : 
                    (N717)? 1'b1 : 
                    (N718)? 1'b0 : 
                    (N719)? 1'b1 : 
                    (N720)? 1'b0 : 
                    (N721)? 1'b0 : 
                    (N722)? 1'b0 : 
                    (N723)? 1'b0 : 
                    (N724)? 1'b1 : 
                    (N725)? 1'b1 : 
                    (N726)? 1'b0 : 
                    (N727)? 1'b0 : 
                    (N728)? 1'b1 : 
                    (N729)? 1'b1 : 
                    (N730)? 1'b0 : 
                    (N731)? 1'b1 : 
                    (N732)? 1'b1 : 
                    (N733)? 1'b1 : 
                    (N734)? 1'b0 : 
                    (N735)? 1'b1 : 
                    (N736)? 1'b0 : 
                    (N737)? 1'b0 : 
                    (N738)? 1'b0 : 
                    (N739)? 1'b0 : 
                    (N740)? 1'b1 : 
                    (N741)? 1'b1 : 
                    (N742)? 1'b0 : 
                    (N743)? 1'b0 : 
                    (N744)? 1'b1 : 
                    (N745)? 1'b1 : 
                    (N746)? 1'b0 : 
                    (N747)? 1'b1 : 
                    (N748)? 1'b1 : 
                    (N749)? 1'b1 : 
                    (N750)? 1'b0 : 
                    (N751)? 1'b0 : 
                    (N752)? 1'b0 : 
                    (N753)? 1'b0 : 
                    (N754)? 1'b0 : 
                    (N755)? 1'b0 : 
                    (N756)? 1'b1 : 
                    (N757)? 1'b1 : 
                    (N758)? 1'b0 : 
                    (N759)? 1'b0 : 
                    (N760)? 1'b1 : 
                    (N761)? 1'b1 : 
                    (N762)? 1'b0 : 
                    (N763)? 1'b1 : 
                    (N764)? 1'b1 : 
                    (N765)? 1'b1 : 
                    (N255)? 1'b0 : 1'b0;
  assign fwd_o[3] = (N511)? 1'b1 : 
                    (N512)? 1'b1 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b1 : 
                    (N515)? 1'b1 : 
                    (N516)? 1'b0 : 
                    (N517)? 1'b0 : 
                    (N518)? 1'b1 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b1 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b1 : 
                    (N523)? 1'b1 : 
                    (N524)? 1'b0 : 
                    (N525)? 1'b0 : 
                    (N526)? 1'b1 : 
                    (N527)? 1'b1 : 
                    (N528)? 1'b0 : 
                    (N529)? 1'b0 : 
                    (N530)? 1'b1 : 
                    (N531)? 1'b0 : 
                    (N532)? 1'b0 : 
                    (N533)? 1'b0 : 
                    (N534)? 1'b1 : 
                    (N535)? 1'b0 : 
                    (N536)? 1'b1 : 
                    (N537)? 1'b1 : 
                    (N538)? 1'b1 : 
                    (N539)? 1'b1 : 
                    (N540)? 1'b0 : 
                    (N541)? 1'b0 : 
                    (N542)? 1'b1 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b1 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b1 : 
                    (N547)? 1'b1 : 
                    (N548)? 1'b0 : 
                    (N549)? 1'b0 : 
                    (N550)? 1'b1 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b1 : 
                    (N553)? 1'b1 : 
                    (N554)? 1'b1 : 
                    (N555)? 1'b1 : 
                    (N556)? 1'b0 : 
                    (N557)? 1'b0 : 
                    (N558)? 1'b1 : 
                    (N559)? 1'b1 : 
                    (N560)? 1'b0 : 
                    (N561)? 1'b0 : 
                    (N562)? 1'b1 : 
                    (N563)? 1'b0 : 
                    (N564)? 1'b0 : 
                    (N565)? 1'b0 : 
                    (N566)? 1'b1 : 
                    (N567)? 1'b0 : 
                    (N568)? 1'b1 : 
                    (N569)? 1'b1 : 
                    (N570)? 1'b1 : 
                    (N571)? 1'b1 : 
                    (N572)? 1'b0 : 
                    (N573)? 1'b0 : 
                    (N574)? 1'b1 : 
                    (N575)? 1'b1 : 
                    (N576)? 1'b0 : 
                    (N577)? 1'b0 : 
                    (N578)? 1'b1 : 
                    (N579)? 1'b0 : 
                    (N580)? 1'b0 : 
                    (N581)? 1'b0 : 
                    (N582)? 1'b1 : 
                    (N583)? 1'b0 : 
                    (N584)? 1'b1 : 
                    (N585)? 1'b1 : 
                    (N586)? 1'b1 : 
                    (N587)? 1'b1 : 
                    (N588)? 1'b0 : 
                    (N589)? 1'b0 : 
                    (N590)? 1'b1 : 
                    (N591)? 1'b0 : 
                    (N592)? 1'b0 : 
                    (N593)? 1'b0 : 
                    (N594)? 1'b1 : 
                    (N595)? 1'b0 : 
                    (N596)? 1'b0 : 
                    (N597)? 1'b0 : 
                    (N598)? 1'b1 : 
                    (N599)? 1'b0 : 
                    (N600)? 1'b1 : 
                    (N601)? 1'b1 : 
                    (N602)? 1'b1 : 
                    (N603)? 1'b1 : 
                    (N604)? 1'b0 : 
                    (N605)? 1'b0 : 
                    (N606)? 1'b1 : 
                    (N607)? 1'b0 : 
                    (N608)? 1'b1 : 
                    (N609)? 1'b1 : 
                    (N610)? 1'b1 : 
                    (N611)? 1'b1 : 
                    (N612)? 1'b0 : 
                    (N613)? 1'b0 : 
                    (N614)? 1'b1 : 
                    (N615)? 1'b1 : 
                    (N616)? 1'b1 : 
                    (N617)? 1'b1 : 
                    (N618)? 1'b1 : 
                    (N619)? 1'b1 : 
                    (N620)? 1'b0 : 
                    (N621)? 1'b0 : 
                    (N622)? 1'b1 : 
                    (N623)? 1'b1 : 
                    (N624)? 1'b0 : 
                    (N625)? 1'b0 : 
                    (N626)? 1'b1 : 
                    (N627)? 1'b0 : 
                    (N628)? 1'b0 : 
                    (N629)? 1'b0 : 
                    (N630)? 1'b1 : 
                    (N631)? 1'b0 : 
                    (N632)? 1'b1 : 
                    (N633)? 1'b1 : 
                    (N634)? 1'b1 : 
                    (N635)? 1'b1 : 
                    (N636)? 1'b0 : 
                    (N637)? 1'b0 : 
                    (N638)? 1'b1 : 
                    (N639)? 1'b0 : 
                    (N640)? 1'b1 : 
                    (N641)? 1'b1 : 
                    (N642)? 1'b1 : 
                    (N643)? 1'b1 : 
                    (N644)? 1'b0 : 
                    (N645)? 1'b0 : 
                    (N646)? 1'b1 : 
                    (N647)? 1'b1 : 
                    (N648)? 1'b1 : 
                    (N649)? 1'b1 : 
                    (N650)? 1'b1 : 
                    (N651)? 1'b1 : 
                    (N652)? 1'b0 : 
                    (N653)? 1'b0 : 
                    (N654)? 1'b1 : 
                    (N655)? 1'b1 : 
                    (N656)? 1'b0 : 
                    (N657)? 1'b0 : 
                    (N658)? 1'b1 : 
                    (N659)? 1'b0 : 
                    (N660)? 1'b0 : 
                    (N661)? 1'b0 : 
                    (N662)? 1'b1 : 
                    (N663)? 1'b0 : 
                    (N664)? 1'b1 : 
                    (N665)? 1'b1 : 
                    (N666)? 1'b1 : 
                    (N667)? 1'b1 : 
                    (N668)? 1'b0 : 
                    (N669)? 1'b0 : 
                    (N670)? 1'b1 : 
                    (N671)? 1'b1 : 
                    (N672)? 1'b1 : 
                    (N673)? 1'b1 : 
                    (N674)? 1'b1 : 
                    (N675)? 1'b1 : 
                    (N676)? 1'b0 : 
                    (N677)? 1'b0 : 
                    (N678)? 1'b1 : 
                    (N679)? 1'b1 : 
                    (N680)? 1'b1 : 
                    (N681)? 1'b1 : 
                    (N682)? 1'b1 : 
                    (N683)? 1'b1 : 
                    (N684)? 1'b0 : 
                    (N685)? 1'b0 : 
                    (N686)? 1'b1 : 
                    (N687)? 1'b1 : 
                    (N688)? 1'b0 : 
                    (N689)? 1'b0 : 
                    (N690)? 1'b1 : 
                    (N691)? 1'b0 : 
                    (N692)? 1'b0 : 
                    (N693)? 1'b0 : 
                    (N694)? 1'b1 : 
                    (N695)? 1'b0 : 
                    (N696)? 1'b1 : 
                    (N697)? 1'b1 : 
                    (N698)? 1'b1 : 
                    (N699)? 1'b1 : 
                    (N700)? 1'b0 : 
                    (N701)? 1'b0 : 
                    (N702)? 1'b1 : 
                    (N703)? 1'b1 : 
                    (N704)? 1'b0 : 
                    (N705)? 1'b0 : 
                    (N706)? 1'b1 : 
                    (N707)? 1'b0 : 
                    (N708)? 1'b0 : 
                    (N709)? 1'b0 : 
                    (N710)? 1'b1 : 
                    (N711)? 1'b0 : 
                    (N712)? 1'b1 : 
                    (N713)? 1'b1 : 
                    (N714)? 1'b1 : 
                    (N715)? 1'b1 : 
                    (N716)? 1'b0 : 
                    (N717)? 1'b0 : 
                    (N718)? 1'b1 : 
                    (N719)? 1'b0 : 
                    (N720)? 1'b0 : 
                    (N721)? 1'b0 : 
                    (N722)? 1'b1 : 
                    (N723)? 1'b0 : 
                    (N724)? 1'b0 : 
                    (N725)? 1'b0 : 
                    (N726)? 1'b1 : 
                    (N727)? 1'b0 : 
                    (N728)? 1'b1 : 
                    (N729)? 1'b1 : 
                    (N730)? 1'b1 : 
                    (N731)? 1'b1 : 
                    (N732)? 1'b0 : 
                    (N733)? 1'b0 : 
                    (N734)? 1'b1 : 
                    (N735)? 1'b0 : 
                    (N736)? 1'b1 : 
                    (N737)? 1'b1 : 
                    (N738)? 1'b1 : 
                    (N739)? 1'b1 : 
                    (N740)? 1'b0 : 
                    (N741)? 1'b0 : 
                    (N742)? 1'b1 : 
                    (N743)? 1'b1 : 
                    (N744)? 1'b1 : 
                    (N745)? 1'b1 : 
                    (N746)? 1'b1 : 
                    (N747)? 1'b1 : 
                    (N748)? 1'b0 : 
                    (N749)? 1'b0 : 
                    (N750)? 1'b1 : 
                    (N751)? 1'b1 : 
                    (N752)? 1'b0 : 
                    (N753)? 1'b0 : 
                    (N754)? 1'b1 : 
                    (N755)? 1'b0 : 
                    (N756)? 1'b0 : 
                    (N757)? 1'b0 : 
                    (N758)? 1'b1 : 
                    (N759)? 1'b0 : 
                    (N760)? 1'b1 : 
                    (N761)? 1'b1 : 
                    (N762)? 1'b1 : 
                    (N763)? 1'b1 : 
                    (N764)? 1'b0 : 
                    (N765)? 1'b0 : 
                    (N255)? 1'b1 : 1'b0;
  assign fwd_o[0] = (N511)? 1'b1 : 
                    (N512)? 1'b0 : 
                    (N513)? 1'b1 : 
                    (N514)? 1'b0 : 
                    (N515)? 1'b0 : 
                    (N516)? 1'b0 : 
                    (N517)? 1'b1 : 
                    (N518)? 1'b0 : 
                    (N519)? 1'b1 : 
                    (N520)? 1'b0 : 
                    (N521)? 1'b1 : 
                    (N522)? 1'b0 : 
                    (N523)? 1'b0 : 
                    (N524)? 1'b0 : 
                    (N525)? 1'b1 : 
                    (N526)? 1'b0 : 
                    (N527)? 1'b0 : 
                    (N528)? 1'b0 : 
                    (N529)? 1'b1 : 
                    (N530)? 1'b0 : 
                    (N531)? 1'b0 : 
                    (N532)? 1'b0 : 
                    (N533)? 1'b1 : 
                    (N534)? 1'b0 : 
                    (N535)? 1'b1 : 
                    (N536)? 1'b0 : 
                    (N537)? 1'b1 : 
                    (N538)? 1'b0 : 
                    (N539)? 1'b0 : 
                    (N540)? 1'b0 : 
                    (N541)? 1'b1 : 
                    (N542)? 1'b0 : 
                    (N543)? 1'b1 : 
                    (N544)? 1'b0 : 
                    (N545)? 1'b1 : 
                    (N546)? 1'b0 : 
                    (N547)? 1'b0 : 
                    (N548)? 1'b0 : 
                    (N549)? 1'b1 : 
                    (N550)? 1'b0 : 
                    (N551)? 1'b1 : 
                    (N552)? 1'b0 : 
                    (N553)? 1'b1 : 
                    (N554)? 1'b0 : 
                    (N555)? 1'b0 : 
                    (N556)? 1'b0 : 
                    (N557)? 1'b1 : 
                    (N558)? 1'b0 : 
                    (N559)? 1'b0 : 
                    (N560)? 1'b0 : 
                    (N561)? 1'b1 : 
                    (N562)? 1'b0 : 
                    (N563)? 1'b0 : 
                    (N564)? 1'b0 : 
                    (N565)? 1'b1 : 
                    (N566)? 1'b0 : 
                    (N567)? 1'b1 : 
                    (N568)? 1'b0 : 
                    (N569)? 1'b1 : 
                    (N570)? 1'b0 : 
                    (N571)? 1'b0 : 
                    (N572)? 1'b0 : 
                    (N573)? 1'b1 : 
                    (N574)? 1'b0 : 
                    (N575)? 1'b0 : 
                    (N576)? 1'b0 : 
                    (N577)? 1'b1 : 
                    (N578)? 1'b0 : 
                    (N579)? 1'b0 : 
                    (N580)? 1'b0 : 
                    (N581)? 1'b1 : 
                    (N582)? 1'b0 : 
                    (N583)? 1'b1 : 
                    (N584)? 1'b0 : 
                    (N585)? 1'b1 : 
                    (N586)? 1'b0 : 
                    (N587)? 1'b0 : 
                    (N588)? 1'b0 : 
                    (N589)? 1'b1 : 
                    (N590)? 1'b0 : 
                    (N591)? 1'b0 : 
                    (N592)? 1'b0 : 
                    (N593)? 1'b1 : 
                    (N594)? 1'b0 : 
                    (N595)? 1'b0 : 
                    (N596)? 1'b0 : 
                    (N597)? 1'b1 : 
                    (N598)? 1'b0 : 
                    (N599)? 1'b1 : 
                    (N600)? 1'b0 : 
                    (N601)? 1'b1 : 
                    (N602)? 1'b0 : 
                    (N603)? 1'b0 : 
                    (N604)? 1'b0 : 
                    (N605)? 1'b1 : 
                    (N606)? 1'b0 : 
                    (N607)? 1'b1 : 
                    (N608)? 1'b0 : 
                    (N609)? 1'b1 : 
                    (N610)? 1'b0 : 
                    (N611)? 1'b0 : 
                    (N612)? 1'b0 : 
                    (N613)? 1'b1 : 
                    (N614)? 1'b0 : 
                    (N615)? 1'b1 : 
                    (N616)? 1'b0 : 
                    (N617)? 1'b1 : 
                    (N618)? 1'b0 : 
                    (N619)? 1'b0 : 
                    (N620)? 1'b0 : 
                    (N621)? 1'b1 : 
                    (N622)? 1'b0 : 
                    (N623)? 1'b0 : 
                    (N624)? 1'b0 : 
                    (N625)? 1'b1 : 
                    (N626)? 1'b0 : 
                    (N627)? 1'b0 : 
                    (N628)? 1'b0 : 
                    (N629)? 1'b1 : 
                    (N630)? 1'b0 : 
                    (N631)? 1'b1 : 
                    (N632)? 1'b0 : 
                    (N633)? 1'b1 : 
                    (N634)? 1'b0 : 
                    (N635)? 1'b0 : 
                    (N636)? 1'b0 : 
                    (N637)? 1'b1 : 
                    (N638)? 1'b0 : 
                    (N639)? 1'b1 : 
                    (N640)? 1'b0 : 
                    (N641)? 1'b1 : 
                    (N642)? 1'b0 : 
                    (N643)? 1'b0 : 
                    (N644)? 1'b0 : 
                    (N645)? 1'b1 : 
                    (N646)? 1'b0 : 
                    (N647)? 1'b1 : 
                    (N648)? 1'b0 : 
                    (N649)? 1'b1 : 
                    (N650)? 1'b0 : 
                    (N651)? 1'b0 : 
                    (N652)? 1'b0 : 
                    (N653)? 1'b1 : 
                    (N654)? 1'b0 : 
                    (N655)? 1'b0 : 
                    (N656)? 1'b0 : 
                    (N657)? 1'b1 : 
                    (N658)? 1'b0 : 
                    (N659)? 1'b0 : 
                    (N660)? 1'b0 : 
                    (N661)? 1'b1 : 
                    (N662)? 1'b0 : 
                    (N663)? 1'b1 : 
                    (N664)? 1'b0 : 
                    (N665)? 1'b1 : 
                    (N666)? 1'b0 : 
                    (N667)? 1'b0 : 
                    (N668)? 1'b0 : 
                    (N669)? 1'b1 : 
                    (N670)? 1'b0 : 
                    (N671)? 1'b1 : 
                    (N672)? 1'b0 : 
                    (N673)? 1'b1 : 
                    (N674)? 1'b0 : 
                    (N675)? 1'b0 : 
                    (N676)? 1'b0 : 
                    (N677)? 1'b1 : 
                    (N678)? 1'b0 : 
                    (N679)? 1'b1 : 
                    (N680)? 1'b0 : 
                    (N681)? 1'b1 : 
                    (N682)? 1'b0 : 
                    (N683)? 1'b0 : 
                    (N684)? 1'b0 : 
                    (N685)? 1'b1 : 
                    (N686)? 1'b0 : 
                    (N687)? 1'b0 : 
                    (N688)? 1'b0 : 
                    (N689)? 1'b1 : 
                    (N690)? 1'b0 : 
                    (N691)? 1'b0 : 
                    (N692)? 1'b0 : 
                    (N693)? 1'b1 : 
                    (N694)? 1'b0 : 
                    (N695)? 1'b1 : 
                    (N696)? 1'b0 : 
                    (N697)? 1'b1 : 
                    (N698)? 1'b0 : 
                    (N699)? 1'b0 : 
                    (N700)? 1'b0 : 
                    (N701)? 1'b1 : 
                    (N702)? 1'b0 : 
                    (N703)? 1'b0 : 
                    (N704)? 1'b0 : 
                    (N705)? 1'b1 : 
                    (N706)? 1'b0 : 
                    (N707)? 1'b0 : 
                    (N708)? 1'b0 : 
                    (N709)? 1'b1 : 
                    (N710)? 1'b0 : 
                    (N711)? 1'b1 : 
                    (N712)? 1'b0 : 
                    (N713)? 1'b1 : 
                    (N714)? 1'b0 : 
                    (N715)? 1'b0 : 
                    (N716)? 1'b0 : 
                    (N717)? 1'b1 : 
                    (N718)? 1'b0 : 
                    (N719)? 1'b0 : 
                    (N720)? 1'b0 : 
                    (N721)? 1'b1 : 
                    (N722)? 1'b0 : 
                    (N723)? 1'b0 : 
                    (N724)? 1'b0 : 
                    (N725)? 1'b1 : 
                    (N726)? 1'b0 : 
                    (N727)? 1'b1 : 
                    (N728)? 1'b0 : 
                    (N729)? 1'b1 : 
                    (N730)? 1'b0 : 
                    (N731)? 1'b0 : 
                    (N732)? 1'b0 : 
                    (N733)? 1'b1 : 
                    (N734)? 1'b0 : 
                    (N735)? 1'b1 : 
                    (N736)? 1'b0 : 
                    (N737)? 1'b1 : 
                    (N738)? 1'b0 : 
                    (N739)? 1'b0 : 
                    (N740)? 1'b0 : 
                    (N741)? 1'b1 : 
                    (N742)? 1'b0 : 
                    (N743)? 1'b1 : 
                    (N744)? 1'b0 : 
                    (N745)? 1'b1 : 
                    (N746)? 1'b0 : 
                    (N747)? 1'b0 : 
                    (N748)? 1'b0 : 
                    (N749)? 1'b1 : 
                    (N750)? 1'b0 : 
                    (N751)? 1'b0 : 
                    (N752)? 1'b0 : 
                    (N753)? 1'b1 : 
                    (N754)? 1'b0 : 
                    (N755)? 1'b0 : 
                    (N756)? 1'b0 : 
                    (N757)? 1'b1 : 
                    (N758)? 1'b0 : 
                    (N759)? 1'b1 : 
                    (N760)? 1'b0 : 
                    (N761)? 1'b1 : 
                    (N762)? 1'b0 : 
                    (N763)? 1'b0 : 
                    (N764)? 1'b0 : 
                    (N765)? 1'b1 : 
                    (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[13] = (N766)? 1'b0 : 
                              (N1)? 1'b0 : 
                              (N767)? 1'b0 : 
                              (N768)? 1'b0 : 
                              (N769)? 1'b0 : 
                              (N770)? 1'b0 : 
                              (N771)? 1'b0 : 
                              (N772)? 1'b0 : 
                              (N773)? 1'b0 : 
                              (N774)? 1'b0 : 
                              (N775)? 1'b0 : 
                              (N776)? 1'b0 : 
                              (N777)? 1'b0 : 
                              (N778)? 1'b0 : 
                              (N779)? 1'b0 : 
                              (N780)? 1'b0 : 
                              (N781)? 1'b0 : 
                              (N782)? 1'b0 : 
                              (N783)? 1'b0 : 
                              (N784)? 1'b0 : 
                              (N785)? 1'b0 : 
                              (N786)? 1'b0 : 
                              (N787)? 1'b0 : 
                              (N788)? 1'b0 : 
                              (N789)? 1'b0 : 
                              (N790)? 1'b0 : 
                              (N791)? 1'b0 : 
                              (N792)? 1'b0 : 
                              (N793)? 1'b0 : 
                              (N794)? 1'b0 : 
                              (N795)? 1'b0 : 
                              (N796)? 1'b0 : 
                              (N797)? 1'b0 : 
                              (N798)? 1'b0 : 
                              (N799)? 1'b0 : 
                              (N800)? 1'b0 : 
                              (N801)? 1'b0 : 
                              (N802)? 1'b0 : 
                              (N803)? 1'b0 : 
                              (N804)? 1'b0 : 
                              (N805)? 1'b0 : 
                              (N806)? 1'b0 : 
                              (N807)? 1'b0 : 
                              (N808)? 1'b0 : 
                              (N809)? 1'b0 : 
                              (N810)? 1'b0 : 
                              (N811)? 1'b0 : 
                              (N812)? 1'b0 : 
                              (N813)? 1'b0 : 
                              (N814)? 1'b0 : 
                              (N815)? 1'b0 : 
                              (N816)? 1'b0 : 
                              (N817)? 1'b0 : 
                              (N818)? 1'b0 : 
                              (N819)? 1'b0 : 
                              (N820)? 1'b0 : 
                              (N821)? 1'b0 : 
                              (N822)? 1'b0 : 
                              (N823)? 1'b0 : 
                              (N824)? 1'b0 : 
                              (N825)? 1'b0 : 
                              (N826)? 1'b0 : 
                              (N827)? 1'b0 : 
                              (N828)? 1'b0 : 
                              (N829)? 1'b0 : 
                              (N830)? 1'b0 : 
                              (N831)? 1'b0 : 
                              (N832)? 1'b0 : 
                              (N833)? 1'b0 : 
                              (N834)? 1'b0 : 
                              (N835)? 1'b0 : 
                              (N836)? 1'b0 : 
                              (N837)? 1'b0 : 
                              (N838)? 1'b0 : 
                              (N839)? 1'b0 : 
                              (N840)? 1'b0 : 
                              (N841)? 1'b0 : 
                              (N842)? 1'b0 : 
                              (N843)? 1'b0 : 
                              (N844)? 1'b1 : 
                              (N845)? 1'b0 : 
                              (N846)? 1'b0 : 
                              (N847)? 1'b0 : 
                              (N848)? 1'b0 : 
                              (N849)? 1'b0 : 
                              (N850)? 1'b0 : 
                              (N851)? 1'b0 : 
                              (N852)? 1'b1 : 
                              (N853)? 1'b0 : 
                              (N854)? 1'b0 : 
                              (N855)? 1'b0 : 
                              (N856)? 1'b1 : 
                              (N857)? 1'b0 : 
                              (N858)? 1'b1 : 
                              (N859)? 1'b1 : 
                              (N860)? 1'b0 : 
                              (N861)? 1'b0 : 
                              (N862)? 1'b0 : 
                              (N863)? 1'b0 : 
                              (N864)? 1'b0 : 
                              (N865)? 1'b0 : 
                              (N866)? 1'b0 : 
                              (N867)? 1'b0 : 
                              (N868)? 1'b1 : 
                              (N869)? 1'b0 : 
                              (N870)? 1'b0 : 
                              (N871)? 1'b0 : 
                              (N872)? 1'b1 : 
                              (N873)? 1'b0 : 
                              (N874)? 1'b1 : 
                              (N875)? 1'b1 : 
                              (N876)? 1'b0 : 
                              (N877)? 1'b0 : 
                              (N878)? 1'b0 : 
                              (N879)? 1'b0 : 
                              (N880)? 1'b1 : 
                              (N881)? 1'b0 : 
                              (N882)? 1'b1 : 
                              (N883)? 1'b1 : 
                              (N884)? 1'b0 : 
                              (N885)? 1'b0 : 
                              (N886)? 1'b1 : 
                              (N887)? 1'b1 : 
                              (N888)? 1'b0 : 
                              (N889)? 1'b1 : 
                              (N890)? 1'b0 : 
                              (N891)? 1'b0 : 
                              (N892)? 1'b0 : 
                              (N893)? 1'b0 : 
                              (N894)? 1'b0 : 
                              (N895)? 1'b0 : 
                              (N896)? 1'b0 : 
                              (N897)? 1'b0 : 
                              (N898)? 1'b0 : 
                              (N899)? 1'b0 : 
                              (N900)? 1'b0 : 
                              (N901)? 1'b0 : 
                              (N902)? 1'b0 : 
                              (N903)? 1'b0 : 
                              (N904)? 1'b0 : 
                              (N905)? 1'b0 : 
                              (N906)? 1'b0 : 
                              (N907)? 1'b0 : 
                              (N908)? 1'b1 : 
                              (N909)? 1'b0 : 
                              (N910)? 1'b0 : 
                              (N911)? 1'b0 : 
                              (N912)? 1'b0 : 
                              (N913)? 1'b0 : 
                              (N914)? 1'b0 : 
                              (N915)? 1'b0 : 
                              (N916)? 1'b1 : 
                              (N917)? 1'b0 : 
                              (N918)? 1'b0 : 
                              (N919)? 1'b0 : 
                              (N920)? 1'b1 : 
                              (N921)? 1'b0 : 
                              (N922)? 1'b1 : 
                              (N923)? 1'b1 : 
                              (N924)? 1'b0 : 
                              (N925)? 1'b0 : 
                              (N926)? 1'b0 : 
                              (N927)? 1'b0 : 
                              (N928)? 1'b0 : 
                              (N929)? 1'b0 : 
                              (N930)? 1'b0 : 
                              (N931)? 1'b0 : 
                              (N932)? 1'b1 : 
                              (N933)? 1'b0 : 
                              (N934)? 1'b0 : 
                              (N935)? 1'b0 : 
                              (N936)? 1'b1 : 
                              (N937)? 1'b0 : 
                              (N938)? 1'b1 : 
                              (N939)? 1'b1 : 
                              (N940)? 1'b0 : 
                              (N941)? 1'b0 : 
                              (N942)? 1'b0 : 
                              (N943)? 1'b0 : 
                              (N944)? 1'b1 : 
                              (N945)? 1'b0 : 
                              (N946)? 1'b1 : 
                              (N947)? 1'b1 : 
                              (N948)? 1'b0 : 
                              (N949)? 1'b0 : 
                              (N950)? 1'b1 : 
                              (N951)? 1'b1 : 
                              (N952)? 1'b0 : 
                              (N953)? 1'b1 : 
                              (N954)? 1'b0 : 
                              (N955)? 1'b0 : 
                              (N956)? 1'b0 : 
                              (N957)? 1'b0 : 
                              (N958)? 1'b0 : 
                              (N959)? 1'b0 : 
                              (N960)? 1'b0 : 
                              (N961)? 1'b0 : 
                              (N962)? 1'b0 : 
                              (N963)? 1'b0 : 
                              (N964)? 1'b1 : 
                              (N965)? 1'b0 : 
                              (N966)? 1'b0 : 
                              (N967)? 1'b0 : 
                              (N968)? 1'b1 : 
                              (N969)? 1'b0 : 
                              (N970)? 1'b1 : 
                              (N971)? 1'b1 : 
                              (N972)? 1'b1 : 
                              (N973)? 1'b0 : 
                              (N974)? 1'b0 : 
                              (N975)? 1'b0 : 
                              (N976)? 1'b1 : 
                              (N977)? 1'b0 : 
                              (N978)? 1'b1 : 
                              (N979)? 1'b1 : 
                              (N980)? 1'b1 : 
                              (N981)? 1'b0 : 
                              (N982)? 1'b1 : 
                              (N983)? 1'b1 : 
                              (N984)? 1'b1 : 
                              (N985)? 1'b1 : 
                              (N986)? 1'b1 : 
                              (N987)? 1'b1 : 
                              (N988)? 1'b0 : 
                              (N989)? 1'b0 : 
                              (N990)? 1'b0 : 
                              (N991)? 1'b0 : 
                              (N992)? 1'b1 : 
                              (N993)? 1'b0 : 
                              (N994)? 1'b1 : 
                              (N995)? 1'b1 : 
                              (N996)? 1'b1 : 
                              (N997)? 1'b0 : 
                              (N998)? 1'b1 : 
                              (N999)? 1'b1 : 
                              (N1000)? 1'b1 : 
                              (N1001)? 1'b1 : 
                              (N1002)? 1'b1 : 
                              (N1003)? 1'b1 : 
                              (N1004)? 1'b0 : 
                              (N1005)? 1'b0 : 
                              (N1006)? 1'b1 : 
                              (N1007)? 1'b1 : 
                              (N1008)? 1'b1 : 
                              (N1009)? 1'b1 : 
                              (N1010)? 1'b1 : 
                              (N1011)? 1'b1 : 
                              (N1012)? 1'b0 : 
                              (N1013)? 1'b1 : 
                              (N1014)? 1'b1 : 
                              (N1015)? 1'b1 : 
                              (N1016)? 1'b0 : 
                              (N1017)? 1'b1 : 
                              (N1018)? 1'b0 : 
                              (N1019)? 1'b0 : 
                              (N255)? 1'b0 : 1'b0;
  assign N766 = N2827;
  assign N767 = N2829;
  assign N768 = N2831;
  assign N769 = N2833;
  assign N770 = N2835;
  assign N771 = N2837;
  assign N772 = N2839;
  assign N773 = N2841;
  assign N774 = N2843;
  assign N775 = N2845;
  assign N776 = N2847;
  assign N777 = N2849;
  assign N778 = N2851;
  assign N779 = N2853;
  assign N780 = N2855;
  assign N781 = N2857;
  assign N782 = N2859;
  assign N783 = N2861;
  assign N784 = N2863;
  assign N785 = N2866;
  assign N786 = N2868;
  assign N787 = N2870;
  assign N788 = N2872;
  assign N789 = N2874;
  assign N790 = N2876;
  assign N791 = N2878;
  assign N792 = N2880;
  assign N793 = N2882;
  assign N794 = N2884;
  assign N795 = N2886;
  assign N796 = N2888;
  assign N797 = N2890;
  assign N798 = N2892;
  assign N799 = N2894;
  assign N800 = N2896;
  assign N801 = N2899;
  assign N802 = N2901;
  assign N803 = N2903;
  assign N804 = N2905;
  assign N805 = N2907;
  assign N806 = N2909;
  assign N807 = N2911;
  assign N808 = N2913;
  assign N809 = N2915;
  assign N810 = N2917;
  assign N811 = N2919;
  assign N812 = N2921;
  assign N813 = N2923;
  assign N814 = N2925;
  assign N815 = N2927;
  assign N816 = N2929;
  assign N817 = N2932;
  assign N818 = N2934;
  assign N819 = N2936;
  assign N820 = N2938;
  assign N821 = N2940;
  assign N822 = N2943;
  assign N823 = N2946;
  assign N824 = N2949;
  assign N825 = N2955;
  assign N826 = N2957;
  assign N827 = N2959;
  assign N828 = N2962;
  assign N829 = N2965;
  assign N830 = N2968;
  assign N831 = N2971;
  assign N832 = N2974;
  assign N833 = N2978;
  assign N834 = N2981;
  assign N835 = N2984;
  assign N836 = N2987;
  assign N837 = N2991;
  assign N838 = N2994;
  assign N839 = N2996;
  assign N840 = N2998;
  assign N841 = N3000;
  assign N842 = N3002;
  assign N843 = N3004;
  assign N844 = N3006;
  assign N845 = N3008;
  assign N846 = N3010;
  assign N847 = N3012;
  assign N848 = N3014;
  assign N849 = N3018;
  assign N850 = N3020;
  assign N851 = N3022;
  assign N852 = N3024;
  assign N853 = N3026;
  assign N854 = N3028;
  assign N855 = N3030;
  assign N856 = N3032;
  assign N857 = N3036;
  assign N858 = N3038;
  assign N859 = N3040;
  assign N860 = N3042;
  assign N861 = N3044;
  assign N862 = N3046;
  assign N863 = N3048;
  assign N864 = N3050;
  assign N865 = N3054;
  assign N866 = N3056;
  assign N867 = N3058;
  assign N868 = N3060;
  assign N869 = N3062;
  assign N870 = N3064;
  assign N871 = N3066;
  assign N872 = N3068;
  assign N873 = N3070;
  assign N874 = N3072;
  assign N875 = N3074;
  assign N876 = N3076;
  assign N877 = N3078;
  assign N878 = N3080;
  assign N879 = N3082;
  assign N880 = N3084;
  assign N881 = N3087;
  assign N882 = N3089;
  assign N883 = N3091;
  assign N884 = N3093;
  assign N885 = N3095;
  assign N886 = N3097;
  assign N887 = N3099;
  assign N888 = N3101;
  assign N889 = N3103;
  assign N890 = N3105;
  assign N891 = N3107;
  assign N892 = N3109;
  assign N893 = N3112;
  assign N894 = N3114;
  assign N895 = N3116;
  assign N896 = N3118;
  assign N897 = N3120;
  assign N898 = N3122;
  assign N899 = N3124;
  assign N900 = N3126;
  assign N901 = N3128;
  assign N902 = N3130;
  assign N903 = N3132;
  assign N904 = N3134;
  assign N905 = N3136;
  assign N906 = N3138;
  assign N907 = N3140;
  assign N908 = N3142;
  assign N909 = N3144;
  assign N910 = N3146;
  assign N911 = N3148;
  assign N912 = N3150;
  assign N913 = N3153;
  assign N914 = N3155;
  assign N915 = N3157;
  assign N916 = N3159;
  assign N917 = N3161;
  assign N918 = N3163;
  assign N919 = N3165;
  assign N920 = N3167;
  assign N921 = N3171;
  assign N922 = N3173;
  assign N923 = N3175;
  assign N924 = N3177;
  assign N925 = N3179;
  assign N926 = N3181;
  assign N927 = N3183;
  assign N928 = N3185;
  assign N929 = N3188;
  assign N930 = N3190;
  assign N931 = N3192;
  assign N932 = N3194;
  assign N933 = N3196;
  assign N934 = N3198;
  assign N935 = N3200;
  assign N936 = N3202;
  assign N937 = N3204;
  assign N938 = N3206;
  assign N939 = N3208;
  assign N940 = N3210;
  assign N941 = N3212;
  assign N942 = N3214;
  assign N943 = N3216;
  assign N944 = N3218;
  assign N945 = N3221;
  assign N946 = N3223;
  assign N947 = N3225;
  assign N948 = N3227;
  assign N949 = N3229;
  assign N950 = N3231;
  assign N951 = N3233;
  assign N952 = N3235;
  assign N953 = N3237;
  assign N954 = N3239;
  assign N955 = N3241;
  assign N956 = N3243;
  assign N957 = N3247;
  assign N958 = N3249;
  assign N959 = N3251;
  assign N960 = N3253;
  assign N961 = N3255;
  assign N962 = N3257;
  assign N963 = N3259;
  assign N964 = N3261;
  assign N965 = N3263;
  assign N966 = N3265;
  assign N967 = N3267;
  assign N968 = N3269;
  assign N969 = N3271;
  assign N970 = N3273;
  assign N971 = N3275;
  assign N972 = N3277;
  assign N973 = N3279;
  assign N974 = N3281;
  assign N975 = N3283;
  assign N976 = N3285;
  assign N977 = N3288;
  assign N978 = N3290;
  assign N979 = N3292;
  assign N980 = N3294;
  assign N981 = N3296;
  assign N982 = N3298;
  assign N983 = N3300;
  assign N984 = N3302;
  assign N985 = N3304;
  assign N986 = N3306;
  assign N987 = N3308;
  assign N988 = N3310;
  assign N989 = N3312;
  assign N990 = N3314;
  assign N991 = N3316;
  assign N992 = N3318;
  assign N993 = N3321;
  assign N994 = N3323;
  assign N995 = N3325;
  assign N996 = N3327;
  assign N997 = N3329;
  assign N998 = N3331;
  assign N999 = N3333;
  assign N1000 = N3335;
  assign N1001 = N3337;
  assign N1002 = N3339;
  assign N1003 = N3341;
  assign N1004 = N3343;
  assign N1005 = N3345;
  assign N1006 = N3347;
  assign N1007 = N3349;
  assign N1008 = N3351;
  assign N1009 = N3354;
  assign N1010 = N3356;
  assign N1011 = N3358;
  assign N1012 = N3360;
  assign N1013 = N3362;
  assign N1014 = N3364;
  assign N1015 = N3368;
  assign N1016 = N3372;
  assign N1017 = N3374;
  assign N1018 = N3378;
  assign N1019 = N3381;
  assign fwd_datapath_o[10] = (N766)? 1'b0 : 
                              (N1)? 1'b0 : 
                              (N767)? 1'b0 : 
                              (N768)? 1'b0 : 
                              (N769)? 1'b0 : 
                              (N770)? 1'b0 : 
                              (N771)? 1'b0 : 
                              (N772)? 1'b0 : 
                              (N773)? 1'b0 : 
                              (N774)? 1'b0 : 
                              (N775)? 1'b0 : 
                              (N776)? 1'b0 : 
                              (N777)? 1'b0 : 
                              (N778)? 1'b0 : 
                              (N779)? 1'b0 : 
                              (N780)? 1'b0 : 
                              (N781)? 1'b0 : 
                              (N782)? 1'b0 : 
                              (N783)? 1'b0 : 
                              (N784)? 1'b0 : 
                              (N785)? 1'b0 : 
                              (N786)? 1'b0 : 
                              (N787)? 1'b0 : 
                              (N788)? 1'b0 : 
                              (N789)? 1'b0 : 
                              (N790)? 1'b0 : 
                              (N791)? 1'b0 : 
                              (N792)? 1'b0 : 
                              (N793)? 1'b0 : 
                              (N794)? 1'b0 : 
                              (N795)? 1'b0 : 
                              (N796)? 1'b0 : 
                              (N797)? 1'b0 : 
                              (N798)? 1'b0 : 
                              (N799)? 1'b0 : 
                              (N800)? 1'b0 : 
                              (N801)? 1'b0 : 
                              (N802)? 1'b0 : 
                              (N803)? 1'b0 : 
                              (N804)? 1'b1 : 
                              (N805)? 1'b0 : 
                              (N806)? 1'b0 : 
                              (N807)? 1'b0 : 
                              (N808)? 1'b1 : 
                              (N809)? 1'b0 : 
                              (N810)? 1'b1 : 
                              (N811)? 1'b1 : 
                              (N812)? 1'b0 : 
                              (N813)? 1'b0 : 
                              (N814)? 1'b0 : 
                              (N815)? 1'b0 : 
                              (N816)? 1'b1 : 
                              (N817)? 1'b0 : 
                              (N818)? 1'b1 : 
                              (N819)? 1'b1 : 
                              (N820)? 1'b0 : 
                              (N821)? 1'b0 : 
                              (N822)? 1'b1 : 
                              (N823)? 1'b1 : 
                              (N824)? 1'b0 : 
                              (N825)? 1'b1 : 
                              (N826)? 1'b0 : 
                              (N827)? 1'b0 : 
                              (N828)? 1'b0 : 
                              (N829)? 1'b0 : 
                              (N830)? 1'b0 : 
                              (N831)? 1'b0 : 
                              (N832)? 1'b0 : 
                              (N833)? 1'b0 : 
                              (N834)? 1'b0 : 
                              (N835)? 1'b0 : 
                              (N836)? 1'b1 : 
                              (N837)? 1'b0 : 
                              (N838)? 1'b0 : 
                              (N839)? 1'b0 : 
                              (N840)? 1'b1 : 
                              (N841)? 1'b0 : 
                              (N842)? 1'b1 : 
                              (N843)? 1'b1 : 
                              (N844)? 1'b0 : 
                              (N845)? 1'b0 : 
                              (N846)? 1'b0 : 
                              (N847)? 1'b0 : 
                              (N848)? 1'b1 : 
                              (N849)? 1'b0 : 
                              (N850)? 1'b1 : 
                              (N851)? 1'b1 : 
                              (N852)? 1'b0 : 
                              (N853)? 1'b0 : 
                              (N854)? 1'b1 : 
                              (N855)? 1'b1 : 
                              (N856)? 1'b0 : 
                              (N857)? 1'b1 : 
                              (N858)? 1'b0 : 
                              (N859)? 1'b0 : 
                              (N860)? 1'b0 : 
                              (N861)? 1'b0 : 
                              (N862)? 1'b0 : 
                              (N863)? 1'b0 : 
                              (N864)? 1'b1 : 
                              (N865)? 1'b0 : 
                              (N866)? 1'b1 : 
                              (N867)? 1'b1 : 
                              (N868)? 1'b1 : 
                              (N869)? 1'b0 : 
                              (N870)? 1'b1 : 
                              (N871)? 1'b1 : 
                              (N872)? 1'b1 : 
                              (N873)? 1'b1 : 
                              (N874)? 1'b1 : 
                              (N875)? 1'b1 : 
                              (N876)? 1'b0 : 
                              (N877)? 1'b0 : 
                              (N878)? 1'b1 : 
                              (N879)? 1'b1 : 
                              (N880)? 1'b1 : 
                              (N881)? 1'b1 : 
                              (N882)? 1'b1 : 
                              (N883)? 1'b1 : 
                              (N884)? 1'b0 : 
                              (N885)? 1'b1 : 
                              (N886)? 1'b1 : 
                              (N887)? 1'b1 : 
                              (N888)? 1'b0 : 
                              (N889)? 1'b1 : 
                              (N890)? 1'b0 : 
                              (N891)? 1'b0 : 
                              (N892)? 1'b0 : 
                              (N893)? 1'b0 : 
                              (N894)? 1'b0 : 
                              (N895)? 1'b0 : 
                              (N896)? 1'b0 : 
                              (N897)? 1'b0 : 
                              (N898)? 1'b0 : 
                              (N899)? 1'b0 : 
                              (N900)? 1'b0 : 
                              (N901)? 1'b0 : 
                              (N902)? 1'b0 : 
                              (N903)? 1'b0 : 
                              (N904)? 1'b0 : 
                              (N905)? 1'b0 : 
                              (N906)? 1'b0 : 
                              (N907)? 1'b0 : 
                              (N908)? 1'b0 : 
                              (N909)? 1'b0 : 
                              (N910)? 1'b0 : 
                              (N911)? 1'b0 : 
                              (N912)? 1'b0 : 
                              (N913)? 1'b0 : 
                              (N914)? 1'b0 : 
                              (N915)? 1'b0 : 
                              (N916)? 1'b0 : 
                              (N917)? 1'b0 : 
                              (N918)? 1'b0 : 
                              (N919)? 1'b0 : 
                              (N920)? 1'b0 : 
                              (N921)? 1'b0 : 
                              (N922)? 1'b0 : 
                              (N923)? 1'b0 : 
                              (N924)? 1'b0 : 
                              (N925)? 1'b0 : 
                              (N926)? 1'b0 : 
                              (N927)? 1'b0 : 
                              (N928)? 1'b0 : 
                              (N929)? 1'b0 : 
                              (N930)? 1'b0 : 
                              (N931)? 1'b0 : 
                              (N932)? 1'b1 : 
                              (N933)? 1'b0 : 
                              (N934)? 1'b0 : 
                              (N935)? 1'b0 : 
                              (N936)? 1'b1 : 
                              (N937)? 1'b0 : 
                              (N938)? 1'b1 : 
                              (N939)? 1'b1 : 
                              (N940)? 1'b0 : 
                              (N941)? 1'b0 : 
                              (N942)? 1'b0 : 
                              (N943)? 1'b0 : 
                              (N944)? 1'b1 : 
                              (N945)? 1'b0 : 
                              (N946)? 1'b1 : 
                              (N947)? 1'b1 : 
                              (N948)? 1'b0 : 
                              (N949)? 1'b0 : 
                              (N950)? 1'b1 : 
                              (N951)? 1'b1 : 
                              (N952)? 1'b0 : 
                              (N953)? 1'b1 : 
                              (N954)? 1'b0 : 
                              (N955)? 1'b0 : 
                              (N956)? 1'b0 : 
                              (N957)? 1'b0 : 
                              (N958)? 1'b0 : 
                              (N959)? 1'b0 : 
                              (N960)? 1'b0 : 
                              (N961)? 1'b0 : 
                              (N962)? 1'b0 : 
                              (N963)? 1'b0 : 
                              (N964)? 1'b1 : 
                              (N965)? 1'b0 : 
                              (N966)? 1'b0 : 
                              (N967)? 1'b0 : 
                              (N968)? 1'b1 : 
                              (N969)? 1'b0 : 
                              (N970)? 1'b1 : 
                              (N971)? 1'b1 : 
                              (N972)? 1'b0 : 
                              (N973)? 1'b0 : 
                              (N974)? 1'b0 : 
                              (N975)? 1'b0 : 
                              (N976)? 1'b1 : 
                              (N977)? 1'b0 : 
                              (N978)? 1'b1 : 
                              (N979)? 1'b1 : 
                              (N980)? 1'b0 : 
                              (N981)? 1'b0 : 
                              (N982)? 1'b1 : 
                              (N983)? 1'b1 : 
                              (N984)? 1'b0 : 
                              (N985)? 1'b1 : 
                              (N986)? 1'b0 : 
                              (N987)? 1'b0 : 
                              (N988)? 1'b0 : 
                              (N989)? 1'b0 : 
                              (N990)? 1'b0 : 
                              (N991)? 1'b0 : 
                              (N992)? 1'b1 : 
                              (N993)? 1'b0 : 
                              (N994)? 1'b1 : 
                              (N995)? 1'b1 : 
                              (N996)? 1'b1 : 
                              (N997)? 1'b0 : 
                              (N998)? 1'b1 : 
                              (N999)? 1'b1 : 
                              (N1000)? 1'b1 : 
                              (N1001)? 1'b1 : 
                              (N1002)? 1'b1 : 
                              (N1003)? 1'b1 : 
                              (N1004)? 1'b0 : 
                              (N1005)? 1'b0 : 
                              (N1006)? 1'b1 : 
                              (N1007)? 1'b1 : 
                              (N1008)? 1'b1 : 
                              (N1009)? 1'b1 : 
                              (N1010)? 1'b1 : 
                              (N1011)? 1'b1 : 
                              (N1012)? 1'b0 : 
                              (N1013)? 1'b1 : 
                              (N1014)? 1'b1 : 
                              (N1015)? 1'b1 : 
                              (N1016)? 1'b0 : 
                              (N1017)? 1'b1 : 
                              (N1018)? 1'b0 : 
                              (N1019)? 1'b0 : 
                              (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[9] = (N766)? 1'b0 : 
                             (N1)? 1'b0 : 
                             (N767)? 1'b0 : 
                             (N768)? 1'b0 : 
                             (N769)? 1'b0 : 
                             (N770)? 1'b0 : 
                             (N771)? 1'b0 : 
                             (N772)? 1'b0 : 
                             (N773)? 1'b0 : 
                             (N774)? 1'b0 : 
                             (N775)? 1'b0 : 
                             (N776)? 1'b0 : 
                             (N777)? 1'b0 : 
                             (N778)? 1'b0 : 
                             (N779)? 1'b0 : 
                             (N780)? 1'b0 : 
                             (N781)? 1'b0 : 
                             (N782)? 1'b0 : 
                             (N783)? 1'b0 : 
                             (N784)? 1'b0 : 
                             (N785)? 1'b0 : 
                             (N786)? 1'b0 : 
                             (N787)? 1'b0 : 
                             (N788)? 1'b1 : 
                             (N789)? 1'b0 : 
                             (N790)? 1'b0 : 
                             (N791)? 1'b0 : 
                             (N792)? 1'b1 : 
                             (N793)? 1'b0 : 
                             (N794)? 1'b1 : 
                             (N795)? 1'b1 : 
                             (N796)? 1'b0 : 
                             (N797)? 1'b0 : 
                             (N798)? 1'b0 : 
                             (N799)? 1'b0 : 
                             (N800)? 1'b0 : 
                             (N801)? 1'b0 : 
                             (N802)? 1'b0 : 
                             (N803)? 1'b0 : 
                             (N804)? 1'b0 : 
                             (N805)? 1'b0 : 
                             (N806)? 1'b0 : 
                             (N807)? 1'b0 : 
                             (N808)? 1'b0 : 
                             (N809)? 1'b0 : 
                             (N810)? 1'b0 : 
                             (N811)? 1'b0 : 
                             (N812)? 1'b0 : 
                             (N813)? 1'b0 : 
                             (N814)? 1'b0 : 
                             (N815)? 1'b0 : 
                             (N816)? 1'b0 : 
                             (N817)? 1'b0 : 
                             (N818)? 1'b0 : 
                             (N819)? 1'b0 : 
                             (N820)? 1'b1 : 
                             (N821)? 1'b0 : 
                             (N822)? 1'b0 : 
                             (N823)? 1'b0 : 
                             (N824)? 1'b1 : 
                             (N825)? 1'b0 : 
                             (N826)? 1'b1 : 
                             (N827)? 1'b1 : 
                             (N828)? 1'b0 : 
                             (N829)? 1'b0 : 
                             (N830)? 1'b0 : 
                             (N831)? 1'b0 : 
                             (N832)? 1'b0 : 
                             (N833)? 1'b0 : 
                             (N834)? 1'b0 : 
                             (N835)? 1'b0 : 
                             (N836)? 1'b1 : 
                             (N837)? 1'b0 : 
                             (N838)? 1'b0 : 
                             (N839)? 1'b0 : 
                             (N840)? 1'b1 : 
                             (N841)? 1'b0 : 
                             (N842)? 1'b1 : 
                             (N843)? 1'b1 : 
                             (N844)? 1'b0 : 
                             (N845)? 1'b0 : 
                             (N846)? 1'b0 : 
                             (N847)? 1'b0 : 
                             (N848)? 1'b1 : 
                             (N849)? 1'b0 : 
                             (N850)? 1'b1 : 
                             (N851)? 1'b1 : 
                             (N852)? 1'b1 : 
                             (N853)? 1'b0 : 
                             (N854)? 1'b1 : 
                             (N855)? 1'b1 : 
                             (N856)? 1'b1 : 
                             (N857)? 1'b1 : 
                             (N858)? 1'b1 : 
                             (N859)? 1'b1 : 
                             (N860)? 1'b0 : 
                             (N861)? 1'b0 : 
                             (N862)? 1'b0 : 
                             (N863)? 1'b0 : 
                             (N864)? 1'b1 : 
                             (N865)? 1'b0 : 
                             (N866)? 1'b1 : 
                             (N867)? 1'b1 : 
                             (N868)? 1'b0 : 
                             (N869)? 1'b0 : 
                             (N870)? 1'b1 : 
                             (N871)? 1'b1 : 
                             (N872)? 1'b0 : 
                             (N873)? 1'b1 : 
                             (N874)? 1'b0 : 
                             (N875)? 1'b0 : 
                             (N876)? 1'b0 : 
                             (N877)? 1'b0 : 
                             (N878)? 1'b1 : 
                             (N879)? 1'b1 : 
                             (N880)? 1'b0 : 
                             (N881)? 1'b1 : 
                             (N882)? 1'b0 : 
                             (N883)? 1'b0 : 
                             (N884)? 1'b1 : 
                             (N885)? 1'b1 : 
                             (N886)? 1'b0 : 
                             (N887)? 1'b0 : 
                             (N888)? 1'b1 : 
                             (N889)? 1'b0 : 
                             (N890)? 1'b1 : 
                             (N891)? 1'b1 : 
                             (N892)? 1'b0 : 
                             (N893)? 1'b0 : 
                             (N894)? 1'b0 : 
                             (N895)? 1'b0 : 
                             (N896)? 1'b0 : 
                             (N897)? 1'b0 : 
                             (N898)? 1'b0 : 
                             (N899)? 1'b0 : 
                             (N900)? 1'b0 : 
                             (N901)? 1'b0 : 
                             (N902)? 1'b0 : 
                             (N903)? 1'b0 : 
                             (N904)? 1'b0 : 
                             (N905)? 1'b0 : 
                             (N906)? 1'b0 : 
                             (N907)? 1'b0 : 
                             (N908)? 1'b0 : 
                             (N909)? 1'b0 : 
                             (N910)? 1'b0 : 
                             (N911)? 1'b0 : 
                             (N912)? 1'b0 : 
                             (N913)? 1'b0 : 
                             (N914)? 1'b0 : 
                             (N915)? 1'b0 : 
                             (N916)? 1'b1 : 
                             (N917)? 1'b0 : 
                             (N918)? 1'b0 : 
                             (N919)? 1'b0 : 
                             (N920)? 1'b1 : 
                             (N921)? 1'b0 : 
                             (N922)? 1'b1 : 
                             (N923)? 1'b1 : 
                             (N924)? 1'b0 : 
                             (N925)? 1'b0 : 
                             (N926)? 1'b0 : 
                             (N927)? 1'b0 : 
                             (N928)? 1'b0 : 
                             (N929)? 1'b0 : 
                             (N930)? 1'b0 : 
                             (N931)? 1'b0 : 
                             (N932)? 1'b0 : 
                             (N933)? 1'b0 : 
                             (N934)? 1'b0 : 
                             (N935)? 1'b0 : 
                             (N936)? 1'b0 : 
                             (N937)? 1'b0 : 
                             (N938)? 1'b0 : 
                             (N939)? 1'b0 : 
                             (N940)? 1'b0 : 
                             (N941)? 1'b0 : 
                             (N942)? 1'b0 : 
                             (N943)? 1'b0 : 
                             (N944)? 1'b0 : 
                             (N945)? 1'b0 : 
                             (N946)? 1'b0 : 
                             (N947)? 1'b0 : 
                             (N948)? 1'b1 : 
                             (N949)? 1'b0 : 
                             (N950)? 1'b0 : 
                             (N951)? 1'b0 : 
                             (N952)? 1'b1 : 
                             (N953)? 1'b0 : 
                             (N954)? 1'b1 : 
                             (N955)? 1'b1 : 
                             (N956)? 1'b0 : 
                             (N957)? 1'b0 : 
                             (N958)? 1'b0 : 
                             (N959)? 1'b0 : 
                             (N960)? 1'b0 : 
                             (N961)? 1'b0 : 
                             (N962)? 1'b0 : 
                             (N963)? 1'b0 : 
                             (N964)? 1'b1 : 
                             (N965)? 1'b0 : 
                             (N966)? 1'b0 : 
                             (N967)? 1'b0 : 
                             (N968)? 1'b1 : 
                             (N969)? 1'b0 : 
                             (N970)? 1'b1 : 
                             (N971)? 1'b1 : 
                             (N972)? 1'b0 : 
                             (N973)? 1'b0 : 
                             (N974)? 1'b0 : 
                             (N975)? 1'b0 : 
                             (N976)? 1'b1 : 
                             (N977)? 1'b0 : 
                             (N978)? 1'b1 : 
                             (N979)? 1'b1 : 
                             (N980)? 1'b1 : 
                             (N981)? 1'b0 : 
                             (N982)? 1'b1 : 
                             (N983)? 1'b1 : 
                             (N984)? 1'b1 : 
                             (N985)? 1'b1 : 
                             (N986)? 1'b1 : 
                             (N987)? 1'b1 : 
                             (N988)? 1'b0 : 
                             (N989)? 1'b0 : 
                             (N990)? 1'b0 : 
                             (N991)? 1'b0 : 
                             (N992)? 1'b1 : 
                             (N993)? 1'b0 : 
                             (N994)? 1'b1 : 
                             (N995)? 1'b1 : 
                             (N996)? 1'b0 : 
                             (N997)? 1'b0 : 
                             (N998)? 1'b1 : 
                             (N999)? 1'b1 : 
                             (N1000)? 1'b0 : 
                             (N1001)? 1'b1 : 
                             (N1002)? 1'b0 : 
                             (N1003)? 1'b0 : 
                             (N1004)? 1'b0 : 
                             (N1005)? 1'b0 : 
                             (N1006)? 1'b1 : 
                             (N1007)? 1'b1 : 
                             (N1008)? 1'b0 : 
                             (N1009)? 1'b1 : 
                             (N1010)? 1'b0 : 
                             (N1011)? 1'b0 : 
                             (N1012)? 1'b1 : 
                             (N1013)? 1'b1 : 
                             (N1014)? 1'b0 : 
                             (N1015)? 1'b0 : 
                             (N1016)? 1'b1 : 
                             (N1017)? 1'b0 : 
                             (N1018)? 1'b1 : 
                             (N1019)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[7] = (N766)? 1'b0 : 
                             (N1)? 1'b0 : 
                             (N767)? 1'b0 : 
                             (N768)? 1'b0 : 
                             (N769)? 1'b0 : 
                             (N770)? 1'b0 : 
                             (N771)? 1'b0 : 
                             (N772)? 1'b0 : 
                             (N773)? 1'b0 : 
                             (N774)? 1'b0 : 
                             (N775)? 1'b0 : 
                             (N776)? 1'b0 : 
                             (N777)? 1'b0 : 
                             (N778)? 1'b0 : 
                             (N779)? 1'b0 : 
                             (N780)? 1'b0 : 
                             (N781)? 1'b0 : 
                             (N782)? 1'b0 : 
                             (N783)? 1'b0 : 
                             (N784)? 1'b1 : 
                             (N785)? 1'b0 : 
                             (N786)? 1'b1 : 
                             (N787)? 1'b1 : 
                             (N788)? 1'b0 : 
                             (N789)? 1'b0 : 
                             (N790)? 1'b1 : 
                             (N791)? 1'b1 : 
                             (N792)? 1'b0 : 
                             (N793)? 1'b1 : 
                             (N794)? 1'b0 : 
                             (N795)? 1'b0 : 
                             (N796)? 1'b0 : 
                             (N797)? 1'b0 : 
                             (N798)? 1'b0 : 
                             (N799)? 1'b0 : 
                             (N800)? 1'b1 : 
                             (N801)? 1'b0 : 
                             (N802)? 1'b1 : 
                             (N803)? 1'b1 : 
                             (N804)? 1'b0 : 
                             (N805)? 1'b0 : 
                             (N806)? 1'b1 : 
                             (N807)? 1'b1 : 
                             (N808)? 1'b0 : 
                             (N809)? 1'b1 : 
                             (N810)? 1'b0 : 
                             (N811)? 1'b0 : 
                             (N812)? 1'b0 : 
                             (N813)? 1'b0 : 
                             (N814)? 1'b1 : 
                             (N815)? 1'b1 : 
                             (N816)? 1'b1 : 
                             (N817)? 1'b1 : 
                             (N818)? 1'b1 : 
                             (N819)? 1'b1 : 
                             (N820)? 1'b0 : 
                             (N821)? 1'b1 : 
                             (N822)? 1'b1 : 
                             (N823)? 1'b1 : 
                             (N824)? 1'b0 : 
                             (N825)? 1'b1 : 
                             (N826)? 1'b0 : 
                             (N827)? 1'b0 : 
                             (N828)? 1'b0 : 
                             (N829)? 1'b0 : 
                             (N830)? 1'b0 : 
                             (N831)? 1'b0 : 
                             (N832)? 1'b0 : 
                             (N833)? 1'b0 : 
                             (N834)? 1'b0 : 
                             (N835)? 1'b0 : 
                             (N836)? 1'b0 : 
                             (N837)? 1'b0 : 
                             (N838)? 1'b0 : 
                             (N839)? 1'b0 : 
                             (N840)? 1'b0 : 
                             (N841)? 1'b0 : 
                             (N842)? 1'b0 : 
                             (N843)? 1'b0 : 
                             (N844)? 1'b0 : 
                             (N845)? 1'b0 : 
                             (N846)? 1'b0 : 
                             (N847)? 1'b0 : 
                             (N848)? 1'b1 : 
                             (N849)? 1'b0 : 
                             (N850)? 1'b1 : 
                             (N851)? 1'b1 : 
                             (N852)? 1'b0 : 
                             (N853)? 1'b0 : 
                             (N854)? 1'b1 : 
                             (N855)? 1'b1 : 
                             (N856)? 1'b0 : 
                             (N857)? 1'b1 : 
                             (N858)? 1'b0 : 
                             (N859)? 1'b0 : 
                             (N860)? 1'b0 : 
                             (N861)? 1'b0 : 
                             (N862)? 1'b0 : 
                             (N863)? 1'b0 : 
                             (N864)? 1'b1 : 
                             (N865)? 1'b0 : 
                             (N866)? 1'b1 : 
                             (N867)? 1'b1 : 
                             (N868)? 1'b0 : 
                             (N869)? 1'b0 : 
                             (N870)? 1'b1 : 
                             (N871)? 1'b1 : 
                             (N872)? 1'b0 : 
                             (N873)? 1'b1 : 
                             (N874)? 1'b0 : 
                             (N875)? 1'b0 : 
                             (N876)? 1'b0 : 
                             (N877)? 1'b0 : 
                             (N878)? 1'b1 : 
                             (N879)? 1'b1 : 
                             (N880)? 1'b1 : 
                             (N881)? 1'b1 : 
                             (N882)? 1'b1 : 
                             (N883)? 1'b1 : 
                             (N884)? 1'b0 : 
                             (N885)? 1'b1 : 
                             (N886)? 1'b1 : 
                             (N887)? 1'b1 : 
                             (N888)? 1'b0 : 
                             (N889)? 1'b1 : 
                             (N890)? 1'b0 : 
                             (N891)? 1'b0 : 
                             (N892)? 1'b0 : 
                             (N893)? 1'b0 : 
                             (N894)? 1'b0 : 
                             (N895)? 1'b0 : 
                             (N896)? 1'b0 : 
                             (N897)? 1'b0 : 
                             (N898)? 1'b0 : 
                             (N899)? 1'b0 : 
                             (N900)? 1'b0 : 
                             (N901)? 1'b0 : 
                             (N902)? 1'b0 : 
                             (N903)? 1'b0 : 
                             (N904)? 1'b0 : 
                             (N905)? 1'b0 : 
                             (N906)? 1'b0 : 
                             (N907)? 1'b0 : 
                             (N908)? 1'b0 : 
                             (N909)? 1'b0 : 
                             (N910)? 1'b0 : 
                             (N911)? 1'b0 : 
                             (N912)? 1'b1 : 
                             (N913)? 1'b0 : 
                             (N914)? 1'b1 : 
                             (N915)? 1'b1 : 
                             (N916)? 1'b0 : 
                             (N917)? 1'b0 : 
                             (N918)? 1'b1 : 
                             (N919)? 1'b1 : 
                             (N920)? 1'b0 : 
                             (N921)? 1'b1 : 
                             (N922)? 1'b0 : 
                             (N923)? 1'b0 : 
                             (N924)? 1'b0 : 
                             (N925)? 1'b0 : 
                             (N926)? 1'b0 : 
                             (N927)? 1'b0 : 
                             (N928)? 1'b1 : 
                             (N929)? 1'b0 : 
                             (N930)? 1'b1 : 
                             (N931)? 1'b1 : 
                             (N932)? 1'b0 : 
                             (N933)? 1'b0 : 
                             (N934)? 1'b1 : 
                             (N935)? 1'b1 : 
                             (N936)? 1'b0 : 
                             (N937)? 1'b1 : 
                             (N938)? 1'b0 : 
                             (N939)? 1'b0 : 
                             (N940)? 1'b0 : 
                             (N941)? 1'b0 : 
                             (N942)? 1'b1 : 
                             (N943)? 1'b1 : 
                             (N944)? 1'b1 : 
                             (N945)? 1'b1 : 
                             (N946)? 1'b1 : 
                             (N947)? 1'b1 : 
                             (N948)? 1'b0 : 
                             (N949)? 1'b1 : 
                             (N950)? 1'b1 : 
                             (N951)? 1'b1 : 
                             (N952)? 1'b0 : 
                             (N953)? 1'b1 : 
                             (N954)? 1'b0 : 
                             (N955)? 1'b0 : 
                             (N956)? 1'b0 : 
                             (N957)? 1'b0 : 
                             (N958)? 1'b0 : 
                             (N959)? 1'b0 : 
                             (N960)? 1'b0 : 
                             (N961)? 1'b0 : 
                             (N962)? 1'b0 : 
                             (N963)? 1'b0 : 
                             (N964)? 1'b0 : 
                             (N965)? 1'b0 : 
                             (N966)? 1'b0 : 
                             (N967)? 1'b0 : 
                             (N968)? 1'b0 : 
                             (N969)? 1'b0 : 
                             (N970)? 1'b0 : 
                             (N971)? 1'b0 : 
                             (N972)? 1'b0 : 
                             (N973)? 1'b0 : 
                             (N974)? 1'b0 : 
                             (N975)? 1'b0 : 
                             (N976)? 1'b1 : 
                             (N977)? 1'b0 : 
                             (N978)? 1'b1 : 
                             (N979)? 1'b1 : 
                             (N980)? 1'b0 : 
                             (N981)? 1'b0 : 
                             (N982)? 1'b1 : 
                             (N983)? 1'b1 : 
                             (N984)? 1'b0 : 
                             (N985)? 1'b1 : 
                             (N986)? 1'b0 : 
                             (N987)? 1'b0 : 
                             (N988)? 1'b0 : 
                             (N989)? 1'b0 : 
                             (N990)? 1'b0 : 
                             (N991)? 1'b0 : 
                             (N992)? 1'b1 : 
                             (N993)? 1'b0 : 
                             (N994)? 1'b1 : 
                             (N995)? 1'b1 : 
                             (N996)? 1'b0 : 
                             (N997)? 1'b0 : 
                             (N998)? 1'b1 : 
                             (N999)? 1'b1 : 
                             (N1000)? 1'b0 : 
                             (N1001)? 1'b1 : 
                             (N1002)? 1'b0 : 
                             (N1003)? 1'b0 : 
                             (N1004)? 1'b0 : 
                             (N1005)? 1'b0 : 
                             (N1006)? 1'b1 : 
                             (N1007)? 1'b1 : 
                             (N1008)? 1'b1 : 
                             (N1009)? 1'b1 : 
                             (N1010)? 1'b1 : 
                             (N1011)? 1'b1 : 
                             (N1012)? 1'b0 : 
                             (N1013)? 1'b1 : 
                             (N1014)? 1'b1 : 
                             (N1015)? 1'b1 : 
                             (N1016)? 1'b0 : 
                             (N1017)? 1'b1 : 
                             (N1018)? 1'b0 : 
                             (N1019)? 1'b0 : 
                             (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[6] = (N766)? 1'b0 : 
                             (N1)? 1'b0 : 
                             (N767)? 1'b0 : 
                             (N768)? 1'b0 : 
                             (N769)? 1'b0 : 
                             (N770)? 1'b0 : 
                             (N771)? 1'b0 : 
                             (N772)? 1'b0 : 
                             (N773)? 1'b0 : 
                             (N774)? 1'b0 : 
                             (N775)? 1'b0 : 
                             (N776)? 1'b1 : 
                             (N777)? 1'b0 : 
                             (N778)? 1'b1 : 
                             (N779)? 1'b1 : 
                             (N780)? 1'b0 : 
                             (N781)? 1'b0 : 
                             (N782)? 1'b0 : 
                             (N783)? 1'b0 : 
                             (N784)? 1'b0 : 
                             (N785)? 1'b0 : 
                             (N786)? 1'b0 : 
                             (N787)? 1'b0 : 
                             (N788)? 1'b0 : 
                             (N789)? 1'b0 : 
                             (N790)? 1'b0 : 
                             (N791)? 1'b0 : 
                             (N792)? 1'b1 : 
                             (N793)? 1'b0 : 
                             (N794)? 1'b1 : 
                             (N795)? 1'b1 : 
                             (N796)? 1'b0 : 
                             (N797)? 1'b0 : 
                             (N798)? 1'b0 : 
                             (N799)? 1'b0 : 
                             (N800)? 1'b1 : 
                             (N801)? 1'b0 : 
                             (N802)? 1'b1 : 
                             (N803)? 1'b1 : 
                             (N804)? 1'b0 : 
                             (N805)? 1'b0 : 
                             (N806)? 1'b1 : 
                             (N807)? 1'b1 : 
                             (N808)? 1'b1 : 
                             (N809)? 1'b1 : 
                             (N810)? 1'b1 : 
                             (N811)? 1'b1 : 
                             (N812)? 1'b0 : 
                             (N813)? 1'b0 : 
                             (N814)? 1'b1 : 
                             (N815)? 1'b1 : 
                             (N816)? 1'b0 : 
                             (N817)? 1'b1 : 
                             (N818)? 1'b0 : 
                             (N819)? 1'b0 : 
                             (N820)? 1'b0 : 
                             (N821)? 1'b1 : 
                             (N822)? 1'b0 : 
                             (N823)? 1'b0 : 
                             (N824)? 1'b1 : 
                             (N825)? 1'b0 : 
                             (N826)? 1'b1 : 
                             (N827)? 1'b1 : 
                             (N828)? 1'b0 : 
                             (N829)? 1'b0 : 
                             (N830)? 1'b0 : 
                             (N831)? 1'b0 : 
                             (N832)? 1'b0 : 
                             (N833)? 1'b0 : 
                             (N834)? 1'b0 : 
                             (N835)? 1'b0 : 
                             (N836)? 1'b0 : 
                             (N837)? 1'b0 : 
                             (N838)? 1'b0 : 
                             (N839)? 1'b0 : 
                             (N840)? 1'b1 : 
                             (N841)? 1'b0 : 
                             (N842)? 1'b1 : 
                             (N843)? 1'b1 : 
                             (N844)? 1'b0 : 
                             (N845)? 1'b0 : 
                             (N846)? 1'b0 : 
                             (N847)? 1'b0 : 
                             (N848)? 1'b0 : 
                             (N849)? 1'b0 : 
                             (N850)? 1'b0 : 
                             (N851)? 1'b0 : 
                             (N852)? 1'b0 : 
                             (N853)? 1'b0 : 
                             (N854)? 1'b0 : 
                             (N855)? 1'b0 : 
                             (N856)? 1'b1 : 
                             (N857)? 1'b0 : 
                             (N858)? 1'b1 : 
                             (N859)? 1'b1 : 
                             (N860)? 1'b0 : 
                             (N861)? 1'b0 : 
                             (N862)? 1'b0 : 
                             (N863)? 1'b0 : 
                             (N864)? 1'b1 : 
                             (N865)? 1'b0 : 
                             (N866)? 1'b1 : 
                             (N867)? 1'b1 : 
                             (N868)? 1'b0 : 
                             (N869)? 1'b0 : 
                             (N870)? 1'b1 : 
                             (N871)? 1'b1 : 
                             (N872)? 1'b1 : 
                             (N873)? 1'b1 : 
                             (N874)? 1'b1 : 
                             (N875)? 1'b1 : 
                             (N876)? 1'b0 : 
                             (N877)? 1'b0 : 
                             (N878)? 1'b1 : 
                             (N879)? 1'b1 : 
                             (N880)? 1'b0 : 
                             (N881)? 1'b1 : 
                             (N882)? 1'b0 : 
                             (N883)? 1'b0 : 
                             (N884)? 1'b0 : 
                             (N885)? 1'b1 : 
                             (N886)? 1'b0 : 
                             (N887)? 1'b0 : 
                             (N888)? 1'b1 : 
                             (N889)? 1'b0 : 
                             (N890)? 1'b1 : 
                             (N891)? 1'b1 : 
                             (N892)? 1'b0 : 
                             (N893)? 1'b0 : 
                             (N894)? 1'b0 : 
                             (N895)? 1'b0 : 
                             (N896)? 1'b1 : 
                             (N897)? 1'b0 : 
                             (N898)? 1'b1 : 
                             (N899)? 1'b1 : 
                             (N900)? 1'b0 : 
                             (N901)? 1'b0 : 
                             (N902)? 1'b1 : 
                             (N903)? 1'b1 : 
                             (N904)? 1'b1 : 
                             (N905)? 1'b1 : 
                             (N906)? 1'b1 : 
                             (N907)? 1'b1 : 
                             (N908)? 1'b0 : 
                             (N909)? 1'b0 : 
                             (N910)? 1'b1 : 
                             (N911)? 1'b1 : 
                             (N912)? 1'b0 : 
                             (N913)? 1'b1 : 
                             (N914)? 1'b0 : 
                             (N915)? 1'b0 : 
                             (N916)? 1'b0 : 
                             (N917)? 1'b1 : 
                             (N918)? 1'b0 : 
                             (N919)? 1'b0 : 
                             (N920)? 1'b1 : 
                             (N921)? 1'b0 : 
                             (N922)? 1'b1 : 
                             (N923)? 1'b1 : 
                             (N924)? 1'b0 : 
                             (N925)? 1'b0 : 
                             (N926)? 1'b1 : 
                             (N927)? 1'b1 : 
                             (N928)? 1'b1 : 
                             (N929)? 1'b1 : 
                             (N930)? 1'b1 : 
                             (N931)? 1'b1 : 
                             (N932)? 1'b0 : 
                             (N933)? 1'b1 : 
                             (N934)? 1'b1 : 
                             (N935)? 1'b1 : 
                             (N936)? 1'b1 : 
                             (N937)? 1'b1 : 
                             (N938)? 1'b1 : 
                             (N939)? 1'b1 : 
                             (N940)? 1'b0 : 
                             (N941)? 1'b1 : 
                             (N942)? 1'b1 : 
                             (N943)? 1'b1 : 
                             (N944)? 1'b0 : 
                             (N945)? 1'b1 : 
                             (N946)? 1'b0 : 
                             (N947)? 1'b0 : 
                             (N948)? 1'b0 : 
                             (N949)? 1'b1 : 
                             (N950)? 1'b0 : 
                             (N951)? 1'b0 : 
                             (N952)? 1'b1 : 
                             (N953)? 1'b0 : 
                             (N954)? 1'b1 : 
                             (N955)? 1'b1 : 
                             (N956)? 1'b0 : 
                             (N957)? 1'b0 : 
                             (N958)? 1'b1 : 
                             (N959)? 1'b1 : 
                             (N960)? 1'b0 : 
                             (N961)? 1'b1 : 
                             (N962)? 1'b0 : 
                             (N963)? 1'b0 : 
                             (N964)? 1'b0 : 
                             (N965)? 1'b1 : 
                             (N966)? 1'b0 : 
                             (N967)? 1'b0 : 
                             (N968)? 1'b1 : 
                             (N969)? 1'b0 : 
                             (N970)? 1'b1 : 
                             (N971)? 1'b1 : 
                             (N972)? 1'b0 : 
                             (N973)? 1'b1 : 
                             (N974)? 1'b0 : 
                             (N975)? 1'b0 : 
                             (N976)? 1'b0 : 
                             (N977)? 1'b0 : 
                             (N978)? 1'b0 : 
                             (N979)? 1'b0 : 
                             (N980)? 1'b0 : 
                             (N981)? 1'b0 : 
                             (N982)? 1'b0 : 
                             (N983)? 1'b0 : 
                             (N984)? 1'b1 : 
                             (N985)? 1'b0 : 
                             (N986)? 1'b1 : 
                             (N987)? 1'b1 : 
                             (N988)? 1'b0 : 
                             (N989)? 1'b1 : 
                             (N990)? 1'b0 : 
                             (N991)? 1'b0 : 
                             (N992)? 1'b1 : 
                             (N993)? 1'b0 : 
                             (N994)? 1'b1 : 
                             (N995)? 1'b1 : 
                             (N996)? 1'b0 : 
                             (N997)? 1'b0 : 
                             (N998)? 1'b1 : 
                             (N999)? 1'b1 : 
                             (N1000)? 1'b1 : 
                             (N1001)? 1'b1 : 
                             (N1002)? 1'b1 : 
                             (N1003)? 1'b1 : 
                             (N1004)? 1'b0 : 
                             (N1005)? 1'b0 : 
                             (N1006)? 1'b1 : 
                             (N1007)? 1'b1 : 
                             (N1008)? 1'b0 : 
                             (N1009)? 1'b1 : 
                             (N1010)? 1'b0 : 
                             (N1011)? 1'b0 : 
                             (N1012)? 1'b0 : 
                             (N1013)? 1'b1 : 
                             (N1014)? 1'b0 : 
                             (N1015)? 1'b0 : 
                             (N1016)? 1'b1 : 
                             (N1017)? 1'b0 : 
                             (N1018)? 1'b1 : 
                             (N1019)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[4] = (N766)? 1'b0 : 
                             (N1)? 1'b0 : 
                             (N767)? 1'b0 : 
                             (N768)? 1'b0 : 
                             (N769)? 1'b0 : 
                             (N770)? 1'b0 : 
                             (N771)? 1'b0 : 
                             (N772)? 1'b0 : 
                             (N773)? 1'b0 : 
                             (N774)? 1'b1 : 
                             (N775)? 1'b1 : 
                             (N776)? 1'b0 : 
                             (N777)? 1'b1 : 
                             (N778)? 1'b0 : 
                             (N779)? 1'b0 : 
                             (N780)? 1'b0 : 
                             (N781)? 1'b0 : 
                             (N782)? 1'b1 : 
                             (N783)? 1'b1 : 
                             (N784)? 1'b0 : 
                             (N785)? 1'b1 : 
                             (N786)? 1'b0 : 
                             (N787)? 1'b0 : 
                             (N788)? 1'b0 : 
                             (N789)? 1'b1 : 
                             (N790)? 1'b1 : 
                             (N791)? 1'b1 : 
                             (N792)? 1'b0 : 
                             (N793)? 1'b1 : 
                             (N794)? 1'b0 : 
                             (N795)? 1'b0 : 
                             (N796)? 1'b0 : 
                             (N797)? 1'b0 : 
                             (N798)? 1'b0 : 
                             (N799)? 1'b0 : 
                             (N800)? 1'b0 : 
                             (N801)? 1'b0 : 
                             (N802)? 1'b0 : 
                             (N803)? 1'b0 : 
                             (N804)? 1'b0 : 
                             (N805)? 1'b0 : 
                             (N806)? 1'b1 : 
                             (N807)? 1'b1 : 
                             (N808)? 1'b0 : 
                             (N809)? 1'b1 : 
                             (N810)? 1'b0 : 
                             (N811)? 1'b0 : 
                             (N812)? 1'b0 : 
                             (N813)? 1'b0 : 
                             (N814)? 1'b1 : 
                             (N815)? 1'b1 : 
                             (N816)? 1'b0 : 
                             (N817)? 1'b1 : 
                             (N818)? 1'b0 : 
                             (N819)? 1'b0 : 
                             (N820)? 1'b0 : 
                             (N821)? 1'b1 : 
                             (N822)? 1'b1 : 
                             (N823)? 1'b1 : 
                             (N824)? 1'b0 : 
                             (N825)? 1'b1 : 
                             (N826)? 1'b0 : 
                             (N827)? 1'b0 : 
                             (N828)? 1'b0 : 
                             (N829)? 1'b0 : 
                             (N830)? 1'b0 : 
                             (N831)? 1'b0 : 
                             (N832)? 1'b0 : 
                             (N833)? 1'b0 : 
                             (N834)? 1'b0 : 
                             (N835)? 1'b0 : 
                             (N836)? 1'b0 : 
                             (N837)? 1'b0 : 
                             (N838)? 1'b1 : 
                             (N839)? 1'b1 : 
                             (N840)? 1'b0 : 
                             (N841)? 1'b1 : 
                             (N842)? 1'b0 : 
                             (N843)? 1'b0 : 
                             (N844)? 1'b0 : 
                             (N845)? 1'b0 : 
                             (N846)? 1'b1 : 
                             (N847)? 1'b1 : 
                             (N848)? 1'b0 : 
                             (N849)? 1'b1 : 
                             (N850)? 1'b0 : 
                             (N851)? 1'b0 : 
                             (N852)? 1'b0 : 
                             (N853)? 1'b1 : 
                             (N854)? 1'b1 : 
                             (N855)? 1'b1 : 
                             (N856)? 1'b0 : 
                             (N857)? 1'b1 : 
                             (N858)? 1'b0 : 
                             (N859)? 1'b0 : 
                             (N860)? 1'b0 : 
                             (N861)? 1'b0 : 
                             (N862)? 1'b0 : 
                             (N863)? 1'b0 : 
                             (N864)? 1'b0 : 
                             (N865)? 1'b0 : 
                             (N866)? 1'b0 : 
                             (N867)? 1'b0 : 
                             (N868)? 1'b0 : 
                             (N869)? 1'b0 : 
                             (N870)? 1'b1 : 
                             (N871)? 1'b1 : 
                             (N872)? 1'b0 : 
                             (N873)? 1'b1 : 
                             (N874)? 1'b0 : 
                             (N875)? 1'b0 : 
                             (N876)? 1'b0 : 
                             (N877)? 1'b0 : 
                             (N878)? 1'b1 : 
                             (N879)? 1'b1 : 
                             (N880)? 1'b0 : 
                             (N881)? 1'b1 : 
                             (N882)? 1'b0 : 
                             (N883)? 1'b0 : 
                             (N884)? 1'b0 : 
                             (N885)? 1'b1 : 
                             (N886)? 1'b1 : 
                             (N887)? 1'b1 : 
                             (N888)? 1'b0 : 
                             (N889)? 1'b1 : 
                             (N890)? 1'b0 : 
                             (N891)? 1'b0 : 
                             (N892)? 1'b0 : 
                             (N893)? 1'b0 : 
                             (N894)? 1'b1 : 
                             (N895)? 1'b1 : 
                             (N896)? 1'b0 : 
                             (N897)? 1'b1 : 
                             (N898)? 1'b0 : 
                             (N899)? 1'b0 : 
                             (N900)? 1'b0 : 
                             (N901)? 1'b1 : 
                             (N902)? 1'b1 : 
                             (N903)? 1'b1 : 
                             (N904)? 1'b0 : 
                             (N905)? 1'b1 : 
                             (N906)? 1'b0 : 
                             (N907)? 1'b0 : 
                             (N908)? 1'b0 : 
                             (N909)? 1'b1 : 
                             (N910)? 1'b1 : 
                             (N911)? 1'b1 : 
                             (N912)? 1'b0 : 
                             (N913)? 1'b1 : 
                             (N914)? 1'b0 : 
                             (N915)? 1'b0 : 
                             (N916)? 1'b0 : 
                             (N917)? 1'b1 : 
                             (N918)? 1'b1 : 
                             (N919)? 1'b1 : 
                             (N920)? 1'b0 : 
                             (N921)? 1'b1 : 
                             (N922)? 1'b0 : 
                             (N923)? 1'b0 : 
                             (N924)? 1'b0 : 
                             (N925)? 1'b1 : 
                             (N926)? 1'b0 : 
                             (N927)? 1'b0 : 
                             (N928)? 1'b0 : 
                             (N929)? 1'b0 : 
                             (N930)? 1'b0 : 
                             (N931)? 1'b0 : 
                             (N932)? 1'b0 : 
                             (N933)? 1'b0 : 
                             (N934)? 1'b1 : 
                             (N935)? 1'b1 : 
                             (N936)? 1'b0 : 
                             (N937)? 1'b1 : 
                             (N938)? 1'b0 : 
                             (N939)? 1'b0 : 
                             (N940)? 1'b0 : 
                             (N941)? 1'b0 : 
                             (N942)? 1'b1 : 
                             (N943)? 1'b1 : 
                             (N944)? 1'b0 : 
                             (N945)? 1'b1 : 
                             (N946)? 1'b0 : 
                             (N947)? 1'b0 : 
                             (N948)? 1'b0 : 
                             (N949)? 1'b1 : 
                             (N950)? 1'b1 : 
                             (N951)? 1'b1 : 
                             (N952)? 1'b0 : 
                             (N953)? 1'b1 : 
                             (N954)? 1'b0 : 
                             (N955)? 1'b0 : 
                             (N956)? 1'b0 : 
                             (N957)? 1'b1 : 
                             (N958)? 1'b0 : 
                             (N959)? 1'b0 : 
                             (N960)? 1'b0 : 
                             (N961)? 1'b0 : 
                             (N962)? 1'b0 : 
                             (N963)? 1'b0 : 
                             (N964)? 1'b0 : 
                             (N965)? 1'b0 : 
                             (N966)? 1'b1 : 
                             (N967)? 1'b1 : 
                             (N968)? 1'b0 : 
                             (N969)? 1'b1 : 
                             (N970)? 1'b0 : 
                             (N971)? 1'b0 : 
                             (N972)? 1'b0 : 
                             (N973)? 1'b0 : 
                             (N974)? 1'b1 : 
                             (N975)? 1'b1 : 
                             (N976)? 1'b0 : 
                             (N977)? 1'b1 : 
                             (N978)? 1'b0 : 
                             (N979)? 1'b0 : 
                             (N980)? 1'b0 : 
                             (N981)? 1'b1 : 
                             (N982)? 1'b1 : 
                             (N983)? 1'b1 : 
                             (N984)? 1'b0 : 
                             (N985)? 1'b1 : 
                             (N986)? 1'b0 : 
                             (N987)? 1'b0 : 
                             (N988)? 1'b0 : 
                             (N989)? 1'b0 : 
                             (N990)? 1'b0 : 
                             (N991)? 1'b0 : 
                             (N992)? 1'b0 : 
                             (N993)? 1'b0 : 
                             (N994)? 1'b0 : 
                             (N995)? 1'b0 : 
                             (N996)? 1'b0 : 
                             (N997)? 1'b0 : 
                             (N998)? 1'b1 : 
                             (N999)? 1'b1 : 
                             (N1000)? 1'b0 : 
                             (N1001)? 1'b1 : 
                             (N1002)? 1'b0 : 
                             (N1003)? 1'b0 : 
                             (N1004)? 1'b0 : 
                             (N1005)? 1'b0 : 
                             (N1006)? 1'b1 : 
                             (N1007)? 1'b1 : 
                             (N1008)? 1'b0 : 
                             (N1009)? 1'b1 : 
                             (N1010)? 1'b0 : 
                             (N1011)? 1'b0 : 
                             (N1012)? 1'b0 : 
                             (N1013)? 1'b1 : 
                             (N1014)? 1'b1 : 
                             (N1015)? 1'b1 : 
                             (N1016)? 1'b0 : 
                             (N1017)? 1'b1 : 
                             (N1018)? 1'b0 : 
                             (N1019)? 1'b0 : 
                             (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[3] = (N766)? 1'b0 : 
                             (N1)? 1'b0 : 
                             (N767)? 1'b0 : 
                             (N768)? 1'b0 : 
                             (N769)? 1'b0 : 
                             (N770)? 1'b1 : 
                             (N771)? 1'b1 : 
                             (N772)? 1'b0 : 
                             (N773)? 1'b0 : 
                             (N774)? 1'b0 : 
                             (N775)? 1'b0 : 
                             (N776)? 1'b0 : 
                             (N777)? 1'b0 : 
                             (N778)? 1'b1 : 
                             (N779)? 1'b1 : 
                             (N780)? 1'b0 : 
                             (N781)? 1'b0 : 
                             (N782)? 1'b1 : 
                             (N783)? 1'b1 : 
                             (N784)? 1'b0 : 
                             (N785)? 1'b1 : 
                             (N786)? 1'b1 : 
                             (N787)? 1'b1 : 
                             (N788)? 1'b0 : 
                             (N789)? 1'b1 : 
                             (N790)? 1'b0 : 
                             (N791)? 1'b0 : 
                             (N792)? 1'b0 : 
                             (N793)? 1'b0 : 
                             (N794)? 1'b1 : 
                             (N795)? 1'b1 : 
                             (N796)? 1'b0 : 
                             (N797)? 1'b0 : 
                             (N798)? 1'b0 : 
                             (N799)? 1'b0 : 
                             (N800)? 1'b0 : 
                             (N801)? 1'b0 : 
                             (N802)? 1'b1 : 
                             (N803)? 1'b1 : 
                             (N804)? 1'b0 : 
                             (N805)? 1'b0 : 
                             (N806)? 1'b0 : 
                             (N807)? 1'b0 : 
                             (N808)? 1'b0 : 
                             (N809)? 1'b0 : 
                             (N810)? 1'b1 : 
                             (N811)? 1'b1 : 
                             (N812)? 1'b0 : 
                             (N813)? 1'b0 : 
                             (N814)? 1'b1 : 
                             (N815)? 1'b1 : 
                             (N816)? 1'b0 : 
                             (N817)? 1'b1 : 
                             (N818)? 1'b1 : 
                             (N819)? 1'b1 : 
                             (N820)? 1'b0 : 
                             (N821)? 1'b1 : 
                             (N822)? 1'b0 : 
                             (N823)? 1'b0 : 
                             (N824)? 1'b0 : 
                             (N825)? 1'b0 : 
                             (N826)? 1'b1 : 
                             (N827)? 1'b1 : 
                             (N828)? 1'b0 : 
                             (N829)? 1'b0 : 
                             (N830)? 1'b1 : 
                             (N831)? 1'b1 : 
                             (N832)? 1'b0 : 
                             (N833)? 1'b1 : 
                             (N834)? 1'b1 : 
                             (N835)? 1'b1 : 
                             (N836)? 1'b0 : 
                             (N837)? 1'b1 : 
                             (N838)? 1'b0 : 
                             (N839)? 1'b0 : 
                             (N840)? 1'b0 : 
                             (N841)? 1'b0 : 
                             (N842)? 1'b1 : 
                             (N843)? 1'b1 : 
                             (N844)? 1'b0 : 
                             (N845)? 1'b1 : 
                             (N846)? 1'b1 : 
                             (N847)? 1'b1 : 
                             (N848)? 1'b0 : 
                             (N849)? 1'b1 : 
                             (N850)? 1'b1 : 
                             (N851)? 1'b1 : 
                             (N852)? 1'b0 : 
                             (N853)? 1'b1 : 
                             (N854)? 1'b0 : 
                             (N855)? 1'b0 : 
                             (N856)? 1'b0 : 
                             (N857)? 1'b0 : 
                             (N858)? 1'b1 : 
                             (N859)? 1'b1 : 
                             (N860)? 1'b0 : 
                             (N861)? 1'b1 : 
                             (N862)? 1'b0 : 
                             (N863)? 1'b0 : 
                             (N864)? 1'b0 : 
                             (N865)? 1'b0 : 
                             (N866)? 1'b1 : 
                             (N867)? 1'b1 : 
                             (N868)? 1'b0 : 
                             (N869)? 1'b0 : 
                             (N870)? 1'b0 : 
                             (N871)? 1'b0 : 
                             (N872)? 1'b0 : 
                             (N873)? 1'b0 : 
                             (N874)? 1'b1 : 
                             (N875)? 1'b1 : 
                             (N876)? 1'b0 : 
                             (N877)? 1'b0 : 
                             (N878)? 1'b1 : 
                             (N879)? 1'b1 : 
                             (N880)? 1'b0 : 
                             (N881)? 1'b1 : 
                             (N882)? 1'b1 : 
                             (N883)? 1'b1 : 
                             (N884)? 1'b0 : 
                             (N885)? 1'b1 : 
                             (N886)? 1'b0 : 
                             (N887)? 1'b0 : 
                             (N888)? 1'b0 : 
                             (N889)? 1'b0 : 
                             (N890)? 1'b1 : 
                             (N891)? 1'b1 : 
                             (N892)? 1'b0 : 
                             (N893)? 1'b0 : 
                             (N894)? 1'b0 : 
                             (N895)? 1'b0 : 
                             (N896)? 1'b0 : 
                             (N897)? 1'b0 : 
                             (N898)? 1'b1 : 
                             (N899)? 1'b1 : 
                             (N900)? 1'b0 : 
                             (N901)? 1'b0 : 
                             (N902)? 1'b0 : 
                             (N903)? 1'b0 : 
                             (N904)? 1'b0 : 
                             (N905)? 1'b0 : 
                             (N906)? 1'b1 : 
                             (N907)? 1'b1 : 
                             (N908)? 1'b0 : 
                             (N909)? 1'b0 : 
                             (N910)? 1'b1 : 
                             (N911)? 1'b1 : 
                             (N912)? 1'b0 : 
                             (N913)? 1'b1 : 
                             (N914)? 1'b1 : 
                             (N915)? 1'b1 : 
                             (N916)? 1'b0 : 
                             (N917)? 1'b1 : 
                             (N918)? 1'b0 : 
                             (N919)? 1'b0 : 
                             (N920)? 1'b0 : 
                             (N921)? 1'b0 : 
                             (N922)? 1'b1 : 
                             (N923)? 1'b1 : 
                             (N924)? 1'b0 : 
                             (N925)? 1'b0 : 
                             (N926)? 1'b0 : 
                             (N927)? 1'b0 : 
                             (N928)? 1'b0 : 
                             (N929)? 1'b0 : 
                             (N930)? 1'b1 : 
                             (N931)? 1'b1 : 
                             (N932)? 1'b0 : 
                             (N933)? 1'b0 : 
                             (N934)? 1'b0 : 
                             (N935)? 1'b0 : 
                             (N936)? 1'b0 : 
                             (N937)? 1'b0 : 
                             (N938)? 1'b1 : 
                             (N939)? 1'b1 : 
                             (N940)? 1'b0 : 
                             (N941)? 1'b0 : 
                             (N942)? 1'b1 : 
                             (N943)? 1'b1 : 
                             (N944)? 1'b0 : 
                             (N945)? 1'b1 : 
                             (N946)? 1'b1 : 
                             (N947)? 1'b1 : 
                             (N948)? 1'b0 : 
                             (N949)? 1'b1 : 
                             (N950)? 1'b0 : 
                             (N951)? 1'b0 : 
                             (N952)? 1'b0 : 
                             (N953)? 1'b0 : 
                             (N954)? 1'b1 : 
                             (N955)? 1'b1 : 
                             (N956)? 1'b0 : 
                             (N957)? 1'b0 : 
                             (N958)? 1'b1 : 
                             (N959)? 1'b1 : 
                             (N960)? 1'b0 : 
                             (N961)? 1'b1 : 
                             (N962)? 1'b1 : 
                             (N963)? 1'b1 : 
                             (N964)? 1'b0 : 
                             (N965)? 1'b1 : 
                             (N966)? 1'b0 : 
                             (N967)? 1'b0 : 
                             (N968)? 1'b0 : 
                             (N969)? 1'b0 : 
                             (N970)? 1'b1 : 
                             (N971)? 1'b1 : 
                             (N972)? 1'b0 : 
                             (N973)? 1'b1 : 
                             (N974)? 1'b1 : 
                             (N975)? 1'b1 : 
                             (N976)? 1'b0 : 
                             (N977)? 1'b1 : 
                             (N978)? 1'b1 : 
                             (N979)? 1'b1 : 
                             (N980)? 1'b0 : 
                             (N981)? 1'b1 : 
                             (N982)? 1'b0 : 
                             (N983)? 1'b0 : 
                             (N984)? 1'b0 : 
                             (N985)? 1'b0 : 
                             (N986)? 1'b1 : 
                             (N987)? 1'b1 : 
                             (N988)? 1'b0 : 
                             (N989)? 1'b1 : 
                             (N990)? 1'b0 : 
                             (N991)? 1'b0 : 
                             (N992)? 1'b0 : 
                             (N993)? 1'b0 : 
                             (N994)? 1'b1 : 
                             (N995)? 1'b1 : 
                             (N996)? 1'b0 : 
                             (N997)? 1'b0 : 
                             (N998)? 1'b0 : 
                             (N999)? 1'b0 : 
                             (N1000)? 1'b0 : 
                             (N1001)? 1'b0 : 
                             (N1002)? 1'b1 : 
                             (N1003)? 1'b1 : 
                             (N1004)? 1'b0 : 
                             (N1005)? 1'b0 : 
                             (N1006)? 1'b1 : 
                             (N1007)? 1'b1 : 
                             (N1008)? 1'b0 : 
                             (N1009)? 1'b1 : 
                             (N1010)? 1'b1 : 
                             (N1011)? 1'b1 : 
                             (N1012)? 1'b0 : 
                             (N1013)? 1'b1 : 
                             (N1014)? 1'b0 : 
                             (N1015)? 1'b0 : 
                             (N1016)? 1'b0 : 
                             (N1017)? 1'b0 : 
                             (N1018)? 1'b1 : 
                             (N1019)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign fwd_datapath_o[0] = (N766)? 1'b0 : 
                             (N1)? 1'b0 : 
                             (N767)? 1'b1 : 
                             (N768)? 1'b0 : 
                             (N769)? 1'b0 : 
                             (N770)? 1'b0 : 
                             (N771)? 1'b1 : 
                             (N772)? 1'b0 : 
                             (N773)? 1'b1 : 
                             (N774)? 1'b0 : 
                             (N775)? 1'b1 : 
                             (N776)? 1'b0 : 
                             (N777)? 1'b0 : 
                             (N778)? 1'b0 : 
                             (N779)? 1'b1 : 
                             (N780)? 1'b0 : 
                             (N781)? 1'b0 : 
                             (N782)? 1'b0 : 
                             (N783)? 1'b1 : 
                             (N784)? 1'b0 : 
                             (N785)? 1'b0 : 
                             (N786)? 1'b0 : 
                             (N787)? 1'b1 : 
                             (N788)? 1'b0 : 
                             (N789)? 1'b1 : 
                             (N790)? 1'b0 : 
                             (N791)? 1'b1 : 
                             (N792)? 1'b0 : 
                             (N793)? 1'b0 : 
                             (N794)? 1'b0 : 
                             (N795)? 1'b1 : 
                             (N796)? 1'b0 : 
                             (N797)? 1'b1 : 
                             (N798)? 1'b0 : 
                             (N799)? 1'b1 : 
                             (N800)? 1'b0 : 
                             (N801)? 1'b0 : 
                             (N802)? 1'b0 : 
                             (N803)? 1'b1 : 
                             (N804)? 1'b0 : 
                             (N805)? 1'b1 : 
                             (N806)? 1'b0 : 
                             (N807)? 1'b1 : 
                             (N808)? 1'b0 : 
                             (N809)? 1'b0 : 
                             (N810)? 1'b0 : 
                             (N811)? 1'b1 : 
                             (N812)? 1'b0 : 
                             (N813)? 1'b0 : 
                             (N814)? 1'b0 : 
                             (N815)? 1'b1 : 
                             (N816)? 1'b0 : 
                             (N817)? 1'b0 : 
                             (N818)? 1'b0 : 
                             (N819)? 1'b1 : 
                             (N820)? 1'b0 : 
                             (N821)? 1'b1 : 
                             (N822)? 1'b0 : 
                             (N823)? 1'b1 : 
                             (N824)? 1'b0 : 
                             (N825)? 1'b0 : 
                             (N826)? 1'b0 : 
                             (N827)? 1'b1 : 
                             (N828)? 1'b0 : 
                             (N829)? 1'b0 : 
                             (N830)? 1'b0 : 
                             (N831)? 1'b1 : 
                             (N832)? 1'b0 : 
                             (N833)? 1'b0 : 
                             (N834)? 1'b0 : 
                             (N835)? 1'b1 : 
                             (N836)? 1'b0 : 
                             (N837)? 1'b1 : 
                             (N838)? 1'b0 : 
                             (N839)? 1'b1 : 
                             (N840)? 1'b0 : 
                             (N841)? 1'b0 : 
                             (N842)? 1'b0 : 
                             (N843)? 1'b1 : 
                             (N844)? 1'b0 : 
                             (N845)? 1'b0 : 
                             (N846)? 1'b0 : 
                             (N847)? 1'b1 : 
                             (N848)? 1'b0 : 
                             (N849)? 1'b0 : 
                             (N850)? 1'b0 : 
                             (N851)? 1'b1 : 
                             (N852)? 1'b0 : 
                             (N853)? 1'b1 : 
                             (N854)? 1'b0 : 
                             (N855)? 1'b1 : 
                             (N856)? 1'b0 : 
                             (N857)? 1'b0 : 
                             (N858)? 1'b0 : 
                             (N859)? 1'b1 : 
                             (N860)? 1'b0 : 
                             (N861)? 1'b1 : 
                             (N862)? 1'b0 : 
                             (N863)? 1'b1 : 
                             (N864)? 1'b0 : 
                             (N865)? 1'b0 : 
                             (N866)? 1'b0 : 
                             (N867)? 1'b1 : 
                             (N868)? 1'b0 : 
                             (N869)? 1'b1 : 
                             (N870)? 1'b0 : 
                             (N871)? 1'b1 : 
                             (N872)? 1'b0 : 
                             (N873)? 1'b0 : 
                             (N874)? 1'b0 : 
                             (N875)? 1'b1 : 
                             (N876)? 1'b0 : 
                             (N877)? 1'b0 : 
                             (N878)? 1'b0 : 
                             (N879)? 1'b1 : 
                             (N880)? 1'b0 : 
                             (N881)? 1'b0 : 
                             (N882)? 1'b0 : 
                             (N883)? 1'b1 : 
                             (N884)? 1'b0 : 
                             (N885)? 1'b1 : 
                             (N886)? 1'b0 : 
                             (N887)? 1'b1 : 
                             (N888)? 1'b0 : 
                             (N889)? 1'b0 : 
                             (N890)? 1'b0 : 
                             (N891)? 1'b1 : 
                             (N892)? 1'b0 : 
                             (N893)? 1'b1 : 
                             (N894)? 1'b0 : 
                             (N895)? 1'b1 : 
                             (N896)? 1'b0 : 
                             (N897)? 1'b0 : 
                             (N898)? 1'b0 : 
                             (N899)? 1'b1 : 
                             (N900)? 1'b0 : 
                             (N901)? 1'b1 : 
                             (N902)? 1'b0 : 
                             (N903)? 1'b1 : 
                             (N904)? 1'b0 : 
                             (N905)? 1'b0 : 
                             (N906)? 1'b0 : 
                             (N907)? 1'b1 : 
                             (N908)? 1'b0 : 
                             (N909)? 1'b0 : 
                             (N910)? 1'b0 : 
                             (N911)? 1'b1 : 
                             (N912)? 1'b0 : 
                             (N913)? 1'b0 : 
                             (N914)? 1'b0 : 
                             (N915)? 1'b1 : 
                             (N916)? 1'b0 : 
                             (N917)? 1'b1 : 
                             (N918)? 1'b0 : 
                             (N919)? 1'b1 : 
                             (N920)? 1'b0 : 
                             (N921)? 1'b0 : 
                             (N922)? 1'b0 : 
                             (N923)? 1'b1 : 
                             (N924)? 1'b0 : 
                             (N925)? 1'b1 : 
                             (N926)? 1'b0 : 
                             (N927)? 1'b1 : 
                             (N928)? 1'b0 : 
                             (N929)? 1'b0 : 
                             (N930)? 1'b0 : 
                             (N931)? 1'b1 : 
                             (N932)? 1'b0 : 
                             (N933)? 1'b1 : 
                             (N934)? 1'b0 : 
                             (N935)? 1'b1 : 
                             (N936)? 1'b0 : 
                             (N937)? 1'b0 : 
                             (N938)? 1'b0 : 
                             (N939)? 1'b1 : 
                             (N940)? 1'b0 : 
                             (N941)? 1'b0 : 
                             (N942)? 1'b0 : 
                             (N943)? 1'b1 : 
                             (N944)? 1'b0 : 
                             (N945)? 1'b0 : 
                             (N946)? 1'b0 : 
                             (N947)? 1'b1 : 
                             (N948)? 1'b0 : 
                             (N949)? 1'b1 : 
                             (N950)? 1'b0 : 
                             (N951)? 1'b1 : 
                             (N952)? 1'b0 : 
                             (N953)? 1'b0 : 
                             (N954)? 1'b0 : 
                             (N955)? 1'b1 : 
                             (N956)? 1'b0 : 
                             (N957)? 1'b0 : 
                             (N958)? 1'b0 : 
                             (N959)? 1'b1 : 
                             (N960)? 1'b0 : 
                             (N961)? 1'b0 : 
                             (N962)? 1'b0 : 
                             (N963)? 1'b1 : 
                             (N964)? 1'b0 : 
                             (N965)? 1'b1 : 
                             (N966)? 1'b0 : 
                             (N967)? 1'b1 : 
                             (N968)? 1'b0 : 
                             (N969)? 1'b0 : 
                             (N970)? 1'b0 : 
                             (N971)? 1'b1 : 
                             (N972)? 1'b0 : 
                             (N973)? 1'b0 : 
                             (N974)? 1'b0 : 
                             (N975)? 1'b1 : 
                             (N976)? 1'b0 : 
                             (N977)? 1'b0 : 
                             (N978)? 1'b0 : 
                             (N979)? 1'b1 : 
                             (N980)? 1'b0 : 
                             (N981)? 1'b1 : 
                             (N982)? 1'b0 : 
                             (N983)? 1'b1 : 
                             (N984)? 1'b0 : 
                             (N985)? 1'b0 : 
                             (N986)? 1'b0 : 
                             (N987)? 1'b1 : 
                             (N988)? 1'b0 : 
                             (N989)? 1'b1 : 
                             (N990)? 1'b0 : 
                             (N991)? 1'b1 : 
                             (N992)? 1'b0 : 
                             (N993)? 1'b0 : 
                             (N994)? 1'b0 : 
                             (N995)? 1'b1 : 
                             (N996)? 1'b0 : 
                             (N997)? 1'b1 : 
                             (N998)? 1'b0 : 
                             (N999)? 1'b1 : 
                             (N1000)? 1'b0 : 
                             (N1001)? 1'b0 : 
                             (N1002)? 1'b0 : 
                             (N1003)? 1'b1 : 
                             (N1004)? 1'b0 : 
                             (N1005)? 1'b0 : 
                             (N1006)? 1'b0 : 
                             (N1007)? 1'b1 : 
                             (N1008)? 1'b0 : 
                             (N1009)? 1'b0 : 
                             (N1010)? 1'b0 : 
                             (N1011)? 1'b1 : 
                             (N1012)? 1'b0 : 
                             (N1013)? 1'b1 : 
                             (N1014)? 1'b0 : 
                             (N1015)? 1'b1 : 
                             (N1016)? 1'b0 : 
                             (N1017)? 1'b0 : 
                             (N1018)? 1'b0 : 
                             (N1019)? 1'b1 : 
                             (N255)? 1'b0 : 1'b0;
  assign N1020 = ~vec_i[7];
  assign N1021 = ~vec_i[6];
  assign N1022 = ~vec_i[5];
  assign N1023 = ~vec_i[4];
  assign N1024 = ~vec_i[3];
  assign N1025 = ~vec_i[2];
  assign N1026 = ~vec_i[1];
  assign N1027 = ~vec_i[0];
  assign N1042 = ~N1041;
  assign N1050 = ~N1049;
  assign N1058 = ~N1057;
  assign N1063 = ~N1062;
  assign N1068 = ~N1067;
  assign N1073 = ~N1072;
  assign N1078 = ~N1077;
  assign N1083 = ~N1082;
  assign N1088 = ~N1087;
  assign N1093 = ~N1092;
  assign N1098 = ~N1097;
  assign N1103 = ~N1102;
  assign N1106 = ~N1105;
  assign N1109 = ~N1108;
  assign N1112 = ~N1111;
  assign N1117 = ~N1116;
  assign N1122 = ~N1121;
  assign N1127 = ~N1126;
  assign N1132 = ~N1131;
  assign N1138 = ~N1137;
  assign N1141 = ~N1140;
  assign N1144 = ~N1143;
  assign N1147 = ~N1146;
  assign N1151 = ~N1150;
  assign N1154 = ~N1153;
  assign N1157 = ~N1156;
  assign N1160 = ~N1159;
  assign N1162 = ~N1161;
  assign N1164 = ~N1163;
  assign N1166 = ~N1165;
  assign N1168 = ~N1167;
  assign N1172 = ~N1171;
  assign N1178 = ~N1177;
  assign N1184 = ~N1183;
  assign N1189 = ~N1188;
  assign N1194 = ~N1193;
  assign N1197 = ~N1196;
  assign N1200 = ~N1199;
  assign N1202 = ~N1201;
  assign N1205 = ~N1204;
  assign N1208 = ~N1207;
  assign N1211 = ~N1210;
  assign N1214 = ~N1213;
  assign N1218 = ~N1217;
  assign N1221 = ~N1220;
  assign N1224 = ~N1223;
  assign N1227 = ~N1226;
  assign N1231 = ~N1230;
  assign N1233 = ~N1232;
  assign N1235 = ~N1234;
  assign N1237 = ~N1236;
  assign N1239 = ~N1238;
  assign N1241 = ~N1240;
  assign N1243 = ~N1242;
  assign N1246 = ~N1245;
  assign N1248 = ~N1247;
  assign N1250 = ~N1249;
  assign N1252 = ~N1251;
  assign N1254 = ~N1253;
  assign N1256 = ~N1255;
  assign N1258 = ~N1257;
  assign N1260 = ~N1259;
  assign N1262 = ~N1261;
  assign N1266 = ~N1265;
  assign N1270 = ~N1269;
  assign N1274 = ~N1273;
  assign N1278 = ~N1277;
  assign N1282 = ~N1281;
  assign N1284 = ~N1283;
  assign N1286 = ~N1285;
  assign N1288 = ~N1287;
  assign N1290 = ~N1289;
  assign N1292 = ~N1291;
  assign N1294 = ~N1293;
  assign N1296 = ~N1295;
  assign N1298 = ~N1297;
  assign N1300 = ~N1299;
  assign N1302 = ~N1301;
  assign N1304 = ~N1303;
  assign N1307 = ~N1306;
  assign N1309 = ~N1308;
  assign N1311 = ~N1310;
  assign N1313 = ~N1312;
  assign N1315 = ~N1314;
  assign N1317 = ~N1316;
  assign N1319 = ~N1318;
  assign N1321 = ~N1320;
  assign N1323 = ~N1322;
  assign N1325 = ~N1324;
  assign N1327 = ~N1326;
  assign N1329 = ~N1328;
  assign N1331 = ~N1330;
  assign N1333 = ~N1332;
  assign N1335 = ~N1334;
  assign N1337 = ~N1336;
  assign N1340 = ~N1339;
  assign N1342 = ~N1341;
  assign N1344 = ~N1343;
  assign N1346 = ~N1345;
  assign N1348 = ~N1347;
  assign N1350 = ~N1349;
  assign N1352 = ~N1351;
  assign N1354 = ~N1353;
  assign N1356 = ~N1355;
  assign N1358 = ~N1357;
  assign N1360 = ~N1359;
  assign N1362 = ~N1361;
  assign N1364 = ~N1363;
  assign N1366 = ~N1365;
  assign N1368 = ~N1367;
  assign N1370 = ~N1369;
  assign N1373 = ~N1372;
  assign N1375 = ~N1374;
  assign N1377 = ~N1376;
  assign N1379 = ~N1378;
  assign N1381 = ~N1380;
  assign N1383 = ~N1382;
  assign N1385 = ~N1384;
  assign N1387 = ~N1386;
  assign N1389 = ~N1388;
  assign N1391 = ~N1390;
  assign N1393 = ~N1392;
  assign N1395 = ~N1394;
  assign N1397 = ~N1396;
  assign N1399 = ~N1398;
  assign N1401 = ~N1400;
  assign N1403 = ~N1402;
  assign N1407 = ~N1406;
  assign N1411 = ~N1410;
  assign N1415 = ~N1414;
  assign N1419 = ~N1418;
  assign N1423 = ~N1422;
  assign N1425 = ~N1424;
  assign N1427 = ~N1426;
  assign N1429 = ~N1428;
  assign N1431 = ~N1430;
  assign N1433 = ~N1432;
  assign N1435 = ~N1434;
  assign N1437 = ~N1436;
  assign N1439 = ~N1438;
  assign N1441 = ~N1440;
  assign N1443 = ~N1442;
  assign N1445 = ~N1444;
  assign N1448 = ~N1447;
  assign N1450 = ~N1449;
  assign N1452 = ~N1451;
  assign N1454 = ~N1453;
  assign N1456 = ~N1455;
  assign N1458 = ~N1457;
  assign N1460 = ~N1459;
  assign N1462 = ~N1461;
  assign N1464 = ~N1463;
  assign N1466 = ~N1465;
  assign N1468 = ~N1467;
  assign N1470 = ~N1469;
  assign N1472 = ~N1471;
  assign N1474 = ~N1473;
  assign N1476 = ~N1475;
  assign N1478 = ~N1477;
  assign N1481 = ~N1480;
  assign N1483 = ~N1482;
  assign N1485 = ~N1484;
  assign N1487 = ~N1486;
  assign N1489 = ~N1488;
  assign N1491 = ~N1490;
  assign N1493 = ~N1492;
  assign N1495 = ~N1494;
  assign N1497 = ~N1496;
  assign N1499 = ~N1498;
  assign N1501 = ~N1500;
  assign N1503 = ~N1502;
  assign N1505 = ~N1504;
  assign N1507 = ~N1506;
  assign N1509 = ~N1508;
  assign N1511 = ~N1510;
  assign N1514 = ~N1513;
  assign N1516 = ~N1515;
  assign N1518 = ~N1517;
  assign N1520 = ~N1519;
  assign N1522 = ~N1521;
  assign N1524 = ~N1523;
  assign N1526 = ~N1525;
  assign N1528 = ~N1527;
  assign N1530 = ~N1529;
  assign N1532 = ~N1531;
  assign N1534 = ~N1533;
  assign N1536 = ~N1535;
  assign N1538 = ~N1537;
  assign N1540 = ~N1539;
  assign N1542 = ~N1541;
  assign N1544 = ~N1543;
  assign N1548 = ~N1547;
  assign N1550 = ~N1549;
  assign N1552 = ~N1551;
  assign N1554 = ~N1553;
  assign N1556 = ~N1555;
  assign N1558 = ~N1557;
  assign N1560 = ~N1559;
  assign N1563 = ~N1562;
  assign N1565 = ~N1564;
  assign N1567 = ~N1566;
  assign N1569 = ~N1568;
  assign N1571 = ~N1570;
  assign N1573 = ~N1572;
  assign N1575 = ~N1574;
  assign N1577 = ~N1576;
  assign N1579 = ~N1578;
  assign N1582 = ~N1581;
  assign N1584 = ~N1583;
  assign N1586 = ~N1585;
  assign N1589 = ~N1588;
  assign N1591 = ~N1590;
  assign N1593 = ~N1592;
  assign N1595 = ~N1594;
  assign N1597 = ~N1596;
  assign N1599 = ~N1598;
  assign N1601 = ~N1600;
  assign N1603 = ~N1602;
  assign N1605 = ~N1604;
  assign N1608 = ~N1607;
  assign N1610 = ~N1609;
  assign N1612 = ~N1611;
  assign N1614 = ~N1613;
  assign N1618 = ~N1617;
  assign N1621 = ~N1620;
  assign N1624 = ~N1623;
  assign N1626 = ~N1625;
  assign N1629 = ~N1628;
  assign N1631 = ~N1630;
  assign N1633 = ~N1632;
  assign N1637 = ~N1636;
  assign N1640 = ~N1639;
  assign N1643 = ~N1642;
  assign N1646 = ~N1645;
  assign N1649 = ~N1648;
  assign N1653 = ~N1652;
  assign N1656 = ~N1655;
  assign N1659 = ~N1658;
  assign N1662 = ~N1661;
  assign N1665 = ~N1664;
  assign N1668 = ~N1667;
  assign N1671 = ~N1670;
  assign N1677 = ~N1676;
  assign N1680 = ~N1679;
  assign N1683 = ~N1682;
  assign N1685 = ~N1684;
  assign N1687 = ~N1686;
  assign N1690 = ~N1689;
  assign N1693 = ~N1692;
  assign N1696 = ~N1695;
  assign N1698 = ~N1697;
  assign N1700 = ~N1699;
  assign N1702 = ~N1701;
  assign N1704 = ~N1703;
  assign N1720 = ~N1719;
  assign N1722 = ~N1721;
  assign N1724 = ~N1723;
  assign N1726 = ~N1725;
  assign N1728 = ~N1727;
  assign N1730 = ~N1729;
  assign N1732 = ~N1731;
  assign N1734 = ~N1733;
  assign N1736 = ~N1735;
  assign N1738 = ~N1737;
  assign N1740 = ~N1739;
  assign N1742 = ~N1741;
  assign N1744 = ~N1743;
  assign N1746 = ~N1745;
  assign N1748 = ~N1747;
  assign N1750 = ~N1749;
  assign N1752 = ~N1751;
  assign N1754 = ~N1753;
  assign N1756 = ~N1755;
  assign N1758 = ~N1757;
  assign N1760 = ~N1759;
  assign N1762 = ~N1761;
  assign N1764 = ~N1763;
  assign N1766 = ~N1765;
  assign N1768 = ~N1767;
  assign N1770 = ~N1769;
  assign N1772 = ~N1771;
  assign N1774 = ~N1773;
  assign N1776 = ~N1775;
  assign N1778 = ~N1777;
  assign N1781 = ~N1780;
  assign N1783 = ~N1782;
  assign N1785 = ~N1784;
  assign N1787 = ~N1786;
  assign N1789 = ~N1788;
  assign N1791 = ~N1790;
  assign N1793 = ~N1792;
  assign N1795 = ~N1794;
  assign N1798 = ~N1797;
  assign N1800 = ~N1799;
  assign N1802 = ~N1801;
  assign N1804 = ~N1803;
  assign N1806 = ~N1805;
  assign N1808 = ~N1807;
  assign N1810 = ~N1809;
  assign N1812 = ~N1811;
  assign N1814 = ~N1813;
  assign N1816 = ~N1815;
  assign N1818 = ~N1817;
  assign N1820 = ~N1819;
  assign N1822 = ~N1821;
  assign N1824 = ~N1823;
  assign N1826 = ~N1825;
  assign N1828 = ~N1827;
  assign N1830 = ~N1829;
  assign N1832 = ~N1831;
  assign N1834 = ~N1833;
  assign N1836 = ~N1835;
  assign N1838 = ~N1837;
  assign N1840 = ~N1839;
  assign N1842 = ~N1841;
  assign N1844 = ~N1843;
  assign N1847 = ~N1846;
  assign N1849 = ~N1848;
  assign N1851 = ~N1850;
  assign N1853 = ~N1852;
  assign N1855 = ~N1854;
  assign N1857 = ~N1856;
  assign N1859 = ~N1858;
  assign N1861 = ~N1860;
  assign N1864 = ~N1863;
  assign N1866 = ~N1865;
  assign N1868 = ~N1867;
  assign N1870 = ~N1869;
  assign N1872 = ~N1871;
  assign N1874 = ~N1873;
  assign N1876 = ~N1875;
  assign N1878 = ~N1877;
  assign N1880 = ~N1879;
  assign N1882 = ~N1881;
  assign N1884 = ~N1883;
  assign N1886 = ~N1885;
  assign N1888 = ~N1887;
  assign N1890 = ~N1889;
  assign N1892 = ~N1891;
  assign N1894 = ~N1893;
  assign N1896 = ~N1895;
  assign N1898 = ~N1897;
  assign N1900 = ~N1899;
  assign N1902 = ~N1901;
  assign N1904 = ~N1903;
  assign N1906 = ~N1905;
  assign N1908 = ~N1907;
  assign N1910 = ~N1909;
  assign N1913 = ~N1912;
  assign N1915 = ~N1914;
  assign N1917 = ~N1916;
  assign N1919 = ~N1918;
  assign N1921 = ~N1920;
  assign N1923 = ~N1922;
  assign N1925 = ~N1924;
  assign N1927 = ~N1926;
  assign N1930 = ~N1929;
  assign N1932 = ~N1931;
  assign N1934 = ~N1933;
  assign N1936 = ~N1935;
  assign N1938 = ~N1937;
  assign N1940 = ~N1939;
  assign N1942 = ~N1941;
  assign N1944 = ~N1943;
  assign N1946 = ~N1945;
  assign N1948 = ~N1947;
  assign N1950 = ~N1949;
  assign N1952 = ~N1951;
  assign N1954 = ~N1953;
  assign N1956 = ~N1955;
  assign N1958 = ~N1957;
  assign N1960 = ~N1959;
  assign N1962 = ~N1961;
  assign N1964 = ~N1963;
  assign N1966 = ~N1965;
  assign N1968 = ~N1967;
  assign N1970 = ~N1969;
  assign N1972 = ~N1971;
  assign N1974 = ~N1973;
  assign N1976 = ~N1975;
  assign N1979 = ~N1978;
  assign N1981 = ~N1980;
  assign N1983 = ~N1982;
  assign N1985 = ~N1984;
  assign N1987 = ~N1986;
  assign N1989 = ~N1988;
  assign N1991 = ~N1990;
  assign N1993 = ~N1992;
  assign N1996 = ~N1995;
  assign N1998 = ~N1997;
  assign N2000 = ~N1999;
  assign N2002 = ~N2001;
  assign N2004 = ~N2003;
  assign N2006 = ~N2005;
  assign N2008 = ~N2007;
  assign N2010 = ~N2009;
  assign N2012 = ~N2011;
  assign N2014 = ~N2013;
  assign N2016 = ~N2015;
  assign N2018 = ~N2017;
  assign N2020 = ~N2019;
  assign N2022 = ~N2021;
  assign N2024 = ~N2023;
  assign N2026 = ~N2025;
  assign N2028 = ~N2027;
  assign N2030 = ~N2029;
  assign N2032 = ~N2031;
  assign N2034 = ~N2033;
  assign N2036 = ~N2035;
  assign N2038 = ~N2037;
  assign N2040 = ~N2039;
  assign N2042 = ~N2041;
  assign N2045 = ~N2044;
  assign N2047 = ~N2046;
  assign N2049 = ~N2048;
  assign N2051 = ~N2050;
  assign N2053 = ~N2052;
  assign N2055 = ~N2054;
  assign N2057 = ~N2056;
  assign N2059 = ~N2058;
  assign N2062 = ~N2061;
  assign N2064 = ~N2063;
  assign N2066 = ~N2065;
  assign N2068 = ~N2067;
  assign N2070 = ~N2069;
  assign N2072 = ~N2071;
  assign N2075 = ~N2074;
  assign N2077 = ~N2076;
  assign N2079 = ~N2078;
  assign N2082 = ~N2081;
  assign N2084 = ~N2083;
  assign N2086 = ~N2085;
  assign N2088 = ~N2087;
  assign N2090 = ~N2089;
  assign N2092 = ~N2091;
  assign N2094 = ~N2093;
  assign N2096 = ~N2095;
  assign N2098 = ~N2097;
  assign N2100 = ~N2099;
  assign N2102 = ~N2101;
  assign N2104 = ~N2103;
  assign N2106 = ~N2105;
  assign N2108 = ~N2107;
  assign N2110 = ~N2109;
  assign N2113 = ~N2112;
  assign N2115 = ~N2114;
  assign N2117 = ~N2116;
  assign N2119 = ~N2118;
  assign N2121 = ~N2120;
  assign N2123 = ~N2122;
  assign N2125 = ~N2124;
  assign N2127 = ~N2126;
  assign N2130 = ~N2129;
  assign N2132 = ~N2131;
  assign N2134 = ~N2133;
  assign N2136 = ~N2135;
  assign N2138 = ~N2137;
  assign N2140 = ~N2139;
  assign N2142 = ~N2141;
  assign N2144 = ~N2143;
  assign N2146 = ~N2145;
  assign N2149 = ~N2148;
  assign N2151 = ~N2150;
  assign N2153 = ~N2152;
  assign N2155 = ~N2154;
  assign N2157 = ~N2156;
  assign N2159 = ~N2158;
  assign N2161 = ~N2160;
  assign N2163 = ~N2162;
  assign N2165 = ~N2164;
  assign N2167 = ~N2166;
  assign N2169 = ~N2168;
  assign N2171 = ~N2170;
  assign N2173 = ~N2172;
  assign N2175 = ~N2174;
  assign N2177 = ~N2176;
  assign N2181 = ~N2180;
  assign N2183 = ~N2182;
  assign N2185 = ~N2184;
  assign N2187 = ~N2186;
  assign N2189 = ~N2188;
  assign N2191 = ~N2190;
  assign N2193 = ~N2192;
  assign N2195 = ~N2194;
  assign N2198 = ~N2197;
  assign N2200 = ~N2199;
  assign N2202 = ~N2201;
  assign N2204 = ~N2203;
  assign N2206 = ~N2205;
  assign N2208 = ~N2207;
  assign N2210 = ~N2209;
  assign N2212 = ~N2211;
  assign N2214 = ~N2213;
  assign N2216 = ~N2215;
  assign N2218 = ~N2217;
  assign N2220 = ~N2219;
  assign N2222 = ~N2221;
  assign N2224 = ~N2223;
  assign N2226 = ~N2225;
  assign N2228 = ~N2227;
  assign N2231 = ~N2230;
  assign N2233 = ~N2232;
  assign N2235 = ~N2234;
  assign N2237 = ~N2236;
  assign N2239 = ~N2238;
  assign N2241 = ~N2240;
  assign N2243 = ~N2242;
  assign N2245 = ~N2244;
  assign N2256 = ~N2255;
  assign N2260 = ~N2259;
  assign N2263 = ~N2262;
  assign N2266 = ~N2265;
  assign N2269 = ~N2268;
  assign N2272 = ~N2271;
  assign N2275 = ~N2274;
  assign N2278 = ~N2277;
  assign N2281 = ~N2280;
  assign N2284 = ~N2283;
  assign N2287 = ~N2286;
  assign N2291 = ~N2290;
  assign N2294 = ~N2293;
  assign N2297 = ~N2296;
  assign N2300 = ~N2299;
  assign N2302 = ~N2301;
  assign N2304 = ~N2303;
  assign N2306 = ~N2305;
  assign N2308 = ~N2307;
  assign N2311 = ~N2310;
  assign N2313 = ~N2312;
  assign N2315 = ~N2314;
  assign N2317 = ~N2316;
  assign N2319 = ~N2318;
  assign N2321 = ~N2320;
  assign N2323 = ~N2322;
  assign N2325 = ~N2324;
  assign N2328 = ~N2327;
  assign N2330 = ~N2329;
  assign N2332 = ~N2331;
  assign N2334 = ~N2333;
  assign N2336 = ~N2335;
  assign N2338 = ~N2337;
  assign N2340 = ~N2339;
  assign N2342 = ~N2341;
  assign N2345 = ~N2344;
  assign N2347 = ~N2346;
  assign N2349 = ~N2348;
  assign N2351 = ~N2350;
  assign N2353 = ~N2352;
  assign N2355 = ~N2354;
  assign N2357 = ~N2356;
  assign N2359 = ~N2358;
  assign N2361 = ~N2360;
  assign N2363 = ~N2362;
  assign N2365 = ~N2364;
  assign N2367 = ~N2366;
  assign N2369 = ~N2368;
  assign N2371 = ~N2370;
  assign N2373 = ~N2372;
  assign N2375 = ~N2374;
  assign N2379 = ~N2378;
  assign N2381 = ~N2380;
  assign N2383 = ~N2382;
  assign N2385 = ~N2384;
  assign N2387 = ~N2386;
  assign N2389 = ~N2388;
  assign N2391 = ~N2390;
  assign N2393 = ~N2392;
  assign N2395 = ~N2394;
  assign N2397 = ~N2396;
  assign N2399 = ~N2398;
  assign N2401 = ~N2400;
  assign N2404 = ~N2403;
  assign N2406 = ~N2405;
  assign N2408 = ~N2407;
  assign N2410 = ~N2409;
  assign N2412 = ~N2411;
  assign N2414 = ~N2413;
  assign N2416 = ~N2415;
  assign N2418 = ~N2417;
  assign N2420 = ~N2419;
  assign N2422 = ~N2421;
  assign N2424 = ~N2423;
  assign N2426 = ~N2425;
  assign N2429 = ~N2428;
  assign N2431 = ~N2430;
  assign N2433 = ~N2432;
  assign N2435 = ~N2434;
  assign N2437 = ~N2436;
  assign N2439 = ~N2438;
  assign N2441 = ~N2440;
  assign N2443 = ~N2442;
  assign N2446 = ~N2445;
  assign N2448 = ~N2447;
  assign N2450 = ~N2449;
  assign N2452 = ~N2451;
  assign N2454 = ~N2453;
  assign N2456 = ~N2455;
  assign N2458 = ~N2457;
  assign N2460 = ~N2459;
  assign N2462 = ~N2461;
  assign N2464 = ~N2463;
  assign N2466 = ~N2465;
  assign N2468 = ~N2467;
  assign N2470 = ~N2469;
  assign N2472 = ~N2471;
  assign N2474 = ~N2473;
  assign N2476 = ~N2475;
  assign N2479 = ~N2478;
  assign N2481 = ~N2480;
  assign N2483 = ~N2482;
  assign N2485 = ~N2484;
  assign N2487 = ~N2486;
  assign N2489 = ~N2488;
  assign N2491 = ~N2490;
  assign N2493 = ~N2492;
  assign N2495 = ~N2494;
  assign N2497 = ~N2496;
  assign N2499 = ~N2498;
  assign N2501 = ~N2500;
  assign N2503 = ~N2502;
  assign N2506 = ~N2505;
  assign N2509 = ~N2508;
  assign N2512 = ~N2511;
  assign N2516 = ~N2515;
  assign N2519 = ~N2518;
  assign N2522 = ~N2521;
  assign N2525 = ~N2524;
  assign N2528 = ~N2527;
  assign N2531 = ~N2530;
  assign N2534 = ~N2533;
  assign N2536 = ~N2535;
  assign N2542 = ~N2541;
  assign N2544 = ~N2543;
  assign N2546 = ~N2545;
  assign N2549 = ~N2548;
  assign N2553 = ~N2552;
  assign N2555 = ~N2554;
  assign N2558 = ~N2557;
  assign N2560 = ~N2559;
  assign N2562 = ~N2561;
  assign N2564 = ~N2563;
  assign N2566 = ~N2565;
  assign N2568 = ~N2567;
  assign N2571 = ~N2570;
  assign N2573 = ~N2572;
  assign N2575 = ~N2574;
  assign N2577 = ~N2576;
  assign N2579 = ~N2578;
  assign N2581 = ~N2580;
  assign N2583 = ~N2582;
  assign N2585 = ~N2584;
  assign N2587 = ~N2586;
  assign N2589 = ~N2588;
  assign N2591 = ~N2590;
  assign N2593 = ~N2592;
  assign N2596 = ~N2595;
  assign N2598 = ~N2597;
  assign N2600 = ~N2599;
  assign N2602 = ~N2601;
  assign N2604 = ~N2603;
  assign N2606 = ~N2605;
  assign N2608 = ~N2607;
  assign N2610 = ~N2609;
  assign N2612 = ~N2611;
  assign N2614 = ~N2613;
  assign N2616 = ~N2615;
  assign N2618 = ~N2617;
  assign N2620 = ~N2619;
  assign N2622 = ~N2621;
  assign N2624 = ~N2623;
  assign N2626 = ~N2625;
  assign N2629 = ~N2628;
  assign N2631 = ~N2630;
  assign N2633 = ~N2632;
  assign N2635 = ~N2634;
  assign N2637 = ~N2636;
  assign N2639 = ~N2638;
  assign N2641 = ~N2640;
  assign N2643 = ~N2642;
  assign N2645 = ~N2644;
  assign N2647 = ~N2646;
  assign N2649 = ~N2648;
  assign N2651 = ~N2650;
  assign N2653 = ~N2652;
  assign N2655 = ~N2654;
  assign N2657 = ~N2656;
  assign N2659 = ~N2658;
  assign N2662 = ~N2661;
  assign N2664 = ~N2663;
  assign N2666 = ~N2665;
  assign N2668 = ~N2667;
  assign N2670 = ~N2669;
  assign N2672 = ~N2671;
  assign N2674 = ~N2673;
  assign N2676 = ~N2675;
  assign N2679 = ~N2678;
  assign N2681 = ~N2680;
  assign N2683 = ~N2682;
  assign N2685 = ~N2684;
  assign N2689 = ~N2688;
  assign N2691 = ~N2690;
  assign N2693 = ~N2692;
  assign N2695 = ~N2694;
  assign N2697 = ~N2696;
  assign N2699 = ~N2698;
  assign N2701 = ~N2700;
  assign N2703 = ~N2702;
  assign N2705 = ~N2704;
  assign N2707 = ~N2706;
  assign N2709 = ~N2708;
  assign N2711 = ~N2710;
  assign N2713 = ~N2712;
  assign N2715 = ~N2714;
  assign N2717 = ~N2716;
  assign N2719 = ~N2718;
  assign N2721 = ~N2720;
  assign N2723 = ~N2722;
  assign N2725 = ~N2724;
  assign N2727 = ~N2726;
  assign N2730 = ~N2729;
  assign N2732 = ~N2731;
  assign N2734 = ~N2733;
  assign N2736 = ~N2735;
  assign N2738 = ~N2737;
  assign N2740 = ~N2739;
  assign N2742 = ~N2741;
  assign N2744 = ~N2743;
  assign N2746 = ~N2745;
  assign N2748 = ~N2747;
  assign N2750 = ~N2749;
  assign N2752 = ~N2751;
  assign N2754 = ~N2753;
  assign N2756 = ~N2755;
  assign N2758 = ~N2757;
  assign N2760 = ~N2759;
  assign N2763 = ~N2762;
  assign N2765 = ~N2764;
  assign N2767 = ~N2766;
  assign N2769 = ~N2768;
  assign N2771 = ~N2770;
  assign N2773 = ~N2772;
  assign N2775 = ~N2774;
  assign N2777 = ~N2776;
  assign N2779 = ~N2778;
  assign N2781 = ~N2780;
  assign N2783 = ~N2782;
  assign N2785 = ~N2784;
  assign N2787 = ~N2786;
  assign N2789 = ~N2788;
  assign N2791 = ~N2790;
  assign N2793 = ~N2792;
  assign N2796 = ~N2795;
  assign N2798 = ~N2797;
  assign N2800 = ~N2799;
  assign N2802 = ~N2801;
  assign N2804 = ~N2803;
  assign N2806 = ~N2805;
  assign N2808 = ~N2807;
  assign N2812 = ~N2811;
  assign N2814 = ~N2813;
  assign N2817 = ~N2816;
  assign N2820 = ~N2819;
  assign N2829 = ~N2828;
  assign N2831 = ~N2830;
  assign N2833 = ~N2832;
  assign N2835 = ~N2834;
  assign N2837 = ~N2836;
  assign N2839 = ~N2838;
  assign N2841 = ~N2840;
  assign N2843 = ~N2842;
  assign N2845 = ~N2844;
  assign N2847 = ~N2846;
  assign N2849 = ~N2848;
  assign N2851 = ~N2850;
  assign N2853 = ~N2852;
  assign N2855 = ~N2854;
  assign N2857 = ~N2856;
  assign N2859 = ~N2858;
  assign N2861 = ~N2860;
  assign N2863 = ~N2862;
  assign N2866 = ~N2865;
  assign N2868 = ~N2867;
  assign N2870 = ~N2869;
  assign N2872 = ~N2871;
  assign N2874 = ~N2873;
  assign N2876 = ~N2875;
  assign N2878 = ~N2877;
  assign N2880 = ~N2879;
  assign N2882 = ~N2881;
  assign N2884 = ~N2883;
  assign N2886 = ~N2885;
  assign N2888 = ~N2887;
  assign N2890 = ~N2889;
  assign N2892 = ~N2891;
  assign N2894 = ~N2893;
  assign N2896 = ~N2895;
  assign N2899 = ~N2898;
  assign N2901 = ~N2900;
  assign N2903 = ~N2902;
  assign N2905 = ~N2904;
  assign N2907 = ~N2906;
  assign N2909 = ~N2908;
  assign N2911 = ~N2910;
  assign N2913 = ~N2912;
  assign N2915 = ~N2914;
  assign N2917 = ~N2916;
  assign N2919 = ~N2918;
  assign N2921 = ~N2920;
  assign N2923 = ~N2922;
  assign N2925 = ~N2924;
  assign N2927 = ~N2926;
  assign N2929 = ~N2928;
  assign N2932 = ~N2931;
  assign N2934 = ~N2933;
  assign N2936 = ~N2935;
  assign N2938 = ~N2937;
  assign N2940 = ~N2939;
  assign N2943 = ~N2942;
  assign N2946 = ~N2945;
  assign N2949 = ~N2948;
  assign N2955 = ~N2954;
  assign N2957 = ~N2956;
  assign N2959 = ~N2958;
  assign N2962 = ~N2961;
  assign N2965 = ~N2964;
  assign N2968 = ~N2967;
  assign N2971 = ~N2970;
  assign N2974 = ~N2973;
  assign N2978 = ~N2977;
  assign N2981 = ~N2980;
  assign N2984 = ~N2983;
  assign N2987 = ~N2986;
  assign N2991 = ~N2990;
  assign N2994 = ~N2993;
  assign N2996 = ~N2995;
  assign N2998 = ~N2997;
  assign N3000 = ~N2999;
  assign N3002 = ~N3001;
  assign N3004 = ~N3003;
  assign N3006 = ~N3005;
  assign N3008 = ~N3007;
  assign N3010 = ~N3009;
  assign N3012 = ~N3011;
  assign N3014 = ~N3013;
  assign N3018 = ~N3017;
  assign N3020 = ~N3019;
  assign N3022 = ~N3021;
  assign N3024 = ~N3023;
  assign N3026 = ~N3025;
  assign N3028 = ~N3027;
  assign N3030 = ~N3029;
  assign N3032 = ~N3031;
  assign N3036 = ~N3035;
  assign N3038 = ~N3037;
  assign N3040 = ~N3039;
  assign N3042 = ~N3041;
  assign N3044 = ~N3043;
  assign N3046 = ~N3045;
  assign N3048 = ~N3047;
  assign N3050 = ~N3049;
  assign N3054 = ~N3053;
  assign N3056 = ~N3055;
  assign N3058 = ~N3057;
  assign N3060 = ~N3059;
  assign N3062 = ~N3061;
  assign N3064 = ~N3063;
  assign N3066 = ~N3065;
  assign N3068 = ~N3067;
  assign N3070 = ~N3069;
  assign N3072 = ~N3071;
  assign N3074 = ~N3073;
  assign N3076 = ~N3075;
  assign N3078 = ~N3077;
  assign N3080 = ~N3079;
  assign N3082 = ~N3081;
  assign N3084 = ~N3083;
  assign N3087 = ~N3086;
  assign N3089 = ~N3088;
  assign N3091 = ~N3090;
  assign N3093 = ~N3092;
  assign N3095 = ~N3094;
  assign N3097 = ~N3096;
  assign N3099 = ~N3098;
  assign N3101 = ~N3100;
  assign N3103 = ~N3102;
  assign N3105 = ~N3104;
  assign N3107 = ~N3106;
  assign N3109 = ~N3108;
  assign N3112 = ~N3111;
  assign N3114 = ~N3113;
  assign N3116 = ~N3115;
  assign N3118 = ~N3117;
  assign N3120 = ~N3119;
  assign N3122 = ~N3121;
  assign N3124 = ~N3123;
  assign N3126 = ~N3125;
  assign N3128 = ~N3127;
  assign N3130 = ~N3129;
  assign N3132 = ~N3131;
  assign N3134 = ~N3133;
  assign N3136 = ~N3135;
  assign N3138 = ~N3137;
  assign N3140 = ~N3139;
  assign N3142 = ~N3141;
  assign N3144 = ~N3143;
  assign N3146 = ~N3145;
  assign N3148 = ~N3147;
  assign N3150 = ~N3149;
  assign N3153 = ~N3152;
  assign N3155 = ~N3154;
  assign N3157 = ~N3156;
  assign N3159 = ~N3158;
  assign N3161 = ~N3160;
  assign N3163 = ~N3162;
  assign N3165 = ~N3164;
  assign N3167 = ~N3166;
  assign N3171 = ~N3170;
  assign N3173 = ~N3172;
  assign N3175 = ~N3174;
  assign N3177 = ~N3176;
  assign N3179 = ~N3178;
  assign N3181 = ~N3180;
  assign N3183 = ~N3182;
  assign N3185 = ~N3184;
  assign N3188 = ~N3187;
  assign N3190 = ~N3189;
  assign N3192 = ~N3191;
  assign N3194 = ~N3193;
  assign N3196 = ~N3195;
  assign N3198 = ~N3197;
  assign N3200 = ~N3199;
  assign N3202 = ~N3201;
  assign N3204 = ~N3203;
  assign N3206 = ~N3205;
  assign N3208 = ~N3207;
  assign N3210 = ~N3209;
  assign N3212 = ~N3211;
  assign N3214 = ~N3213;
  assign N3216 = ~N3215;
  assign N3218 = ~N3217;
  assign N3221 = ~N3220;
  assign N3223 = ~N3222;
  assign N3225 = ~N3224;
  assign N3227 = ~N3226;
  assign N3229 = ~N3228;
  assign N3231 = ~N3230;
  assign N3233 = ~N3232;
  assign N3235 = ~N3234;
  assign N3237 = ~N3236;
  assign N3239 = ~N3238;
  assign N3241 = ~N3240;
  assign N3243 = ~N3242;
  assign N3247 = ~N3246;
  assign N3249 = ~N3248;
  assign N3251 = ~N3250;
  assign N3253 = ~N3252;
  assign N3255 = ~N3254;
  assign N3257 = ~N3256;
  assign N3259 = ~N3258;
  assign N3261 = ~N3260;
  assign N3263 = ~N3262;
  assign N3265 = ~N3264;
  assign N3267 = ~N3266;
  assign N3269 = ~N3268;
  assign N3271 = ~N3270;
  assign N3273 = ~N3272;
  assign N3275 = ~N3274;
  assign N3277 = ~N3276;
  assign N3279 = ~N3278;
  assign N3281 = ~N3280;
  assign N3283 = ~N3282;
  assign N3285 = ~N3284;
  assign N3288 = ~N3287;
  assign N3290 = ~N3289;
  assign N3292 = ~N3291;
  assign N3294 = ~N3293;
  assign N3296 = ~N3295;
  assign N3298 = ~N3297;
  assign N3300 = ~N3299;
  assign N3302 = ~N3301;
  assign N3304 = ~N3303;
  assign N3306 = ~N3305;
  assign N3308 = ~N3307;
  assign N3310 = ~N3309;
  assign N3312 = ~N3311;
  assign N3314 = ~N3313;
  assign N3316 = ~N3315;
  assign N3318 = ~N3317;
  assign N3321 = ~N3320;
  assign N3323 = ~N3322;
  assign N3325 = ~N3324;
  assign N3327 = ~N3326;
  assign N3329 = ~N3328;
  assign N3331 = ~N3330;
  assign N3333 = ~N3332;
  assign N3335 = ~N3334;
  assign N3337 = ~N3336;
  assign N3339 = ~N3338;
  assign N3341 = ~N3340;
  assign N3343 = ~N3342;
  assign N3345 = ~N3344;
  assign N3347 = ~N3346;
  assign N3349 = ~N3348;
  assign N3351 = ~N3350;
  assign N3354 = ~N3353;
  assign N3356 = ~N3355;
  assign N3358 = ~N3357;
  assign N3360 = ~N3359;
  assign N3362 = ~N3361;
  assign N3364 = ~N3363;
  assign N3368 = ~N3367;
  assign N3372 = ~N3371;
  assign N3374 = ~N3373;
  assign N3378 = ~N3377;
  assign N3381 = ~N3380;

endmodule

