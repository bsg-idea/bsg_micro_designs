

module top
(
  clk,
  reset,
  calibration_done_i,
  valid_i,
  data_i,
  ready_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [1279:0] data_i;
  input [3:0] in_top_channel_i;
  input [3:0] out_top_channel_i;
  output [9:0] valid_o;
  output [1279:0] data_o;
  input [9:0] ready_i;
  input clk;
  input reset;
  input calibration_done_i;
  input valid_i;
  output ready_o;

  bsg_assembler_out
  wrapper
  (
    .data_i(data_i),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .ready_i(ready_i),
    .clk(clk),
    .reset(reset),
    .calibration_done_i(calibration_done_i),
    .valid_i(valid_i),
    .ready_o(ready_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p128_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [127:0] w_data_i;
  input [0:0] r_addr_i;
  output [127:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [127:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10;
  reg [255:0] mem;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[255] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[254] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[253] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[252] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[251] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[250] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[249] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[248] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[247] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[246] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[245] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[244] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[243] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[242] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[241] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[240] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[239] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[238] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[237] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[236] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[235] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[234] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[233] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[232] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[231] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[230] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[229] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[228] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[227] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[226] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[225] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[224] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[223] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[222] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[221] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[220] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[219] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[218] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[217] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[216] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[215] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[214] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[213] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[212] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[211] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[210] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[209] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[208] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[207] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[206] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[205] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[204] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[203] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[202] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[201] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[200] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[199] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[198] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[197] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[196] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[195] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[194] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[193] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[192] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[191] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[190] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[189] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[188] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[187] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[186] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[185] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[184] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[183] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[182] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[181] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[180] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[179] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[178] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[177] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[176] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[175] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[174] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[173] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[172] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[171] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[170] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[169] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[168] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[167] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[166] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[165] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[164] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[163] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[162] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[161] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[160] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[159] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[158] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[157] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[156] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[155] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[154] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[153] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[152] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[151] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[150] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[149] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[148] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[147] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[146] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[145] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[144] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[143] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[142] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[141] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[140] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[139] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[138] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[137] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[136] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[135] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[134] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[133] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[132] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[131] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[130] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[129] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[128] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], N5, N5 } : 
                               (N2)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N9) begin
      { mem[255:157], mem[128:128] } <= { w_data_i[127:29], w_data_i[0:0] };
    end 
    if(N10) begin
      { mem[156:129] } <= { w_data_i[28:1] };
    end 
    if(N7) begin
      { mem[127:29], mem[0:0] } <= { w_data_i[127:29], w_data_i[0:0] };
    end 
    if(N8) begin
      { mem[28:1] } <= { w_data_i[28:1] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p128_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [127:0] w_data_i;
  input [0:0] r_addr_i;
  output [127:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [127:0] r_data_o;

  bsg_mem_1r1w_synth_width_p128_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p128_ready_THEN_valid_p1
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [127:0] data_o;
  wire ready_o,v_o,N0,N1,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p128_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(v_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = v_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N16 | N19;
  assign N16 = empty_r & N15;
  assign N15 = ~v_i;
  assign N19 = N18 & N15;
  assign N18 = N17 & yumi_i;
  assign N17 = ~full_r;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & v_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_make_2D_array_width_p128_items_p10
(
  i,
  o
);

  input [1279:0] i;
  output [1279:0] o;
  wire [1279:0] o;
  assign o[1279] = i[1279];
  assign o[1278] = i[1278];
  assign o[1277] = i[1277];
  assign o[1276] = i[1276];
  assign o[1275] = i[1275];
  assign o[1274] = i[1274];
  assign o[1273] = i[1273];
  assign o[1272] = i[1272];
  assign o[1271] = i[1271];
  assign o[1270] = i[1270];
  assign o[1269] = i[1269];
  assign o[1268] = i[1268];
  assign o[1267] = i[1267];
  assign o[1266] = i[1266];
  assign o[1265] = i[1265];
  assign o[1264] = i[1264];
  assign o[1263] = i[1263];
  assign o[1262] = i[1262];
  assign o[1261] = i[1261];
  assign o[1260] = i[1260];
  assign o[1259] = i[1259];
  assign o[1258] = i[1258];
  assign o[1257] = i[1257];
  assign o[1256] = i[1256];
  assign o[1255] = i[1255];
  assign o[1254] = i[1254];
  assign o[1253] = i[1253];
  assign o[1252] = i[1252];
  assign o[1251] = i[1251];
  assign o[1250] = i[1250];
  assign o[1249] = i[1249];
  assign o[1248] = i[1248];
  assign o[1247] = i[1247];
  assign o[1246] = i[1246];
  assign o[1245] = i[1245];
  assign o[1244] = i[1244];
  assign o[1243] = i[1243];
  assign o[1242] = i[1242];
  assign o[1241] = i[1241];
  assign o[1240] = i[1240];
  assign o[1239] = i[1239];
  assign o[1238] = i[1238];
  assign o[1237] = i[1237];
  assign o[1236] = i[1236];
  assign o[1235] = i[1235];
  assign o[1234] = i[1234];
  assign o[1233] = i[1233];
  assign o[1232] = i[1232];
  assign o[1231] = i[1231];
  assign o[1230] = i[1230];
  assign o[1229] = i[1229];
  assign o[1228] = i[1228];
  assign o[1227] = i[1227];
  assign o[1226] = i[1226];
  assign o[1225] = i[1225];
  assign o[1224] = i[1224];
  assign o[1223] = i[1223];
  assign o[1222] = i[1222];
  assign o[1221] = i[1221];
  assign o[1220] = i[1220];
  assign o[1219] = i[1219];
  assign o[1218] = i[1218];
  assign o[1217] = i[1217];
  assign o[1216] = i[1216];
  assign o[1215] = i[1215];
  assign o[1214] = i[1214];
  assign o[1213] = i[1213];
  assign o[1212] = i[1212];
  assign o[1211] = i[1211];
  assign o[1210] = i[1210];
  assign o[1209] = i[1209];
  assign o[1208] = i[1208];
  assign o[1207] = i[1207];
  assign o[1206] = i[1206];
  assign o[1205] = i[1205];
  assign o[1204] = i[1204];
  assign o[1203] = i[1203];
  assign o[1202] = i[1202];
  assign o[1201] = i[1201];
  assign o[1200] = i[1200];
  assign o[1199] = i[1199];
  assign o[1198] = i[1198];
  assign o[1197] = i[1197];
  assign o[1196] = i[1196];
  assign o[1195] = i[1195];
  assign o[1194] = i[1194];
  assign o[1193] = i[1193];
  assign o[1192] = i[1192];
  assign o[1191] = i[1191];
  assign o[1190] = i[1190];
  assign o[1189] = i[1189];
  assign o[1188] = i[1188];
  assign o[1187] = i[1187];
  assign o[1186] = i[1186];
  assign o[1185] = i[1185];
  assign o[1184] = i[1184];
  assign o[1183] = i[1183];
  assign o[1182] = i[1182];
  assign o[1181] = i[1181];
  assign o[1180] = i[1180];
  assign o[1179] = i[1179];
  assign o[1178] = i[1178];
  assign o[1177] = i[1177];
  assign o[1176] = i[1176];
  assign o[1175] = i[1175];
  assign o[1174] = i[1174];
  assign o[1173] = i[1173];
  assign o[1172] = i[1172];
  assign o[1171] = i[1171];
  assign o[1170] = i[1170];
  assign o[1169] = i[1169];
  assign o[1168] = i[1168];
  assign o[1167] = i[1167];
  assign o[1166] = i[1166];
  assign o[1165] = i[1165];
  assign o[1164] = i[1164];
  assign o[1163] = i[1163];
  assign o[1162] = i[1162];
  assign o[1161] = i[1161];
  assign o[1160] = i[1160];
  assign o[1159] = i[1159];
  assign o[1158] = i[1158];
  assign o[1157] = i[1157];
  assign o[1156] = i[1156];
  assign o[1155] = i[1155];
  assign o[1154] = i[1154];
  assign o[1153] = i[1153];
  assign o[1152] = i[1152];
  assign o[1151] = i[1151];
  assign o[1150] = i[1150];
  assign o[1149] = i[1149];
  assign o[1148] = i[1148];
  assign o[1147] = i[1147];
  assign o[1146] = i[1146];
  assign o[1145] = i[1145];
  assign o[1144] = i[1144];
  assign o[1143] = i[1143];
  assign o[1142] = i[1142];
  assign o[1141] = i[1141];
  assign o[1140] = i[1140];
  assign o[1139] = i[1139];
  assign o[1138] = i[1138];
  assign o[1137] = i[1137];
  assign o[1136] = i[1136];
  assign o[1135] = i[1135];
  assign o[1134] = i[1134];
  assign o[1133] = i[1133];
  assign o[1132] = i[1132];
  assign o[1131] = i[1131];
  assign o[1130] = i[1130];
  assign o[1129] = i[1129];
  assign o[1128] = i[1128];
  assign o[1127] = i[1127];
  assign o[1126] = i[1126];
  assign o[1125] = i[1125];
  assign o[1124] = i[1124];
  assign o[1123] = i[1123];
  assign o[1122] = i[1122];
  assign o[1121] = i[1121];
  assign o[1120] = i[1120];
  assign o[1119] = i[1119];
  assign o[1118] = i[1118];
  assign o[1117] = i[1117];
  assign o[1116] = i[1116];
  assign o[1115] = i[1115];
  assign o[1114] = i[1114];
  assign o[1113] = i[1113];
  assign o[1112] = i[1112];
  assign o[1111] = i[1111];
  assign o[1110] = i[1110];
  assign o[1109] = i[1109];
  assign o[1108] = i[1108];
  assign o[1107] = i[1107];
  assign o[1106] = i[1106];
  assign o[1105] = i[1105];
  assign o[1104] = i[1104];
  assign o[1103] = i[1103];
  assign o[1102] = i[1102];
  assign o[1101] = i[1101];
  assign o[1100] = i[1100];
  assign o[1099] = i[1099];
  assign o[1098] = i[1098];
  assign o[1097] = i[1097];
  assign o[1096] = i[1096];
  assign o[1095] = i[1095];
  assign o[1094] = i[1094];
  assign o[1093] = i[1093];
  assign o[1092] = i[1092];
  assign o[1091] = i[1091];
  assign o[1090] = i[1090];
  assign o[1089] = i[1089];
  assign o[1088] = i[1088];
  assign o[1087] = i[1087];
  assign o[1086] = i[1086];
  assign o[1085] = i[1085];
  assign o[1084] = i[1084];
  assign o[1083] = i[1083];
  assign o[1082] = i[1082];
  assign o[1081] = i[1081];
  assign o[1080] = i[1080];
  assign o[1079] = i[1079];
  assign o[1078] = i[1078];
  assign o[1077] = i[1077];
  assign o[1076] = i[1076];
  assign o[1075] = i[1075];
  assign o[1074] = i[1074];
  assign o[1073] = i[1073];
  assign o[1072] = i[1072];
  assign o[1071] = i[1071];
  assign o[1070] = i[1070];
  assign o[1069] = i[1069];
  assign o[1068] = i[1068];
  assign o[1067] = i[1067];
  assign o[1066] = i[1066];
  assign o[1065] = i[1065];
  assign o[1064] = i[1064];
  assign o[1063] = i[1063];
  assign o[1062] = i[1062];
  assign o[1061] = i[1061];
  assign o[1060] = i[1060];
  assign o[1059] = i[1059];
  assign o[1058] = i[1058];
  assign o[1057] = i[1057];
  assign o[1056] = i[1056];
  assign o[1055] = i[1055];
  assign o[1054] = i[1054];
  assign o[1053] = i[1053];
  assign o[1052] = i[1052];
  assign o[1051] = i[1051];
  assign o[1050] = i[1050];
  assign o[1049] = i[1049];
  assign o[1048] = i[1048];
  assign o[1047] = i[1047];
  assign o[1046] = i[1046];
  assign o[1045] = i[1045];
  assign o[1044] = i[1044];
  assign o[1043] = i[1043];
  assign o[1042] = i[1042];
  assign o[1041] = i[1041];
  assign o[1040] = i[1040];
  assign o[1039] = i[1039];
  assign o[1038] = i[1038];
  assign o[1037] = i[1037];
  assign o[1036] = i[1036];
  assign o[1035] = i[1035];
  assign o[1034] = i[1034];
  assign o[1033] = i[1033];
  assign o[1032] = i[1032];
  assign o[1031] = i[1031];
  assign o[1030] = i[1030];
  assign o[1029] = i[1029];
  assign o[1028] = i[1028];
  assign o[1027] = i[1027];
  assign o[1026] = i[1026];
  assign o[1025] = i[1025];
  assign o[1024] = i[1024];
  assign o[1023] = i[1023];
  assign o[1022] = i[1022];
  assign o[1021] = i[1021];
  assign o[1020] = i[1020];
  assign o[1019] = i[1019];
  assign o[1018] = i[1018];
  assign o[1017] = i[1017];
  assign o[1016] = i[1016];
  assign o[1015] = i[1015];
  assign o[1014] = i[1014];
  assign o[1013] = i[1013];
  assign o[1012] = i[1012];
  assign o[1011] = i[1011];
  assign o[1010] = i[1010];
  assign o[1009] = i[1009];
  assign o[1008] = i[1008];
  assign o[1007] = i[1007];
  assign o[1006] = i[1006];
  assign o[1005] = i[1005];
  assign o[1004] = i[1004];
  assign o[1003] = i[1003];
  assign o[1002] = i[1002];
  assign o[1001] = i[1001];
  assign o[1000] = i[1000];
  assign o[999] = i[999];
  assign o[998] = i[998];
  assign o[997] = i[997];
  assign o[996] = i[996];
  assign o[995] = i[995];
  assign o[994] = i[994];
  assign o[993] = i[993];
  assign o[992] = i[992];
  assign o[991] = i[991];
  assign o[990] = i[990];
  assign o[989] = i[989];
  assign o[988] = i[988];
  assign o[987] = i[987];
  assign o[986] = i[986];
  assign o[985] = i[985];
  assign o[984] = i[984];
  assign o[983] = i[983];
  assign o[982] = i[982];
  assign o[981] = i[981];
  assign o[980] = i[980];
  assign o[979] = i[979];
  assign o[978] = i[978];
  assign o[977] = i[977];
  assign o[976] = i[976];
  assign o[975] = i[975];
  assign o[974] = i[974];
  assign o[973] = i[973];
  assign o[972] = i[972];
  assign o[971] = i[971];
  assign o[970] = i[970];
  assign o[969] = i[969];
  assign o[968] = i[968];
  assign o[967] = i[967];
  assign o[966] = i[966];
  assign o[965] = i[965];
  assign o[964] = i[964];
  assign o[963] = i[963];
  assign o[962] = i[962];
  assign o[961] = i[961];
  assign o[960] = i[960];
  assign o[959] = i[959];
  assign o[958] = i[958];
  assign o[957] = i[957];
  assign o[956] = i[956];
  assign o[955] = i[955];
  assign o[954] = i[954];
  assign o[953] = i[953];
  assign o[952] = i[952];
  assign o[951] = i[951];
  assign o[950] = i[950];
  assign o[949] = i[949];
  assign o[948] = i[948];
  assign o[947] = i[947];
  assign o[946] = i[946];
  assign o[945] = i[945];
  assign o[944] = i[944];
  assign o[943] = i[943];
  assign o[942] = i[942];
  assign o[941] = i[941];
  assign o[940] = i[940];
  assign o[939] = i[939];
  assign o[938] = i[938];
  assign o[937] = i[937];
  assign o[936] = i[936];
  assign o[935] = i[935];
  assign o[934] = i[934];
  assign o[933] = i[933];
  assign o[932] = i[932];
  assign o[931] = i[931];
  assign o[930] = i[930];
  assign o[929] = i[929];
  assign o[928] = i[928];
  assign o[927] = i[927];
  assign o[926] = i[926];
  assign o[925] = i[925];
  assign o[924] = i[924];
  assign o[923] = i[923];
  assign o[922] = i[922];
  assign o[921] = i[921];
  assign o[920] = i[920];
  assign o[919] = i[919];
  assign o[918] = i[918];
  assign o[917] = i[917];
  assign o[916] = i[916];
  assign o[915] = i[915];
  assign o[914] = i[914];
  assign o[913] = i[913];
  assign o[912] = i[912];
  assign o[911] = i[911];
  assign o[910] = i[910];
  assign o[909] = i[909];
  assign o[908] = i[908];
  assign o[907] = i[907];
  assign o[906] = i[906];
  assign o[905] = i[905];
  assign o[904] = i[904];
  assign o[903] = i[903];
  assign o[902] = i[902];
  assign o[901] = i[901];
  assign o[900] = i[900];
  assign o[899] = i[899];
  assign o[898] = i[898];
  assign o[897] = i[897];
  assign o[896] = i[896];
  assign o[895] = i[895];
  assign o[894] = i[894];
  assign o[893] = i[893];
  assign o[892] = i[892];
  assign o[891] = i[891];
  assign o[890] = i[890];
  assign o[889] = i[889];
  assign o[888] = i[888];
  assign o[887] = i[887];
  assign o[886] = i[886];
  assign o[885] = i[885];
  assign o[884] = i[884];
  assign o[883] = i[883];
  assign o[882] = i[882];
  assign o[881] = i[881];
  assign o[880] = i[880];
  assign o[879] = i[879];
  assign o[878] = i[878];
  assign o[877] = i[877];
  assign o[876] = i[876];
  assign o[875] = i[875];
  assign o[874] = i[874];
  assign o[873] = i[873];
  assign o[872] = i[872];
  assign o[871] = i[871];
  assign o[870] = i[870];
  assign o[869] = i[869];
  assign o[868] = i[868];
  assign o[867] = i[867];
  assign o[866] = i[866];
  assign o[865] = i[865];
  assign o[864] = i[864];
  assign o[863] = i[863];
  assign o[862] = i[862];
  assign o[861] = i[861];
  assign o[860] = i[860];
  assign o[859] = i[859];
  assign o[858] = i[858];
  assign o[857] = i[857];
  assign o[856] = i[856];
  assign o[855] = i[855];
  assign o[854] = i[854];
  assign o[853] = i[853];
  assign o[852] = i[852];
  assign o[851] = i[851];
  assign o[850] = i[850];
  assign o[849] = i[849];
  assign o[848] = i[848];
  assign o[847] = i[847];
  assign o[846] = i[846];
  assign o[845] = i[845];
  assign o[844] = i[844];
  assign o[843] = i[843];
  assign o[842] = i[842];
  assign o[841] = i[841];
  assign o[840] = i[840];
  assign o[839] = i[839];
  assign o[838] = i[838];
  assign o[837] = i[837];
  assign o[836] = i[836];
  assign o[835] = i[835];
  assign o[834] = i[834];
  assign o[833] = i[833];
  assign o[832] = i[832];
  assign o[831] = i[831];
  assign o[830] = i[830];
  assign o[829] = i[829];
  assign o[828] = i[828];
  assign o[827] = i[827];
  assign o[826] = i[826];
  assign o[825] = i[825];
  assign o[824] = i[824];
  assign o[823] = i[823];
  assign o[822] = i[822];
  assign o[821] = i[821];
  assign o[820] = i[820];
  assign o[819] = i[819];
  assign o[818] = i[818];
  assign o[817] = i[817];
  assign o[816] = i[816];
  assign o[815] = i[815];
  assign o[814] = i[814];
  assign o[813] = i[813];
  assign o[812] = i[812];
  assign o[811] = i[811];
  assign o[810] = i[810];
  assign o[809] = i[809];
  assign o[808] = i[808];
  assign o[807] = i[807];
  assign o[806] = i[806];
  assign o[805] = i[805];
  assign o[804] = i[804];
  assign o[803] = i[803];
  assign o[802] = i[802];
  assign o[801] = i[801];
  assign o[800] = i[800];
  assign o[799] = i[799];
  assign o[798] = i[798];
  assign o[797] = i[797];
  assign o[796] = i[796];
  assign o[795] = i[795];
  assign o[794] = i[794];
  assign o[793] = i[793];
  assign o[792] = i[792];
  assign o[791] = i[791];
  assign o[790] = i[790];
  assign o[789] = i[789];
  assign o[788] = i[788];
  assign o[787] = i[787];
  assign o[786] = i[786];
  assign o[785] = i[785];
  assign o[784] = i[784];
  assign o[783] = i[783];
  assign o[782] = i[782];
  assign o[781] = i[781];
  assign o[780] = i[780];
  assign o[779] = i[779];
  assign o[778] = i[778];
  assign o[777] = i[777];
  assign o[776] = i[776];
  assign o[775] = i[775];
  assign o[774] = i[774];
  assign o[773] = i[773];
  assign o[772] = i[772];
  assign o[771] = i[771];
  assign o[770] = i[770];
  assign o[769] = i[769];
  assign o[768] = i[768];
  assign o[767] = i[767];
  assign o[766] = i[766];
  assign o[765] = i[765];
  assign o[764] = i[764];
  assign o[763] = i[763];
  assign o[762] = i[762];
  assign o[761] = i[761];
  assign o[760] = i[760];
  assign o[759] = i[759];
  assign o[758] = i[758];
  assign o[757] = i[757];
  assign o[756] = i[756];
  assign o[755] = i[755];
  assign o[754] = i[754];
  assign o[753] = i[753];
  assign o[752] = i[752];
  assign o[751] = i[751];
  assign o[750] = i[750];
  assign o[749] = i[749];
  assign o[748] = i[748];
  assign o[747] = i[747];
  assign o[746] = i[746];
  assign o[745] = i[745];
  assign o[744] = i[744];
  assign o[743] = i[743];
  assign o[742] = i[742];
  assign o[741] = i[741];
  assign o[740] = i[740];
  assign o[739] = i[739];
  assign o[738] = i[738];
  assign o[737] = i[737];
  assign o[736] = i[736];
  assign o[735] = i[735];
  assign o[734] = i[734];
  assign o[733] = i[733];
  assign o[732] = i[732];
  assign o[731] = i[731];
  assign o[730] = i[730];
  assign o[729] = i[729];
  assign o[728] = i[728];
  assign o[727] = i[727];
  assign o[726] = i[726];
  assign o[725] = i[725];
  assign o[724] = i[724];
  assign o[723] = i[723];
  assign o[722] = i[722];
  assign o[721] = i[721];
  assign o[720] = i[720];
  assign o[719] = i[719];
  assign o[718] = i[718];
  assign o[717] = i[717];
  assign o[716] = i[716];
  assign o[715] = i[715];
  assign o[714] = i[714];
  assign o[713] = i[713];
  assign o[712] = i[712];
  assign o[711] = i[711];
  assign o[710] = i[710];
  assign o[709] = i[709];
  assign o[708] = i[708];
  assign o[707] = i[707];
  assign o[706] = i[706];
  assign o[705] = i[705];
  assign o[704] = i[704];
  assign o[703] = i[703];
  assign o[702] = i[702];
  assign o[701] = i[701];
  assign o[700] = i[700];
  assign o[699] = i[699];
  assign o[698] = i[698];
  assign o[697] = i[697];
  assign o[696] = i[696];
  assign o[695] = i[695];
  assign o[694] = i[694];
  assign o[693] = i[693];
  assign o[692] = i[692];
  assign o[691] = i[691];
  assign o[690] = i[690];
  assign o[689] = i[689];
  assign o[688] = i[688];
  assign o[687] = i[687];
  assign o[686] = i[686];
  assign o[685] = i[685];
  assign o[684] = i[684];
  assign o[683] = i[683];
  assign o[682] = i[682];
  assign o[681] = i[681];
  assign o[680] = i[680];
  assign o[679] = i[679];
  assign o[678] = i[678];
  assign o[677] = i[677];
  assign o[676] = i[676];
  assign o[675] = i[675];
  assign o[674] = i[674];
  assign o[673] = i[673];
  assign o[672] = i[672];
  assign o[671] = i[671];
  assign o[670] = i[670];
  assign o[669] = i[669];
  assign o[668] = i[668];
  assign o[667] = i[667];
  assign o[666] = i[666];
  assign o[665] = i[665];
  assign o[664] = i[664];
  assign o[663] = i[663];
  assign o[662] = i[662];
  assign o[661] = i[661];
  assign o[660] = i[660];
  assign o[659] = i[659];
  assign o[658] = i[658];
  assign o[657] = i[657];
  assign o[656] = i[656];
  assign o[655] = i[655];
  assign o[654] = i[654];
  assign o[653] = i[653];
  assign o[652] = i[652];
  assign o[651] = i[651];
  assign o[650] = i[650];
  assign o[649] = i[649];
  assign o[648] = i[648];
  assign o[647] = i[647];
  assign o[646] = i[646];
  assign o[645] = i[645];
  assign o[644] = i[644];
  assign o[643] = i[643];
  assign o[642] = i[642];
  assign o[641] = i[641];
  assign o[640] = i[640];
  assign o[639] = i[639];
  assign o[638] = i[638];
  assign o[637] = i[637];
  assign o[636] = i[636];
  assign o[635] = i[635];
  assign o[634] = i[634];
  assign o[633] = i[633];
  assign o[632] = i[632];
  assign o[631] = i[631];
  assign o[630] = i[630];
  assign o[629] = i[629];
  assign o[628] = i[628];
  assign o[627] = i[627];
  assign o[626] = i[626];
  assign o[625] = i[625];
  assign o[624] = i[624];
  assign o[623] = i[623];
  assign o[622] = i[622];
  assign o[621] = i[621];
  assign o[620] = i[620];
  assign o[619] = i[619];
  assign o[618] = i[618];
  assign o[617] = i[617];
  assign o[616] = i[616];
  assign o[615] = i[615];
  assign o[614] = i[614];
  assign o[613] = i[613];
  assign o[612] = i[612];
  assign o[611] = i[611];
  assign o[610] = i[610];
  assign o[609] = i[609];
  assign o[608] = i[608];
  assign o[607] = i[607];
  assign o[606] = i[606];
  assign o[605] = i[605];
  assign o[604] = i[604];
  assign o[603] = i[603];
  assign o[602] = i[602];
  assign o[601] = i[601];
  assign o[600] = i[600];
  assign o[599] = i[599];
  assign o[598] = i[598];
  assign o[597] = i[597];
  assign o[596] = i[596];
  assign o[595] = i[595];
  assign o[594] = i[594];
  assign o[593] = i[593];
  assign o[592] = i[592];
  assign o[591] = i[591];
  assign o[590] = i[590];
  assign o[589] = i[589];
  assign o[588] = i[588];
  assign o[587] = i[587];
  assign o[586] = i[586];
  assign o[585] = i[585];
  assign o[584] = i[584];
  assign o[583] = i[583];
  assign o[582] = i[582];
  assign o[581] = i[581];
  assign o[580] = i[580];
  assign o[579] = i[579];
  assign o[578] = i[578];
  assign o[577] = i[577];
  assign o[576] = i[576];
  assign o[575] = i[575];
  assign o[574] = i[574];
  assign o[573] = i[573];
  assign o[572] = i[572];
  assign o[571] = i[571];
  assign o[570] = i[570];
  assign o[569] = i[569];
  assign o[568] = i[568];
  assign o[567] = i[567];
  assign o[566] = i[566];
  assign o[565] = i[565];
  assign o[564] = i[564];
  assign o[563] = i[563];
  assign o[562] = i[562];
  assign o[561] = i[561];
  assign o[560] = i[560];
  assign o[559] = i[559];
  assign o[558] = i[558];
  assign o[557] = i[557];
  assign o[556] = i[556];
  assign o[555] = i[555];
  assign o[554] = i[554];
  assign o[553] = i[553];
  assign o[552] = i[552];
  assign o[551] = i[551];
  assign o[550] = i[550];
  assign o[549] = i[549];
  assign o[548] = i[548];
  assign o[547] = i[547];
  assign o[546] = i[546];
  assign o[545] = i[545];
  assign o[544] = i[544];
  assign o[543] = i[543];
  assign o[542] = i[542];
  assign o[541] = i[541];
  assign o[540] = i[540];
  assign o[539] = i[539];
  assign o[538] = i[538];
  assign o[537] = i[537];
  assign o[536] = i[536];
  assign o[535] = i[535];
  assign o[534] = i[534];
  assign o[533] = i[533];
  assign o[532] = i[532];
  assign o[531] = i[531];
  assign o[530] = i[530];
  assign o[529] = i[529];
  assign o[528] = i[528];
  assign o[527] = i[527];
  assign o[526] = i[526];
  assign o[525] = i[525];
  assign o[524] = i[524];
  assign o[523] = i[523];
  assign o[522] = i[522];
  assign o[521] = i[521];
  assign o[520] = i[520];
  assign o[519] = i[519];
  assign o[518] = i[518];
  assign o[517] = i[517];
  assign o[516] = i[516];
  assign o[515] = i[515];
  assign o[514] = i[514];
  assign o[513] = i[513];
  assign o[512] = i[512];
  assign o[511] = i[511];
  assign o[510] = i[510];
  assign o[509] = i[509];
  assign o[508] = i[508];
  assign o[507] = i[507];
  assign o[506] = i[506];
  assign o[505] = i[505];
  assign o[504] = i[504];
  assign o[503] = i[503];
  assign o[502] = i[502];
  assign o[501] = i[501];
  assign o[500] = i[500];
  assign o[499] = i[499];
  assign o[498] = i[498];
  assign o[497] = i[497];
  assign o[496] = i[496];
  assign o[495] = i[495];
  assign o[494] = i[494];
  assign o[493] = i[493];
  assign o[492] = i[492];
  assign o[491] = i[491];
  assign o[490] = i[490];
  assign o[489] = i[489];
  assign o[488] = i[488];
  assign o[487] = i[487];
  assign o[486] = i[486];
  assign o[485] = i[485];
  assign o[484] = i[484];
  assign o[483] = i[483];
  assign o[482] = i[482];
  assign o[481] = i[481];
  assign o[480] = i[480];
  assign o[479] = i[479];
  assign o[478] = i[478];
  assign o[477] = i[477];
  assign o[476] = i[476];
  assign o[475] = i[475];
  assign o[474] = i[474];
  assign o[473] = i[473];
  assign o[472] = i[472];
  assign o[471] = i[471];
  assign o[470] = i[470];
  assign o[469] = i[469];
  assign o[468] = i[468];
  assign o[467] = i[467];
  assign o[466] = i[466];
  assign o[465] = i[465];
  assign o[464] = i[464];
  assign o[463] = i[463];
  assign o[462] = i[462];
  assign o[461] = i[461];
  assign o[460] = i[460];
  assign o[459] = i[459];
  assign o[458] = i[458];
  assign o[457] = i[457];
  assign o[456] = i[456];
  assign o[455] = i[455];
  assign o[454] = i[454];
  assign o[453] = i[453];
  assign o[452] = i[452];
  assign o[451] = i[451];
  assign o[450] = i[450];
  assign o[449] = i[449];
  assign o[448] = i[448];
  assign o[447] = i[447];
  assign o[446] = i[446];
  assign o[445] = i[445];
  assign o[444] = i[444];
  assign o[443] = i[443];
  assign o[442] = i[442];
  assign o[441] = i[441];
  assign o[440] = i[440];
  assign o[439] = i[439];
  assign o[438] = i[438];
  assign o[437] = i[437];
  assign o[436] = i[436];
  assign o[435] = i[435];
  assign o[434] = i[434];
  assign o[433] = i[433];
  assign o[432] = i[432];
  assign o[431] = i[431];
  assign o[430] = i[430];
  assign o[429] = i[429];
  assign o[428] = i[428];
  assign o[427] = i[427];
  assign o[426] = i[426];
  assign o[425] = i[425];
  assign o[424] = i[424];
  assign o[423] = i[423];
  assign o[422] = i[422];
  assign o[421] = i[421];
  assign o[420] = i[420];
  assign o[419] = i[419];
  assign o[418] = i[418];
  assign o[417] = i[417];
  assign o[416] = i[416];
  assign o[415] = i[415];
  assign o[414] = i[414];
  assign o[413] = i[413];
  assign o[412] = i[412];
  assign o[411] = i[411];
  assign o[410] = i[410];
  assign o[409] = i[409];
  assign o[408] = i[408];
  assign o[407] = i[407];
  assign o[406] = i[406];
  assign o[405] = i[405];
  assign o[404] = i[404];
  assign o[403] = i[403];
  assign o[402] = i[402];
  assign o[401] = i[401];
  assign o[400] = i[400];
  assign o[399] = i[399];
  assign o[398] = i[398];
  assign o[397] = i[397];
  assign o[396] = i[396];
  assign o[395] = i[395];
  assign o[394] = i[394];
  assign o[393] = i[393];
  assign o[392] = i[392];
  assign o[391] = i[391];
  assign o[390] = i[390];
  assign o[389] = i[389];
  assign o[388] = i[388];
  assign o[387] = i[387];
  assign o[386] = i[386];
  assign o[385] = i[385];
  assign o[384] = i[384];
  assign o[383] = i[383];
  assign o[382] = i[382];
  assign o[381] = i[381];
  assign o[380] = i[380];
  assign o[379] = i[379];
  assign o[378] = i[378];
  assign o[377] = i[377];
  assign o[376] = i[376];
  assign o[375] = i[375];
  assign o[374] = i[374];
  assign o[373] = i[373];
  assign o[372] = i[372];
  assign o[371] = i[371];
  assign o[370] = i[370];
  assign o[369] = i[369];
  assign o[368] = i[368];
  assign o[367] = i[367];
  assign o[366] = i[366];
  assign o[365] = i[365];
  assign o[364] = i[364];
  assign o[363] = i[363];
  assign o[362] = i[362];
  assign o[361] = i[361];
  assign o[360] = i[360];
  assign o[359] = i[359];
  assign o[358] = i[358];
  assign o[357] = i[357];
  assign o[356] = i[356];
  assign o[355] = i[355];
  assign o[354] = i[354];
  assign o[353] = i[353];
  assign o[352] = i[352];
  assign o[351] = i[351];
  assign o[350] = i[350];
  assign o[349] = i[349];
  assign o[348] = i[348];
  assign o[347] = i[347];
  assign o[346] = i[346];
  assign o[345] = i[345];
  assign o[344] = i[344];
  assign o[343] = i[343];
  assign o[342] = i[342];
  assign o[341] = i[341];
  assign o[340] = i[340];
  assign o[339] = i[339];
  assign o[338] = i[338];
  assign o[337] = i[337];
  assign o[336] = i[336];
  assign o[335] = i[335];
  assign o[334] = i[334];
  assign o[333] = i[333];
  assign o[332] = i[332];
  assign o[331] = i[331];
  assign o[330] = i[330];
  assign o[329] = i[329];
  assign o[328] = i[328];
  assign o[327] = i[327];
  assign o[326] = i[326];
  assign o[325] = i[325];
  assign o[324] = i[324];
  assign o[323] = i[323];
  assign o[322] = i[322];
  assign o[321] = i[321];
  assign o[320] = i[320];
  assign o[319] = i[319];
  assign o[318] = i[318];
  assign o[317] = i[317];
  assign o[316] = i[316];
  assign o[315] = i[315];
  assign o[314] = i[314];
  assign o[313] = i[313];
  assign o[312] = i[312];
  assign o[311] = i[311];
  assign o[310] = i[310];
  assign o[309] = i[309];
  assign o[308] = i[308];
  assign o[307] = i[307];
  assign o[306] = i[306];
  assign o[305] = i[305];
  assign o[304] = i[304];
  assign o[303] = i[303];
  assign o[302] = i[302];
  assign o[301] = i[301];
  assign o[300] = i[300];
  assign o[299] = i[299];
  assign o[298] = i[298];
  assign o[297] = i[297];
  assign o[296] = i[296];
  assign o[295] = i[295];
  assign o[294] = i[294];
  assign o[293] = i[293];
  assign o[292] = i[292];
  assign o[291] = i[291];
  assign o[290] = i[290];
  assign o[289] = i[289];
  assign o[288] = i[288];
  assign o[287] = i[287];
  assign o[286] = i[286];
  assign o[285] = i[285];
  assign o[284] = i[284];
  assign o[283] = i[283];
  assign o[282] = i[282];
  assign o[281] = i[281];
  assign o[280] = i[280];
  assign o[279] = i[279];
  assign o[278] = i[278];
  assign o[277] = i[277];
  assign o[276] = i[276];
  assign o[275] = i[275];
  assign o[274] = i[274];
  assign o[273] = i[273];
  assign o[272] = i[272];
  assign o[271] = i[271];
  assign o[270] = i[270];
  assign o[269] = i[269];
  assign o[268] = i[268];
  assign o[267] = i[267];
  assign o[266] = i[266];
  assign o[265] = i[265];
  assign o[264] = i[264];
  assign o[263] = i[263];
  assign o[262] = i[262];
  assign o[261] = i[261];
  assign o[260] = i[260];
  assign o[259] = i[259];
  assign o[258] = i[258];
  assign o[257] = i[257];
  assign o[256] = i[256];
  assign o[255] = i[255];
  assign o[254] = i[254];
  assign o[253] = i[253];
  assign o[252] = i[252];
  assign o[251] = i[251];
  assign o[250] = i[250];
  assign o[249] = i[249];
  assign o[248] = i[248];
  assign o[247] = i[247];
  assign o[246] = i[246];
  assign o[245] = i[245];
  assign o[244] = i[244];
  assign o[243] = i[243];
  assign o[242] = i[242];
  assign o[241] = i[241];
  assign o[240] = i[240];
  assign o[239] = i[239];
  assign o[238] = i[238];
  assign o[237] = i[237];
  assign o[236] = i[236];
  assign o[235] = i[235];
  assign o[234] = i[234];
  assign o[233] = i[233];
  assign o[232] = i[232];
  assign o[231] = i[231];
  assign o[230] = i[230];
  assign o[229] = i[229];
  assign o[228] = i[228];
  assign o[227] = i[227];
  assign o[226] = i[226];
  assign o[225] = i[225];
  assign o[224] = i[224];
  assign o[223] = i[223];
  assign o[222] = i[222];
  assign o[221] = i[221];
  assign o[220] = i[220];
  assign o[219] = i[219];
  assign o[218] = i[218];
  assign o[217] = i[217];
  assign o[216] = i[216];
  assign o[215] = i[215];
  assign o[214] = i[214];
  assign o[213] = i[213];
  assign o[212] = i[212];
  assign o[211] = i[211];
  assign o[210] = i[210];
  assign o[209] = i[209];
  assign o[208] = i[208];
  assign o[207] = i[207];
  assign o[206] = i[206];
  assign o[205] = i[205];
  assign o[204] = i[204];
  assign o[203] = i[203];
  assign o[202] = i[202];
  assign o[201] = i[201];
  assign o[200] = i[200];
  assign o[199] = i[199];
  assign o[198] = i[198];
  assign o[197] = i[197];
  assign o[196] = i[196];
  assign o[195] = i[195];
  assign o[194] = i[194];
  assign o[193] = i[193];
  assign o[192] = i[192];
  assign o[191] = i[191];
  assign o[190] = i[190];
  assign o[189] = i[189];
  assign o[188] = i[188];
  assign o[187] = i[187];
  assign o[186] = i[186];
  assign o[185] = i[185];
  assign o[184] = i[184];
  assign o[183] = i[183];
  assign o[182] = i[182];
  assign o[181] = i[181];
  assign o[180] = i[180];
  assign o[179] = i[179];
  assign o[178] = i[178];
  assign o[177] = i[177];
  assign o[176] = i[176];
  assign o[175] = i[175];
  assign o[174] = i[174];
  assign o[173] = i[173];
  assign o[172] = i[172];
  assign o[171] = i[171];
  assign o[170] = i[170];
  assign o[169] = i[169];
  assign o[168] = i[168];
  assign o[167] = i[167];
  assign o[166] = i[166];
  assign o[165] = i[165];
  assign o[164] = i[164];
  assign o[163] = i[163];
  assign o[162] = i[162];
  assign o[161] = i[161];
  assign o[160] = i[160];
  assign o[159] = i[159];
  assign o[158] = i[158];
  assign o[157] = i[157];
  assign o[156] = i[156];
  assign o[155] = i[155];
  assign o[154] = i[154];
  assign o[153] = i[153];
  assign o[152] = i[152];
  assign o[151] = i[151];
  assign o[150] = i[150];
  assign o[149] = i[149];
  assign o[148] = i[148];
  assign o[147] = i[147];
  assign o[146] = i[146];
  assign o[145] = i[145];
  assign o[144] = i[144];
  assign o[143] = i[143];
  assign o[142] = i[142];
  assign o[141] = i[141];
  assign o[140] = i[140];
  assign o[139] = i[139];
  assign o[138] = i[138];
  assign o[137] = i[137];
  assign o[136] = i[136];
  assign o[135] = i[135];
  assign o[134] = i[134];
  assign o[133] = i[133];
  assign o[132] = i[132];
  assign o[131] = i[131];
  assign o[130] = i[130];
  assign o[129] = i[129];
  assign o[128] = i[128];
  assign o[127] = i[127];
  assign o[126] = i[126];
  assign o[125] = i[125];
  assign o[124] = i[124];
  assign o[123] = i[123];
  assign o[122] = i[122];
  assign o[121] = i[121];
  assign o[120] = i[120];
  assign o[119] = i[119];
  assign o[118] = i[118];
  assign o[117] = i[117];
  assign o[116] = i[116];
  assign o[115] = i[115];
  assign o[114] = i[114];
  assign o[113] = i[113];
  assign o[112] = i[112];
  assign o[111] = i[111];
  assign o[110] = i[110];
  assign o[109] = i[109];
  assign o[108] = i[108];
  assign o[107] = i[107];
  assign o[106] = i[106];
  assign o[105] = i[105];
  assign o[104] = i[104];
  assign o[103] = i[103];
  assign o[102] = i[102];
  assign o[101] = i[101];
  assign o[100] = i[100];
  assign o[99] = i[99];
  assign o[98] = i[98];
  assign o[97] = i[97];
  assign o[96] = i[96];
  assign o[95] = i[95];
  assign o[94] = i[94];
  assign o[93] = i[93];
  assign o[92] = i[92];
  assign o[91] = i[91];
  assign o[90] = i[90];
  assign o[89] = i[89];
  assign o[88] = i[88];
  assign o[87] = i[87];
  assign o[86] = i[86];
  assign o[85] = i[85];
  assign o[84] = i[84];
  assign o[83] = i[83];
  assign o[82] = i[82];
  assign o[81] = i[81];
  assign o[80] = i[80];
  assign o[79] = i[79];
  assign o[78] = i[78];
  assign o[77] = i[77];
  assign o[76] = i[76];
  assign o[75] = i[75];
  assign o[74] = i[74];
  assign o[73] = i[73];
  assign o[72] = i[72];
  assign o[71] = i[71];
  assign o[70] = i[70];
  assign o[69] = i[69];
  assign o[68] = i[68];
  assign o[67] = i[67];
  assign o[66] = i[66];
  assign o[65] = i[65];
  assign o[64] = i[64];
  assign o[63] = i[63];
  assign o[62] = i[62];
  assign o[61] = i[61];
  assign o[60] = i[60];
  assign o[59] = i[59];
  assign o[58] = i[58];
  assign o[57] = i[57];
  assign o[56] = i[56];
  assign o[55] = i[55];
  assign o[54] = i[54];
  assign o[53] = i[53];
  assign o[52] = i[52];
  assign o[51] = i[51];
  assign o[50] = i[50];
  assign o[49] = i[49];
  assign o[48] = i[48];
  assign o[47] = i[47];
  assign o[46] = i[46];
  assign o[45] = i[45];
  assign o[44] = i[44];
  assign o[43] = i[43];
  assign o[42] = i[42];
  assign o[41] = i[41];
  assign o[40] = i[40];
  assign o[39] = i[39];
  assign o[38] = i[38];
  assign o[37] = i[37];
  assign o[36] = i[36];
  assign o[35] = i[35];
  assign o[34] = i[34];
  assign o[33] = i[33];
  assign o[32] = i[32];
  assign o[31] = i[31];
  assign o[30] = i[30];
  assign o[29] = i[29];
  assign o[28] = i[28];
  assign o[27] = i[27];
  assign o[26] = i[26];
  assign o[25] = i[25];
  assign o[24] = i[24];
  assign o[23] = i[23];
  assign o[22] = i[22];
  assign o[21] = i[21];
  assign o[20] = i[20];
  assign o[19] = i[19];
  assign o[18] = i[18];
  assign o[17] = i[17];
  assign o[16] = i[16];
  assign o[15] = i[15];
  assign o[14] = i[14];
  assign o[13] = i[13];
  assign o[12] = i[12];
  assign o[11] = i[11];
  assign o[10] = i[10];
  assign o[9] = i[9];
  assign o[8] = i[8];
  assign o[7] = i[7];
  assign o[6] = i[6];
  assign o[5] = i[5];
  assign o[4] = i[4];
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_rotate_right_width_p10
(
  data_i,
  rot_i,
  o
);

  input [9:0] data_i;
  input [3:0] rot_i;
  output [9:0] o;
  wire [9:0] o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10;
  assign { SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, o } = { data_i, data_i } >> rot_i;

endmodule



module bsg_circular_ptr_slots_p10_max_add_p10
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [3:0] add_i;
  output [3:0] o;
  output [3:0] n_o;
  input clk;
  input reset_i;
  wire [3:0] n_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  wire [4:0] ptr_wrap;
  reg [3:0] o;
  assign { N17, N16, N15, N14 } = o + add_i;
  assign { N13, N12, N11, N10, N9 } = o - { 1'b1, 1'b0, 1'b1, 1'b0 };
  assign ptr_wrap = { N13, N12, N11, N10, N9 } + add_i;
  assign { N8, N7, N6, N5 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N1)? n_o : 1'b0;
  assign N0 = reset_i;
  assign N1 = N4;
  assign n_o = (N2)? ptr_wrap[3:0] : 
               (N3)? { N17, N16, N15, N14 } : 1'b0;
  assign N2 = N18;
  assign N3 = ptr_wrap[4];
  assign N4 = ~reset_i;
  assign N18 = ~ptr_wrap[4];

  always @(posedge clk) begin
    if(1'b1) begin
      { o[3:0] } <= { N8, N7, N6, N5 };
    end 
  end


endmodule



module bsg_rr_f2f_input_width_p128_num_in_p10_middle_meet_p10
(
  clk,
  reset,
  valid_i,
  data_i,
  data_head_o,
  valid_head_o,
  go_channels_i,
  go_cnt_i,
  yumi_o
);

  input [9:0] valid_i;
  input [1279:0] data_i;
  output [1279:0] data_head_o;
  output [9:0] valid_head_o;
  input [9:0] go_channels_i;
  input [3:0] go_cnt_i;
  output [9:0] yumi_o;
  input clk;
  input reset;
  wire [1279:0] data_head_o,data_head_o_flat_pretrunc;
  wire [9:0] valid_head_o,yumi_o;
  wire SYNOPSYS_UNCONNECTED_1,SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,
  SYNOPSYS_UNCONNECTED_4,SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,
  SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,
  SYNOPSYS_UNCONNECTED_11,SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13,
  SYNOPSYS_UNCONNECTED_14,SYNOPSYS_UNCONNECTED_15,SYNOPSYS_UNCONNECTED_16,SYNOPSYS_UNCONNECTED_17,
  SYNOPSYS_UNCONNECTED_18,SYNOPSYS_UNCONNECTED_19,SYNOPSYS_UNCONNECTED_20,
  SYNOPSYS_UNCONNECTED_21,SYNOPSYS_UNCONNECTED_22,SYNOPSYS_UNCONNECTED_23,
  SYNOPSYS_UNCONNECTED_24,SYNOPSYS_UNCONNECTED_25,SYNOPSYS_UNCONNECTED_26,SYNOPSYS_UNCONNECTED_27,
  SYNOPSYS_UNCONNECTED_28,SYNOPSYS_UNCONNECTED_29,SYNOPSYS_UNCONNECTED_30,
  SYNOPSYS_UNCONNECTED_31,SYNOPSYS_UNCONNECTED_32,SYNOPSYS_UNCONNECTED_33,
  SYNOPSYS_UNCONNECTED_34,SYNOPSYS_UNCONNECTED_35,SYNOPSYS_UNCONNECTED_36,SYNOPSYS_UNCONNECTED_37,
  SYNOPSYS_UNCONNECTED_38,SYNOPSYS_UNCONNECTED_39,SYNOPSYS_UNCONNECTED_40,
  SYNOPSYS_UNCONNECTED_41,SYNOPSYS_UNCONNECTED_42,SYNOPSYS_UNCONNECTED_43,
  SYNOPSYS_UNCONNECTED_44,SYNOPSYS_UNCONNECTED_45,SYNOPSYS_UNCONNECTED_46,SYNOPSYS_UNCONNECTED_47,
  SYNOPSYS_UNCONNECTED_48,SYNOPSYS_UNCONNECTED_49,SYNOPSYS_UNCONNECTED_50,
  SYNOPSYS_UNCONNECTED_51,SYNOPSYS_UNCONNECTED_52,SYNOPSYS_UNCONNECTED_53,
  SYNOPSYS_UNCONNECTED_54,SYNOPSYS_UNCONNECTED_55,SYNOPSYS_UNCONNECTED_56,SYNOPSYS_UNCONNECTED_57,
  SYNOPSYS_UNCONNECTED_58,SYNOPSYS_UNCONNECTED_59,SYNOPSYS_UNCONNECTED_60,
  SYNOPSYS_UNCONNECTED_61,SYNOPSYS_UNCONNECTED_62,SYNOPSYS_UNCONNECTED_63,
  SYNOPSYS_UNCONNECTED_64,SYNOPSYS_UNCONNECTED_65,SYNOPSYS_UNCONNECTED_66,SYNOPSYS_UNCONNECTED_67,
  SYNOPSYS_UNCONNECTED_68,SYNOPSYS_UNCONNECTED_69,SYNOPSYS_UNCONNECTED_70,
  SYNOPSYS_UNCONNECTED_71,SYNOPSYS_UNCONNECTED_72,SYNOPSYS_UNCONNECTED_73,
  SYNOPSYS_UNCONNECTED_74,SYNOPSYS_UNCONNECTED_75,SYNOPSYS_UNCONNECTED_76,SYNOPSYS_UNCONNECTED_77,
  SYNOPSYS_UNCONNECTED_78,SYNOPSYS_UNCONNECTED_79,SYNOPSYS_UNCONNECTED_80,
  SYNOPSYS_UNCONNECTED_81,SYNOPSYS_UNCONNECTED_82,SYNOPSYS_UNCONNECTED_83,
  SYNOPSYS_UNCONNECTED_84,SYNOPSYS_UNCONNECTED_85,SYNOPSYS_UNCONNECTED_86,SYNOPSYS_UNCONNECTED_87,
  SYNOPSYS_UNCONNECTED_88,SYNOPSYS_UNCONNECTED_89,SYNOPSYS_UNCONNECTED_90,
  SYNOPSYS_UNCONNECTED_91,SYNOPSYS_UNCONNECTED_92,SYNOPSYS_UNCONNECTED_93,
  SYNOPSYS_UNCONNECTED_94,SYNOPSYS_UNCONNECTED_95,SYNOPSYS_UNCONNECTED_96,SYNOPSYS_UNCONNECTED_97,
  SYNOPSYS_UNCONNECTED_98,SYNOPSYS_UNCONNECTED_99,SYNOPSYS_UNCONNECTED_100,
  SYNOPSYS_UNCONNECTED_101,SYNOPSYS_UNCONNECTED_102,SYNOPSYS_UNCONNECTED_103,
  SYNOPSYS_UNCONNECTED_104,SYNOPSYS_UNCONNECTED_105,SYNOPSYS_UNCONNECTED_106,
  SYNOPSYS_UNCONNECTED_107,SYNOPSYS_UNCONNECTED_108,SYNOPSYS_UNCONNECTED_109,
  SYNOPSYS_UNCONNECTED_110,SYNOPSYS_UNCONNECTED_111,SYNOPSYS_UNCONNECTED_112,SYNOPSYS_UNCONNECTED_113,
  SYNOPSYS_UNCONNECTED_114,SYNOPSYS_UNCONNECTED_115,SYNOPSYS_UNCONNECTED_116,
  SYNOPSYS_UNCONNECTED_117,SYNOPSYS_UNCONNECTED_118,SYNOPSYS_UNCONNECTED_119,
  SYNOPSYS_UNCONNECTED_120,SYNOPSYS_UNCONNECTED_121,SYNOPSYS_UNCONNECTED_122,
  SYNOPSYS_UNCONNECTED_123,SYNOPSYS_UNCONNECTED_124,SYNOPSYS_UNCONNECTED_125,
  SYNOPSYS_UNCONNECTED_126,SYNOPSYS_UNCONNECTED_127,SYNOPSYS_UNCONNECTED_128,SYNOPSYS_UNCONNECTED_129,
  SYNOPSYS_UNCONNECTED_130,SYNOPSYS_UNCONNECTED_131,SYNOPSYS_UNCONNECTED_132,
  SYNOPSYS_UNCONNECTED_133,SYNOPSYS_UNCONNECTED_134,SYNOPSYS_UNCONNECTED_135,
  SYNOPSYS_UNCONNECTED_136,SYNOPSYS_UNCONNECTED_137,SYNOPSYS_UNCONNECTED_138,
  SYNOPSYS_UNCONNECTED_139,SYNOPSYS_UNCONNECTED_140,SYNOPSYS_UNCONNECTED_141,
  SYNOPSYS_UNCONNECTED_142,SYNOPSYS_UNCONNECTED_143,SYNOPSYS_UNCONNECTED_144,SYNOPSYS_UNCONNECTED_145,
  SYNOPSYS_UNCONNECTED_146,SYNOPSYS_UNCONNECTED_147,SYNOPSYS_UNCONNECTED_148,
  SYNOPSYS_UNCONNECTED_149,SYNOPSYS_UNCONNECTED_150,SYNOPSYS_UNCONNECTED_151,
  SYNOPSYS_UNCONNECTED_152,SYNOPSYS_UNCONNECTED_153,SYNOPSYS_UNCONNECTED_154,
  SYNOPSYS_UNCONNECTED_155,SYNOPSYS_UNCONNECTED_156,SYNOPSYS_UNCONNECTED_157,
  SYNOPSYS_UNCONNECTED_158,SYNOPSYS_UNCONNECTED_159,SYNOPSYS_UNCONNECTED_160,SYNOPSYS_UNCONNECTED_161,
  SYNOPSYS_UNCONNECTED_162,SYNOPSYS_UNCONNECTED_163,SYNOPSYS_UNCONNECTED_164,
  SYNOPSYS_UNCONNECTED_165,SYNOPSYS_UNCONNECTED_166,SYNOPSYS_UNCONNECTED_167,
  SYNOPSYS_UNCONNECTED_168,SYNOPSYS_UNCONNECTED_169,SYNOPSYS_UNCONNECTED_170,
  SYNOPSYS_UNCONNECTED_171,SYNOPSYS_UNCONNECTED_172,SYNOPSYS_UNCONNECTED_173,
  SYNOPSYS_UNCONNECTED_174,SYNOPSYS_UNCONNECTED_175,SYNOPSYS_UNCONNECTED_176,SYNOPSYS_UNCONNECTED_177,
  SYNOPSYS_UNCONNECTED_178,SYNOPSYS_UNCONNECTED_179,SYNOPSYS_UNCONNECTED_180,
  SYNOPSYS_UNCONNECTED_181,SYNOPSYS_UNCONNECTED_182,SYNOPSYS_UNCONNECTED_183,
  SYNOPSYS_UNCONNECTED_184,SYNOPSYS_UNCONNECTED_185,SYNOPSYS_UNCONNECTED_186,
  SYNOPSYS_UNCONNECTED_187,SYNOPSYS_UNCONNECTED_188,SYNOPSYS_UNCONNECTED_189,
  SYNOPSYS_UNCONNECTED_190,SYNOPSYS_UNCONNECTED_191,SYNOPSYS_UNCONNECTED_192,SYNOPSYS_UNCONNECTED_193,
  SYNOPSYS_UNCONNECTED_194,SYNOPSYS_UNCONNECTED_195,SYNOPSYS_UNCONNECTED_196,
  SYNOPSYS_UNCONNECTED_197,SYNOPSYS_UNCONNECTED_198,SYNOPSYS_UNCONNECTED_199,
  SYNOPSYS_UNCONNECTED_200,SYNOPSYS_UNCONNECTED_201,SYNOPSYS_UNCONNECTED_202,
  SYNOPSYS_UNCONNECTED_203,SYNOPSYS_UNCONNECTED_204,SYNOPSYS_UNCONNECTED_205,
  SYNOPSYS_UNCONNECTED_206,SYNOPSYS_UNCONNECTED_207,SYNOPSYS_UNCONNECTED_208,SYNOPSYS_UNCONNECTED_209,
  SYNOPSYS_UNCONNECTED_210,SYNOPSYS_UNCONNECTED_211,SYNOPSYS_UNCONNECTED_212,
  SYNOPSYS_UNCONNECTED_213,SYNOPSYS_UNCONNECTED_214,SYNOPSYS_UNCONNECTED_215,
  SYNOPSYS_UNCONNECTED_216,SYNOPSYS_UNCONNECTED_217,SYNOPSYS_UNCONNECTED_218,
  SYNOPSYS_UNCONNECTED_219,SYNOPSYS_UNCONNECTED_220,SYNOPSYS_UNCONNECTED_221,
  SYNOPSYS_UNCONNECTED_222,SYNOPSYS_UNCONNECTED_223,SYNOPSYS_UNCONNECTED_224,SYNOPSYS_UNCONNECTED_225,
  SYNOPSYS_UNCONNECTED_226,SYNOPSYS_UNCONNECTED_227,SYNOPSYS_UNCONNECTED_228,
  SYNOPSYS_UNCONNECTED_229,SYNOPSYS_UNCONNECTED_230,SYNOPSYS_UNCONNECTED_231,
  SYNOPSYS_UNCONNECTED_232,SYNOPSYS_UNCONNECTED_233,SYNOPSYS_UNCONNECTED_234,
  SYNOPSYS_UNCONNECTED_235,SYNOPSYS_UNCONNECTED_236,SYNOPSYS_UNCONNECTED_237,
  SYNOPSYS_UNCONNECTED_238,SYNOPSYS_UNCONNECTED_239,SYNOPSYS_UNCONNECTED_240,SYNOPSYS_UNCONNECTED_241,
  SYNOPSYS_UNCONNECTED_242,SYNOPSYS_UNCONNECTED_243,SYNOPSYS_UNCONNECTED_244,
  SYNOPSYS_UNCONNECTED_245,SYNOPSYS_UNCONNECTED_246,SYNOPSYS_UNCONNECTED_247,
  SYNOPSYS_UNCONNECTED_248,SYNOPSYS_UNCONNECTED_249,SYNOPSYS_UNCONNECTED_250,
  SYNOPSYS_UNCONNECTED_251,SYNOPSYS_UNCONNECTED_252,SYNOPSYS_UNCONNECTED_253,
  SYNOPSYS_UNCONNECTED_254,SYNOPSYS_UNCONNECTED_255,SYNOPSYS_UNCONNECTED_256,SYNOPSYS_UNCONNECTED_257,
  SYNOPSYS_UNCONNECTED_258,SYNOPSYS_UNCONNECTED_259,SYNOPSYS_UNCONNECTED_260,
  SYNOPSYS_UNCONNECTED_261,SYNOPSYS_UNCONNECTED_262,SYNOPSYS_UNCONNECTED_263,
  SYNOPSYS_UNCONNECTED_264,SYNOPSYS_UNCONNECTED_265,SYNOPSYS_UNCONNECTED_266,
  SYNOPSYS_UNCONNECTED_267,SYNOPSYS_UNCONNECTED_268,SYNOPSYS_UNCONNECTED_269,
  SYNOPSYS_UNCONNECTED_270,SYNOPSYS_UNCONNECTED_271,SYNOPSYS_UNCONNECTED_272,SYNOPSYS_UNCONNECTED_273,
  SYNOPSYS_UNCONNECTED_274,SYNOPSYS_UNCONNECTED_275,SYNOPSYS_UNCONNECTED_276,
  SYNOPSYS_UNCONNECTED_277,SYNOPSYS_UNCONNECTED_278,SYNOPSYS_UNCONNECTED_279,
  SYNOPSYS_UNCONNECTED_280,SYNOPSYS_UNCONNECTED_281,SYNOPSYS_UNCONNECTED_282,
  SYNOPSYS_UNCONNECTED_283,SYNOPSYS_UNCONNECTED_284,SYNOPSYS_UNCONNECTED_285,
  SYNOPSYS_UNCONNECTED_286,SYNOPSYS_UNCONNECTED_287,SYNOPSYS_UNCONNECTED_288,SYNOPSYS_UNCONNECTED_289,
  SYNOPSYS_UNCONNECTED_290,SYNOPSYS_UNCONNECTED_291,SYNOPSYS_UNCONNECTED_292,
  SYNOPSYS_UNCONNECTED_293,SYNOPSYS_UNCONNECTED_294,SYNOPSYS_UNCONNECTED_295,
  SYNOPSYS_UNCONNECTED_296,SYNOPSYS_UNCONNECTED_297,SYNOPSYS_UNCONNECTED_298,
  SYNOPSYS_UNCONNECTED_299,SYNOPSYS_UNCONNECTED_300,SYNOPSYS_UNCONNECTED_301,
  SYNOPSYS_UNCONNECTED_302,SYNOPSYS_UNCONNECTED_303,SYNOPSYS_UNCONNECTED_304,SYNOPSYS_UNCONNECTED_305,
  SYNOPSYS_UNCONNECTED_306,SYNOPSYS_UNCONNECTED_307,SYNOPSYS_UNCONNECTED_308,
  SYNOPSYS_UNCONNECTED_309,SYNOPSYS_UNCONNECTED_310,SYNOPSYS_UNCONNECTED_311,
  SYNOPSYS_UNCONNECTED_312,SYNOPSYS_UNCONNECTED_313,SYNOPSYS_UNCONNECTED_314,
  SYNOPSYS_UNCONNECTED_315,SYNOPSYS_UNCONNECTED_316,SYNOPSYS_UNCONNECTED_317,
  SYNOPSYS_UNCONNECTED_318,SYNOPSYS_UNCONNECTED_319,SYNOPSYS_UNCONNECTED_320,SYNOPSYS_UNCONNECTED_321,
  SYNOPSYS_UNCONNECTED_322,SYNOPSYS_UNCONNECTED_323,SYNOPSYS_UNCONNECTED_324,
  SYNOPSYS_UNCONNECTED_325,SYNOPSYS_UNCONNECTED_326,SYNOPSYS_UNCONNECTED_327,
  SYNOPSYS_UNCONNECTED_328,SYNOPSYS_UNCONNECTED_329,SYNOPSYS_UNCONNECTED_330,
  SYNOPSYS_UNCONNECTED_331,SYNOPSYS_UNCONNECTED_332,SYNOPSYS_UNCONNECTED_333,
  SYNOPSYS_UNCONNECTED_334,SYNOPSYS_UNCONNECTED_335,SYNOPSYS_UNCONNECTED_336,SYNOPSYS_UNCONNECTED_337,
  SYNOPSYS_UNCONNECTED_338,SYNOPSYS_UNCONNECTED_339,SYNOPSYS_UNCONNECTED_340,
  SYNOPSYS_UNCONNECTED_341,SYNOPSYS_UNCONNECTED_342,SYNOPSYS_UNCONNECTED_343,
  SYNOPSYS_UNCONNECTED_344,SYNOPSYS_UNCONNECTED_345,SYNOPSYS_UNCONNECTED_346,
  SYNOPSYS_UNCONNECTED_347,SYNOPSYS_UNCONNECTED_348,SYNOPSYS_UNCONNECTED_349,
  SYNOPSYS_UNCONNECTED_350,SYNOPSYS_UNCONNECTED_351,SYNOPSYS_UNCONNECTED_352,SYNOPSYS_UNCONNECTED_353,
  SYNOPSYS_UNCONNECTED_354,SYNOPSYS_UNCONNECTED_355,SYNOPSYS_UNCONNECTED_356,
  SYNOPSYS_UNCONNECTED_357,SYNOPSYS_UNCONNECTED_358,SYNOPSYS_UNCONNECTED_359,
  SYNOPSYS_UNCONNECTED_360,SYNOPSYS_UNCONNECTED_361,SYNOPSYS_UNCONNECTED_362,
  SYNOPSYS_UNCONNECTED_363,SYNOPSYS_UNCONNECTED_364,SYNOPSYS_UNCONNECTED_365,
  SYNOPSYS_UNCONNECTED_366,SYNOPSYS_UNCONNECTED_367,SYNOPSYS_UNCONNECTED_368,SYNOPSYS_UNCONNECTED_369,
  SYNOPSYS_UNCONNECTED_370,SYNOPSYS_UNCONNECTED_371,SYNOPSYS_UNCONNECTED_372,
  SYNOPSYS_UNCONNECTED_373,SYNOPSYS_UNCONNECTED_374,SYNOPSYS_UNCONNECTED_375,
  SYNOPSYS_UNCONNECTED_376,SYNOPSYS_UNCONNECTED_377,SYNOPSYS_UNCONNECTED_378,
  SYNOPSYS_UNCONNECTED_379,SYNOPSYS_UNCONNECTED_380,SYNOPSYS_UNCONNECTED_381,
  SYNOPSYS_UNCONNECTED_382,SYNOPSYS_UNCONNECTED_383,SYNOPSYS_UNCONNECTED_384,SYNOPSYS_UNCONNECTED_385,
  SYNOPSYS_UNCONNECTED_386,SYNOPSYS_UNCONNECTED_387,SYNOPSYS_UNCONNECTED_388,
  SYNOPSYS_UNCONNECTED_389,SYNOPSYS_UNCONNECTED_390,SYNOPSYS_UNCONNECTED_391,
  SYNOPSYS_UNCONNECTED_392,SYNOPSYS_UNCONNECTED_393,SYNOPSYS_UNCONNECTED_394,
  SYNOPSYS_UNCONNECTED_395,SYNOPSYS_UNCONNECTED_396,SYNOPSYS_UNCONNECTED_397,
  SYNOPSYS_UNCONNECTED_398,SYNOPSYS_UNCONNECTED_399,SYNOPSYS_UNCONNECTED_400,SYNOPSYS_UNCONNECTED_401,
  SYNOPSYS_UNCONNECTED_402,SYNOPSYS_UNCONNECTED_403,SYNOPSYS_UNCONNECTED_404,
  SYNOPSYS_UNCONNECTED_405,SYNOPSYS_UNCONNECTED_406,SYNOPSYS_UNCONNECTED_407,
  SYNOPSYS_UNCONNECTED_408,SYNOPSYS_UNCONNECTED_409,SYNOPSYS_UNCONNECTED_410,
  SYNOPSYS_UNCONNECTED_411,SYNOPSYS_UNCONNECTED_412,SYNOPSYS_UNCONNECTED_413,
  SYNOPSYS_UNCONNECTED_414,SYNOPSYS_UNCONNECTED_415,SYNOPSYS_UNCONNECTED_416,SYNOPSYS_UNCONNECTED_417,
  SYNOPSYS_UNCONNECTED_418,SYNOPSYS_UNCONNECTED_419,SYNOPSYS_UNCONNECTED_420,
  SYNOPSYS_UNCONNECTED_421,SYNOPSYS_UNCONNECTED_422,SYNOPSYS_UNCONNECTED_423,
  SYNOPSYS_UNCONNECTED_424,SYNOPSYS_UNCONNECTED_425,SYNOPSYS_UNCONNECTED_426,
  SYNOPSYS_UNCONNECTED_427,SYNOPSYS_UNCONNECTED_428,SYNOPSYS_UNCONNECTED_429,
  SYNOPSYS_UNCONNECTED_430,SYNOPSYS_UNCONNECTED_431,SYNOPSYS_UNCONNECTED_432,SYNOPSYS_UNCONNECTED_433,
  SYNOPSYS_UNCONNECTED_434,SYNOPSYS_UNCONNECTED_435,SYNOPSYS_UNCONNECTED_436,
  SYNOPSYS_UNCONNECTED_437,SYNOPSYS_UNCONNECTED_438,SYNOPSYS_UNCONNECTED_439,
  SYNOPSYS_UNCONNECTED_440,SYNOPSYS_UNCONNECTED_441,SYNOPSYS_UNCONNECTED_442,
  SYNOPSYS_UNCONNECTED_443,SYNOPSYS_UNCONNECTED_444,SYNOPSYS_UNCONNECTED_445,
  SYNOPSYS_UNCONNECTED_446,SYNOPSYS_UNCONNECTED_447,SYNOPSYS_UNCONNECTED_448,SYNOPSYS_UNCONNECTED_449,
  SYNOPSYS_UNCONNECTED_450,SYNOPSYS_UNCONNECTED_451,SYNOPSYS_UNCONNECTED_452,
  SYNOPSYS_UNCONNECTED_453,SYNOPSYS_UNCONNECTED_454,SYNOPSYS_UNCONNECTED_455,
  SYNOPSYS_UNCONNECTED_456,SYNOPSYS_UNCONNECTED_457,SYNOPSYS_UNCONNECTED_458,
  SYNOPSYS_UNCONNECTED_459,SYNOPSYS_UNCONNECTED_460,SYNOPSYS_UNCONNECTED_461,
  SYNOPSYS_UNCONNECTED_462,SYNOPSYS_UNCONNECTED_463,SYNOPSYS_UNCONNECTED_464,SYNOPSYS_UNCONNECTED_465,
  SYNOPSYS_UNCONNECTED_466,SYNOPSYS_UNCONNECTED_467,SYNOPSYS_UNCONNECTED_468,
  SYNOPSYS_UNCONNECTED_469,SYNOPSYS_UNCONNECTED_470,SYNOPSYS_UNCONNECTED_471,
  SYNOPSYS_UNCONNECTED_472,SYNOPSYS_UNCONNECTED_473,SYNOPSYS_UNCONNECTED_474,
  SYNOPSYS_UNCONNECTED_475,SYNOPSYS_UNCONNECTED_476,SYNOPSYS_UNCONNECTED_477,
  SYNOPSYS_UNCONNECTED_478,SYNOPSYS_UNCONNECTED_479,SYNOPSYS_UNCONNECTED_480,SYNOPSYS_UNCONNECTED_481,
  SYNOPSYS_UNCONNECTED_482,SYNOPSYS_UNCONNECTED_483,SYNOPSYS_UNCONNECTED_484,
  SYNOPSYS_UNCONNECTED_485,SYNOPSYS_UNCONNECTED_486,SYNOPSYS_UNCONNECTED_487,
  SYNOPSYS_UNCONNECTED_488,SYNOPSYS_UNCONNECTED_489,SYNOPSYS_UNCONNECTED_490,
  SYNOPSYS_UNCONNECTED_491,SYNOPSYS_UNCONNECTED_492,SYNOPSYS_UNCONNECTED_493,
  SYNOPSYS_UNCONNECTED_494,SYNOPSYS_UNCONNECTED_495,SYNOPSYS_UNCONNECTED_496,SYNOPSYS_UNCONNECTED_497,
  SYNOPSYS_UNCONNECTED_498,SYNOPSYS_UNCONNECTED_499,SYNOPSYS_UNCONNECTED_500,
  SYNOPSYS_UNCONNECTED_501,SYNOPSYS_UNCONNECTED_502,SYNOPSYS_UNCONNECTED_503,
  SYNOPSYS_UNCONNECTED_504,SYNOPSYS_UNCONNECTED_505,SYNOPSYS_UNCONNECTED_506,
  SYNOPSYS_UNCONNECTED_507,SYNOPSYS_UNCONNECTED_508,SYNOPSYS_UNCONNECTED_509,
  SYNOPSYS_UNCONNECTED_510,SYNOPSYS_UNCONNECTED_511,SYNOPSYS_UNCONNECTED_512,SYNOPSYS_UNCONNECTED_513,
  SYNOPSYS_UNCONNECTED_514,SYNOPSYS_UNCONNECTED_515,SYNOPSYS_UNCONNECTED_516,
  SYNOPSYS_UNCONNECTED_517,SYNOPSYS_UNCONNECTED_518,SYNOPSYS_UNCONNECTED_519,
  SYNOPSYS_UNCONNECTED_520,SYNOPSYS_UNCONNECTED_521,SYNOPSYS_UNCONNECTED_522,
  SYNOPSYS_UNCONNECTED_523,SYNOPSYS_UNCONNECTED_524,SYNOPSYS_UNCONNECTED_525,
  SYNOPSYS_UNCONNECTED_526,SYNOPSYS_UNCONNECTED_527,SYNOPSYS_UNCONNECTED_528,SYNOPSYS_UNCONNECTED_529,
  SYNOPSYS_UNCONNECTED_530,SYNOPSYS_UNCONNECTED_531,SYNOPSYS_UNCONNECTED_532,
  SYNOPSYS_UNCONNECTED_533,SYNOPSYS_UNCONNECTED_534,SYNOPSYS_UNCONNECTED_535,
  SYNOPSYS_UNCONNECTED_536,SYNOPSYS_UNCONNECTED_537,SYNOPSYS_UNCONNECTED_538,
  SYNOPSYS_UNCONNECTED_539,SYNOPSYS_UNCONNECTED_540,SYNOPSYS_UNCONNECTED_541,
  SYNOPSYS_UNCONNECTED_542,SYNOPSYS_UNCONNECTED_543,SYNOPSYS_UNCONNECTED_544,SYNOPSYS_UNCONNECTED_545,
  SYNOPSYS_UNCONNECTED_546,SYNOPSYS_UNCONNECTED_547,SYNOPSYS_UNCONNECTED_548,
  SYNOPSYS_UNCONNECTED_549,SYNOPSYS_UNCONNECTED_550,SYNOPSYS_UNCONNECTED_551,
  SYNOPSYS_UNCONNECTED_552,SYNOPSYS_UNCONNECTED_553,SYNOPSYS_UNCONNECTED_554,
  SYNOPSYS_UNCONNECTED_555,SYNOPSYS_UNCONNECTED_556,SYNOPSYS_UNCONNECTED_557,
  SYNOPSYS_UNCONNECTED_558,SYNOPSYS_UNCONNECTED_559,SYNOPSYS_UNCONNECTED_560,SYNOPSYS_UNCONNECTED_561,
  SYNOPSYS_UNCONNECTED_562,SYNOPSYS_UNCONNECTED_563,SYNOPSYS_UNCONNECTED_564,
  SYNOPSYS_UNCONNECTED_565,SYNOPSYS_UNCONNECTED_566,SYNOPSYS_UNCONNECTED_567,
  SYNOPSYS_UNCONNECTED_568,SYNOPSYS_UNCONNECTED_569,SYNOPSYS_UNCONNECTED_570,
  SYNOPSYS_UNCONNECTED_571,SYNOPSYS_UNCONNECTED_572,SYNOPSYS_UNCONNECTED_573,
  SYNOPSYS_UNCONNECTED_574,SYNOPSYS_UNCONNECTED_575,SYNOPSYS_UNCONNECTED_576,SYNOPSYS_UNCONNECTED_577,
  SYNOPSYS_UNCONNECTED_578,SYNOPSYS_UNCONNECTED_579,SYNOPSYS_UNCONNECTED_580,
  SYNOPSYS_UNCONNECTED_581,SYNOPSYS_UNCONNECTED_582,SYNOPSYS_UNCONNECTED_583,
  SYNOPSYS_UNCONNECTED_584,SYNOPSYS_UNCONNECTED_585,SYNOPSYS_UNCONNECTED_586,
  SYNOPSYS_UNCONNECTED_587,SYNOPSYS_UNCONNECTED_588,SYNOPSYS_UNCONNECTED_589,
  SYNOPSYS_UNCONNECTED_590,SYNOPSYS_UNCONNECTED_591,SYNOPSYS_UNCONNECTED_592,SYNOPSYS_UNCONNECTED_593,
  SYNOPSYS_UNCONNECTED_594,SYNOPSYS_UNCONNECTED_595,SYNOPSYS_UNCONNECTED_596,
  SYNOPSYS_UNCONNECTED_597,SYNOPSYS_UNCONNECTED_598,SYNOPSYS_UNCONNECTED_599,
  SYNOPSYS_UNCONNECTED_600,SYNOPSYS_UNCONNECTED_601,SYNOPSYS_UNCONNECTED_602,
  SYNOPSYS_UNCONNECTED_603,SYNOPSYS_UNCONNECTED_604,SYNOPSYS_UNCONNECTED_605,
  SYNOPSYS_UNCONNECTED_606,SYNOPSYS_UNCONNECTED_607,SYNOPSYS_UNCONNECTED_608,SYNOPSYS_UNCONNECTED_609,
  SYNOPSYS_UNCONNECTED_610,SYNOPSYS_UNCONNECTED_611,SYNOPSYS_UNCONNECTED_612,
  SYNOPSYS_UNCONNECTED_613,SYNOPSYS_UNCONNECTED_614,SYNOPSYS_UNCONNECTED_615,
  SYNOPSYS_UNCONNECTED_616,SYNOPSYS_UNCONNECTED_617,SYNOPSYS_UNCONNECTED_618,
  SYNOPSYS_UNCONNECTED_619,SYNOPSYS_UNCONNECTED_620,SYNOPSYS_UNCONNECTED_621,
  SYNOPSYS_UNCONNECTED_622,SYNOPSYS_UNCONNECTED_623,SYNOPSYS_UNCONNECTED_624,SYNOPSYS_UNCONNECTED_625,
  SYNOPSYS_UNCONNECTED_626,SYNOPSYS_UNCONNECTED_627,SYNOPSYS_UNCONNECTED_628,
  SYNOPSYS_UNCONNECTED_629,SYNOPSYS_UNCONNECTED_630,SYNOPSYS_UNCONNECTED_631,
  SYNOPSYS_UNCONNECTED_632,SYNOPSYS_UNCONNECTED_633,SYNOPSYS_UNCONNECTED_634,
  SYNOPSYS_UNCONNECTED_635,SYNOPSYS_UNCONNECTED_636,SYNOPSYS_UNCONNECTED_637,
  SYNOPSYS_UNCONNECTED_638,SYNOPSYS_UNCONNECTED_639,SYNOPSYS_UNCONNECTED_640,SYNOPSYS_UNCONNECTED_641,
  SYNOPSYS_UNCONNECTED_642,SYNOPSYS_UNCONNECTED_643,SYNOPSYS_UNCONNECTED_644,
  SYNOPSYS_UNCONNECTED_645,SYNOPSYS_UNCONNECTED_646,SYNOPSYS_UNCONNECTED_647,
  SYNOPSYS_UNCONNECTED_648,SYNOPSYS_UNCONNECTED_649,SYNOPSYS_UNCONNECTED_650,
  SYNOPSYS_UNCONNECTED_651,SYNOPSYS_UNCONNECTED_652,SYNOPSYS_UNCONNECTED_653,
  SYNOPSYS_UNCONNECTED_654,SYNOPSYS_UNCONNECTED_655,SYNOPSYS_UNCONNECTED_656,SYNOPSYS_UNCONNECTED_657,
  SYNOPSYS_UNCONNECTED_658,SYNOPSYS_UNCONNECTED_659,SYNOPSYS_UNCONNECTED_660,
  SYNOPSYS_UNCONNECTED_661,SYNOPSYS_UNCONNECTED_662,SYNOPSYS_UNCONNECTED_663,
  SYNOPSYS_UNCONNECTED_664,SYNOPSYS_UNCONNECTED_665,SYNOPSYS_UNCONNECTED_666,
  SYNOPSYS_UNCONNECTED_667,SYNOPSYS_UNCONNECTED_668,SYNOPSYS_UNCONNECTED_669,
  SYNOPSYS_UNCONNECTED_670,SYNOPSYS_UNCONNECTED_671,SYNOPSYS_UNCONNECTED_672,SYNOPSYS_UNCONNECTED_673,
  SYNOPSYS_UNCONNECTED_674,SYNOPSYS_UNCONNECTED_675,SYNOPSYS_UNCONNECTED_676,
  SYNOPSYS_UNCONNECTED_677,SYNOPSYS_UNCONNECTED_678,SYNOPSYS_UNCONNECTED_679,
  SYNOPSYS_UNCONNECTED_680,SYNOPSYS_UNCONNECTED_681,SYNOPSYS_UNCONNECTED_682,
  SYNOPSYS_UNCONNECTED_683,SYNOPSYS_UNCONNECTED_684,SYNOPSYS_UNCONNECTED_685,
  SYNOPSYS_UNCONNECTED_686,SYNOPSYS_UNCONNECTED_687,SYNOPSYS_UNCONNECTED_688,SYNOPSYS_UNCONNECTED_689,
  SYNOPSYS_UNCONNECTED_690,SYNOPSYS_UNCONNECTED_691,SYNOPSYS_UNCONNECTED_692,
  SYNOPSYS_UNCONNECTED_693,SYNOPSYS_UNCONNECTED_694,SYNOPSYS_UNCONNECTED_695,
  SYNOPSYS_UNCONNECTED_696,SYNOPSYS_UNCONNECTED_697,SYNOPSYS_UNCONNECTED_698,
  SYNOPSYS_UNCONNECTED_699,SYNOPSYS_UNCONNECTED_700,SYNOPSYS_UNCONNECTED_701,
  SYNOPSYS_UNCONNECTED_702,SYNOPSYS_UNCONNECTED_703,SYNOPSYS_UNCONNECTED_704,SYNOPSYS_UNCONNECTED_705,
  SYNOPSYS_UNCONNECTED_706,SYNOPSYS_UNCONNECTED_707,SYNOPSYS_UNCONNECTED_708,
  SYNOPSYS_UNCONNECTED_709,SYNOPSYS_UNCONNECTED_710,SYNOPSYS_UNCONNECTED_711,
  SYNOPSYS_UNCONNECTED_712,SYNOPSYS_UNCONNECTED_713,SYNOPSYS_UNCONNECTED_714,
  SYNOPSYS_UNCONNECTED_715,SYNOPSYS_UNCONNECTED_716,SYNOPSYS_UNCONNECTED_717,
  SYNOPSYS_UNCONNECTED_718,SYNOPSYS_UNCONNECTED_719,SYNOPSYS_UNCONNECTED_720,SYNOPSYS_UNCONNECTED_721,
  SYNOPSYS_UNCONNECTED_722,SYNOPSYS_UNCONNECTED_723,SYNOPSYS_UNCONNECTED_724,
  SYNOPSYS_UNCONNECTED_725,SYNOPSYS_UNCONNECTED_726,SYNOPSYS_UNCONNECTED_727,
  SYNOPSYS_UNCONNECTED_728,SYNOPSYS_UNCONNECTED_729,SYNOPSYS_UNCONNECTED_730,
  SYNOPSYS_UNCONNECTED_731,SYNOPSYS_UNCONNECTED_732,SYNOPSYS_UNCONNECTED_733,
  SYNOPSYS_UNCONNECTED_734,SYNOPSYS_UNCONNECTED_735,SYNOPSYS_UNCONNECTED_736,SYNOPSYS_UNCONNECTED_737,
  SYNOPSYS_UNCONNECTED_738,SYNOPSYS_UNCONNECTED_739,SYNOPSYS_UNCONNECTED_740,
  SYNOPSYS_UNCONNECTED_741,SYNOPSYS_UNCONNECTED_742,SYNOPSYS_UNCONNECTED_743,
  SYNOPSYS_UNCONNECTED_744,SYNOPSYS_UNCONNECTED_745,SYNOPSYS_UNCONNECTED_746,
  SYNOPSYS_UNCONNECTED_747,SYNOPSYS_UNCONNECTED_748,SYNOPSYS_UNCONNECTED_749,
  SYNOPSYS_UNCONNECTED_750,SYNOPSYS_UNCONNECTED_751,SYNOPSYS_UNCONNECTED_752,SYNOPSYS_UNCONNECTED_753,
  SYNOPSYS_UNCONNECTED_754,SYNOPSYS_UNCONNECTED_755,SYNOPSYS_UNCONNECTED_756,
  SYNOPSYS_UNCONNECTED_757,SYNOPSYS_UNCONNECTED_758,SYNOPSYS_UNCONNECTED_759,
  SYNOPSYS_UNCONNECTED_760,SYNOPSYS_UNCONNECTED_761,SYNOPSYS_UNCONNECTED_762,
  SYNOPSYS_UNCONNECTED_763,SYNOPSYS_UNCONNECTED_764,SYNOPSYS_UNCONNECTED_765,
  SYNOPSYS_UNCONNECTED_766,SYNOPSYS_UNCONNECTED_767,SYNOPSYS_UNCONNECTED_768,SYNOPSYS_UNCONNECTED_769,
  SYNOPSYS_UNCONNECTED_770,SYNOPSYS_UNCONNECTED_771,SYNOPSYS_UNCONNECTED_772,
  SYNOPSYS_UNCONNECTED_773,SYNOPSYS_UNCONNECTED_774,SYNOPSYS_UNCONNECTED_775,
  SYNOPSYS_UNCONNECTED_776,SYNOPSYS_UNCONNECTED_777,SYNOPSYS_UNCONNECTED_778,
  SYNOPSYS_UNCONNECTED_779,SYNOPSYS_UNCONNECTED_780,SYNOPSYS_UNCONNECTED_781,
  SYNOPSYS_UNCONNECTED_782,SYNOPSYS_UNCONNECTED_783,SYNOPSYS_UNCONNECTED_784,SYNOPSYS_UNCONNECTED_785,
  SYNOPSYS_UNCONNECTED_786,SYNOPSYS_UNCONNECTED_787,SYNOPSYS_UNCONNECTED_788,
  SYNOPSYS_UNCONNECTED_789,SYNOPSYS_UNCONNECTED_790,SYNOPSYS_UNCONNECTED_791,
  SYNOPSYS_UNCONNECTED_792,SYNOPSYS_UNCONNECTED_793,SYNOPSYS_UNCONNECTED_794,
  SYNOPSYS_UNCONNECTED_795,SYNOPSYS_UNCONNECTED_796,SYNOPSYS_UNCONNECTED_797,
  SYNOPSYS_UNCONNECTED_798,SYNOPSYS_UNCONNECTED_799,SYNOPSYS_UNCONNECTED_800,SYNOPSYS_UNCONNECTED_801,
  SYNOPSYS_UNCONNECTED_802,SYNOPSYS_UNCONNECTED_803,SYNOPSYS_UNCONNECTED_804,
  SYNOPSYS_UNCONNECTED_805,SYNOPSYS_UNCONNECTED_806,SYNOPSYS_UNCONNECTED_807,
  SYNOPSYS_UNCONNECTED_808,SYNOPSYS_UNCONNECTED_809,SYNOPSYS_UNCONNECTED_810,
  SYNOPSYS_UNCONNECTED_811,SYNOPSYS_UNCONNECTED_812,SYNOPSYS_UNCONNECTED_813,
  SYNOPSYS_UNCONNECTED_814,SYNOPSYS_UNCONNECTED_815,SYNOPSYS_UNCONNECTED_816,SYNOPSYS_UNCONNECTED_817,
  SYNOPSYS_UNCONNECTED_818,SYNOPSYS_UNCONNECTED_819,SYNOPSYS_UNCONNECTED_820,
  SYNOPSYS_UNCONNECTED_821,SYNOPSYS_UNCONNECTED_822,SYNOPSYS_UNCONNECTED_823,
  SYNOPSYS_UNCONNECTED_824,SYNOPSYS_UNCONNECTED_825,SYNOPSYS_UNCONNECTED_826,
  SYNOPSYS_UNCONNECTED_827,SYNOPSYS_UNCONNECTED_828,SYNOPSYS_UNCONNECTED_829,
  SYNOPSYS_UNCONNECTED_830,SYNOPSYS_UNCONNECTED_831,SYNOPSYS_UNCONNECTED_832,SYNOPSYS_UNCONNECTED_833,
  SYNOPSYS_UNCONNECTED_834,SYNOPSYS_UNCONNECTED_835,SYNOPSYS_UNCONNECTED_836,
  SYNOPSYS_UNCONNECTED_837,SYNOPSYS_UNCONNECTED_838,SYNOPSYS_UNCONNECTED_839,
  SYNOPSYS_UNCONNECTED_840,SYNOPSYS_UNCONNECTED_841,SYNOPSYS_UNCONNECTED_842,
  SYNOPSYS_UNCONNECTED_843,SYNOPSYS_UNCONNECTED_844,SYNOPSYS_UNCONNECTED_845,
  SYNOPSYS_UNCONNECTED_846,SYNOPSYS_UNCONNECTED_847,SYNOPSYS_UNCONNECTED_848,SYNOPSYS_UNCONNECTED_849,
  SYNOPSYS_UNCONNECTED_850,SYNOPSYS_UNCONNECTED_851,SYNOPSYS_UNCONNECTED_852,
  SYNOPSYS_UNCONNECTED_853,SYNOPSYS_UNCONNECTED_854,SYNOPSYS_UNCONNECTED_855,
  SYNOPSYS_UNCONNECTED_856,SYNOPSYS_UNCONNECTED_857,SYNOPSYS_UNCONNECTED_858,
  SYNOPSYS_UNCONNECTED_859,SYNOPSYS_UNCONNECTED_860,SYNOPSYS_UNCONNECTED_861,
  SYNOPSYS_UNCONNECTED_862,SYNOPSYS_UNCONNECTED_863,SYNOPSYS_UNCONNECTED_864,SYNOPSYS_UNCONNECTED_865,
  SYNOPSYS_UNCONNECTED_866,SYNOPSYS_UNCONNECTED_867,SYNOPSYS_UNCONNECTED_868,
  SYNOPSYS_UNCONNECTED_869,SYNOPSYS_UNCONNECTED_870,SYNOPSYS_UNCONNECTED_871,
  SYNOPSYS_UNCONNECTED_872,SYNOPSYS_UNCONNECTED_873,SYNOPSYS_UNCONNECTED_874,
  SYNOPSYS_UNCONNECTED_875,SYNOPSYS_UNCONNECTED_876,SYNOPSYS_UNCONNECTED_877,
  SYNOPSYS_UNCONNECTED_878,SYNOPSYS_UNCONNECTED_879,SYNOPSYS_UNCONNECTED_880,SYNOPSYS_UNCONNECTED_881,
  SYNOPSYS_UNCONNECTED_882,SYNOPSYS_UNCONNECTED_883,SYNOPSYS_UNCONNECTED_884,
  SYNOPSYS_UNCONNECTED_885,SYNOPSYS_UNCONNECTED_886,SYNOPSYS_UNCONNECTED_887,
  SYNOPSYS_UNCONNECTED_888,SYNOPSYS_UNCONNECTED_889,SYNOPSYS_UNCONNECTED_890,
  SYNOPSYS_UNCONNECTED_891,SYNOPSYS_UNCONNECTED_892,SYNOPSYS_UNCONNECTED_893,
  SYNOPSYS_UNCONNECTED_894,SYNOPSYS_UNCONNECTED_895,SYNOPSYS_UNCONNECTED_896,SYNOPSYS_UNCONNECTED_897,
  SYNOPSYS_UNCONNECTED_898,SYNOPSYS_UNCONNECTED_899,SYNOPSYS_UNCONNECTED_900,
  SYNOPSYS_UNCONNECTED_901,SYNOPSYS_UNCONNECTED_902,SYNOPSYS_UNCONNECTED_903,
  SYNOPSYS_UNCONNECTED_904,SYNOPSYS_UNCONNECTED_905,SYNOPSYS_UNCONNECTED_906,
  SYNOPSYS_UNCONNECTED_907,SYNOPSYS_UNCONNECTED_908,SYNOPSYS_UNCONNECTED_909,
  SYNOPSYS_UNCONNECTED_910,SYNOPSYS_UNCONNECTED_911,SYNOPSYS_UNCONNECTED_912,SYNOPSYS_UNCONNECTED_913,
  SYNOPSYS_UNCONNECTED_914,SYNOPSYS_UNCONNECTED_915,SYNOPSYS_UNCONNECTED_916,
  SYNOPSYS_UNCONNECTED_917,SYNOPSYS_UNCONNECTED_918,SYNOPSYS_UNCONNECTED_919,
  SYNOPSYS_UNCONNECTED_920,SYNOPSYS_UNCONNECTED_921,SYNOPSYS_UNCONNECTED_922,
  SYNOPSYS_UNCONNECTED_923,SYNOPSYS_UNCONNECTED_924,SYNOPSYS_UNCONNECTED_925,
  SYNOPSYS_UNCONNECTED_926,SYNOPSYS_UNCONNECTED_927,SYNOPSYS_UNCONNECTED_928,SYNOPSYS_UNCONNECTED_929,
  SYNOPSYS_UNCONNECTED_930,SYNOPSYS_UNCONNECTED_931,SYNOPSYS_UNCONNECTED_932,
  SYNOPSYS_UNCONNECTED_933,SYNOPSYS_UNCONNECTED_934,SYNOPSYS_UNCONNECTED_935,
  SYNOPSYS_UNCONNECTED_936,SYNOPSYS_UNCONNECTED_937,SYNOPSYS_UNCONNECTED_938,
  SYNOPSYS_UNCONNECTED_939,SYNOPSYS_UNCONNECTED_940,SYNOPSYS_UNCONNECTED_941,
  SYNOPSYS_UNCONNECTED_942,SYNOPSYS_UNCONNECTED_943,SYNOPSYS_UNCONNECTED_944,SYNOPSYS_UNCONNECTED_945,
  SYNOPSYS_UNCONNECTED_946,SYNOPSYS_UNCONNECTED_947,SYNOPSYS_UNCONNECTED_948,
  SYNOPSYS_UNCONNECTED_949,SYNOPSYS_UNCONNECTED_950,SYNOPSYS_UNCONNECTED_951,
  SYNOPSYS_UNCONNECTED_952,SYNOPSYS_UNCONNECTED_953,SYNOPSYS_UNCONNECTED_954,
  SYNOPSYS_UNCONNECTED_955,SYNOPSYS_UNCONNECTED_956,SYNOPSYS_UNCONNECTED_957,
  SYNOPSYS_UNCONNECTED_958,SYNOPSYS_UNCONNECTED_959,SYNOPSYS_UNCONNECTED_960,SYNOPSYS_UNCONNECTED_961,
  SYNOPSYS_UNCONNECTED_962,SYNOPSYS_UNCONNECTED_963,SYNOPSYS_UNCONNECTED_964,
  SYNOPSYS_UNCONNECTED_965,SYNOPSYS_UNCONNECTED_966,SYNOPSYS_UNCONNECTED_967,
  SYNOPSYS_UNCONNECTED_968,SYNOPSYS_UNCONNECTED_969,SYNOPSYS_UNCONNECTED_970,
  SYNOPSYS_UNCONNECTED_971,SYNOPSYS_UNCONNECTED_972,SYNOPSYS_UNCONNECTED_973,
  SYNOPSYS_UNCONNECTED_974,SYNOPSYS_UNCONNECTED_975,SYNOPSYS_UNCONNECTED_976,SYNOPSYS_UNCONNECTED_977,
  SYNOPSYS_UNCONNECTED_978,SYNOPSYS_UNCONNECTED_979,SYNOPSYS_UNCONNECTED_980,
  SYNOPSYS_UNCONNECTED_981,SYNOPSYS_UNCONNECTED_982,SYNOPSYS_UNCONNECTED_983,
  SYNOPSYS_UNCONNECTED_984,SYNOPSYS_UNCONNECTED_985,SYNOPSYS_UNCONNECTED_986,
  SYNOPSYS_UNCONNECTED_987,SYNOPSYS_UNCONNECTED_988,SYNOPSYS_UNCONNECTED_989,
  SYNOPSYS_UNCONNECTED_990,SYNOPSYS_UNCONNECTED_991,SYNOPSYS_UNCONNECTED_992,SYNOPSYS_UNCONNECTED_993,
  SYNOPSYS_UNCONNECTED_994,SYNOPSYS_UNCONNECTED_995,SYNOPSYS_UNCONNECTED_996,
  SYNOPSYS_UNCONNECTED_997,SYNOPSYS_UNCONNECTED_998,SYNOPSYS_UNCONNECTED_999,
  SYNOPSYS_UNCONNECTED_1000,SYNOPSYS_UNCONNECTED_1001,SYNOPSYS_UNCONNECTED_1002,
  SYNOPSYS_UNCONNECTED_1003,SYNOPSYS_UNCONNECTED_1004,SYNOPSYS_UNCONNECTED_1005,
  SYNOPSYS_UNCONNECTED_1006,SYNOPSYS_UNCONNECTED_1007,SYNOPSYS_UNCONNECTED_1008,
  SYNOPSYS_UNCONNECTED_1009,SYNOPSYS_UNCONNECTED_1010,SYNOPSYS_UNCONNECTED_1011,
  SYNOPSYS_UNCONNECTED_1012,SYNOPSYS_UNCONNECTED_1013,SYNOPSYS_UNCONNECTED_1014,
  SYNOPSYS_UNCONNECTED_1015,SYNOPSYS_UNCONNECTED_1016,SYNOPSYS_UNCONNECTED_1017,
  SYNOPSYS_UNCONNECTED_1018,SYNOPSYS_UNCONNECTED_1019,SYNOPSYS_UNCONNECTED_1020,SYNOPSYS_UNCONNECTED_1021,
  SYNOPSYS_UNCONNECTED_1022,SYNOPSYS_UNCONNECTED_1023,SYNOPSYS_UNCONNECTED_1024,
  SYNOPSYS_UNCONNECTED_1025,SYNOPSYS_UNCONNECTED_1026,SYNOPSYS_UNCONNECTED_1027,
  SYNOPSYS_UNCONNECTED_1028,SYNOPSYS_UNCONNECTED_1029,SYNOPSYS_UNCONNECTED_1030,
  SYNOPSYS_UNCONNECTED_1031,SYNOPSYS_UNCONNECTED_1032,SYNOPSYS_UNCONNECTED_1033,
  SYNOPSYS_UNCONNECTED_1034,SYNOPSYS_UNCONNECTED_1035,SYNOPSYS_UNCONNECTED_1036,
  SYNOPSYS_UNCONNECTED_1037,SYNOPSYS_UNCONNECTED_1038,SYNOPSYS_UNCONNECTED_1039,
  SYNOPSYS_UNCONNECTED_1040,SYNOPSYS_UNCONNECTED_1041,SYNOPSYS_UNCONNECTED_1042,
  SYNOPSYS_UNCONNECTED_1043,SYNOPSYS_UNCONNECTED_1044,SYNOPSYS_UNCONNECTED_1045,
  SYNOPSYS_UNCONNECTED_1046,SYNOPSYS_UNCONNECTED_1047,SYNOPSYS_UNCONNECTED_1048,
  SYNOPSYS_UNCONNECTED_1049,SYNOPSYS_UNCONNECTED_1050,SYNOPSYS_UNCONNECTED_1051,
  SYNOPSYS_UNCONNECTED_1052,SYNOPSYS_UNCONNECTED_1053,SYNOPSYS_UNCONNECTED_1054,
  SYNOPSYS_UNCONNECTED_1055,SYNOPSYS_UNCONNECTED_1056,SYNOPSYS_UNCONNECTED_1057,
  SYNOPSYS_UNCONNECTED_1058,SYNOPSYS_UNCONNECTED_1059,SYNOPSYS_UNCONNECTED_1060,SYNOPSYS_UNCONNECTED_1061,
  SYNOPSYS_UNCONNECTED_1062,SYNOPSYS_UNCONNECTED_1063,SYNOPSYS_UNCONNECTED_1064,
  SYNOPSYS_UNCONNECTED_1065,SYNOPSYS_UNCONNECTED_1066,SYNOPSYS_UNCONNECTED_1067,
  SYNOPSYS_UNCONNECTED_1068,SYNOPSYS_UNCONNECTED_1069,SYNOPSYS_UNCONNECTED_1070,
  SYNOPSYS_UNCONNECTED_1071,SYNOPSYS_UNCONNECTED_1072,SYNOPSYS_UNCONNECTED_1073,
  SYNOPSYS_UNCONNECTED_1074,SYNOPSYS_UNCONNECTED_1075,SYNOPSYS_UNCONNECTED_1076,
  SYNOPSYS_UNCONNECTED_1077,SYNOPSYS_UNCONNECTED_1078,SYNOPSYS_UNCONNECTED_1079,
  SYNOPSYS_UNCONNECTED_1080,SYNOPSYS_UNCONNECTED_1081,SYNOPSYS_UNCONNECTED_1082,
  SYNOPSYS_UNCONNECTED_1083,SYNOPSYS_UNCONNECTED_1084,SYNOPSYS_UNCONNECTED_1085,
  SYNOPSYS_UNCONNECTED_1086,SYNOPSYS_UNCONNECTED_1087,SYNOPSYS_UNCONNECTED_1088,
  SYNOPSYS_UNCONNECTED_1089,SYNOPSYS_UNCONNECTED_1090,SYNOPSYS_UNCONNECTED_1091,
  SYNOPSYS_UNCONNECTED_1092,SYNOPSYS_UNCONNECTED_1093,SYNOPSYS_UNCONNECTED_1094,
  SYNOPSYS_UNCONNECTED_1095,SYNOPSYS_UNCONNECTED_1096,SYNOPSYS_UNCONNECTED_1097,
  SYNOPSYS_UNCONNECTED_1098,SYNOPSYS_UNCONNECTED_1099,SYNOPSYS_UNCONNECTED_1100,SYNOPSYS_UNCONNECTED_1101,
  SYNOPSYS_UNCONNECTED_1102,SYNOPSYS_UNCONNECTED_1103,SYNOPSYS_UNCONNECTED_1104,
  SYNOPSYS_UNCONNECTED_1105,SYNOPSYS_UNCONNECTED_1106,SYNOPSYS_UNCONNECTED_1107,
  SYNOPSYS_UNCONNECTED_1108,SYNOPSYS_UNCONNECTED_1109,SYNOPSYS_UNCONNECTED_1110,
  SYNOPSYS_UNCONNECTED_1111,SYNOPSYS_UNCONNECTED_1112,SYNOPSYS_UNCONNECTED_1113,
  SYNOPSYS_UNCONNECTED_1114,SYNOPSYS_UNCONNECTED_1115,SYNOPSYS_UNCONNECTED_1116,
  SYNOPSYS_UNCONNECTED_1117,SYNOPSYS_UNCONNECTED_1118,SYNOPSYS_UNCONNECTED_1119,
  SYNOPSYS_UNCONNECTED_1120,SYNOPSYS_UNCONNECTED_1121,SYNOPSYS_UNCONNECTED_1122,
  SYNOPSYS_UNCONNECTED_1123,SYNOPSYS_UNCONNECTED_1124,SYNOPSYS_UNCONNECTED_1125,
  SYNOPSYS_UNCONNECTED_1126,SYNOPSYS_UNCONNECTED_1127,SYNOPSYS_UNCONNECTED_1128,
  SYNOPSYS_UNCONNECTED_1129,SYNOPSYS_UNCONNECTED_1130,SYNOPSYS_UNCONNECTED_1131,
  SYNOPSYS_UNCONNECTED_1132,SYNOPSYS_UNCONNECTED_1133,SYNOPSYS_UNCONNECTED_1134,
  SYNOPSYS_UNCONNECTED_1135,SYNOPSYS_UNCONNECTED_1136,SYNOPSYS_UNCONNECTED_1137,
  SYNOPSYS_UNCONNECTED_1138,SYNOPSYS_UNCONNECTED_1139,SYNOPSYS_UNCONNECTED_1140,SYNOPSYS_UNCONNECTED_1141,
  SYNOPSYS_UNCONNECTED_1142,SYNOPSYS_UNCONNECTED_1143,SYNOPSYS_UNCONNECTED_1144,
  SYNOPSYS_UNCONNECTED_1145,SYNOPSYS_UNCONNECTED_1146,SYNOPSYS_UNCONNECTED_1147,
  SYNOPSYS_UNCONNECTED_1148,SYNOPSYS_UNCONNECTED_1149,SYNOPSYS_UNCONNECTED_1150,
  SYNOPSYS_UNCONNECTED_1151,SYNOPSYS_UNCONNECTED_1152,SYNOPSYS_UNCONNECTED_1153,
  SYNOPSYS_UNCONNECTED_1154,SYNOPSYS_UNCONNECTED_1155,SYNOPSYS_UNCONNECTED_1156,
  SYNOPSYS_UNCONNECTED_1157,SYNOPSYS_UNCONNECTED_1158,SYNOPSYS_UNCONNECTED_1159,
  SYNOPSYS_UNCONNECTED_1160,SYNOPSYS_UNCONNECTED_1161,SYNOPSYS_UNCONNECTED_1162,
  SYNOPSYS_UNCONNECTED_1163,SYNOPSYS_UNCONNECTED_1164,SYNOPSYS_UNCONNECTED_1165,
  SYNOPSYS_UNCONNECTED_1166,SYNOPSYS_UNCONNECTED_1167,SYNOPSYS_UNCONNECTED_1168,
  SYNOPSYS_UNCONNECTED_1169,SYNOPSYS_UNCONNECTED_1170,SYNOPSYS_UNCONNECTED_1171,
  SYNOPSYS_UNCONNECTED_1172,SYNOPSYS_UNCONNECTED_1173,SYNOPSYS_UNCONNECTED_1174,
  SYNOPSYS_UNCONNECTED_1175,SYNOPSYS_UNCONNECTED_1176,SYNOPSYS_UNCONNECTED_1177,
  SYNOPSYS_UNCONNECTED_1178,SYNOPSYS_UNCONNECTED_1179,SYNOPSYS_UNCONNECTED_1180,SYNOPSYS_UNCONNECTED_1181,
  SYNOPSYS_UNCONNECTED_1182,SYNOPSYS_UNCONNECTED_1183,SYNOPSYS_UNCONNECTED_1184,
  SYNOPSYS_UNCONNECTED_1185,SYNOPSYS_UNCONNECTED_1186,SYNOPSYS_UNCONNECTED_1187,
  SYNOPSYS_UNCONNECTED_1188,SYNOPSYS_UNCONNECTED_1189,SYNOPSYS_UNCONNECTED_1190,
  SYNOPSYS_UNCONNECTED_1191,SYNOPSYS_UNCONNECTED_1192,SYNOPSYS_UNCONNECTED_1193,
  SYNOPSYS_UNCONNECTED_1194,SYNOPSYS_UNCONNECTED_1195,SYNOPSYS_UNCONNECTED_1196,
  SYNOPSYS_UNCONNECTED_1197,SYNOPSYS_UNCONNECTED_1198,SYNOPSYS_UNCONNECTED_1199,
  SYNOPSYS_UNCONNECTED_1200,SYNOPSYS_UNCONNECTED_1201,SYNOPSYS_UNCONNECTED_1202,
  SYNOPSYS_UNCONNECTED_1203,SYNOPSYS_UNCONNECTED_1204,SYNOPSYS_UNCONNECTED_1205,
  SYNOPSYS_UNCONNECTED_1206,SYNOPSYS_UNCONNECTED_1207,SYNOPSYS_UNCONNECTED_1208,
  SYNOPSYS_UNCONNECTED_1209,SYNOPSYS_UNCONNECTED_1210,SYNOPSYS_UNCONNECTED_1211,
  SYNOPSYS_UNCONNECTED_1212,SYNOPSYS_UNCONNECTED_1213,SYNOPSYS_UNCONNECTED_1214,
  SYNOPSYS_UNCONNECTED_1215,SYNOPSYS_UNCONNECTED_1216,SYNOPSYS_UNCONNECTED_1217,
  SYNOPSYS_UNCONNECTED_1218,SYNOPSYS_UNCONNECTED_1219,SYNOPSYS_UNCONNECTED_1220,SYNOPSYS_UNCONNECTED_1221,
  SYNOPSYS_UNCONNECTED_1222,SYNOPSYS_UNCONNECTED_1223,SYNOPSYS_UNCONNECTED_1224,
  SYNOPSYS_UNCONNECTED_1225,SYNOPSYS_UNCONNECTED_1226,SYNOPSYS_UNCONNECTED_1227,
  SYNOPSYS_UNCONNECTED_1228,SYNOPSYS_UNCONNECTED_1229,SYNOPSYS_UNCONNECTED_1230,
  SYNOPSYS_UNCONNECTED_1231,SYNOPSYS_UNCONNECTED_1232,SYNOPSYS_UNCONNECTED_1233,
  SYNOPSYS_UNCONNECTED_1234,SYNOPSYS_UNCONNECTED_1235,SYNOPSYS_UNCONNECTED_1236,
  SYNOPSYS_UNCONNECTED_1237,SYNOPSYS_UNCONNECTED_1238,SYNOPSYS_UNCONNECTED_1239,
  SYNOPSYS_UNCONNECTED_1240,SYNOPSYS_UNCONNECTED_1241,SYNOPSYS_UNCONNECTED_1242,
  SYNOPSYS_UNCONNECTED_1243,SYNOPSYS_UNCONNECTED_1244,SYNOPSYS_UNCONNECTED_1245,
  SYNOPSYS_UNCONNECTED_1246,SYNOPSYS_UNCONNECTED_1247,SYNOPSYS_UNCONNECTED_1248,
  SYNOPSYS_UNCONNECTED_1249,SYNOPSYS_UNCONNECTED_1250,SYNOPSYS_UNCONNECTED_1251,
  SYNOPSYS_UNCONNECTED_1252,SYNOPSYS_UNCONNECTED_1253,SYNOPSYS_UNCONNECTED_1254,
  SYNOPSYS_UNCONNECTED_1255,SYNOPSYS_UNCONNECTED_1256,SYNOPSYS_UNCONNECTED_1257,
  SYNOPSYS_UNCONNECTED_1258,SYNOPSYS_UNCONNECTED_1259,SYNOPSYS_UNCONNECTED_1260,SYNOPSYS_UNCONNECTED_1261,
  SYNOPSYS_UNCONNECTED_1262,SYNOPSYS_UNCONNECTED_1263,SYNOPSYS_UNCONNECTED_1264,
  SYNOPSYS_UNCONNECTED_1265,SYNOPSYS_UNCONNECTED_1266,SYNOPSYS_UNCONNECTED_1267,
  SYNOPSYS_UNCONNECTED_1268,SYNOPSYS_UNCONNECTED_1269,SYNOPSYS_UNCONNECTED_1270,
  SYNOPSYS_UNCONNECTED_1271,SYNOPSYS_UNCONNECTED_1272,SYNOPSYS_UNCONNECTED_1273,
  SYNOPSYS_UNCONNECTED_1274,SYNOPSYS_UNCONNECTED_1275,SYNOPSYS_UNCONNECTED_1276,
  SYNOPSYS_UNCONNECTED_1277,SYNOPSYS_UNCONNECTED_1278,SYNOPSYS_UNCONNECTED_1279,
  SYNOPSYS_UNCONNECTED_1280,SYNOPSYS_UNCONNECTED_1281,SYNOPSYS_UNCONNECTED_1282,
  SYNOPSYS_UNCONNECTED_1283,SYNOPSYS_UNCONNECTED_1284,SYNOPSYS_UNCONNECTED_1285,
  SYNOPSYS_UNCONNECTED_1286,SYNOPSYS_UNCONNECTED_1287,SYNOPSYS_UNCONNECTED_1288,
  SYNOPSYS_UNCONNECTED_1289,SYNOPSYS_UNCONNECTED_1290,SYNOPSYS_UNCONNECTED_1291,
  SYNOPSYS_UNCONNECTED_1292,SYNOPSYS_UNCONNECTED_1293,SYNOPSYS_UNCONNECTED_1294,
  SYNOPSYS_UNCONNECTED_1295,SYNOPSYS_UNCONNECTED_1296,SYNOPSYS_UNCONNECTED_1297,
  SYNOPSYS_UNCONNECTED_1298;
  wire [3:0] iptr_r,iptr_r_data;

  bsg_make_2D_array_width_p128_items_p10
  bm2Da
  (
    .i(data_head_o_flat_pretrunc),
    .o(data_head_o)
  );


  bsg_rotate_right_width_p10
  valid_rr
  (
    .data_i(valid_i),
    .rot_i(iptr_r),
    .o(valid_head_o)
  );

  assign { SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18, SYNOPSYS_UNCONNECTED_19, SYNOPSYS_UNCONNECTED_20, SYNOPSYS_UNCONNECTED_21, SYNOPSYS_UNCONNECTED_22, SYNOPSYS_UNCONNECTED_23, SYNOPSYS_UNCONNECTED_24, SYNOPSYS_UNCONNECTED_25, SYNOPSYS_UNCONNECTED_26, SYNOPSYS_UNCONNECTED_27, SYNOPSYS_UNCONNECTED_28, SYNOPSYS_UNCONNECTED_29, SYNOPSYS_UNCONNECTED_30, SYNOPSYS_UNCONNECTED_31, SYNOPSYS_UNCONNECTED_32, SYNOPSYS_UNCONNECTED_33, SYNOPSYS_UNCONNECTED_34, SYNOPSYS_UNCONNECTED_35, SYNOPSYS_UNCONNECTED_36, SYNOPSYS_UNCONNECTED_37, SYNOPSYS_UNCONNECTED_38, SYNOPSYS_UNCONNECTED_39, SYNOPSYS_UNCONNECTED_40, SYNOPSYS_UNCONNECTED_41, SYNOPSYS_UNCONNECTED_42, SYNOPSYS_UNCONNECTED_43, SYNOPSYS_UNCONNECTED_44, SYNOPSYS_UNCONNECTED_45, SYNOPSYS_UNCONNECTED_46, SYNOPSYS_UNCONNECTED_47, SYNOPSYS_UNCONNECTED_48, SYNOPSYS_UNCONNECTED_49, SYNOPSYS_UNCONNECTED_50, SYNOPSYS_UNCONNECTED_51, SYNOPSYS_UNCONNECTED_52, SYNOPSYS_UNCONNECTED_53, SYNOPSYS_UNCONNECTED_54, SYNOPSYS_UNCONNECTED_55, SYNOPSYS_UNCONNECTED_56, SYNOPSYS_UNCONNECTED_57, SYNOPSYS_UNCONNECTED_58, SYNOPSYS_UNCONNECTED_59, SYNOPSYS_UNCONNECTED_60, SYNOPSYS_UNCONNECTED_61, SYNOPSYS_UNCONNECTED_62, SYNOPSYS_UNCONNECTED_63, SYNOPSYS_UNCONNECTED_64, SYNOPSYS_UNCONNECTED_65, SYNOPSYS_UNCONNECTED_66, SYNOPSYS_UNCONNECTED_67, SYNOPSYS_UNCONNECTED_68, SYNOPSYS_UNCONNECTED_69, SYNOPSYS_UNCONNECTED_70, SYNOPSYS_UNCONNECTED_71, SYNOPSYS_UNCONNECTED_72, SYNOPSYS_UNCONNECTED_73, SYNOPSYS_UNCONNECTED_74, SYNOPSYS_UNCONNECTED_75, SYNOPSYS_UNCONNECTED_76, SYNOPSYS_UNCONNECTED_77, SYNOPSYS_UNCONNECTED_78, SYNOPSYS_UNCONNECTED_79, SYNOPSYS_UNCONNECTED_80, SYNOPSYS_UNCONNECTED_81, SYNOPSYS_UNCONNECTED_82, SYNOPSYS_UNCONNECTED_83, SYNOPSYS_UNCONNECTED_84, SYNOPSYS_UNCONNECTED_85, SYNOPSYS_UNCONNECTED_86, SYNOPSYS_UNCONNECTED_87, SYNOPSYS_UNCONNECTED_88, SYNOPSYS_UNCONNECTED_89, SYNOPSYS_UNCONNECTED_90, SYNOPSYS_UNCONNECTED_91, SYNOPSYS_UNCONNECTED_92, SYNOPSYS_UNCONNECTED_93, SYNOPSYS_UNCONNECTED_94, SYNOPSYS_UNCONNECTED_95, SYNOPSYS_UNCONNECTED_96, SYNOPSYS_UNCONNECTED_97, SYNOPSYS_UNCONNECTED_98, SYNOPSYS_UNCONNECTED_99, SYNOPSYS_UNCONNECTED_100, SYNOPSYS_UNCONNECTED_101, SYNOPSYS_UNCONNECTED_102, SYNOPSYS_UNCONNECTED_103, SYNOPSYS_UNCONNECTED_104, SYNOPSYS_UNCONNECTED_105, SYNOPSYS_UNCONNECTED_106, SYNOPSYS_UNCONNECTED_107, SYNOPSYS_UNCONNECTED_108, SYNOPSYS_UNCONNECTED_109, SYNOPSYS_UNCONNECTED_110, SYNOPSYS_UNCONNECTED_111, SYNOPSYS_UNCONNECTED_112, SYNOPSYS_UNCONNECTED_113, SYNOPSYS_UNCONNECTED_114, SYNOPSYS_UNCONNECTED_115, SYNOPSYS_UNCONNECTED_116, SYNOPSYS_UNCONNECTED_117, SYNOPSYS_UNCONNECTED_118, SYNOPSYS_UNCONNECTED_119, SYNOPSYS_UNCONNECTED_120, SYNOPSYS_UNCONNECTED_121, SYNOPSYS_UNCONNECTED_122, SYNOPSYS_UNCONNECTED_123, SYNOPSYS_UNCONNECTED_124, SYNOPSYS_UNCONNECTED_125, SYNOPSYS_UNCONNECTED_126, SYNOPSYS_UNCONNECTED_127, SYNOPSYS_UNCONNECTED_128, SYNOPSYS_UNCONNECTED_129, SYNOPSYS_UNCONNECTED_130, SYNOPSYS_UNCONNECTED_131, SYNOPSYS_UNCONNECTED_132, SYNOPSYS_UNCONNECTED_133, SYNOPSYS_UNCONNECTED_134, SYNOPSYS_UNCONNECTED_135, SYNOPSYS_UNCONNECTED_136, SYNOPSYS_UNCONNECTED_137, SYNOPSYS_UNCONNECTED_138, SYNOPSYS_UNCONNECTED_139, SYNOPSYS_UNCONNECTED_140, SYNOPSYS_UNCONNECTED_141, SYNOPSYS_UNCONNECTED_142, SYNOPSYS_UNCONNECTED_143, SYNOPSYS_UNCONNECTED_144, SYNOPSYS_UNCONNECTED_145, SYNOPSYS_UNCONNECTED_146, SYNOPSYS_UNCONNECTED_147, SYNOPSYS_UNCONNECTED_148, SYNOPSYS_UNCONNECTED_149, SYNOPSYS_UNCONNECTED_150, SYNOPSYS_UNCONNECTED_151, SYNOPSYS_UNCONNECTED_152, SYNOPSYS_UNCONNECTED_153, SYNOPSYS_UNCONNECTED_154, SYNOPSYS_UNCONNECTED_155, SYNOPSYS_UNCONNECTED_156, SYNOPSYS_UNCONNECTED_157, SYNOPSYS_UNCONNECTED_158, SYNOPSYS_UNCONNECTED_159, SYNOPSYS_UNCONNECTED_160, SYNOPSYS_UNCONNECTED_161, SYNOPSYS_UNCONNECTED_162, SYNOPSYS_UNCONNECTED_163, SYNOPSYS_UNCONNECTED_164, SYNOPSYS_UNCONNECTED_165, SYNOPSYS_UNCONNECTED_166, SYNOPSYS_UNCONNECTED_167, SYNOPSYS_UNCONNECTED_168, SYNOPSYS_UNCONNECTED_169, SYNOPSYS_UNCONNECTED_170, SYNOPSYS_UNCONNECTED_171, SYNOPSYS_UNCONNECTED_172, SYNOPSYS_UNCONNECTED_173, SYNOPSYS_UNCONNECTED_174, SYNOPSYS_UNCONNECTED_175, SYNOPSYS_UNCONNECTED_176, SYNOPSYS_UNCONNECTED_177, SYNOPSYS_UNCONNECTED_178, SYNOPSYS_UNCONNECTED_179, SYNOPSYS_UNCONNECTED_180, SYNOPSYS_UNCONNECTED_181, SYNOPSYS_UNCONNECTED_182, SYNOPSYS_UNCONNECTED_183, SYNOPSYS_UNCONNECTED_184, SYNOPSYS_UNCONNECTED_185, SYNOPSYS_UNCONNECTED_186, SYNOPSYS_UNCONNECTED_187, SYNOPSYS_UNCONNECTED_188, SYNOPSYS_UNCONNECTED_189, SYNOPSYS_UNCONNECTED_190, SYNOPSYS_UNCONNECTED_191, SYNOPSYS_UNCONNECTED_192, SYNOPSYS_UNCONNECTED_193, SYNOPSYS_UNCONNECTED_194, SYNOPSYS_UNCONNECTED_195, SYNOPSYS_UNCONNECTED_196, SYNOPSYS_UNCONNECTED_197, SYNOPSYS_UNCONNECTED_198, SYNOPSYS_UNCONNECTED_199, SYNOPSYS_UNCONNECTED_200, SYNOPSYS_UNCONNECTED_201, SYNOPSYS_UNCONNECTED_202, SYNOPSYS_UNCONNECTED_203, SYNOPSYS_UNCONNECTED_204, SYNOPSYS_UNCONNECTED_205, SYNOPSYS_UNCONNECTED_206, SYNOPSYS_UNCONNECTED_207, SYNOPSYS_UNCONNECTED_208, SYNOPSYS_UNCONNECTED_209, SYNOPSYS_UNCONNECTED_210, SYNOPSYS_UNCONNECTED_211, SYNOPSYS_UNCONNECTED_212, SYNOPSYS_UNCONNECTED_213, SYNOPSYS_UNCONNECTED_214, SYNOPSYS_UNCONNECTED_215, SYNOPSYS_UNCONNECTED_216, SYNOPSYS_UNCONNECTED_217, SYNOPSYS_UNCONNECTED_218, SYNOPSYS_UNCONNECTED_219, SYNOPSYS_UNCONNECTED_220, SYNOPSYS_UNCONNECTED_221, SYNOPSYS_UNCONNECTED_222, SYNOPSYS_UNCONNECTED_223, SYNOPSYS_UNCONNECTED_224, SYNOPSYS_UNCONNECTED_225, SYNOPSYS_UNCONNECTED_226, SYNOPSYS_UNCONNECTED_227, SYNOPSYS_UNCONNECTED_228, SYNOPSYS_UNCONNECTED_229, SYNOPSYS_UNCONNECTED_230, SYNOPSYS_UNCONNECTED_231, SYNOPSYS_UNCONNECTED_232, SYNOPSYS_UNCONNECTED_233, SYNOPSYS_UNCONNECTED_234, SYNOPSYS_UNCONNECTED_235, SYNOPSYS_UNCONNECTED_236, SYNOPSYS_UNCONNECTED_237, SYNOPSYS_UNCONNECTED_238, SYNOPSYS_UNCONNECTED_239, SYNOPSYS_UNCONNECTED_240, SYNOPSYS_UNCONNECTED_241, SYNOPSYS_UNCONNECTED_242, SYNOPSYS_UNCONNECTED_243, SYNOPSYS_UNCONNECTED_244, SYNOPSYS_UNCONNECTED_245, SYNOPSYS_UNCONNECTED_246, SYNOPSYS_UNCONNECTED_247, SYNOPSYS_UNCONNECTED_248, SYNOPSYS_UNCONNECTED_249, SYNOPSYS_UNCONNECTED_250, SYNOPSYS_UNCONNECTED_251, SYNOPSYS_UNCONNECTED_252, SYNOPSYS_UNCONNECTED_253, SYNOPSYS_UNCONNECTED_254, SYNOPSYS_UNCONNECTED_255, SYNOPSYS_UNCONNECTED_256, SYNOPSYS_UNCONNECTED_257, SYNOPSYS_UNCONNECTED_258, SYNOPSYS_UNCONNECTED_259, SYNOPSYS_UNCONNECTED_260, SYNOPSYS_UNCONNECTED_261, SYNOPSYS_UNCONNECTED_262, SYNOPSYS_UNCONNECTED_263, SYNOPSYS_UNCONNECTED_264, SYNOPSYS_UNCONNECTED_265, SYNOPSYS_UNCONNECTED_266, SYNOPSYS_UNCONNECTED_267, SYNOPSYS_UNCONNECTED_268, SYNOPSYS_UNCONNECTED_269, SYNOPSYS_UNCONNECTED_270, SYNOPSYS_UNCONNECTED_271, SYNOPSYS_UNCONNECTED_272, SYNOPSYS_UNCONNECTED_273, SYNOPSYS_UNCONNECTED_274, SYNOPSYS_UNCONNECTED_275, SYNOPSYS_UNCONNECTED_276, SYNOPSYS_UNCONNECTED_277, SYNOPSYS_UNCONNECTED_278, SYNOPSYS_UNCONNECTED_279, SYNOPSYS_UNCONNECTED_280, SYNOPSYS_UNCONNECTED_281, SYNOPSYS_UNCONNECTED_282, SYNOPSYS_UNCONNECTED_283, SYNOPSYS_UNCONNECTED_284, SYNOPSYS_UNCONNECTED_285, SYNOPSYS_UNCONNECTED_286, SYNOPSYS_UNCONNECTED_287, SYNOPSYS_UNCONNECTED_288, SYNOPSYS_UNCONNECTED_289, SYNOPSYS_UNCONNECTED_290, SYNOPSYS_UNCONNECTED_291, SYNOPSYS_UNCONNECTED_292, SYNOPSYS_UNCONNECTED_293, SYNOPSYS_UNCONNECTED_294, SYNOPSYS_UNCONNECTED_295, SYNOPSYS_UNCONNECTED_296, SYNOPSYS_UNCONNECTED_297, SYNOPSYS_UNCONNECTED_298, SYNOPSYS_UNCONNECTED_299, SYNOPSYS_UNCONNECTED_300, SYNOPSYS_UNCONNECTED_301, SYNOPSYS_UNCONNECTED_302, SYNOPSYS_UNCONNECTED_303, SYNOPSYS_UNCONNECTED_304, SYNOPSYS_UNCONNECTED_305, SYNOPSYS_UNCONNECTED_306, SYNOPSYS_UNCONNECTED_307, SYNOPSYS_UNCONNECTED_308, SYNOPSYS_UNCONNECTED_309, SYNOPSYS_UNCONNECTED_310, SYNOPSYS_UNCONNECTED_311, SYNOPSYS_UNCONNECTED_312, SYNOPSYS_UNCONNECTED_313, SYNOPSYS_UNCONNECTED_314, SYNOPSYS_UNCONNECTED_315, SYNOPSYS_UNCONNECTED_316, SYNOPSYS_UNCONNECTED_317, SYNOPSYS_UNCONNECTED_318, SYNOPSYS_UNCONNECTED_319, SYNOPSYS_UNCONNECTED_320, SYNOPSYS_UNCONNECTED_321, SYNOPSYS_UNCONNECTED_322, SYNOPSYS_UNCONNECTED_323, SYNOPSYS_UNCONNECTED_324, SYNOPSYS_UNCONNECTED_325, SYNOPSYS_UNCONNECTED_326, SYNOPSYS_UNCONNECTED_327, SYNOPSYS_UNCONNECTED_328, SYNOPSYS_UNCONNECTED_329, SYNOPSYS_UNCONNECTED_330, SYNOPSYS_UNCONNECTED_331, SYNOPSYS_UNCONNECTED_332, SYNOPSYS_UNCONNECTED_333, SYNOPSYS_UNCONNECTED_334, SYNOPSYS_UNCONNECTED_335, SYNOPSYS_UNCONNECTED_336, SYNOPSYS_UNCONNECTED_337, SYNOPSYS_UNCONNECTED_338, SYNOPSYS_UNCONNECTED_339, SYNOPSYS_UNCONNECTED_340, SYNOPSYS_UNCONNECTED_341, SYNOPSYS_UNCONNECTED_342, SYNOPSYS_UNCONNECTED_343, SYNOPSYS_UNCONNECTED_344, SYNOPSYS_UNCONNECTED_345, SYNOPSYS_UNCONNECTED_346, SYNOPSYS_UNCONNECTED_347, SYNOPSYS_UNCONNECTED_348, SYNOPSYS_UNCONNECTED_349, SYNOPSYS_UNCONNECTED_350, SYNOPSYS_UNCONNECTED_351, SYNOPSYS_UNCONNECTED_352, SYNOPSYS_UNCONNECTED_353, SYNOPSYS_UNCONNECTED_354, SYNOPSYS_UNCONNECTED_355, SYNOPSYS_UNCONNECTED_356, SYNOPSYS_UNCONNECTED_357, SYNOPSYS_UNCONNECTED_358, SYNOPSYS_UNCONNECTED_359, SYNOPSYS_UNCONNECTED_360, SYNOPSYS_UNCONNECTED_361, SYNOPSYS_UNCONNECTED_362, SYNOPSYS_UNCONNECTED_363, SYNOPSYS_UNCONNECTED_364, SYNOPSYS_UNCONNECTED_365, SYNOPSYS_UNCONNECTED_366, SYNOPSYS_UNCONNECTED_367, SYNOPSYS_UNCONNECTED_368, SYNOPSYS_UNCONNECTED_369, SYNOPSYS_UNCONNECTED_370, SYNOPSYS_UNCONNECTED_371, SYNOPSYS_UNCONNECTED_372, SYNOPSYS_UNCONNECTED_373, SYNOPSYS_UNCONNECTED_374, SYNOPSYS_UNCONNECTED_375, SYNOPSYS_UNCONNECTED_376, SYNOPSYS_UNCONNECTED_377, SYNOPSYS_UNCONNECTED_378, SYNOPSYS_UNCONNECTED_379, SYNOPSYS_UNCONNECTED_380, SYNOPSYS_UNCONNECTED_381, SYNOPSYS_UNCONNECTED_382, SYNOPSYS_UNCONNECTED_383, SYNOPSYS_UNCONNECTED_384, SYNOPSYS_UNCONNECTED_385, SYNOPSYS_UNCONNECTED_386, SYNOPSYS_UNCONNECTED_387, SYNOPSYS_UNCONNECTED_388, SYNOPSYS_UNCONNECTED_389, SYNOPSYS_UNCONNECTED_390, SYNOPSYS_UNCONNECTED_391, SYNOPSYS_UNCONNECTED_392, SYNOPSYS_UNCONNECTED_393, SYNOPSYS_UNCONNECTED_394, SYNOPSYS_UNCONNECTED_395, SYNOPSYS_UNCONNECTED_396, SYNOPSYS_UNCONNECTED_397, SYNOPSYS_UNCONNECTED_398, SYNOPSYS_UNCONNECTED_399, SYNOPSYS_UNCONNECTED_400, SYNOPSYS_UNCONNECTED_401, SYNOPSYS_UNCONNECTED_402, SYNOPSYS_UNCONNECTED_403, SYNOPSYS_UNCONNECTED_404, SYNOPSYS_UNCONNECTED_405, SYNOPSYS_UNCONNECTED_406, SYNOPSYS_UNCONNECTED_407, SYNOPSYS_UNCONNECTED_408, SYNOPSYS_UNCONNECTED_409, SYNOPSYS_UNCONNECTED_410, SYNOPSYS_UNCONNECTED_411, SYNOPSYS_UNCONNECTED_412, SYNOPSYS_UNCONNECTED_413, SYNOPSYS_UNCONNECTED_414, SYNOPSYS_UNCONNECTED_415, SYNOPSYS_UNCONNECTED_416, SYNOPSYS_UNCONNECTED_417, SYNOPSYS_UNCONNECTED_418, SYNOPSYS_UNCONNECTED_419, SYNOPSYS_UNCONNECTED_420, SYNOPSYS_UNCONNECTED_421, SYNOPSYS_UNCONNECTED_422, SYNOPSYS_UNCONNECTED_423, SYNOPSYS_UNCONNECTED_424, SYNOPSYS_UNCONNECTED_425, SYNOPSYS_UNCONNECTED_426, SYNOPSYS_UNCONNECTED_427, SYNOPSYS_UNCONNECTED_428, SYNOPSYS_UNCONNECTED_429, SYNOPSYS_UNCONNECTED_430, SYNOPSYS_UNCONNECTED_431, SYNOPSYS_UNCONNECTED_432, SYNOPSYS_UNCONNECTED_433, SYNOPSYS_UNCONNECTED_434, SYNOPSYS_UNCONNECTED_435, SYNOPSYS_UNCONNECTED_436, SYNOPSYS_UNCONNECTED_437, SYNOPSYS_UNCONNECTED_438, SYNOPSYS_UNCONNECTED_439, SYNOPSYS_UNCONNECTED_440, SYNOPSYS_UNCONNECTED_441, SYNOPSYS_UNCONNECTED_442, SYNOPSYS_UNCONNECTED_443, SYNOPSYS_UNCONNECTED_444, SYNOPSYS_UNCONNECTED_445, SYNOPSYS_UNCONNECTED_446, SYNOPSYS_UNCONNECTED_447, SYNOPSYS_UNCONNECTED_448, SYNOPSYS_UNCONNECTED_449, SYNOPSYS_UNCONNECTED_450, SYNOPSYS_UNCONNECTED_451, SYNOPSYS_UNCONNECTED_452, SYNOPSYS_UNCONNECTED_453, SYNOPSYS_UNCONNECTED_454, SYNOPSYS_UNCONNECTED_455, SYNOPSYS_UNCONNECTED_456, SYNOPSYS_UNCONNECTED_457, SYNOPSYS_UNCONNECTED_458, SYNOPSYS_UNCONNECTED_459, SYNOPSYS_UNCONNECTED_460, SYNOPSYS_UNCONNECTED_461, SYNOPSYS_UNCONNECTED_462, SYNOPSYS_UNCONNECTED_463, SYNOPSYS_UNCONNECTED_464, SYNOPSYS_UNCONNECTED_465, SYNOPSYS_UNCONNECTED_466, SYNOPSYS_UNCONNECTED_467, SYNOPSYS_UNCONNECTED_468, SYNOPSYS_UNCONNECTED_469, SYNOPSYS_UNCONNECTED_470, SYNOPSYS_UNCONNECTED_471, SYNOPSYS_UNCONNECTED_472, SYNOPSYS_UNCONNECTED_473, SYNOPSYS_UNCONNECTED_474, SYNOPSYS_UNCONNECTED_475, SYNOPSYS_UNCONNECTED_476, SYNOPSYS_UNCONNECTED_477, SYNOPSYS_UNCONNECTED_478, SYNOPSYS_UNCONNECTED_479, SYNOPSYS_UNCONNECTED_480, SYNOPSYS_UNCONNECTED_481, SYNOPSYS_UNCONNECTED_482, SYNOPSYS_UNCONNECTED_483, SYNOPSYS_UNCONNECTED_484, SYNOPSYS_UNCONNECTED_485, SYNOPSYS_UNCONNECTED_486, SYNOPSYS_UNCONNECTED_487, SYNOPSYS_UNCONNECTED_488, SYNOPSYS_UNCONNECTED_489, SYNOPSYS_UNCONNECTED_490, SYNOPSYS_UNCONNECTED_491, SYNOPSYS_UNCONNECTED_492, SYNOPSYS_UNCONNECTED_493, SYNOPSYS_UNCONNECTED_494, SYNOPSYS_UNCONNECTED_495, SYNOPSYS_UNCONNECTED_496, SYNOPSYS_UNCONNECTED_497, SYNOPSYS_UNCONNECTED_498, SYNOPSYS_UNCONNECTED_499, SYNOPSYS_UNCONNECTED_500, SYNOPSYS_UNCONNECTED_501, SYNOPSYS_UNCONNECTED_502, SYNOPSYS_UNCONNECTED_503, SYNOPSYS_UNCONNECTED_504, SYNOPSYS_UNCONNECTED_505, SYNOPSYS_UNCONNECTED_506, SYNOPSYS_UNCONNECTED_507, SYNOPSYS_UNCONNECTED_508, SYNOPSYS_UNCONNECTED_509, SYNOPSYS_UNCONNECTED_510, SYNOPSYS_UNCONNECTED_511, SYNOPSYS_UNCONNECTED_512, SYNOPSYS_UNCONNECTED_513, SYNOPSYS_UNCONNECTED_514, SYNOPSYS_UNCONNECTED_515, SYNOPSYS_UNCONNECTED_516, SYNOPSYS_UNCONNECTED_517, SYNOPSYS_UNCONNECTED_518, SYNOPSYS_UNCONNECTED_519, SYNOPSYS_UNCONNECTED_520, SYNOPSYS_UNCONNECTED_521, SYNOPSYS_UNCONNECTED_522, SYNOPSYS_UNCONNECTED_523, SYNOPSYS_UNCONNECTED_524, SYNOPSYS_UNCONNECTED_525, SYNOPSYS_UNCONNECTED_526, SYNOPSYS_UNCONNECTED_527, SYNOPSYS_UNCONNECTED_528, SYNOPSYS_UNCONNECTED_529, SYNOPSYS_UNCONNECTED_530, SYNOPSYS_UNCONNECTED_531, SYNOPSYS_UNCONNECTED_532, SYNOPSYS_UNCONNECTED_533, SYNOPSYS_UNCONNECTED_534, SYNOPSYS_UNCONNECTED_535, SYNOPSYS_UNCONNECTED_536, SYNOPSYS_UNCONNECTED_537, SYNOPSYS_UNCONNECTED_538, SYNOPSYS_UNCONNECTED_539, SYNOPSYS_UNCONNECTED_540, SYNOPSYS_UNCONNECTED_541, SYNOPSYS_UNCONNECTED_542, SYNOPSYS_UNCONNECTED_543, SYNOPSYS_UNCONNECTED_544, SYNOPSYS_UNCONNECTED_545, SYNOPSYS_UNCONNECTED_546, SYNOPSYS_UNCONNECTED_547, SYNOPSYS_UNCONNECTED_548, SYNOPSYS_UNCONNECTED_549, SYNOPSYS_UNCONNECTED_550, SYNOPSYS_UNCONNECTED_551, SYNOPSYS_UNCONNECTED_552, SYNOPSYS_UNCONNECTED_553, SYNOPSYS_UNCONNECTED_554, SYNOPSYS_UNCONNECTED_555, SYNOPSYS_UNCONNECTED_556, SYNOPSYS_UNCONNECTED_557, SYNOPSYS_UNCONNECTED_558, SYNOPSYS_UNCONNECTED_559, SYNOPSYS_UNCONNECTED_560, SYNOPSYS_UNCONNECTED_561, SYNOPSYS_UNCONNECTED_562, SYNOPSYS_UNCONNECTED_563, SYNOPSYS_UNCONNECTED_564, SYNOPSYS_UNCONNECTED_565, SYNOPSYS_UNCONNECTED_566, SYNOPSYS_UNCONNECTED_567, SYNOPSYS_UNCONNECTED_568, SYNOPSYS_UNCONNECTED_569, SYNOPSYS_UNCONNECTED_570, SYNOPSYS_UNCONNECTED_571, SYNOPSYS_UNCONNECTED_572, SYNOPSYS_UNCONNECTED_573, SYNOPSYS_UNCONNECTED_574, SYNOPSYS_UNCONNECTED_575, SYNOPSYS_UNCONNECTED_576, SYNOPSYS_UNCONNECTED_577, SYNOPSYS_UNCONNECTED_578, SYNOPSYS_UNCONNECTED_579, SYNOPSYS_UNCONNECTED_580, SYNOPSYS_UNCONNECTED_581, SYNOPSYS_UNCONNECTED_582, SYNOPSYS_UNCONNECTED_583, SYNOPSYS_UNCONNECTED_584, SYNOPSYS_UNCONNECTED_585, SYNOPSYS_UNCONNECTED_586, SYNOPSYS_UNCONNECTED_587, SYNOPSYS_UNCONNECTED_588, SYNOPSYS_UNCONNECTED_589, SYNOPSYS_UNCONNECTED_590, SYNOPSYS_UNCONNECTED_591, SYNOPSYS_UNCONNECTED_592, SYNOPSYS_UNCONNECTED_593, SYNOPSYS_UNCONNECTED_594, SYNOPSYS_UNCONNECTED_595, SYNOPSYS_UNCONNECTED_596, SYNOPSYS_UNCONNECTED_597, SYNOPSYS_UNCONNECTED_598, SYNOPSYS_UNCONNECTED_599, SYNOPSYS_UNCONNECTED_600, SYNOPSYS_UNCONNECTED_601, SYNOPSYS_UNCONNECTED_602, SYNOPSYS_UNCONNECTED_603, SYNOPSYS_UNCONNECTED_604, SYNOPSYS_UNCONNECTED_605, SYNOPSYS_UNCONNECTED_606, SYNOPSYS_UNCONNECTED_607, SYNOPSYS_UNCONNECTED_608, SYNOPSYS_UNCONNECTED_609, SYNOPSYS_UNCONNECTED_610, SYNOPSYS_UNCONNECTED_611, SYNOPSYS_UNCONNECTED_612, SYNOPSYS_UNCONNECTED_613, SYNOPSYS_UNCONNECTED_614, SYNOPSYS_UNCONNECTED_615, SYNOPSYS_UNCONNECTED_616, SYNOPSYS_UNCONNECTED_617, SYNOPSYS_UNCONNECTED_618, SYNOPSYS_UNCONNECTED_619, SYNOPSYS_UNCONNECTED_620, SYNOPSYS_UNCONNECTED_621, SYNOPSYS_UNCONNECTED_622, SYNOPSYS_UNCONNECTED_623, SYNOPSYS_UNCONNECTED_624, SYNOPSYS_UNCONNECTED_625, SYNOPSYS_UNCONNECTED_626, SYNOPSYS_UNCONNECTED_627, SYNOPSYS_UNCONNECTED_628, SYNOPSYS_UNCONNECTED_629, SYNOPSYS_UNCONNECTED_630, SYNOPSYS_UNCONNECTED_631, SYNOPSYS_UNCONNECTED_632, SYNOPSYS_UNCONNECTED_633, SYNOPSYS_UNCONNECTED_634, SYNOPSYS_UNCONNECTED_635, SYNOPSYS_UNCONNECTED_636, SYNOPSYS_UNCONNECTED_637, SYNOPSYS_UNCONNECTED_638, SYNOPSYS_UNCONNECTED_639, SYNOPSYS_UNCONNECTED_640, SYNOPSYS_UNCONNECTED_641, SYNOPSYS_UNCONNECTED_642, SYNOPSYS_UNCONNECTED_643, SYNOPSYS_UNCONNECTED_644, SYNOPSYS_UNCONNECTED_645, SYNOPSYS_UNCONNECTED_646, SYNOPSYS_UNCONNECTED_647, SYNOPSYS_UNCONNECTED_648, SYNOPSYS_UNCONNECTED_649, SYNOPSYS_UNCONNECTED_650, SYNOPSYS_UNCONNECTED_651, SYNOPSYS_UNCONNECTED_652, SYNOPSYS_UNCONNECTED_653, SYNOPSYS_UNCONNECTED_654, SYNOPSYS_UNCONNECTED_655, SYNOPSYS_UNCONNECTED_656, SYNOPSYS_UNCONNECTED_657, SYNOPSYS_UNCONNECTED_658, SYNOPSYS_UNCONNECTED_659, SYNOPSYS_UNCONNECTED_660, SYNOPSYS_UNCONNECTED_661, SYNOPSYS_UNCONNECTED_662, SYNOPSYS_UNCONNECTED_663, SYNOPSYS_UNCONNECTED_664, SYNOPSYS_UNCONNECTED_665, SYNOPSYS_UNCONNECTED_666, SYNOPSYS_UNCONNECTED_667, SYNOPSYS_UNCONNECTED_668, SYNOPSYS_UNCONNECTED_669, SYNOPSYS_UNCONNECTED_670, SYNOPSYS_UNCONNECTED_671, SYNOPSYS_UNCONNECTED_672, SYNOPSYS_UNCONNECTED_673, SYNOPSYS_UNCONNECTED_674, SYNOPSYS_UNCONNECTED_675, SYNOPSYS_UNCONNECTED_676, SYNOPSYS_UNCONNECTED_677, SYNOPSYS_UNCONNECTED_678, SYNOPSYS_UNCONNECTED_679, SYNOPSYS_UNCONNECTED_680, SYNOPSYS_UNCONNECTED_681, SYNOPSYS_UNCONNECTED_682, SYNOPSYS_UNCONNECTED_683, SYNOPSYS_UNCONNECTED_684, SYNOPSYS_UNCONNECTED_685, SYNOPSYS_UNCONNECTED_686, SYNOPSYS_UNCONNECTED_687, SYNOPSYS_UNCONNECTED_688, SYNOPSYS_UNCONNECTED_689, SYNOPSYS_UNCONNECTED_690, SYNOPSYS_UNCONNECTED_691, SYNOPSYS_UNCONNECTED_692, SYNOPSYS_UNCONNECTED_693, SYNOPSYS_UNCONNECTED_694, SYNOPSYS_UNCONNECTED_695, SYNOPSYS_UNCONNECTED_696, SYNOPSYS_UNCONNECTED_697, SYNOPSYS_UNCONNECTED_698, SYNOPSYS_UNCONNECTED_699, SYNOPSYS_UNCONNECTED_700, SYNOPSYS_UNCONNECTED_701, SYNOPSYS_UNCONNECTED_702, SYNOPSYS_UNCONNECTED_703, SYNOPSYS_UNCONNECTED_704, SYNOPSYS_UNCONNECTED_705, SYNOPSYS_UNCONNECTED_706, SYNOPSYS_UNCONNECTED_707, SYNOPSYS_UNCONNECTED_708, SYNOPSYS_UNCONNECTED_709, SYNOPSYS_UNCONNECTED_710, SYNOPSYS_UNCONNECTED_711, SYNOPSYS_UNCONNECTED_712, SYNOPSYS_UNCONNECTED_713, SYNOPSYS_UNCONNECTED_714, SYNOPSYS_UNCONNECTED_715, SYNOPSYS_UNCONNECTED_716, SYNOPSYS_UNCONNECTED_717, SYNOPSYS_UNCONNECTED_718, SYNOPSYS_UNCONNECTED_719, SYNOPSYS_UNCONNECTED_720, SYNOPSYS_UNCONNECTED_721, SYNOPSYS_UNCONNECTED_722, SYNOPSYS_UNCONNECTED_723, SYNOPSYS_UNCONNECTED_724, SYNOPSYS_UNCONNECTED_725, SYNOPSYS_UNCONNECTED_726, SYNOPSYS_UNCONNECTED_727, SYNOPSYS_UNCONNECTED_728, SYNOPSYS_UNCONNECTED_729, SYNOPSYS_UNCONNECTED_730, SYNOPSYS_UNCONNECTED_731, SYNOPSYS_UNCONNECTED_732, SYNOPSYS_UNCONNECTED_733, SYNOPSYS_UNCONNECTED_734, SYNOPSYS_UNCONNECTED_735, SYNOPSYS_UNCONNECTED_736, SYNOPSYS_UNCONNECTED_737, SYNOPSYS_UNCONNECTED_738, SYNOPSYS_UNCONNECTED_739, SYNOPSYS_UNCONNECTED_740, SYNOPSYS_UNCONNECTED_741, SYNOPSYS_UNCONNECTED_742, SYNOPSYS_UNCONNECTED_743, SYNOPSYS_UNCONNECTED_744, SYNOPSYS_UNCONNECTED_745, SYNOPSYS_UNCONNECTED_746, SYNOPSYS_UNCONNECTED_747, SYNOPSYS_UNCONNECTED_748, SYNOPSYS_UNCONNECTED_749, SYNOPSYS_UNCONNECTED_750, SYNOPSYS_UNCONNECTED_751, SYNOPSYS_UNCONNECTED_752, SYNOPSYS_UNCONNECTED_753, SYNOPSYS_UNCONNECTED_754, SYNOPSYS_UNCONNECTED_755, SYNOPSYS_UNCONNECTED_756, SYNOPSYS_UNCONNECTED_757, SYNOPSYS_UNCONNECTED_758, SYNOPSYS_UNCONNECTED_759, SYNOPSYS_UNCONNECTED_760, SYNOPSYS_UNCONNECTED_761, SYNOPSYS_UNCONNECTED_762, SYNOPSYS_UNCONNECTED_763, SYNOPSYS_UNCONNECTED_764, SYNOPSYS_UNCONNECTED_765, SYNOPSYS_UNCONNECTED_766, SYNOPSYS_UNCONNECTED_767, SYNOPSYS_UNCONNECTED_768, SYNOPSYS_UNCONNECTED_769, SYNOPSYS_UNCONNECTED_770, SYNOPSYS_UNCONNECTED_771, SYNOPSYS_UNCONNECTED_772, SYNOPSYS_UNCONNECTED_773, SYNOPSYS_UNCONNECTED_774, SYNOPSYS_UNCONNECTED_775, SYNOPSYS_UNCONNECTED_776, SYNOPSYS_UNCONNECTED_777, SYNOPSYS_UNCONNECTED_778, SYNOPSYS_UNCONNECTED_779, SYNOPSYS_UNCONNECTED_780, SYNOPSYS_UNCONNECTED_781, SYNOPSYS_UNCONNECTED_782, SYNOPSYS_UNCONNECTED_783, SYNOPSYS_UNCONNECTED_784, SYNOPSYS_UNCONNECTED_785, SYNOPSYS_UNCONNECTED_786, SYNOPSYS_UNCONNECTED_787, SYNOPSYS_UNCONNECTED_788, SYNOPSYS_UNCONNECTED_789, SYNOPSYS_UNCONNECTED_790, SYNOPSYS_UNCONNECTED_791, SYNOPSYS_UNCONNECTED_792, SYNOPSYS_UNCONNECTED_793, SYNOPSYS_UNCONNECTED_794, SYNOPSYS_UNCONNECTED_795, SYNOPSYS_UNCONNECTED_796, SYNOPSYS_UNCONNECTED_797, SYNOPSYS_UNCONNECTED_798, SYNOPSYS_UNCONNECTED_799, SYNOPSYS_UNCONNECTED_800, SYNOPSYS_UNCONNECTED_801, SYNOPSYS_UNCONNECTED_802, SYNOPSYS_UNCONNECTED_803, SYNOPSYS_UNCONNECTED_804, SYNOPSYS_UNCONNECTED_805, SYNOPSYS_UNCONNECTED_806, SYNOPSYS_UNCONNECTED_807, SYNOPSYS_UNCONNECTED_808, SYNOPSYS_UNCONNECTED_809, SYNOPSYS_UNCONNECTED_810, SYNOPSYS_UNCONNECTED_811, SYNOPSYS_UNCONNECTED_812, SYNOPSYS_UNCONNECTED_813, SYNOPSYS_UNCONNECTED_814, SYNOPSYS_UNCONNECTED_815, SYNOPSYS_UNCONNECTED_816, SYNOPSYS_UNCONNECTED_817, SYNOPSYS_UNCONNECTED_818, SYNOPSYS_UNCONNECTED_819, SYNOPSYS_UNCONNECTED_820, SYNOPSYS_UNCONNECTED_821, SYNOPSYS_UNCONNECTED_822, SYNOPSYS_UNCONNECTED_823, SYNOPSYS_UNCONNECTED_824, SYNOPSYS_UNCONNECTED_825, SYNOPSYS_UNCONNECTED_826, SYNOPSYS_UNCONNECTED_827, SYNOPSYS_UNCONNECTED_828, SYNOPSYS_UNCONNECTED_829, SYNOPSYS_UNCONNECTED_830, SYNOPSYS_UNCONNECTED_831, SYNOPSYS_UNCONNECTED_832, SYNOPSYS_UNCONNECTED_833, SYNOPSYS_UNCONNECTED_834, SYNOPSYS_UNCONNECTED_835, SYNOPSYS_UNCONNECTED_836, SYNOPSYS_UNCONNECTED_837, SYNOPSYS_UNCONNECTED_838, SYNOPSYS_UNCONNECTED_839, SYNOPSYS_UNCONNECTED_840, SYNOPSYS_UNCONNECTED_841, SYNOPSYS_UNCONNECTED_842, SYNOPSYS_UNCONNECTED_843, SYNOPSYS_UNCONNECTED_844, SYNOPSYS_UNCONNECTED_845, SYNOPSYS_UNCONNECTED_846, SYNOPSYS_UNCONNECTED_847, SYNOPSYS_UNCONNECTED_848, SYNOPSYS_UNCONNECTED_849, SYNOPSYS_UNCONNECTED_850, SYNOPSYS_UNCONNECTED_851, SYNOPSYS_UNCONNECTED_852, SYNOPSYS_UNCONNECTED_853, SYNOPSYS_UNCONNECTED_854, SYNOPSYS_UNCONNECTED_855, SYNOPSYS_UNCONNECTED_856, SYNOPSYS_UNCONNECTED_857, SYNOPSYS_UNCONNECTED_858, SYNOPSYS_UNCONNECTED_859, SYNOPSYS_UNCONNECTED_860, SYNOPSYS_UNCONNECTED_861, SYNOPSYS_UNCONNECTED_862, SYNOPSYS_UNCONNECTED_863, SYNOPSYS_UNCONNECTED_864, SYNOPSYS_UNCONNECTED_865, SYNOPSYS_UNCONNECTED_866, SYNOPSYS_UNCONNECTED_867, SYNOPSYS_UNCONNECTED_868, SYNOPSYS_UNCONNECTED_869, SYNOPSYS_UNCONNECTED_870, SYNOPSYS_UNCONNECTED_871, SYNOPSYS_UNCONNECTED_872, SYNOPSYS_UNCONNECTED_873, SYNOPSYS_UNCONNECTED_874, SYNOPSYS_UNCONNECTED_875, SYNOPSYS_UNCONNECTED_876, SYNOPSYS_UNCONNECTED_877, SYNOPSYS_UNCONNECTED_878, SYNOPSYS_UNCONNECTED_879, SYNOPSYS_UNCONNECTED_880, SYNOPSYS_UNCONNECTED_881, SYNOPSYS_UNCONNECTED_882, SYNOPSYS_UNCONNECTED_883, SYNOPSYS_UNCONNECTED_884, SYNOPSYS_UNCONNECTED_885, SYNOPSYS_UNCONNECTED_886, SYNOPSYS_UNCONNECTED_887, SYNOPSYS_UNCONNECTED_888, SYNOPSYS_UNCONNECTED_889, SYNOPSYS_UNCONNECTED_890, SYNOPSYS_UNCONNECTED_891, SYNOPSYS_UNCONNECTED_892, SYNOPSYS_UNCONNECTED_893, SYNOPSYS_UNCONNECTED_894, SYNOPSYS_UNCONNECTED_895, SYNOPSYS_UNCONNECTED_896, SYNOPSYS_UNCONNECTED_897, SYNOPSYS_UNCONNECTED_898, SYNOPSYS_UNCONNECTED_899, SYNOPSYS_UNCONNECTED_900, SYNOPSYS_UNCONNECTED_901, SYNOPSYS_UNCONNECTED_902, SYNOPSYS_UNCONNECTED_903, SYNOPSYS_UNCONNECTED_904, SYNOPSYS_UNCONNECTED_905, SYNOPSYS_UNCONNECTED_906, SYNOPSYS_UNCONNECTED_907, SYNOPSYS_UNCONNECTED_908, SYNOPSYS_UNCONNECTED_909, SYNOPSYS_UNCONNECTED_910, SYNOPSYS_UNCONNECTED_911, SYNOPSYS_UNCONNECTED_912, SYNOPSYS_UNCONNECTED_913, SYNOPSYS_UNCONNECTED_914, SYNOPSYS_UNCONNECTED_915, SYNOPSYS_UNCONNECTED_916, SYNOPSYS_UNCONNECTED_917, SYNOPSYS_UNCONNECTED_918, SYNOPSYS_UNCONNECTED_919, SYNOPSYS_UNCONNECTED_920, SYNOPSYS_UNCONNECTED_921, SYNOPSYS_UNCONNECTED_922, SYNOPSYS_UNCONNECTED_923, SYNOPSYS_UNCONNECTED_924, SYNOPSYS_UNCONNECTED_925, SYNOPSYS_UNCONNECTED_926, SYNOPSYS_UNCONNECTED_927, SYNOPSYS_UNCONNECTED_928, SYNOPSYS_UNCONNECTED_929, SYNOPSYS_UNCONNECTED_930, SYNOPSYS_UNCONNECTED_931, SYNOPSYS_UNCONNECTED_932, SYNOPSYS_UNCONNECTED_933, SYNOPSYS_UNCONNECTED_934, SYNOPSYS_UNCONNECTED_935, SYNOPSYS_UNCONNECTED_936, SYNOPSYS_UNCONNECTED_937, SYNOPSYS_UNCONNECTED_938, SYNOPSYS_UNCONNECTED_939, SYNOPSYS_UNCONNECTED_940, SYNOPSYS_UNCONNECTED_941, SYNOPSYS_UNCONNECTED_942, SYNOPSYS_UNCONNECTED_943, SYNOPSYS_UNCONNECTED_944, SYNOPSYS_UNCONNECTED_945, SYNOPSYS_UNCONNECTED_946, SYNOPSYS_UNCONNECTED_947, SYNOPSYS_UNCONNECTED_948, SYNOPSYS_UNCONNECTED_949, SYNOPSYS_UNCONNECTED_950, SYNOPSYS_UNCONNECTED_951, SYNOPSYS_UNCONNECTED_952, SYNOPSYS_UNCONNECTED_953, SYNOPSYS_UNCONNECTED_954, SYNOPSYS_UNCONNECTED_955, SYNOPSYS_UNCONNECTED_956, SYNOPSYS_UNCONNECTED_957, SYNOPSYS_UNCONNECTED_958, SYNOPSYS_UNCONNECTED_959, SYNOPSYS_UNCONNECTED_960, SYNOPSYS_UNCONNECTED_961, SYNOPSYS_UNCONNECTED_962, SYNOPSYS_UNCONNECTED_963, SYNOPSYS_UNCONNECTED_964, SYNOPSYS_UNCONNECTED_965, SYNOPSYS_UNCONNECTED_966, SYNOPSYS_UNCONNECTED_967, SYNOPSYS_UNCONNECTED_968, SYNOPSYS_UNCONNECTED_969, SYNOPSYS_UNCONNECTED_970, SYNOPSYS_UNCONNECTED_971, SYNOPSYS_UNCONNECTED_972, SYNOPSYS_UNCONNECTED_973, SYNOPSYS_UNCONNECTED_974, SYNOPSYS_UNCONNECTED_975, SYNOPSYS_UNCONNECTED_976, SYNOPSYS_UNCONNECTED_977, SYNOPSYS_UNCONNECTED_978, SYNOPSYS_UNCONNECTED_979, SYNOPSYS_UNCONNECTED_980, SYNOPSYS_UNCONNECTED_981, SYNOPSYS_UNCONNECTED_982, SYNOPSYS_UNCONNECTED_983, SYNOPSYS_UNCONNECTED_984, SYNOPSYS_UNCONNECTED_985, SYNOPSYS_UNCONNECTED_986, SYNOPSYS_UNCONNECTED_987, SYNOPSYS_UNCONNECTED_988, SYNOPSYS_UNCONNECTED_989, SYNOPSYS_UNCONNECTED_990, SYNOPSYS_UNCONNECTED_991, SYNOPSYS_UNCONNECTED_992, SYNOPSYS_UNCONNECTED_993, SYNOPSYS_UNCONNECTED_994, SYNOPSYS_UNCONNECTED_995, SYNOPSYS_UNCONNECTED_996, SYNOPSYS_UNCONNECTED_997, SYNOPSYS_UNCONNECTED_998, SYNOPSYS_UNCONNECTED_999, SYNOPSYS_UNCONNECTED_1000, SYNOPSYS_UNCONNECTED_1001, SYNOPSYS_UNCONNECTED_1002, SYNOPSYS_UNCONNECTED_1003, SYNOPSYS_UNCONNECTED_1004, SYNOPSYS_UNCONNECTED_1005, SYNOPSYS_UNCONNECTED_1006, SYNOPSYS_UNCONNECTED_1007, SYNOPSYS_UNCONNECTED_1008, SYNOPSYS_UNCONNECTED_1009, SYNOPSYS_UNCONNECTED_1010, SYNOPSYS_UNCONNECTED_1011, SYNOPSYS_UNCONNECTED_1012, SYNOPSYS_UNCONNECTED_1013, SYNOPSYS_UNCONNECTED_1014, SYNOPSYS_UNCONNECTED_1015, SYNOPSYS_UNCONNECTED_1016, SYNOPSYS_UNCONNECTED_1017, SYNOPSYS_UNCONNECTED_1018, SYNOPSYS_UNCONNECTED_1019, SYNOPSYS_UNCONNECTED_1020, SYNOPSYS_UNCONNECTED_1021, SYNOPSYS_UNCONNECTED_1022, SYNOPSYS_UNCONNECTED_1023, SYNOPSYS_UNCONNECTED_1024, SYNOPSYS_UNCONNECTED_1025, SYNOPSYS_UNCONNECTED_1026, SYNOPSYS_UNCONNECTED_1027, SYNOPSYS_UNCONNECTED_1028, SYNOPSYS_UNCONNECTED_1029, SYNOPSYS_UNCONNECTED_1030, SYNOPSYS_UNCONNECTED_1031, SYNOPSYS_UNCONNECTED_1032, SYNOPSYS_UNCONNECTED_1033, SYNOPSYS_UNCONNECTED_1034, SYNOPSYS_UNCONNECTED_1035, SYNOPSYS_UNCONNECTED_1036, SYNOPSYS_UNCONNECTED_1037, SYNOPSYS_UNCONNECTED_1038, SYNOPSYS_UNCONNECTED_1039, SYNOPSYS_UNCONNECTED_1040, SYNOPSYS_UNCONNECTED_1041, SYNOPSYS_UNCONNECTED_1042, SYNOPSYS_UNCONNECTED_1043, SYNOPSYS_UNCONNECTED_1044, SYNOPSYS_UNCONNECTED_1045, SYNOPSYS_UNCONNECTED_1046, SYNOPSYS_UNCONNECTED_1047, SYNOPSYS_UNCONNECTED_1048, SYNOPSYS_UNCONNECTED_1049, SYNOPSYS_UNCONNECTED_1050, SYNOPSYS_UNCONNECTED_1051, SYNOPSYS_UNCONNECTED_1052, SYNOPSYS_UNCONNECTED_1053, SYNOPSYS_UNCONNECTED_1054, SYNOPSYS_UNCONNECTED_1055, SYNOPSYS_UNCONNECTED_1056, SYNOPSYS_UNCONNECTED_1057, SYNOPSYS_UNCONNECTED_1058, SYNOPSYS_UNCONNECTED_1059, SYNOPSYS_UNCONNECTED_1060, SYNOPSYS_UNCONNECTED_1061, SYNOPSYS_UNCONNECTED_1062, SYNOPSYS_UNCONNECTED_1063, SYNOPSYS_UNCONNECTED_1064, SYNOPSYS_UNCONNECTED_1065, SYNOPSYS_UNCONNECTED_1066, SYNOPSYS_UNCONNECTED_1067, SYNOPSYS_UNCONNECTED_1068, SYNOPSYS_UNCONNECTED_1069, SYNOPSYS_UNCONNECTED_1070, SYNOPSYS_UNCONNECTED_1071, SYNOPSYS_UNCONNECTED_1072, SYNOPSYS_UNCONNECTED_1073, SYNOPSYS_UNCONNECTED_1074, SYNOPSYS_UNCONNECTED_1075, SYNOPSYS_UNCONNECTED_1076, SYNOPSYS_UNCONNECTED_1077, SYNOPSYS_UNCONNECTED_1078, SYNOPSYS_UNCONNECTED_1079, SYNOPSYS_UNCONNECTED_1080, SYNOPSYS_UNCONNECTED_1081, SYNOPSYS_UNCONNECTED_1082, SYNOPSYS_UNCONNECTED_1083, SYNOPSYS_UNCONNECTED_1084, SYNOPSYS_UNCONNECTED_1085, SYNOPSYS_UNCONNECTED_1086, SYNOPSYS_UNCONNECTED_1087, SYNOPSYS_UNCONNECTED_1088, SYNOPSYS_UNCONNECTED_1089, SYNOPSYS_UNCONNECTED_1090, SYNOPSYS_UNCONNECTED_1091, SYNOPSYS_UNCONNECTED_1092, SYNOPSYS_UNCONNECTED_1093, SYNOPSYS_UNCONNECTED_1094, SYNOPSYS_UNCONNECTED_1095, SYNOPSYS_UNCONNECTED_1096, SYNOPSYS_UNCONNECTED_1097, SYNOPSYS_UNCONNECTED_1098, SYNOPSYS_UNCONNECTED_1099, SYNOPSYS_UNCONNECTED_1100, SYNOPSYS_UNCONNECTED_1101, SYNOPSYS_UNCONNECTED_1102, SYNOPSYS_UNCONNECTED_1103, SYNOPSYS_UNCONNECTED_1104, SYNOPSYS_UNCONNECTED_1105, SYNOPSYS_UNCONNECTED_1106, SYNOPSYS_UNCONNECTED_1107, SYNOPSYS_UNCONNECTED_1108, SYNOPSYS_UNCONNECTED_1109, SYNOPSYS_UNCONNECTED_1110, SYNOPSYS_UNCONNECTED_1111, SYNOPSYS_UNCONNECTED_1112, SYNOPSYS_UNCONNECTED_1113, SYNOPSYS_UNCONNECTED_1114, SYNOPSYS_UNCONNECTED_1115, SYNOPSYS_UNCONNECTED_1116, SYNOPSYS_UNCONNECTED_1117, SYNOPSYS_UNCONNECTED_1118, SYNOPSYS_UNCONNECTED_1119, SYNOPSYS_UNCONNECTED_1120, SYNOPSYS_UNCONNECTED_1121, SYNOPSYS_UNCONNECTED_1122, SYNOPSYS_UNCONNECTED_1123, SYNOPSYS_UNCONNECTED_1124, SYNOPSYS_UNCONNECTED_1125, SYNOPSYS_UNCONNECTED_1126, SYNOPSYS_UNCONNECTED_1127, SYNOPSYS_UNCONNECTED_1128, SYNOPSYS_UNCONNECTED_1129, SYNOPSYS_UNCONNECTED_1130, SYNOPSYS_UNCONNECTED_1131, SYNOPSYS_UNCONNECTED_1132, SYNOPSYS_UNCONNECTED_1133, SYNOPSYS_UNCONNECTED_1134, SYNOPSYS_UNCONNECTED_1135, SYNOPSYS_UNCONNECTED_1136, SYNOPSYS_UNCONNECTED_1137, SYNOPSYS_UNCONNECTED_1138, SYNOPSYS_UNCONNECTED_1139, SYNOPSYS_UNCONNECTED_1140, SYNOPSYS_UNCONNECTED_1141, SYNOPSYS_UNCONNECTED_1142, SYNOPSYS_UNCONNECTED_1143, SYNOPSYS_UNCONNECTED_1144, SYNOPSYS_UNCONNECTED_1145, SYNOPSYS_UNCONNECTED_1146, SYNOPSYS_UNCONNECTED_1147, SYNOPSYS_UNCONNECTED_1148, SYNOPSYS_UNCONNECTED_1149, SYNOPSYS_UNCONNECTED_1150, SYNOPSYS_UNCONNECTED_1151, SYNOPSYS_UNCONNECTED_1152, SYNOPSYS_UNCONNECTED_1153, SYNOPSYS_UNCONNECTED_1154, SYNOPSYS_UNCONNECTED_1155, SYNOPSYS_UNCONNECTED_1156, SYNOPSYS_UNCONNECTED_1157, SYNOPSYS_UNCONNECTED_1158, SYNOPSYS_UNCONNECTED_1159, SYNOPSYS_UNCONNECTED_1160, SYNOPSYS_UNCONNECTED_1161, SYNOPSYS_UNCONNECTED_1162, SYNOPSYS_UNCONNECTED_1163, SYNOPSYS_UNCONNECTED_1164, SYNOPSYS_UNCONNECTED_1165, SYNOPSYS_UNCONNECTED_1166, SYNOPSYS_UNCONNECTED_1167, SYNOPSYS_UNCONNECTED_1168, SYNOPSYS_UNCONNECTED_1169, SYNOPSYS_UNCONNECTED_1170, SYNOPSYS_UNCONNECTED_1171, SYNOPSYS_UNCONNECTED_1172, SYNOPSYS_UNCONNECTED_1173, SYNOPSYS_UNCONNECTED_1174, SYNOPSYS_UNCONNECTED_1175, SYNOPSYS_UNCONNECTED_1176, SYNOPSYS_UNCONNECTED_1177, SYNOPSYS_UNCONNECTED_1178, SYNOPSYS_UNCONNECTED_1179, SYNOPSYS_UNCONNECTED_1180, SYNOPSYS_UNCONNECTED_1181, SYNOPSYS_UNCONNECTED_1182, SYNOPSYS_UNCONNECTED_1183, SYNOPSYS_UNCONNECTED_1184, SYNOPSYS_UNCONNECTED_1185, SYNOPSYS_UNCONNECTED_1186, SYNOPSYS_UNCONNECTED_1187, SYNOPSYS_UNCONNECTED_1188, SYNOPSYS_UNCONNECTED_1189, SYNOPSYS_UNCONNECTED_1190, SYNOPSYS_UNCONNECTED_1191, SYNOPSYS_UNCONNECTED_1192, SYNOPSYS_UNCONNECTED_1193, SYNOPSYS_UNCONNECTED_1194, SYNOPSYS_UNCONNECTED_1195, SYNOPSYS_UNCONNECTED_1196, SYNOPSYS_UNCONNECTED_1197, SYNOPSYS_UNCONNECTED_1198, SYNOPSYS_UNCONNECTED_1199, SYNOPSYS_UNCONNECTED_1200, SYNOPSYS_UNCONNECTED_1201, SYNOPSYS_UNCONNECTED_1202, SYNOPSYS_UNCONNECTED_1203, SYNOPSYS_UNCONNECTED_1204, SYNOPSYS_UNCONNECTED_1205, SYNOPSYS_UNCONNECTED_1206, SYNOPSYS_UNCONNECTED_1207, SYNOPSYS_UNCONNECTED_1208, SYNOPSYS_UNCONNECTED_1209, SYNOPSYS_UNCONNECTED_1210, SYNOPSYS_UNCONNECTED_1211, SYNOPSYS_UNCONNECTED_1212, SYNOPSYS_UNCONNECTED_1213, SYNOPSYS_UNCONNECTED_1214, SYNOPSYS_UNCONNECTED_1215, SYNOPSYS_UNCONNECTED_1216, SYNOPSYS_UNCONNECTED_1217, SYNOPSYS_UNCONNECTED_1218, SYNOPSYS_UNCONNECTED_1219, SYNOPSYS_UNCONNECTED_1220, SYNOPSYS_UNCONNECTED_1221, SYNOPSYS_UNCONNECTED_1222, SYNOPSYS_UNCONNECTED_1223, SYNOPSYS_UNCONNECTED_1224, SYNOPSYS_UNCONNECTED_1225, SYNOPSYS_UNCONNECTED_1226, SYNOPSYS_UNCONNECTED_1227, SYNOPSYS_UNCONNECTED_1228, SYNOPSYS_UNCONNECTED_1229, SYNOPSYS_UNCONNECTED_1230, SYNOPSYS_UNCONNECTED_1231, SYNOPSYS_UNCONNECTED_1232, SYNOPSYS_UNCONNECTED_1233, SYNOPSYS_UNCONNECTED_1234, SYNOPSYS_UNCONNECTED_1235, SYNOPSYS_UNCONNECTED_1236, SYNOPSYS_UNCONNECTED_1237, SYNOPSYS_UNCONNECTED_1238, SYNOPSYS_UNCONNECTED_1239, SYNOPSYS_UNCONNECTED_1240, SYNOPSYS_UNCONNECTED_1241, SYNOPSYS_UNCONNECTED_1242, SYNOPSYS_UNCONNECTED_1243, SYNOPSYS_UNCONNECTED_1244, SYNOPSYS_UNCONNECTED_1245, SYNOPSYS_UNCONNECTED_1246, SYNOPSYS_UNCONNECTED_1247, SYNOPSYS_UNCONNECTED_1248, SYNOPSYS_UNCONNECTED_1249, SYNOPSYS_UNCONNECTED_1250, SYNOPSYS_UNCONNECTED_1251, SYNOPSYS_UNCONNECTED_1252, SYNOPSYS_UNCONNECTED_1253, SYNOPSYS_UNCONNECTED_1254, SYNOPSYS_UNCONNECTED_1255, SYNOPSYS_UNCONNECTED_1256, SYNOPSYS_UNCONNECTED_1257, SYNOPSYS_UNCONNECTED_1258, SYNOPSYS_UNCONNECTED_1259, SYNOPSYS_UNCONNECTED_1260, SYNOPSYS_UNCONNECTED_1261, SYNOPSYS_UNCONNECTED_1262, SYNOPSYS_UNCONNECTED_1263, SYNOPSYS_UNCONNECTED_1264, SYNOPSYS_UNCONNECTED_1265, SYNOPSYS_UNCONNECTED_1266, SYNOPSYS_UNCONNECTED_1267, SYNOPSYS_UNCONNECTED_1268, SYNOPSYS_UNCONNECTED_1269, SYNOPSYS_UNCONNECTED_1270, SYNOPSYS_UNCONNECTED_1271, SYNOPSYS_UNCONNECTED_1272, SYNOPSYS_UNCONNECTED_1273, SYNOPSYS_UNCONNECTED_1274, SYNOPSYS_UNCONNECTED_1275, SYNOPSYS_UNCONNECTED_1276, SYNOPSYS_UNCONNECTED_1277, SYNOPSYS_UNCONNECTED_1278, SYNOPSYS_UNCONNECTED_1279, SYNOPSYS_UNCONNECTED_1280, data_head_o_flat_pretrunc } = { data_i, data_i } >> { iptr_r_data, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 };
  assign { yumi_o, SYNOPSYS_UNCONNECTED_1281, SYNOPSYS_UNCONNECTED_1282, SYNOPSYS_UNCONNECTED_1283, SYNOPSYS_UNCONNECTED_1284, SYNOPSYS_UNCONNECTED_1285, SYNOPSYS_UNCONNECTED_1286, SYNOPSYS_UNCONNECTED_1287, SYNOPSYS_UNCONNECTED_1288, SYNOPSYS_UNCONNECTED_1289, SYNOPSYS_UNCONNECTED_1290 } = { go_channels_i, go_channels_i } << iptr_r;

  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r),
    .n_o({ SYNOPSYS_UNCONNECTED_1291, SYNOPSYS_UNCONNECTED_1292, SYNOPSYS_UNCONNECTED_1293, SYNOPSYS_UNCONNECTED_1294 })
  );


  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(iptr_r_data),
    .n_o({ SYNOPSYS_UNCONNECTED_1295, SYNOPSYS_UNCONNECTED_1296, SYNOPSYS_UNCONNECTED_1297, SYNOPSYS_UNCONNECTED_1298 })
  );


endmodule



module bsg_scan_width_p10_and_p1_lo_to_hi_p1
(
  i,
  o
);

  input [9:0] i;
  output [9:0] o;
  wire [9:0] o;
  wire t_3__9_,t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,
  t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,
  t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__9_ = i[0] & 1'b1;
  assign t_1__8_ = i[1] & i[0];
  assign t_1__7_ = i[2] & i[1];
  assign t_1__6_ = i[3] & i[2];
  assign t_1__5_ = i[4] & i[3];
  assign t_1__4_ = i[5] & i[4];
  assign t_1__3_ = i[6] & i[5];
  assign t_1__2_ = i[7] & i[6];
  assign t_1__1_ = i[8] & i[7];
  assign t_1__0_ = i[9] & i[8];
  assign t_2__9_ = t_1__9_ & 1'b1;
  assign t_2__8_ = t_1__8_ & 1'b1;
  assign t_2__7_ = t_1__7_ & t_1__9_;
  assign t_2__6_ = t_1__6_ & t_1__8_;
  assign t_2__5_ = t_1__5_ & t_1__7_;
  assign t_2__4_ = t_1__4_ & t_1__6_;
  assign t_2__3_ = t_1__3_ & t_1__5_;
  assign t_2__2_ = t_1__2_ & t_1__4_;
  assign t_2__1_ = t_1__1_ & t_1__3_;
  assign t_2__0_ = t_1__0_ & t_1__2_;
  assign t_3__9_ = t_2__9_ & 1'b1;
  assign t_3__8_ = t_2__8_ & 1'b1;
  assign t_3__7_ = t_2__7_ & 1'b1;
  assign t_3__6_ = t_2__6_ & 1'b1;
  assign t_3__5_ = t_2__5_ & t_2__9_;
  assign t_3__4_ = t_2__4_ & t_2__8_;
  assign t_3__3_ = t_2__3_ & t_2__7_;
  assign t_3__2_ = t_2__2_ & t_2__6_;
  assign t_3__1_ = t_2__1_ & t_2__5_;
  assign t_3__0_ = t_2__0_ & t_2__4_;
  assign o[0] = t_3__9_ & 1'b1;
  assign o[1] = t_3__8_ & 1'b1;
  assign o[2] = t_3__7_ & 1'b1;
  assign o[3] = t_3__6_ & 1'b1;
  assign o[4] = t_3__5_ & 1'b1;
  assign o[5] = t_3__4_ & 1'b1;
  assign o[6] = t_3__3_ & 1'b1;
  assign o[7] = t_3__2_ & 1'b1;
  assign o[8] = t_3__1_ & t_3__9_;
  assign o[9] = t_3__0_ & t_3__8_;

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_width_p16
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [5:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p8
  aligned_left
  (
    .i(i[7:0]),
    .addr_o(aligned_addrs[2:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p8
  aligned_right
  (
    .i(i[15:8]),
    .addr_o(aligned_addrs[5:3]),
    .v_o(addr_o[3])
  );

  assign v_o = addr_o[3] | aligned_vs[0];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[5];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[4];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[3];

endmodule



module bsg_encode_one_hot_width_p11
(
  i,
  addr_o,
  v_o
);

  input [10:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;

  bsg_encode_one_hot_width_p16
  unaligned_align
  (
    .i({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, i }),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_thermometer_count_width_p10
(
  i,
  o
);

  input [9:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  wire [9:0] big_one_hot;

  bsg_encode_one_hot_width_p11
  big_encode_one_hot
  (
    .i({ i[9:9], big_one_hot }),
    .addr_o(o)
  );

  assign big_one_hot[9] = N0 & i[8];
  assign N0 = ~i[9];
  assign big_one_hot[8] = N1 & i[7];
  assign N1 = ~i[8];
  assign big_one_hot[7] = N2 & i[6];
  assign N2 = ~i[7];
  assign big_one_hot[6] = N3 & i[5];
  assign N3 = ~i[6];
  assign big_one_hot[5] = N4 & i[4];
  assign N4 = ~i[5];
  assign big_one_hot[4] = N5 & i[3];
  assign N5 = ~i[4];
  assign big_one_hot[3] = N6 & i[2];
  assign N6 = ~i[3];
  assign big_one_hot[2] = N7 & i[1];
  assign N7 = ~i[2];
  assign big_one_hot[1] = N8 & i[0];
  assign N8 = ~i[1];
  assign big_one_hot[0] = ~i[0];

endmodule



module bsg_rr_f2f_middle_width_p128_middle_meet_p10
(
  valid_head_i,
  ready_head_i,
  go_channels_o,
  go_cnt_o
);

  input [9:0] valid_head_i;
  input [9:0] ready_head_i;
  output [9:0] go_channels_o;
  output [3:0] go_cnt_o;
  wire [9:0] go_channels_o,happy_channels;
  wire [3:0] go_cnt_o;

  bsg_scan_width_p10_and_p1_lo_to_hi_p1
  and_scan
  (
    .i(happy_channels),
    .o(go_channels_o)
  );


  bsg_thermometer_count_width_p10
  genblk1_genblk1_thermo
  (
    .i(go_channels_o),
    .o(go_cnt_o)
  );

  assign happy_channels[9] = valid_head_i[9] & ready_head_i[9];
  assign happy_channels[8] = valid_head_i[8] & ready_head_i[8];
  assign happy_channels[7] = valid_head_i[7] & ready_head_i[7];
  assign happy_channels[6] = valid_head_i[6] & ready_head_i[6];
  assign happy_channels[5] = valid_head_i[5] & ready_head_i[5];
  assign happy_channels[4] = valid_head_i[4] & ready_head_i[4];
  assign happy_channels[3] = valid_head_i[3] & ready_head_i[3];
  assign happy_channels[2] = valid_head_i[2] & ready_head_i[2];
  assign happy_channels[1] = valid_head_i[1] & ready_head_i[1];
  assign happy_channels[0] = valid_head_i[0] & ready_head_i[0];

endmodule



module bsg_rr_f2f_output_width_p128_num_out_p10_middle_meet_p10
(
  clk,
  reset,
  ready_i,
  ready_head_o,
  go_channels_i,
  go_cnt_i,
  data_head_i,
  valid_o,
  data_o
);

  input [9:0] ready_i;
  output [9:0] ready_head_o;
  input [9:0] go_channels_i;
  input [3:0] go_cnt_i;
  input [1279:0] data_head_i;
  output [9:0] valid_o;
  output [1279:0] data_o;
  input clk;
  input reset;
  wire [9:0] ready_head_o,valid_o;
  wire [1279:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,SYNOPSYS_UNCONNECTED_1,
  SYNOPSYS_UNCONNECTED_2,SYNOPSYS_UNCONNECTED_3,SYNOPSYS_UNCONNECTED_4,
  SYNOPSYS_UNCONNECTED_5,SYNOPSYS_UNCONNECTED_6,SYNOPSYS_UNCONNECTED_7,SYNOPSYS_UNCONNECTED_8,
  SYNOPSYS_UNCONNECTED_9,SYNOPSYS_UNCONNECTED_10,SYNOPSYS_UNCONNECTED_11,
  SYNOPSYS_UNCONNECTED_12,SYNOPSYS_UNCONNECTED_13,SYNOPSYS_UNCONNECTED_14,
  SYNOPSYS_UNCONNECTED_15,SYNOPSYS_UNCONNECTED_16,SYNOPSYS_UNCONNECTED_17,SYNOPSYS_UNCONNECTED_18;
  wire [3:0] optr_r,optr_r_data;

  bsg_rotate_right_width_p10
  ready_rr
  (
    .data_i(ready_i),
    .rot_i(optr_r),
    .o(ready_head_o)
  );

  assign { valid_o, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10 } = { go_channels_i, go_channels_i } << optr_r;

  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r),
    .n_o({ SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14 })
  );


  bsg_circular_ptr_slots_p10_max_add_p10
  c_ptr_data
  (
    .clk(clk),
    .reset_i(reset),
    .add_i(go_cnt_i),
    .o(optr_r_data),
    .n_o({ SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16, SYNOPSYS_UNCONNECTED_17, SYNOPSYS_UNCONNECTED_18 })
  );

  assign N370 = N0 & optr_r_data[3];
  assign N0 = ~optr_r_data[2];
  assign N371 = optr_r_data[2] & N1;
  assign N1 = ~optr_r_data[3];
  assign N372 = N2 & N3;
  assign N2 = ~optr_r_data[2];
  assign N3 = ~optr_r_data[3];
  assign N373 = optr_r_data[0] & optr_r_data[1];
  assign N374 = N4 & optr_r_data[1];
  assign N4 = ~optr_r_data[0];
  assign N375 = optr_r_data[0] & N5;
  assign N5 = ~optr_r_data[1];
  assign N376 = N6 & N7;
  assign N6 = ~optr_r_data[0];
  assign N7 = ~optr_r_data[1];
  assign N235 = N370 & N374;
  assign N234 = N370 & N375;
  assign N233 = N370 & N376;
  assign N232 = N371 & N373;
  assign N231 = N371 & N374;
  assign N230 = N371 & N375;
  assign N229 = N371 & N376;
  assign N228 = N372 & N373;
  assign N227 = N372 & N374;
  assign N226 = N372 & N375;
  assign N225 = N372 & N376;
  assign N377 = N8 & optr_r_data[3];
  assign N8 = ~optr_r_data[2];
  assign N378 = optr_r_data[2] & N9;
  assign N9 = ~optr_r_data[3];
  assign N379 = N10 & N11;
  assign N10 = ~optr_r_data[2];
  assign N11 = ~optr_r_data[3];
  assign N380 = optr_r_data[0] & optr_r_data[1];
  assign N381 = N12 & optr_r_data[1];
  assign N12 = ~optr_r_data[0];
  assign N382 = optr_r_data[0] & N13;
  assign N13 = ~optr_r_data[1];
  assign N383 = N14 & N15;
  assign N14 = ~optr_r_data[0];
  assign N15 = ~optr_r_data[1];
  assign N247 = N377 & N380;
  assign N246 = N377 & N381;
  assign N245 = N377 & N382;
  assign N244 = N377 & N383;
  assign N243 = N378 & N380;
  assign N242 = N378 & N381;
  assign N241 = N378 & N382;
  assign N240 = N378 & N383;
  assign N239 = N379 & N380;
  assign N238 = N379 & N381;
  assign N237 = N379 & N382;
  assign N236 = N379 & N383;
  assign N384 = optr_r_data[2] & optr_r_data[3];
  assign N385 = N16 & optr_r_data[3];
  assign N16 = ~optr_r_data[2];
  assign N386 = optr_r_data[2] & N17;
  assign N17 = ~optr_r_data[3];
  assign N387 = N18 & N19;
  assign N18 = ~optr_r_data[2];
  assign N19 = ~optr_r_data[3];
  assign N388 = optr_r_data[0] & optr_r_data[1];
  assign N389 = N20 & optr_r_data[1];
  assign N20 = ~optr_r_data[0];
  assign N390 = optr_r_data[0] & N21;
  assign N21 = ~optr_r_data[1];
  assign N391 = N22 & N23;
  assign N22 = ~optr_r_data[0];
  assign N23 = ~optr_r_data[1];
  assign N260 = N384 & N391;
  assign N259 = N385 & N388;
  assign N258 = N385 & N389;
  assign N257 = N385 & N390;
  assign N256 = N385 & N391;
  assign N255 = N386 & N388;
  assign N254 = N386 & N389;
  assign N253 = N386 & N390;
  assign N252 = N386 & N391;
  assign N251 = N387 & N388;
  assign N250 = N387 & N389;
  assign N249 = N387 & N390;
  assign N248 = N387 & N391;
  assign N392 = optr_r_data[2] & optr_r_data[3];
  assign N393 = N24 & optr_r_data[3];
  assign N24 = ~optr_r_data[2];
  assign N394 = optr_r_data[2] & N25;
  assign N25 = ~optr_r_data[3];
  assign N395 = N26 & N27;
  assign N26 = ~optr_r_data[2];
  assign N27 = ~optr_r_data[3];
  assign N396 = optr_r_data[0] & optr_r_data[1];
  assign N397 = N28 & optr_r_data[1];
  assign N28 = ~optr_r_data[0];
  assign N398 = optr_r_data[0] & N29;
  assign N29 = ~optr_r_data[1];
  assign N399 = N30 & N31;
  assign N30 = ~optr_r_data[0];
  assign N31 = ~optr_r_data[1];
  assign N274 = N392 & N398;
  assign N273 = N392 & N399;
  assign N272 = N393 & N396;
  assign N271 = N393 & N397;
  assign N270 = N393 & N398;
  assign N269 = N393 & N399;
  assign N268 = N394 & N396;
  assign N267 = N394 & N397;
  assign N266 = N394 & N398;
  assign N265 = N394 & N399;
  assign N264 = N395 & N396;
  assign N263 = N395 & N397;
  assign N262 = N395 & N398;
  assign N261 = N395 & N399;
  assign N400 = optr_r_data[2] & optr_r_data[3];
  assign N401 = N32 & optr_r_data[3];
  assign N32 = ~optr_r_data[2];
  assign N402 = optr_r_data[2] & N33;
  assign N33 = ~optr_r_data[3];
  assign N403 = N34 & N35;
  assign N34 = ~optr_r_data[2];
  assign N35 = ~optr_r_data[3];
  assign N404 = optr_r_data[0] & optr_r_data[1];
  assign N405 = N36 & optr_r_data[1];
  assign N36 = ~optr_r_data[0];
  assign N406 = optr_r_data[0] & N37;
  assign N37 = ~optr_r_data[1];
  assign N407 = N38 & N39;
  assign N38 = ~optr_r_data[0];
  assign N39 = ~optr_r_data[1];
  assign N289 = N400 & N405;
  assign N288 = N400 & N406;
  assign N287 = N400 & N407;
  assign N286 = N401 & N404;
  assign N285 = N401 & N405;
  assign N284 = N401 & N406;
  assign N283 = N401 & N407;
  assign N282 = N402 & N404;
  assign N281 = N402 & N405;
  assign N280 = N402 & N406;
  assign N279 = N402 & N407;
  assign N278 = N403 & N404;
  assign N277 = N403 & N405;
  assign N276 = N403 & N406;
  assign N275 = N403 & N407;
  assign N408 = optr_r_data[2] & optr_r_data[3];
  assign N409 = N40 & optr_r_data[3];
  assign N40 = ~optr_r_data[2];
  assign N410 = optr_r_data[2] & N41;
  assign N41 = ~optr_r_data[3];
  assign N411 = N42 & N43;
  assign N42 = ~optr_r_data[2];
  assign N43 = ~optr_r_data[3];
  assign N412 = optr_r_data[0] & optr_r_data[1];
  assign N413 = N44 & optr_r_data[1];
  assign N44 = ~optr_r_data[0];
  assign N414 = optr_r_data[0] & N45;
  assign N45 = ~optr_r_data[1];
  assign N415 = N46 & N47;
  assign N46 = ~optr_r_data[0];
  assign N47 = ~optr_r_data[1];
  assign N305 = N408 & N412;
  assign N304 = N408 & N413;
  assign N303 = N408 & N414;
  assign N302 = N408 & N415;
  assign N301 = N409 & N412;
  assign N300 = N409 & N413;
  assign N299 = N409 & N414;
  assign N298 = N409 & N415;
  assign N297 = N410 & N412;
  assign N296 = N410 & N413;
  assign N295 = N410 & N414;
  assign N294 = N410 & N415;
  assign N293 = N411 & N412;
  assign N292 = N411 & N413;
  assign N291 = N411 & N414;
  assign N290 = N411 & N415;
  assign N416 = optr_r_data[2] & optr_r_data[3];
  assign N417 = N48 & optr_r_data[3];
  assign N48 = ~optr_r_data[2];
  assign N418 = optr_r_data[2] & N49;
  assign N49 = ~optr_r_data[3];
  assign N419 = N50 & N51;
  assign N50 = ~optr_r_data[2];
  assign N51 = ~optr_r_data[3];
  assign N420 = optr_r_data[0] & optr_r_data[1];
  assign N421 = N52 & optr_r_data[1];
  assign N52 = ~optr_r_data[0];
  assign N422 = optr_r_data[0] & N53;
  assign N53 = ~optr_r_data[1];
  assign N423 = N54 & N55;
  assign N54 = ~optr_r_data[0];
  assign N55 = ~optr_r_data[1];
  assign N321 = N416 & N420;
  assign N320 = N416 & N421;
  assign N319 = N416 & N422;
  assign N318 = N416 & N423;
  assign N317 = N417 & N420;
  assign N316 = N417 & N421;
  assign N315 = N417 & N422;
  assign N314 = N417 & N423;
  assign N313 = N418 & N420;
  assign N312 = N418 & N421;
  assign N311 = N418 & N422;
  assign N310 = N418 & N423;
  assign N309 = N419 & N420;
  assign N308 = N419 & N421;
  assign N307 = N419 & N422;
  assign N306 = N419 & N423;
  assign N424 = optr_r_data[2] & optr_r_data[3];
  assign N425 = N56 & optr_r_data[3];
  assign N56 = ~optr_r_data[2];
  assign N426 = optr_r_data[2] & N57;
  assign N57 = ~optr_r_data[3];
  assign N427 = N58 & N59;
  assign N58 = ~optr_r_data[2];
  assign N59 = ~optr_r_data[3];
  assign N428 = optr_r_data[0] & optr_r_data[1];
  assign N429 = N60 & optr_r_data[1];
  assign N60 = ~optr_r_data[0];
  assign N430 = optr_r_data[0] & N61;
  assign N61 = ~optr_r_data[1];
  assign N431 = N62 & N63;
  assign N62 = ~optr_r_data[0];
  assign N63 = ~optr_r_data[1];
  assign N337 = N424 & N428;
  assign N336 = N424 & N429;
  assign N335 = N424 & N430;
  assign N334 = N424 & N431;
  assign N333 = N425 & N428;
  assign N332 = N425 & N429;
  assign N331 = N425 & N430;
  assign N330 = N425 & N431;
  assign N329 = N426 & N428;
  assign N328 = N426 & N429;
  assign N327 = N426 & N430;
  assign N326 = N426 & N431;
  assign N325 = N427 & N428;
  assign N324 = N427 & N429;
  assign N323 = N427 & N430;
  assign N322 = N427 & N431;
  assign N432 = optr_r_data[2] & optr_r_data[3];
  assign N433 = N64 & optr_r_data[3];
  assign N64 = ~optr_r_data[2];
  assign N434 = optr_r_data[2] & N65;
  assign N65 = ~optr_r_data[3];
  assign N435 = N66 & N67;
  assign N66 = ~optr_r_data[2];
  assign N67 = ~optr_r_data[3];
  assign N436 = optr_r_data[0] & optr_r_data[1];
  assign N437 = N68 & optr_r_data[1];
  assign N68 = ~optr_r_data[0];
  assign N438 = optr_r_data[0] & N69;
  assign N69 = ~optr_r_data[1];
  assign N439 = N70 & N71;
  assign N70 = ~optr_r_data[0];
  assign N71 = ~optr_r_data[1];
  assign N353 = N432 & N436;
  assign N352 = N432 & N437;
  assign N351 = N432 & N438;
  assign N350 = N432 & N439;
  assign N349 = N433 & N436;
  assign N348 = N433 & N437;
  assign N347 = N433 & N438;
  assign N346 = N433 & N439;
  assign N345 = N434 & N436;
  assign N344 = N434 & N437;
  assign N343 = N434 & N438;
  assign N342 = N434 & N439;
  assign N341 = N435 & N436;
  assign N340 = N435 & N437;
  assign N339 = N435 & N438;
  assign N338 = N435 & N439;
  assign N440 = optr_r_data[2] & optr_r_data[3];
  assign N441 = N72 & optr_r_data[3];
  assign N72 = ~optr_r_data[2];
  assign N442 = optr_r_data[2] & N73;
  assign N73 = ~optr_r_data[3];
  assign N443 = N74 & N75;
  assign N74 = ~optr_r_data[2];
  assign N75 = ~optr_r_data[3];
  assign N444 = optr_r_data[0] & optr_r_data[1];
  assign N445 = N76 & optr_r_data[1];
  assign N76 = ~optr_r_data[0];
  assign N446 = optr_r_data[0] & N77;
  assign N77 = ~optr_r_data[1];
  assign N447 = N78 & N79;
  assign N78 = ~optr_r_data[0];
  assign N79 = ~optr_r_data[1];
  assign N369 = N440 & N444;
  assign N368 = N440 & N445;
  assign N367 = N440 & N446;
  assign N366 = N440 & N447;
  assign N365 = N441 & N444;
  assign N364 = N441 & N445;
  assign N363 = N441 & N446;
  assign N362 = N441 & N447;
  assign N361 = N442 & N444;
  assign N360 = N442 & N445;
  assign N359 = N442 & N446;
  assign N358 = N442 & N447;
  assign N357 = N443 & N444;
  assign N356 = N443 & N445;
  assign N355 = N443 & N446;
  assign N354 = N443 & N447;
  assign data_o[127:0] = (N80)? data_head_i[127:0] : 
                         (N81)? data_head_i[255:128] : 
                         (N82)? data_head_i[383:256] : 
                         (N83)? data_head_i[511:384] : 
                         (N84)? data_head_i[639:512] : 
                         (N85)? data_head_i[767:640] : 
                         (N86)? data_head_i[895:768] : 
                         (N87)? data_head_i[1023:896] : 
                         (N88)? data_head_i[1151:1024] : 
                         (N89)? data_head_i[1279:1152] : 
                         (N90)? data_head_i[127:0] : 1'b0;
  assign N80 = N235;
  assign N81 = N234;
  assign N82 = N233;
  assign N83 = N232;
  assign N84 = N231;
  assign N85 = N230;
  assign N86 = N229;
  assign N87 = N228;
  assign N88 = N227;
  assign N89 = N226;
  assign N90 = N225;
  assign data_o[255:128] = (N91)? data_head_i[127:0] : 
                           (N92)? data_head_i[255:128] : 
                           (N93)? data_head_i[383:256] : 
                           (N94)? data_head_i[511:384] : 
                           (N95)? data_head_i[639:512] : 
                           (N96)? data_head_i[767:640] : 
                           (N97)? data_head_i[895:768] : 
                           (N98)? data_head_i[1023:896] : 
                           (N99)? data_head_i[1151:1024] : 
                           (N100)? data_head_i[1279:1152] : 
                           (N101)? data_head_i[127:0] : 
                           (N102)? data_head_i[255:128] : 1'b0;
  assign N91 = N247;
  assign N92 = N246;
  assign N93 = N245;
  assign N94 = N244;
  assign N95 = N243;
  assign N96 = N242;
  assign N97 = N241;
  assign N98 = N240;
  assign N99 = N239;
  assign N100 = N238;
  assign N101 = N237;
  assign N102 = N236;
  assign data_o[383:256] = (N103)? data_head_i[127:0] : 
                           (N104)? data_head_i[255:128] : 
                           (N105)? data_head_i[383:256] : 
                           (N106)? data_head_i[511:384] : 
                           (N107)? data_head_i[639:512] : 
                           (N108)? data_head_i[767:640] : 
                           (N109)? data_head_i[895:768] : 
                           (N110)? data_head_i[1023:896] : 
                           (N111)? data_head_i[1151:1024] : 
                           (N112)? data_head_i[1279:1152] : 
                           (N113)? data_head_i[127:0] : 
                           (N114)? data_head_i[255:128] : 
                           (N115)? data_head_i[383:256] : 1'b0;
  assign N103 = N260;
  assign N104 = N259;
  assign N105 = N258;
  assign N106 = N257;
  assign N107 = N256;
  assign N108 = N255;
  assign N109 = N254;
  assign N110 = N253;
  assign N111 = N252;
  assign N112 = N251;
  assign N113 = N250;
  assign N114 = N249;
  assign N115 = N248;
  assign data_o[511:384] = (N116)? data_head_i[127:0] : 
                           (N117)? data_head_i[255:128] : 
                           (N118)? data_head_i[383:256] : 
                           (N119)? data_head_i[511:384] : 
                           (N120)? data_head_i[639:512] : 
                           (N121)? data_head_i[767:640] : 
                           (N122)? data_head_i[895:768] : 
                           (N123)? data_head_i[1023:896] : 
                           (N124)? data_head_i[1151:1024] : 
                           (N125)? data_head_i[1279:1152] : 
                           (N126)? data_head_i[127:0] : 
                           (N127)? data_head_i[255:128] : 
                           (N128)? data_head_i[383:256] : 
                           (N129)? data_head_i[511:384] : 1'b0;
  assign N116 = N274;
  assign N117 = N273;
  assign N118 = N272;
  assign N119 = N271;
  assign N120 = N270;
  assign N121 = N269;
  assign N122 = N268;
  assign N123 = N267;
  assign N124 = N266;
  assign N125 = N265;
  assign N126 = N264;
  assign N127 = N263;
  assign N128 = N262;
  assign N129 = N261;
  assign data_o[639:512] = (N130)? data_head_i[127:0] : 
                           (N131)? data_head_i[255:128] : 
                           (N132)? data_head_i[383:256] : 
                           (N133)? data_head_i[511:384] : 
                           (N134)? data_head_i[639:512] : 
                           (N135)? data_head_i[767:640] : 
                           (N136)? data_head_i[895:768] : 
                           (N137)? data_head_i[1023:896] : 
                           (N138)? data_head_i[1151:1024] : 
                           (N139)? data_head_i[1279:1152] : 
                           (N140)? data_head_i[127:0] : 
                           (N141)? data_head_i[255:128] : 
                           (N142)? data_head_i[383:256] : 
                           (N143)? data_head_i[511:384] : 
                           (N144)? data_head_i[639:512] : 1'b0;
  assign N130 = N289;
  assign N131 = N288;
  assign N132 = N287;
  assign N133 = N286;
  assign N134 = N285;
  assign N135 = N284;
  assign N136 = N283;
  assign N137 = N282;
  assign N138 = N281;
  assign N139 = N280;
  assign N140 = N279;
  assign N141 = N278;
  assign N142 = N277;
  assign N143 = N276;
  assign N144 = N275;
  assign data_o[767:640] = (N145)? data_head_i[127:0] : 
                           (N146)? data_head_i[255:128] : 
                           (N147)? data_head_i[383:256] : 
                           (N148)? data_head_i[511:384] : 
                           (N149)? data_head_i[639:512] : 
                           (N150)? data_head_i[767:640] : 
                           (N151)? data_head_i[895:768] : 
                           (N152)? data_head_i[1023:896] : 
                           (N153)? data_head_i[1151:1024] : 
                           (N154)? data_head_i[1279:1152] : 
                           (N155)? data_head_i[127:0] : 
                           (N156)? data_head_i[255:128] : 
                           (N157)? data_head_i[383:256] : 
                           (N158)? data_head_i[511:384] : 
                           (N159)? data_head_i[639:512] : 
                           (N160)? data_head_i[767:640] : 1'b0;
  assign N145 = N305;
  assign N146 = N304;
  assign N147 = N303;
  assign N148 = N302;
  assign N149 = N301;
  assign N150 = N300;
  assign N151 = N299;
  assign N152 = N298;
  assign N153 = N297;
  assign N154 = N296;
  assign N155 = N295;
  assign N156 = N294;
  assign N157 = N293;
  assign N158 = N292;
  assign N159 = N291;
  assign N160 = N290;
  assign data_o[895:768] = (N161)? data_head_i[255:128] : 
                           (N162)? data_head_i[383:256] : 
                           (N163)? data_head_i[511:384] : 
                           (N164)? data_head_i[639:512] : 
                           (N165)? data_head_i[767:640] : 
                           (N166)? data_head_i[895:768] : 
                           (N167)? data_head_i[1023:896] : 
                           (N168)? data_head_i[1151:1024] : 
                           (N169)? data_head_i[1279:1152] : 
                           (N170)? data_head_i[127:0] : 
                           (N171)? data_head_i[255:128] : 
                           (N172)? data_head_i[383:256] : 
                           (N173)? data_head_i[511:384] : 
                           (N174)? data_head_i[639:512] : 
                           (N175)? data_head_i[767:640] : 
                           (N176)? data_head_i[895:768] : 1'b0;
  assign N161 = N321;
  assign N162 = N320;
  assign N163 = N319;
  assign N164 = N318;
  assign N165 = N317;
  assign N166 = N316;
  assign N167 = N315;
  assign N168 = N314;
  assign N169 = N313;
  assign N170 = N312;
  assign N171 = N311;
  assign N172 = N310;
  assign N173 = N309;
  assign N174 = N308;
  assign N175 = N307;
  assign N176 = N306;
  assign data_o[1023:896] = (N177)? data_head_i[383:256] : 
                            (N178)? data_head_i[511:384] : 
                            (N179)? data_head_i[639:512] : 
                            (N180)? data_head_i[767:640] : 
                            (N181)? data_head_i[895:768] : 
                            (N182)? data_head_i[1023:896] : 
                            (N183)? data_head_i[1151:1024] : 
                            (N184)? data_head_i[1279:1152] : 
                            (N185)? data_head_i[127:0] : 
                            (N186)? data_head_i[255:128] : 
                            (N187)? data_head_i[383:256] : 
                            (N188)? data_head_i[511:384] : 
                            (N189)? data_head_i[639:512] : 
                            (N190)? data_head_i[767:640] : 
                            (N191)? data_head_i[895:768] : 
                            (N192)? data_head_i[1023:896] : 1'b0;
  assign N177 = N337;
  assign N178 = N336;
  assign N179 = N335;
  assign N180 = N334;
  assign N181 = N333;
  assign N182 = N332;
  assign N183 = N331;
  assign N184 = N330;
  assign N185 = N329;
  assign N186 = N328;
  assign N187 = N327;
  assign N188 = N326;
  assign N189 = N325;
  assign N190 = N324;
  assign N191 = N323;
  assign N192 = N322;
  assign data_o[1151:1024] = (N193)? data_head_i[511:384] : 
                             (N194)? data_head_i[639:512] : 
                             (N195)? data_head_i[767:640] : 
                             (N196)? data_head_i[895:768] : 
                             (N197)? data_head_i[1023:896] : 
                             (N198)? data_head_i[1151:1024] : 
                             (N199)? data_head_i[1279:1152] : 
                             (N200)? data_head_i[127:0] : 
                             (N201)? data_head_i[255:128] : 
                             (N202)? data_head_i[383:256] : 
                             (N203)? data_head_i[511:384] : 
                             (N204)? data_head_i[639:512] : 
                             (N205)? data_head_i[767:640] : 
                             (N206)? data_head_i[895:768] : 
                             (N207)? data_head_i[1023:896] : 
                             (N208)? data_head_i[1151:1024] : 1'b0;
  assign N193 = N353;
  assign N194 = N352;
  assign N195 = N351;
  assign N196 = N350;
  assign N197 = N349;
  assign N198 = N348;
  assign N199 = N347;
  assign N200 = N346;
  assign N201 = N345;
  assign N202 = N344;
  assign N203 = N343;
  assign N204 = N342;
  assign N205 = N341;
  assign N206 = N340;
  assign N207 = N339;
  assign N208 = N338;
  assign data_o[1279:1152] = (N209)? data_head_i[639:512] : 
                             (N210)? data_head_i[767:640] : 
                             (N211)? data_head_i[895:768] : 
                             (N212)? data_head_i[1023:896] : 
                             (N213)? data_head_i[1151:1024] : 
                             (N214)? data_head_i[1279:1152] : 
                             (N215)? data_head_i[127:0] : 
                             (N216)? data_head_i[255:128] : 
                             (N217)? data_head_i[383:256] : 
                             (N218)? data_head_i[511:384] : 
                             (N219)? data_head_i[639:512] : 
                             (N220)? data_head_i[767:640] : 
                             (N221)? data_head_i[895:768] : 
                             (N222)? data_head_i[1023:896] : 
                             (N223)? data_head_i[1151:1024] : 
                             (N224)? data_head_i[1279:1152] : 1'b0;
  assign N209 = N369;
  assign N210 = N368;
  assign N211 = N367;
  assign N212 = N366;
  assign N213 = N365;
  assign N214 = N364;
  assign N215 = N363;
  assign N216 = N362;
  assign N217 = N361;
  assign N218 = N360;
  assign N219 = N359;
  assign N220 = N358;
  assign N221 = N357;
  assign N222 = N356;
  assign N223 = N355;
  assign N224 = N354;

endmodule



module bsg_round_robin_fifo_to_fifo_width_p128_num_in_p10_num_out_p10_out_channel_count_mask_p512
(
  clk,
  reset,
  valid_i,
  data_i,
  yumi_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [9:0] valid_i;
  input [1279:0] data_i;
  output [9:0] yumi_o;
  input [3:0] in_top_channel_i;
  input [3:0] out_top_channel_i;
  output [9:0] valid_o;
  output [1279:0] data_o;
  input [9:0] ready_i;
  input clk;
  input reset;
  wire [9:0] yumi_o,valid_o,go_channels;
  wire [1279:0] data_o,data_o_flat,oc_9__out_chan_data_head_array;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,yumi_int_o_9__9_,yumi_int_o_9__8_,
  yumi_int_o_9__7_,yumi_int_o_9__6_,yumi_int_o_9__5_,yumi_int_o_9__4_,yumi_int_o_9__3_,
  yumi_int_o_9__2_,yumi_int_o_9__1_,yumi_int_o_9__0_,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,valid_int_o_9__9_,valid_int_o_9__8_,valid_int_o_9__7_,
  valid_int_o_9__6_,valid_int_o_9__5_,valid_int_o_9__4_,valid_int_o_9__3_,valid_int_o_9__2_,
  valid_int_o_9__1_,valid_int_o_9__0_,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,data_int_o_9__1279_,data_int_o_9__1278_,data_int_o_9__1277_,
  data_int_o_9__1276_,data_int_o_9__1275_,data_int_o_9__1274_,data_int_o_9__1273_,
  data_int_o_9__1272_,data_int_o_9__1271_,data_int_o_9__1270_,data_int_o_9__1269_,
  data_int_o_9__1268_,data_int_o_9__1267_,data_int_o_9__1266_,data_int_o_9__1265_,
  data_int_o_9__1264_,data_int_o_9__1263_,data_int_o_9__1262_,data_int_o_9__1261_,
  data_int_o_9__1260_,data_int_o_9__1259_,data_int_o_9__1258_,data_int_o_9__1257_,
  data_int_o_9__1256_,data_int_o_9__1255_,data_int_o_9__1254_,data_int_o_9__1253_,
  data_int_o_9__1252_,data_int_o_9__1251_,data_int_o_9__1250_,data_int_o_9__1249_,
  data_int_o_9__1248_,data_int_o_9__1247_,data_int_o_9__1246_,data_int_o_9__1245_,
  data_int_o_9__1244_,data_int_o_9__1243_,data_int_o_9__1242_,data_int_o_9__1241_,
  data_int_o_9__1240_,data_int_o_9__1239_,data_int_o_9__1238_,data_int_o_9__1237_,
  data_int_o_9__1236_,data_int_o_9__1235_,data_int_o_9__1234_,data_int_o_9__1233_,
  data_int_o_9__1232_,data_int_o_9__1231_,data_int_o_9__1230_,data_int_o_9__1229_,
  data_int_o_9__1228_,data_int_o_9__1227_,data_int_o_9__1226_,data_int_o_9__1225_,
  data_int_o_9__1224_,data_int_o_9__1223_,data_int_o_9__1222_,data_int_o_9__1221_,
  data_int_o_9__1220_,data_int_o_9__1219_,data_int_o_9__1218_,data_int_o_9__1217_,
  data_int_o_9__1216_,data_int_o_9__1215_,data_int_o_9__1214_,data_int_o_9__1213_,
  data_int_o_9__1212_,data_int_o_9__1211_,data_int_o_9__1210_,data_int_o_9__1209_,
  data_int_o_9__1208_,data_int_o_9__1207_,data_int_o_9__1206_,data_int_o_9__1205_,
  data_int_o_9__1204_,data_int_o_9__1203_,data_int_o_9__1202_,data_int_o_9__1201_,
  data_int_o_9__1200_,data_int_o_9__1199_,data_int_o_9__1198_,data_int_o_9__1197_,
  data_int_o_9__1196_,data_int_o_9__1195_,data_int_o_9__1194_,data_int_o_9__1193_,
  data_int_o_9__1192_,data_int_o_9__1191_,data_int_o_9__1190_,data_int_o_9__1189_,
  data_int_o_9__1188_,data_int_o_9__1187_,data_int_o_9__1186_,data_int_o_9__1185_,
  data_int_o_9__1184_,data_int_o_9__1183_,data_int_o_9__1182_,data_int_o_9__1181_,
  data_int_o_9__1180_,data_int_o_9__1179_,data_int_o_9__1178_,data_int_o_9__1177_,
  data_int_o_9__1176_,data_int_o_9__1175_,data_int_o_9__1174_,data_int_o_9__1173_,
  data_int_o_9__1172_,data_int_o_9__1171_,data_int_o_9__1170_,data_int_o_9__1169_,
  data_int_o_9__1168_,data_int_o_9__1167_,data_int_o_9__1166_,data_int_o_9__1165_,
  data_int_o_9__1164_,data_int_o_9__1163_,data_int_o_9__1162_,data_int_o_9__1161_,
  data_int_o_9__1160_,data_int_o_9__1159_,data_int_o_9__1158_,data_int_o_9__1157_,
  data_int_o_9__1156_,data_int_o_9__1155_,data_int_o_9__1154_,data_int_o_9__1153_,
  data_int_o_9__1152_,data_int_o_9__1151_,data_int_o_9__1150_,data_int_o_9__1149_,
  data_int_o_9__1148_,data_int_o_9__1147_,data_int_o_9__1146_,data_int_o_9__1145_,
  data_int_o_9__1144_,data_int_o_9__1143_,data_int_o_9__1142_,data_int_o_9__1141_,
  data_int_o_9__1140_,data_int_o_9__1139_,data_int_o_9__1138_,data_int_o_9__1137_,
  data_int_o_9__1136_,data_int_o_9__1135_,data_int_o_9__1134_,data_int_o_9__1133_,
  data_int_o_9__1132_,data_int_o_9__1131_,data_int_o_9__1130_,data_int_o_9__1129_,
  data_int_o_9__1128_,data_int_o_9__1127_,data_int_o_9__1126_,data_int_o_9__1125_,
  data_int_o_9__1124_,data_int_o_9__1123_,data_int_o_9__1122_,data_int_o_9__1121_,
  data_int_o_9__1120_,data_int_o_9__1119_,data_int_o_9__1118_,data_int_o_9__1117_,
  data_int_o_9__1116_,data_int_o_9__1115_,data_int_o_9__1114_,data_int_o_9__1113_,
  data_int_o_9__1112_,data_int_o_9__1111_,data_int_o_9__1110_,data_int_o_9__1109_,
  data_int_o_9__1108_,data_int_o_9__1107_,data_int_o_9__1106_,data_int_o_9__1105_,
  data_int_o_9__1104_,data_int_o_9__1103_,data_int_o_9__1102_,data_int_o_9__1101_,
  data_int_o_9__1100_,data_int_o_9__1099_,data_int_o_9__1098_,data_int_o_9__1097_,
  data_int_o_9__1096_,data_int_o_9__1095_,data_int_o_9__1094_,data_int_o_9__1093_,
  data_int_o_9__1092_,data_int_o_9__1091_,data_int_o_9__1090_,data_int_o_9__1089_,
  data_int_o_9__1088_,data_int_o_9__1087_,data_int_o_9__1086_,data_int_o_9__1085_,
  data_int_o_9__1084_,data_int_o_9__1083_,data_int_o_9__1082_,data_int_o_9__1081_,
  data_int_o_9__1080_,data_int_o_9__1079_,data_int_o_9__1078_,data_int_o_9__1077_,
  data_int_o_9__1076_,data_int_o_9__1075_,data_int_o_9__1074_,data_int_o_9__1073_,
  data_int_o_9__1072_,data_int_o_9__1071_,data_int_o_9__1070_,data_int_o_9__1069_,
  data_int_o_9__1068_,data_int_o_9__1067_,data_int_o_9__1066_,data_int_o_9__1065_,
  data_int_o_9__1064_,data_int_o_9__1063_,data_int_o_9__1062_,data_int_o_9__1061_,
  data_int_o_9__1060_,data_int_o_9__1059_,data_int_o_9__1058_,data_int_o_9__1057_,
  data_int_o_9__1056_,data_int_o_9__1055_,data_int_o_9__1054_,data_int_o_9__1053_,
  data_int_o_9__1052_,data_int_o_9__1051_,data_int_o_9__1050_,data_int_o_9__1049_,
  data_int_o_9__1048_,data_int_o_9__1047_,data_int_o_9__1046_,data_int_o_9__1045_,
  data_int_o_9__1044_,data_int_o_9__1043_,data_int_o_9__1042_,data_int_o_9__1041_,
  data_int_o_9__1040_,data_int_o_9__1039_,data_int_o_9__1038_,data_int_o_9__1037_,
  data_int_o_9__1036_,data_int_o_9__1035_,data_int_o_9__1034_,data_int_o_9__1033_,
  data_int_o_9__1032_,data_int_o_9__1031_,data_int_o_9__1030_,data_int_o_9__1029_,
  data_int_o_9__1028_,data_int_o_9__1027_,data_int_o_9__1026_,data_int_o_9__1025_,
  data_int_o_9__1024_,data_int_o_9__1023_,data_int_o_9__1022_,data_int_o_9__1021_,
  data_int_o_9__1020_,data_int_o_9__1019_,data_int_o_9__1018_,data_int_o_9__1017_,
  data_int_o_9__1016_,data_int_o_9__1015_,data_int_o_9__1014_,data_int_o_9__1013_,
  data_int_o_9__1012_,data_int_o_9__1011_,data_int_o_9__1010_,data_int_o_9__1009_,
  data_int_o_9__1008_,data_int_o_9__1007_,data_int_o_9__1006_,data_int_o_9__1005_,
  data_int_o_9__1004_,data_int_o_9__1003_,data_int_o_9__1002_,data_int_o_9__1001_,
  data_int_o_9__1000_,data_int_o_9__999_,data_int_o_9__998_,data_int_o_9__997_,
  data_int_o_9__996_,data_int_o_9__995_,data_int_o_9__994_,data_int_o_9__993_,data_int_o_9__992_,
  data_int_o_9__991_,data_int_o_9__990_,data_int_o_9__989_,data_int_o_9__988_,
  data_int_o_9__987_,data_int_o_9__986_,data_int_o_9__985_,data_int_o_9__984_,
  data_int_o_9__983_,data_int_o_9__982_,data_int_o_9__981_,data_int_o_9__980_,
  data_int_o_9__979_,data_int_o_9__978_,data_int_o_9__977_,data_int_o_9__976_,data_int_o_9__975_,
  data_int_o_9__974_,data_int_o_9__973_,data_int_o_9__972_,data_int_o_9__971_,
  data_int_o_9__970_,data_int_o_9__969_,data_int_o_9__968_,data_int_o_9__967_,
  data_int_o_9__966_,data_int_o_9__965_,data_int_o_9__964_,data_int_o_9__963_,
  data_int_o_9__962_,data_int_o_9__961_,data_int_o_9__960_,data_int_o_9__959_,
  data_int_o_9__958_,data_int_o_9__957_,data_int_o_9__956_,data_int_o_9__955_,data_int_o_9__954_,
  data_int_o_9__953_,data_int_o_9__952_,data_int_o_9__951_,data_int_o_9__950_,
  data_int_o_9__949_,data_int_o_9__948_,data_int_o_9__947_,data_int_o_9__946_,
  data_int_o_9__945_,data_int_o_9__944_,data_int_o_9__943_,data_int_o_9__942_,
  data_int_o_9__941_,data_int_o_9__940_,data_int_o_9__939_,data_int_o_9__938_,
  data_int_o_9__937_,data_int_o_9__936_,data_int_o_9__935_,data_int_o_9__934_,data_int_o_9__933_,
  data_int_o_9__932_,data_int_o_9__931_,data_int_o_9__930_,data_int_o_9__929_,
  data_int_o_9__928_,data_int_o_9__927_,data_int_o_9__926_,data_int_o_9__925_,
  data_int_o_9__924_,data_int_o_9__923_,data_int_o_9__922_,data_int_o_9__921_,
  data_int_o_9__920_,data_int_o_9__919_,data_int_o_9__918_,data_int_o_9__917_,
  data_int_o_9__916_,data_int_o_9__915_,data_int_o_9__914_,data_int_o_9__913_,data_int_o_9__912_,
  data_int_o_9__911_,data_int_o_9__910_,data_int_o_9__909_,data_int_o_9__908_,
  data_int_o_9__907_,data_int_o_9__906_,data_int_o_9__905_,data_int_o_9__904_,
  data_int_o_9__903_,data_int_o_9__902_,data_int_o_9__901_,data_int_o_9__900_,
  data_int_o_9__899_,data_int_o_9__898_,data_int_o_9__897_,data_int_o_9__896_,data_int_o_9__895_,
  data_int_o_9__894_,data_int_o_9__893_,data_int_o_9__892_,data_int_o_9__891_,
  data_int_o_9__890_,data_int_o_9__889_,data_int_o_9__888_,data_int_o_9__887_,
  data_int_o_9__886_,data_int_o_9__885_,data_int_o_9__884_,data_int_o_9__883_,
  data_int_o_9__882_,data_int_o_9__881_,data_int_o_9__880_,data_int_o_9__879_,
  data_int_o_9__878_,data_int_o_9__877_,data_int_o_9__876_,data_int_o_9__875_,data_int_o_9__874_,
  data_int_o_9__873_,data_int_o_9__872_,data_int_o_9__871_,data_int_o_9__870_,
  data_int_o_9__869_,data_int_o_9__868_,data_int_o_9__867_,data_int_o_9__866_,
  data_int_o_9__865_,data_int_o_9__864_,data_int_o_9__863_,data_int_o_9__862_,
  data_int_o_9__861_,data_int_o_9__860_,data_int_o_9__859_,data_int_o_9__858_,
  data_int_o_9__857_,data_int_o_9__856_,data_int_o_9__855_,data_int_o_9__854_,data_int_o_9__853_,
  data_int_o_9__852_,data_int_o_9__851_,data_int_o_9__850_,data_int_o_9__849_,
  data_int_o_9__848_,data_int_o_9__847_,data_int_o_9__846_,data_int_o_9__845_,
  data_int_o_9__844_,data_int_o_9__843_,data_int_o_9__842_,data_int_o_9__841_,
  data_int_o_9__840_,data_int_o_9__839_,data_int_o_9__838_,data_int_o_9__837_,
  data_int_o_9__836_,data_int_o_9__835_,data_int_o_9__834_,data_int_o_9__833_,data_int_o_9__832_,
  data_int_o_9__831_,data_int_o_9__830_,data_int_o_9__829_,data_int_o_9__828_,
  data_int_o_9__827_,data_int_o_9__826_,data_int_o_9__825_,data_int_o_9__824_,
  data_int_o_9__823_,data_int_o_9__822_,data_int_o_9__821_,data_int_o_9__820_,
  data_int_o_9__819_,data_int_o_9__818_,data_int_o_9__817_,data_int_o_9__816_,data_int_o_9__815_,
  data_int_o_9__814_,data_int_o_9__813_,data_int_o_9__812_,data_int_o_9__811_,
  data_int_o_9__810_,data_int_o_9__809_,data_int_o_9__808_,data_int_o_9__807_,
  data_int_o_9__806_,data_int_o_9__805_,data_int_o_9__804_,data_int_o_9__803_,
  data_int_o_9__802_,data_int_o_9__801_,data_int_o_9__800_,data_int_o_9__799_,
  data_int_o_9__798_,data_int_o_9__797_,data_int_o_9__796_,data_int_o_9__795_,data_int_o_9__794_,
  data_int_o_9__793_,data_int_o_9__792_,data_int_o_9__791_,data_int_o_9__790_,
  data_int_o_9__789_,data_int_o_9__788_,data_int_o_9__787_,data_int_o_9__786_,
  data_int_o_9__785_,data_int_o_9__784_,data_int_o_9__783_,data_int_o_9__782_,
  data_int_o_9__781_,data_int_o_9__780_,data_int_o_9__779_,data_int_o_9__778_,
  data_int_o_9__777_,data_int_o_9__776_,data_int_o_9__775_,data_int_o_9__774_,data_int_o_9__773_,
  data_int_o_9__772_,data_int_o_9__771_,data_int_o_9__770_,data_int_o_9__769_,
  data_int_o_9__768_,data_int_o_9__767_,data_int_o_9__766_,data_int_o_9__765_,
  data_int_o_9__764_,data_int_o_9__763_,data_int_o_9__762_,data_int_o_9__761_,
  data_int_o_9__760_,data_int_o_9__759_,data_int_o_9__758_,data_int_o_9__757_,
  data_int_o_9__756_,data_int_o_9__755_,data_int_o_9__754_,data_int_o_9__753_,data_int_o_9__752_,
  data_int_o_9__751_,data_int_o_9__750_,data_int_o_9__749_,data_int_o_9__748_,
  data_int_o_9__747_,data_int_o_9__746_,data_int_o_9__745_,data_int_o_9__744_,
  data_int_o_9__743_,data_int_o_9__742_,data_int_o_9__741_,data_int_o_9__740_,
  data_int_o_9__739_,data_int_o_9__738_,data_int_o_9__737_,data_int_o_9__736_,data_int_o_9__735_,
  data_int_o_9__734_,data_int_o_9__733_,data_int_o_9__732_,data_int_o_9__731_,
  data_int_o_9__730_,data_int_o_9__729_,data_int_o_9__728_,data_int_o_9__727_,
  data_int_o_9__726_,data_int_o_9__725_,data_int_o_9__724_,data_int_o_9__723_,
  data_int_o_9__722_,data_int_o_9__721_,data_int_o_9__720_,data_int_o_9__719_,
  data_int_o_9__718_,data_int_o_9__717_,data_int_o_9__716_,data_int_o_9__715_,data_int_o_9__714_,
  data_int_o_9__713_,data_int_o_9__712_,data_int_o_9__711_,data_int_o_9__710_,
  data_int_o_9__709_,data_int_o_9__708_,data_int_o_9__707_,data_int_o_9__706_,
  data_int_o_9__705_,data_int_o_9__704_,data_int_o_9__703_,data_int_o_9__702_,
  data_int_o_9__701_,data_int_o_9__700_,data_int_o_9__699_,data_int_o_9__698_,
  data_int_o_9__697_,data_int_o_9__696_,data_int_o_9__695_,data_int_o_9__694_,data_int_o_9__693_,
  data_int_o_9__692_,data_int_o_9__691_,data_int_o_9__690_,data_int_o_9__689_,
  data_int_o_9__688_,data_int_o_9__687_,data_int_o_9__686_,data_int_o_9__685_,
  data_int_o_9__684_,data_int_o_9__683_,data_int_o_9__682_,data_int_o_9__681_,
  data_int_o_9__680_,data_int_o_9__679_,data_int_o_9__678_,data_int_o_9__677_,
  data_int_o_9__676_,data_int_o_9__675_,data_int_o_9__674_,data_int_o_9__673_,data_int_o_9__672_,
  data_int_o_9__671_,data_int_o_9__670_,data_int_o_9__669_,data_int_o_9__668_,
  data_int_o_9__667_,data_int_o_9__666_,data_int_o_9__665_,data_int_o_9__664_,
  data_int_o_9__663_,data_int_o_9__662_,data_int_o_9__661_,data_int_o_9__660_,
  data_int_o_9__659_,data_int_o_9__658_,data_int_o_9__657_,data_int_o_9__656_,data_int_o_9__655_,
  data_int_o_9__654_,data_int_o_9__653_,data_int_o_9__652_,data_int_o_9__651_,
  data_int_o_9__650_,data_int_o_9__649_,data_int_o_9__648_,data_int_o_9__647_,
  data_int_o_9__646_,data_int_o_9__645_,data_int_o_9__644_,data_int_o_9__643_,
  data_int_o_9__642_,data_int_o_9__641_,data_int_o_9__640_,data_int_o_9__639_,
  data_int_o_9__638_,data_int_o_9__637_,data_int_o_9__636_,data_int_o_9__635_,data_int_o_9__634_,
  data_int_o_9__633_,data_int_o_9__632_,data_int_o_9__631_,data_int_o_9__630_,
  data_int_o_9__629_,data_int_o_9__628_,data_int_o_9__627_,data_int_o_9__626_,
  data_int_o_9__625_,data_int_o_9__624_,data_int_o_9__623_,data_int_o_9__622_,
  data_int_o_9__621_,data_int_o_9__620_,data_int_o_9__619_,data_int_o_9__618_,
  data_int_o_9__617_,data_int_o_9__616_,data_int_o_9__615_,data_int_o_9__614_,data_int_o_9__613_,
  data_int_o_9__612_,data_int_o_9__611_,data_int_o_9__610_,data_int_o_9__609_,
  data_int_o_9__608_,data_int_o_9__607_,data_int_o_9__606_,data_int_o_9__605_,
  data_int_o_9__604_,data_int_o_9__603_,data_int_o_9__602_,data_int_o_9__601_,
  data_int_o_9__600_,data_int_o_9__599_,data_int_o_9__598_,data_int_o_9__597_,
  data_int_o_9__596_,data_int_o_9__595_,data_int_o_9__594_,data_int_o_9__593_,data_int_o_9__592_,
  data_int_o_9__591_,data_int_o_9__590_,data_int_o_9__589_,data_int_o_9__588_,
  data_int_o_9__587_,data_int_o_9__586_,data_int_o_9__585_,data_int_o_9__584_,
  data_int_o_9__583_,data_int_o_9__582_,data_int_o_9__581_,data_int_o_9__580_,
  data_int_o_9__579_,data_int_o_9__578_,data_int_o_9__577_,data_int_o_9__576_,data_int_o_9__575_,
  data_int_o_9__574_,data_int_o_9__573_,data_int_o_9__572_,data_int_o_9__571_,
  data_int_o_9__570_,data_int_o_9__569_,data_int_o_9__568_,data_int_o_9__567_,
  data_int_o_9__566_,data_int_o_9__565_,data_int_o_9__564_,data_int_o_9__563_,
  data_int_o_9__562_,data_int_o_9__561_,data_int_o_9__560_,data_int_o_9__559_,
  data_int_o_9__558_,data_int_o_9__557_,data_int_o_9__556_,data_int_o_9__555_,data_int_o_9__554_,
  data_int_o_9__553_,data_int_o_9__552_,data_int_o_9__551_,data_int_o_9__550_,
  data_int_o_9__549_,data_int_o_9__548_,data_int_o_9__547_,data_int_o_9__546_,
  data_int_o_9__545_,data_int_o_9__544_,data_int_o_9__543_,data_int_o_9__542_,
  data_int_o_9__541_,data_int_o_9__540_,data_int_o_9__539_,data_int_o_9__538_,
  data_int_o_9__537_,data_int_o_9__536_,data_int_o_9__535_,data_int_o_9__534_,data_int_o_9__533_,
  data_int_o_9__532_,data_int_o_9__531_,data_int_o_9__530_,data_int_o_9__529_,
  data_int_o_9__528_,data_int_o_9__527_,data_int_o_9__526_,data_int_o_9__525_,
  data_int_o_9__524_,data_int_o_9__523_,data_int_o_9__522_,data_int_o_9__521_,
  data_int_o_9__520_,data_int_o_9__519_,data_int_o_9__518_,data_int_o_9__517_,
  data_int_o_9__516_,data_int_o_9__515_,data_int_o_9__514_,data_int_o_9__513_,data_int_o_9__512_,
  data_int_o_9__511_,data_int_o_9__510_,data_int_o_9__509_,data_int_o_9__508_,
  data_int_o_9__507_,data_int_o_9__506_,data_int_o_9__505_,data_int_o_9__504_,
  data_int_o_9__503_,data_int_o_9__502_,data_int_o_9__501_,data_int_o_9__500_,
  data_int_o_9__499_,data_int_o_9__498_,data_int_o_9__497_,data_int_o_9__496_,data_int_o_9__495_,
  data_int_o_9__494_,data_int_o_9__493_,data_int_o_9__492_,data_int_o_9__491_,
  data_int_o_9__490_,data_int_o_9__489_,data_int_o_9__488_,data_int_o_9__487_,
  data_int_o_9__486_,data_int_o_9__485_,data_int_o_9__484_,data_int_o_9__483_,
  data_int_o_9__482_,data_int_o_9__481_,data_int_o_9__480_,data_int_o_9__479_,
  data_int_o_9__478_,data_int_o_9__477_,data_int_o_9__476_,data_int_o_9__475_,data_int_o_9__474_,
  data_int_o_9__473_,data_int_o_9__472_,data_int_o_9__471_,data_int_o_9__470_,
  data_int_o_9__469_,data_int_o_9__468_,data_int_o_9__467_,data_int_o_9__466_,
  data_int_o_9__465_,data_int_o_9__464_,data_int_o_9__463_,data_int_o_9__462_,
  data_int_o_9__461_,data_int_o_9__460_,data_int_o_9__459_,data_int_o_9__458_,
  data_int_o_9__457_,data_int_o_9__456_,data_int_o_9__455_,data_int_o_9__454_,data_int_o_9__453_,
  data_int_o_9__452_,data_int_o_9__451_,data_int_o_9__450_,data_int_o_9__449_,
  data_int_o_9__448_,data_int_o_9__447_,data_int_o_9__446_,data_int_o_9__445_,
  data_int_o_9__444_,data_int_o_9__443_,data_int_o_9__442_,data_int_o_9__441_,
  data_int_o_9__440_,data_int_o_9__439_,data_int_o_9__438_,data_int_o_9__437_,
  data_int_o_9__436_,data_int_o_9__435_,data_int_o_9__434_,data_int_o_9__433_,data_int_o_9__432_,
  data_int_o_9__431_,data_int_o_9__430_,data_int_o_9__429_,data_int_o_9__428_,
  data_int_o_9__427_,data_int_o_9__426_,data_int_o_9__425_,data_int_o_9__424_,
  data_int_o_9__423_,data_int_o_9__422_,data_int_o_9__421_,data_int_o_9__420_,
  data_int_o_9__419_,data_int_o_9__418_,data_int_o_9__417_,data_int_o_9__416_,data_int_o_9__415_,
  data_int_o_9__414_,data_int_o_9__413_,data_int_o_9__412_,data_int_o_9__411_,
  data_int_o_9__410_,data_int_o_9__409_,data_int_o_9__408_,data_int_o_9__407_,
  data_int_o_9__406_,data_int_o_9__405_,data_int_o_9__404_,data_int_o_9__403_,
  data_int_o_9__402_,data_int_o_9__401_,data_int_o_9__400_,data_int_o_9__399_,
  data_int_o_9__398_,data_int_o_9__397_,data_int_o_9__396_,data_int_o_9__395_,data_int_o_9__394_,
  data_int_o_9__393_,data_int_o_9__392_,data_int_o_9__391_,data_int_o_9__390_,
  data_int_o_9__389_,data_int_o_9__388_,data_int_o_9__387_,data_int_o_9__386_,
  data_int_o_9__385_,data_int_o_9__384_,data_int_o_9__383_,data_int_o_9__382_,
  data_int_o_9__381_,data_int_o_9__380_,data_int_o_9__379_,data_int_o_9__378_,
  data_int_o_9__377_,data_int_o_9__376_,data_int_o_9__375_,data_int_o_9__374_,data_int_o_9__373_,
  data_int_o_9__372_,data_int_o_9__371_,data_int_o_9__370_,data_int_o_9__369_,
  data_int_o_9__368_,data_int_o_9__367_,data_int_o_9__366_,data_int_o_9__365_,
  data_int_o_9__364_,data_int_o_9__363_,data_int_o_9__362_,data_int_o_9__361_,
  data_int_o_9__360_,data_int_o_9__359_,data_int_o_9__358_,data_int_o_9__357_,
  data_int_o_9__356_,data_int_o_9__355_,data_int_o_9__354_,data_int_o_9__353_,data_int_o_9__352_,
  data_int_o_9__351_,data_int_o_9__350_,data_int_o_9__349_,data_int_o_9__348_,
  data_int_o_9__347_,data_int_o_9__346_,data_int_o_9__345_,data_int_o_9__344_,
  data_int_o_9__343_,data_int_o_9__342_,data_int_o_9__341_,data_int_o_9__340_,
  data_int_o_9__339_,data_int_o_9__338_,data_int_o_9__337_,data_int_o_9__336_,data_int_o_9__335_,
  data_int_o_9__334_,data_int_o_9__333_,data_int_o_9__332_,data_int_o_9__331_,
  data_int_o_9__330_,data_int_o_9__329_,data_int_o_9__328_,data_int_o_9__327_,
  data_int_o_9__326_,data_int_o_9__325_,data_int_o_9__324_,data_int_o_9__323_,
  data_int_o_9__322_,data_int_o_9__321_,data_int_o_9__320_,data_int_o_9__319_,
  data_int_o_9__318_,data_int_o_9__317_,data_int_o_9__316_,data_int_o_9__315_,data_int_o_9__314_,
  data_int_o_9__313_,data_int_o_9__312_,data_int_o_9__311_,data_int_o_9__310_,
  data_int_o_9__309_,data_int_o_9__308_,data_int_o_9__307_,data_int_o_9__306_,
  data_int_o_9__305_,data_int_o_9__304_,data_int_o_9__303_,data_int_o_9__302_,
  data_int_o_9__301_,data_int_o_9__300_,data_int_o_9__299_,data_int_o_9__298_,
  data_int_o_9__297_,data_int_o_9__296_,data_int_o_9__295_,data_int_o_9__294_,data_int_o_9__293_,
  data_int_o_9__292_,data_int_o_9__291_,data_int_o_9__290_,data_int_o_9__289_,
  data_int_o_9__288_,data_int_o_9__287_,data_int_o_9__286_,data_int_o_9__285_,
  data_int_o_9__284_,data_int_o_9__283_,data_int_o_9__282_,data_int_o_9__281_,
  data_int_o_9__280_,data_int_o_9__279_,data_int_o_9__278_,data_int_o_9__277_,
  data_int_o_9__276_,data_int_o_9__275_,data_int_o_9__274_,data_int_o_9__273_,data_int_o_9__272_,
  data_int_o_9__271_,data_int_o_9__270_,data_int_o_9__269_,data_int_o_9__268_,
  data_int_o_9__267_,data_int_o_9__266_,data_int_o_9__265_,data_int_o_9__264_,
  data_int_o_9__263_,data_int_o_9__262_,data_int_o_9__261_,data_int_o_9__260_,
  data_int_o_9__259_,data_int_o_9__258_,data_int_o_9__257_,data_int_o_9__256_,data_int_o_9__255_,
  data_int_o_9__254_,data_int_o_9__253_,data_int_o_9__252_,data_int_o_9__251_,
  data_int_o_9__250_,data_int_o_9__249_,data_int_o_9__248_,data_int_o_9__247_,
  data_int_o_9__246_,data_int_o_9__245_,data_int_o_9__244_,data_int_o_9__243_,
  data_int_o_9__242_,data_int_o_9__241_,data_int_o_9__240_,data_int_o_9__239_,
  data_int_o_9__238_,data_int_o_9__237_,data_int_o_9__236_,data_int_o_9__235_,data_int_o_9__234_,
  data_int_o_9__233_,data_int_o_9__232_,data_int_o_9__231_,data_int_o_9__230_,
  data_int_o_9__229_,data_int_o_9__228_,data_int_o_9__227_,data_int_o_9__226_,
  data_int_o_9__225_,data_int_o_9__224_,data_int_o_9__223_,data_int_o_9__222_,
  data_int_o_9__221_,data_int_o_9__220_,data_int_o_9__219_,data_int_o_9__218_,
  data_int_o_9__217_,data_int_o_9__216_,data_int_o_9__215_,data_int_o_9__214_,data_int_o_9__213_,
  data_int_o_9__212_,data_int_o_9__211_,data_int_o_9__210_,data_int_o_9__209_,
  data_int_o_9__208_,data_int_o_9__207_,data_int_o_9__206_,data_int_o_9__205_,
  data_int_o_9__204_,data_int_o_9__203_,data_int_o_9__202_,data_int_o_9__201_,
  data_int_o_9__200_,data_int_o_9__199_,data_int_o_9__198_,data_int_o_9__197_,
  data_int_o_9__196_,data_int_o_9__195_,data_int_o_9__194_,data_int_o_9__193_,data_int_o_9__192_,
  data_int_o_9__191_,data_int_o_9__190_,data_int_o_9__189_,data_int_o_9__188_,
  data_int_o_9__187_,data_int_o_9__186_,data_int_o_9__185_,data_int_o_9__184_,
  data_int_o_9__183_,data_int_o_9__182_,data_int_o_9__181_,data_int_o_9__180_,
  data_int_o_9__179_,data_int_o_9__178_,data_int_o_9__177_,data_int_o_9__176_,data_int_o_9__175_,
  data_int_o_9__174_,data_int_o_9__173_,data_int_o_9__172_,data_int_o_9__171_,
  data_int_o_9__170_,data_int_o_9__169_,data_int_o_9__168_,data_int_o_9__167_,
  data_int_o_9__166_,data_int_o_9__165_,data_int_o_9__164_,data_int_o_9__163_,
  data_int_o_9__162_,data_int_o_9__161_,data_int_o_9__160_,data_int_o_9__159_,
  data_int_o_9__158_,data_int_o_9__157_,data_int_o_9__156_,data_int_o_9__155_,data_int_o_9__154_,
  data_int_o_9__153_,data_int_o_9__152_,data_int_o_9__151_,data_int_o_9__150_,
  data_int_o_9__149_,data_int_o_9__148_,data_int_o_9__147_,data_int_o_9__146_,
  data_int_o_9__145_,data_int_o_9__144_,data_int_o_9__143_,data_int_o_9__142_,
  data_int_o_9__141_,data_int_o_9__140_,data_int_o_9__139_,data_int_o_9__138_,
  data_int_o_9__137_,data_int_o_9__136_,data_int_o_9__135_,data_int_o_9__134_,data_int_o_9__133_,
  data_int_o_9__132_,data_int_o_9__131_,data_int_o_9__130_,data_int_o_9__129_,
  data_int_o_9__128_,data_int_o_9__127_,data_int_o_9__126_,data_int_o_9__125_,
  data_int_o_9__124_,data_int_o_9__123_,data_int_o_9__122_,data_int_o_9__121_,
  data_int_o_9__120_,data_int_o_9__119_,data_int_o_9__118_,data_int_o_9__117_,
  data_int_o_9__116_,data_int_o_9__115_,data_int_o_9__114_,data_int_o_9__113_,data_int_o_9__112_,
  data_int_o_9__111_,data_int_o_9__110_,data_int_o_9__109_,data_int_o_9__108_,
  data_int_o_9__107_,data_int_o_9__106_,data_int_o_9__105_,data_int_o_9__104_,
  data_int_o_9__103_,data_int_o_9__102_,data_int_o_9__101_,data_int_o_9__100_,
  data_int_o_9__99_,data_int_o_9__98_,data_int_o_9__97_,data_int_o_9__96_,data_int_o_9__95_,
  data_int_o_9__94_,data_int_o_9__93_,data_int_o_9__92_,data_int_o_9__91_,
  data_int_o_9__90_,data_int_o_9__89_,data_int_o_9__88_,data_int_o_9__87_,data_int_o_9__86_,
  data_int_o_9__85_,data_int_o_9__84_,data_int_o_9__83_,data_int_o_9__82_,
  data_int_o_9__81_,data_int_o_9__80_,data_int_o_9__79_,data_int_o_9__78_,data_int_o_9__77_,
  data_int_o_9__76_,data_int_o_9__75_,data_int_o_9__74_,data_int_o_9__73_,
  data_int_o_9__72_,data_int_o_9__71_,data_int_o_9__70_,data_int_o_9__69_,
  data_int_o_9__68_,data_int_o_9__67_,data_int_o_9__66_,data_int_o_9__65_,data_int_o_9__64_,
  data_int_o_9__63_,data_int_o_9__62_,data_int_o_9__61_,data_int_o_9__60_,
  data_int_o_9__59_,data_int_o_9__58_,data_int_o_9__57_,data_int_o_9__56_,data_int_o_9__55_,
  data_int_o_9__54_,data_int_o_9__53_,data_int_o_9__52_,data_int_o_9__51_,
  data_int_o_9__50_,data_int_o_9__49_,data_int_o_9__48_,data_int_o_9__47_,data_int_o_9__46_,
  data_int_o_9__45_,data_int_o_9__44_,data_int_o_9__43_,data_int_o_9__42_,
  data_int_o_9__41_,data_int_o_9__40_,data_int_o_9__39_,data_int_o_9__38_,data_int_o_9__37_,
  data_int_o_9__36_,data_int_o_9__35_,data_int_o_9__34_,data_int_o_9__33_,
  data_int_o_9__32_,data_int_o_9__31_,data_int_o_9__30_,data_int_o_9__29_,
  data_int_o_9__28_,data_int_o_9__27_,data_int_o_9__26_,data_int_o_9__25_,data_int_o_9__24_,
  data_int_o_9__23_,data_int_o_9__22_,data_int_o_9__21_,data_int_o_9__20_,
  data_int_o_9__19_,data_int_o_9__18_,data_int_o_9__17_,data_int_o_9__16_,data_int_o_9__15_,
  data_int_o_9__14_,data_int_o_9__13_,data_int_o_9__12_,data_int_o_9__11_,
  data_int_o_9__10_,data_int_o_9__9_,data_int_o_9__8_,data_int_o_9__7_,data_int_o_9__6_,
  data_int_o_9__5_,data_int_o_9__4_,data_int_o_9__3_,data_int_o_9__2_,data_int_o_9__1_,
  data_int_o_9__0_,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  data_head_9__1279_,data_head_9__1278_,data_head_9__1277_,data_head_9__1276_,data_head_9__1275_,
  data_head_9__1274_,data_head_9__1273_,data_head_9__1272_,data_head_9__1271_,
  data_head_9__1270_,data_head_9__1269_,data_head_9__1268_,data_head_9__1267_,
  data_head_9__1266_,data_head_9__1265_,data_head_9__1264_,data_head_9__1263_,
  data_head_9__1262_,data_head_9__1261_,data_head_9__1260_,data_head_9__1259_,
  data_head_9__1258_,data_head_9__1257_,data_head_9__1256_,data_head_9__1255_,data_head_9__1254_,
  data_head_9__1253_,data_head_9__1252_,data_head_9__1251_,data_head_9__1250_,
  data_head_9__1249_,data_head_9__1248_,data_head_9__1247_,data_head_9__1246_,
  data_head_9__1245_,data_head_9__1244_,data_head_9__1243_,data_head_9__1242_,
  data_head_9__1241_,data_head_9__1240_,data_head_9__1239_,data_head_9__1238_,
  data_head_9__1237_,data_head_9__1236_,data_head_9__1235_,data_head_9__1234_,data_head_9__1233_,
  data_head_9__1232_,data_head_9__1231_,data_head_9__1230_,data_head_9__1229_,
  data_head_9__1228_,data_head_9__1227_,data_head_9__1226_,data_head_9__1225_,
  data_head_9__1224_,data_head_9__1223_,data_head_9__1222_,data_head_9__1221_,
  data_head_9__1220_,data_head_9__1219_,data_head_9__1218_,data_head_9__1217_,
  data_head_9__1216_,data_head_9__1215_,data_head_9__1214_,data_head_9__1213_,data_head_9__1212_,
  data_head_9__1211_,data_head_9__1210_,data_head_9__1209_,data_head_9__1208_,
  data_head_9__1207_,data_head_9__1206_,data_head_9__1205_,data_head_9__1204_,
  data_head_9__1203_,data_head_9__1202_,data_head_9__1201_,data_head_9__1200_,
  data_head_9__1199_,data_head_9__1198_,data_head_9__1197_,data_head_9__1196_,data_head_9__1195_,
  data_head_9__1194_,data_head_9__1193_,data_head_9__1192_,data_head_9__1191_,
  data_head_9__1190_,data_head_9__1189_,data_head_9__1188_,data_head_9__1187_,
  data_head_9__1186_,data_head_9__1185_,data_head_9__1184_,data_head_9__1183_,
  data_head_9__1182_,data_head_9__1181_,data_head_9__1180_,data_head_9__1179_,
  data_head_9__1178_,data_head_9__1177_,data_head_9__1176_,data_head_9__1175_,data_head_9__1174_,
  data_head_9__1173_,data_head_9__1172_,data_head_9__1171_,data_head_9__1170_,
  data_head_9__1169_,data_head_9__1168_,data_head_9__1167_,data_head_9__1166_,
  data_head_9__1165_,data_head_9__1164_,data_head_9__1163_,data_head_9__1162_,
  data_head_9__1161_,data_head_9__1160_,data_head_9__1159_,data_head_9__1158_,
  data_head_9__1157_,data_head_9__1156_,data_head_9__1155_,data_head_9__1154_,data_head_9__1153_,
  data_head_9__1152_,data_head_9__1151_,data_head_9__1150_,data_head_9__1149_,
  data_head_9__1148_,data_head_9__1147_,data_head_9__1146_,data_head_9__1145_,
  data_head_9__1144_,data_head_9__1143_,data_head_9__1142_,data_head_9__1141_,
  data_head_9__1140_,data_head_9__1139_,data_head_9__1138_,data_head_9__1137_,
  data_head_9__1136_,data_head_9__1135_,data_head_9__1134_,data_head_9__1133_,data_head_9__1132_,
  data_head_9__1131_,data_head_9__1130_,data_head_9__1129_,data_head_9__1128_,
  data_head_9__1127_,data_head_9__1126_,data_head_9__1125_,data_head_9__1124_,
  data_head_9__1123_,data_head_9__1122_,data_head_9__1121_,data_head_9__1120_,
  data_head_9__1119_,data_head_9__1118_,data_head_9__1117_,data_head_9__1116_,data_head_9__1115_,
  data_head_9__1114_,data_head_9__1113_,data_head_9__1112_,data_head_9__1111_,
  data_head_9__1110_,data_head_9__1109_,data_head_9__1108_,data_head_9__1107_,
  data_head_9__1106_,data_head_9__1105_,data_head_9__1104_,data_head_9__1103_,
  data_head_9__1102_,data_head_9__1101_,data_head_9__1100_,data_head_9__1099_,
  data_head_9__1098_,data_head_9__1097_,data_head_9__1096_,data_head_9__1095_,data_head_9__1094_,
  data_head_9__1093_,data_head_9__1092_,data_head_9__1091_,data_head_9__1090_,
  data_head_9__1089_,data_head_9__1088_,data_head_9__1087_,data_head_9__1086_,
  data_head_9__1085_,data_head_9__1084_,data_head_9__1083_,data_head_9__1082_,
  data_head_9__1081_,data_head_9__1080_,data_head_9__1079_,data_head_9__1078_,
  data_head_9__1077_,data_head_9__1076_,data_head_9__1075_,data_head_9__1074_,data_head_9__1073_,
  data_head_9__1072_,data_head_9__1071_,data_head_9__1070_,data_head_9__1069_,
  data_head_9__1068_,data_head_9__1067_,data_head_9__1066_,data_head_9__1065_,
  data_head_9__1064_,data_head_9__1063_,data_head_9__1062_,data_head_9__1061_,
  data_head_9__1060_,data_head_9__1059_,data_head_9__1058_,data_head_9__1057_,
  data_head_9__1056_,data_head_9__1055_,data_head_9__1054_,data_head_9__1053_,data_head_9__1052_,
  data_head_9__1051_,data_head_9__1050_,data_head_9__1049_,data_head_9__1048_,
  data_head_9__1047_,data_head_9__1046_,data_head_9__1045_,data_head_9__1044_,
  data_head_9__1043_,data_head_9__1042_,data_head_9__1041_,data_head_9__1040_,
  data_head_9__1039_,data_head_9__1038_,data_head_9__1037_,data_head_9__1036_,data_head_9__1035_,
  data_head_9__1034_,data_head_9__1033_,data_head_9__1032_,data_head_9__1031_,
  data_head_9__1030_,data_head_9__1029_,data_head_9__1028_,data_head_9__1027_,
  data_head_9__1026_,data_head_9__1025_,data_head_9__1024_,data_head_9__1023_,
  data_head_9__1022_,data_head_9__1021_,data_head_9__1020_,data_head_9__1019_,
  data_head_9__1018_,data_head_9__1017_,data_head_9__1016_,data_head_9__1015_,data_head_9__1014_,
  data_head_9__1013_,data_head_9__1012_,data_head_9__1011_,data_head_9__1010_,
  data_head_9__1009_,data_head_9__1008_,data_head_9__1007_,data_head_9__1006_,
  data_head_9__1005_,data_head_9__1004_,data_head_9__1003_,data_head_9__1002_,
  data_head_9__1001_,data_head_9__1000_,data_head_9__999_,data_head_9__998_,data_head_9__997_,
  data_head_9__996_,data_head_9__995_,data_head_9__994_,data_head_9__993_,
  data_head_9__992_,data_head_9__991_,data_head_9__990_,data_head_9__989_,
  data_head_9__988_,data_head_9__987_,data_head_9__986_,data_head_9__985_,data_head_9__984_,
  data_head_9__983_,data_head_9__982_,data_head_9__981_,data_head_9__980_,
  data_head_9__979_,data_head_9__978_,data_head_9__977_,data_head_9__976_,data_head_9__975_,
  data_head_9__974_,data_head_9__973_,data_head_9__972_,data_head_9__971_,
  data_head_9__970_,data_head_9__969_,data_head_9__968_,data_head_9__967_,data_head_9__966_,
  data_head_9__965_,data_head_9__964_,data_head_9__963_,data_head_9__962_,
  data_head_9__961_,data_head_9__960_,data_head_9__959_,data_head_9__958_,data_head_9__957_,
  data_head_9__956_,data_head_9__955_,data_head_9__954_,data_head_9__953_,
  data_head_9__952_,data_head_9__951_,data_head_9__950_,data_head_9__949_,
  data_head_9__948_,data_head_9__947_,data_head_9__946_,data_head_9__945_,data_head_9__944_,
  data_head_9__943_,data_head_9__942_,data_head_9__941_,data_head_9__940_,
  data_head_9__939_,data_head_9__938_,data_head_9__937_,data_head_9__936_,data_head_9__935_,
  data_head_9__934_,data_head_9__933_,data_head_9__932_,data_head_9__931_,
  data_head_9__930_,data_head_9__929_,data_head_9__928_,data_head_9__927_,data_head_9__926_,
  data_head_9__925_,data_head_9__924_,data_head_9__923_,data_head_9__922_,
  data_head_9__921_,data_head_9__920_,data_head_9__919_,data_head_9__918_,data_head_9__917_,
  data_head_9__916_,data_head_9__915_,data_head_9__914_,data_head_9__913_,
  data_head_9__912_,data_head_9__911_,data_head_9__910_,data_head_9__909_,
  data_head_9__908_,data_head_9__907_,data_head_9__906_,data_head_9__905_,data_head_9__904_,
  data_head_9__903_,data_head_9__902_,data_head_9__901_,data_head_9__900_,
  data_head_9__899_,data_head_9__898_,data_head_9__897_,data_head_9__896_,data_head_9__895_,
  data_head_9__894_,data_head_9__893_,data_head_9__892_,data_head_9__891_,
  data_head_9__890_,data_head_9__889_,data_head_9__888_,data_head_9__887_,data_head_9__886_,
  data_head_9__885_,data_head_9__884_,data_head_9__883_,data_head_9__882_,
  data_head_9__881_,data_head_9__880_,data_head_9__879_,data_head_9__878_,data_head_9__877_,
  data_head_9__876_,data_head_9__875_,data_head_9__874_,data_head_9__873_,
  data_head_9__872_,data_head_9__871_,data_head_9__870_,data_head_9__869_,
  data_head_9__868_,data_head_9__867_,data_head_9__866_,data_head_9__865_,data_head_9__864_,
  data_head_9__863_,data_head_9__862_,data_head_9__861_,data_head_9__860_,
  data_head_9__859_,data_head_9__858_,data_head_9__857_,data_head_9__856_,data_head_9__855_,
  data_head_9__854_,data_head_9__853_,data_head_9__852_,data_head_9__851_,
  data_head_9__850_,data_head_9__849_,data_head_9__848_,data_head_9__847_,data_head_9__846_,
  data_head_9__845_,data_head_9__844_,data_head_9__843_,data_head_9__842_,
  data_head_9__841_,data_head_9__840_,data_head_9__839_,data_head_9__838_,data_head_9__837_,
  data_head_9__836_,data_head_9__835_,data_head_9__834_,data_head_9__833_,
  data_head_9__832_,data_head_9__831_,data_head_9__830_,data_head_9__829_,
  data_head_9__828_,data_head_9__827_,data_head_9__826_,data_head_9__825_,data_head_9__824_,
  data_head_9__823_,data_head_9__822_,data_head_9__821_,data_head_9__820_,
  data_head_9__819_,data_head_9__818_,data_head_9__817_,data_head_9__816_,data_head_9__815_,
  data_head_9__814_,data_head_9__813_,data_head_9__812_,data_head_9__811_,
  data_head_9__810_,data_head_9__809_,data_head_9__808_,data_head_9__807_,data_head_9__806_,
  data_head_9__805_,data_head_9__804_,data_head_9__803_,data_head_9__802_,
  data_head_9__801_,data_head_9__800_,data_head_9__799_,data_head_9__798_,data_head_9__797_,
  data_head_9__796_,data_head_9__795_,data_head_9__794_,data_head_9__793_,
  data_head_9__792_,data_head_9__791_,data_head_9__790_,data_head_9__789_,
  data_head_9__788_,data_head_9__787_,data_head_9__786_,data_head_9__785_,data_head_9__784_,
  data_head_9__783_,data_head_9__782_,data_head_9__781_,data_head_9__780_,
  data_head_9__779_,data_head_9__778_,data_head_9__777_,data_head_9__776_,data_head_9__775_,
  data_head_9__774_,data_head_9__773_,data_head_9__772_,data_head_9__771_,
  data_head_9__770_,data_head_9__769_,data_head_9__768_,data_head_9__767_,data_head_9__766_,
  data_head_9__765_,data_head_9__764_,data_head_9__763_,data_head_9__762_,
  data_head_9__761_,data_head_9__760_,data_head_9__759_,data_head_9__758_,data_head_9__757_,
  data_head_9__756_,data_head_9__755_,data_head_9__754_,data_head_9__753_,
  data_head_9__752_,data_head_9__751_,data_head_9__750_,data_head_9__749_,
  data_head_9__748_,data_head_9__747_,data_head_9__746_,data_head_9__745_,data_head_9__744_,
  data_head_9__743_,data_head_9__742_,data_head_9__741_,data_head_9__740_,
  data_head_9__739_,data_head_9__738_,data_head_9__737_,data_head_9__736_,data_head_9__735_,
  data_head_9__734_,data_head_9__733_,data_head_9__732_,data_head_9__731_,
  data_head_9__730_,data_head_9__729_,data_head_9__728_,data_head_9__727_,data_head_9__726_,
  data_head_9__725_,data_head_9__724_,data_head_9__723_,data_head_9__722_,
  data_head_9__721_,data_head_9__720_,data_head_9__719_,data_head_9__718_,data_head_9__717_,
  data_head_9__716_,data_head_9__715_,data_head_9__714_,data_head_9__713_,
  data_head_9__712_,data_head_9__711_,data_head_9__710_,data_head_9__709_,
  data_head_9__708_,data_head_9__707_,data_head_9__706_,data_head_9__705_,data_head_9__704_,
  data_head_9__703_,data_head_9__702_,data_head_9__701_,data_head_9__700_,
  data_head_9__699_,data_head_9__698_,data_head_9__697_,data_head_9__696_,data_head_9__695_,
  data_head_9__694_,data_head_9__693_,data_head_9__692_,data_head_9__691_,
  data_head_9__690_,data_head_9__689_,data_head_9__688_,data_head_9__687_,data_head_9__686_,
  data_head_9__685_,data_head_9__684_,data_head_9__683_,data_head_9__682_,
  data_head_9__681_,data_head_9__680_,data_head_9__679_,data_head_9__678_,data_head_9__677_,
  data_head_9__676_,data_head_9__675_,data_head_9__674_,data_head_9__673_,
  data_head_9__672_,data_head_9__671_,data_head_9__670_,data_head_9__669_,
  data_head_9__668_,data_head_9__667_,data_head_9__666_,data_head_9__665_,data_head_9__664_,
  data_head_9__663_,data_head_9__662_,data_head_9__661_,data_head_9__660_,
  data_head_9__659_,data_head_9__658_,data_head_9__657_,data_head_9__656_,data_head_9__655_,
  data_head_9__654_,data_head_9__653_,data_head_9__652_,data_head_9__651_,
  data_head_9__650_,data_head_9__649_,data_head_9__648_,data_head_9__647_,data_head_9__646_,
  data_head_9__645_,data_head_9__644_,data_head_9__643_,data_head_9__642_,
  data_head_9__641_,data_head_9__640_,data_head_9__639_,data_head_9__638_,data_head_9__637_,
  data_head_9__636_,data_head_9__635_,data_head_9__634_,data_head_9__633_,
  data_head_9__632_,data_head_9__631_,data_head_9__630_,data_head_9__629_,
  data_head_9__628_,data_head_9__627_,data_head_9__626_,data_head_9__625_,data_head_9__624_,
  data_head_9__623_,data_head_9__622_,data_head_9__621_,data_head_9__620_,
  data_head_9__619_,data_head_9__618_,data_head_9__617_,data_head_9__616_,data_head_9__615_,
  data_head_9__614_,data_head_9__613_,data_head_9__612_,data_head_9__611_,
  data_head_9__610_,data_head_9__609_,data_head_9__608_,data_head_9__607_,data_head_9__606_,
  data_head_9__605_,data_head_9__604_,data_head_9__603_,data_head_9__602_,
  data_head_9__601_,data_head_9__600_,data_head_9__599_,data_head_9__598_,data_head_9__597_,
  data_head_9__596_,data_head_9__595_,data_head_9__594_,data_head_9__593_,
  data_head_9__592_,data_head_9__591_,data_head_9__590_,data_head_9__589_,
  data_head_9__588_,data_head_9__587_,data_head_9__586_,data_head_9__585_,data_head_9__584_,
  data_head_9__583_,data_head_9__582_,data_head_9__581_,data_head_9__580_,
  data_head_9__579_,data_head_9__578_,data_head_9__577_,data_head_9__576_,data_head_9__575_,
  data_head_9__574_,data_head_9__573_,data_head_9__572_,data_head_9__571_,
  data_head_9__570_,data_head_9__569_,data_head_9__568_,data_head_9__567_,data_head_9__566_,
  data_head_9__565_,data_head_9__564_,data_head_9__563_,data_head_9__562_,
  data_head_9__561_,data_head_9__560_,data_head_9__559_,data_head_9__558_,data_head_9__557_,
  data_head_9__556_,data_head_9__555_,data_head_9__554_,data_head_9__553_,
  data_head_9__552_,data_head_9__551_,data_head_9__550_,data_head_9__549_,
  data_head_9__548_,data_head_9__547_,data_head_9__546_,data_head_9__545_,data_head_9__544_,
  data_head_9__543_,data_head_9__542_,data_head_9__541_,data_head_9__540_,
  data_head_9__539_,data_head_9__538_,data_head_9__537_,data_head_9__536_,data_head_9__535_,
  data_head_9__534_,data_head_9__533_,data_head_9__532_,data_head_9__531_,
  data_head_9__530_,data_head_9__529_,data_head_9__528_,data_head_9__527_,data_head_9__526_,
  data_head_9__525_,data_head_9__524_,data_head_9__523_,data_head_9__522_,
  data_head_9__521_,data_head_9__520_,data_head_9__519_,data_head_9__518_,data_head_9__517_,
  data_head_9__516_,data_head_9__515_,data_head_9__514_,data_head_9__513_,
  data_head_9__512_,data_head_9__511_,data_head_9__510_,data_head_9__509_,
  data_head_9__508_,data_head_9__507_,data_head_9__506_,data_head_9__505_,data_head_9__504_,
  data_head_9__503_,data_head_9__502_,data_head_9__501_,data_head_9__500_,
  data_head_9__499_,data_head_9__498_,data_head_9__497_,data_head_9__496_,data_head_9__495_,
  data_head_9__494_,data_head_9__493_,data_head_9__492_,data_head_9__491_,
  data_head_9__490_,data_head_9__489_,data_head_9__488_,data_head_9__487_,data_head_9__486_,
  data_head_9__485_,data_head_9__484_,data_head_9__483_,data_head_9__482_,
  data_head_9__481_,data_head_9__480_,data_head_9__479_,data_head_9__478_,data_head_9__477_,
  data_head_9__476_,data_head_9__475_,data_head_9__474_,data_head_9__473_,
  data_head_9__472_,data_head_9__471_,data_head_9__470_,data_head_9__469_,
  data_head_9__468_,data_head_9__467_,data_head_9__466_,data_head_9__465_,data_head_9__464_,
  data_head_9__463_,data_head_9__462_,data_head_9__461_,data_head_9__460_,
  data_head_9__459_,data_head_9__458_,data_head_9__457_,data_head_9__456_,data_head_9__455_,
  data_head_9__454_,data_head_9__453_,data_head_9__452_,data_head_9__451_,
  data_head_9__450_,data_head_9__449_,data_head_9__448_,data_head_9__447_,data_head_9__446_,
  data_head_9__445_,data_head_9__444_,data_head_9__443_,data_head_9__442_,
  data_head_9__441_,data_head_9__440_,data_head_9__439_,data_head_9__438_,data_head_9__437_,
  data_head_9__436_,data_head_9__435_,data_head_9__434_,data_head_9__433_,
  data_head_9__432_,data_head_9__431_,data_head_9__430_,data_head_9__429_,
  data_head_9__428_,data_head_9__427_,data_head_9__426_,data_head_9__425_,data_head_9__424_,
  data_head_9__423_,data_head_9__422_,data_head_9__421_,data_head_9__420_,
  data_head_9__419_,data_head_9__418_,data_head_9__417_,data_head_9__416_,data_head_9__415_,
  data_head_9__414_,data_head_9__413_,data_head_9__412_,data_head_9__411_,
  data_head_9__410_,data_head_9__409_,data_head_9__408_,data_head_9__407_,data_head_9__406_,
  data_head_9__405_,data_head_9__404_,data_head_9__403_,data_head_9__402_,
  data_head_9__401_,data_head_9__400_,data_head_9__399_,data_head_9__398_,data_head_9__397_,
  data_head_9__396_,data_head_9__395_,data_head_9__394_,data_head_9__393_,
  data_head_9__392_,data_head_9__391_,data_head_9__390_,data_head_9__389_,
  data_head_9__388_,data_head_9__387_,data_head_9__386_,data_head_9__385_,data_head_9__384_,
  data_head_9__383_,data_head_9__382_,data_head_9__381_,data_head_9__380_,
  data_head_9__379_,data_head_9__378_,data_head_9__377_,data_head_9__376_,data_head_9__375_,
  data_head_9__374_,data_head_9__373_,data_head_9__372_,data_head_9__371_,
  data_head_9__370_,data_head_9__369_,data_head_9__368_,data_head_9__367_,data_head_9__366_,
  data_head_9__365_,data_head_9__364_,data_head_9__363_,data_head_9__362_,
  data_head_9__361_,data_head_9__360_,data_head_9__359_,data_head_9__358_,data_head_9__357_,
  data_head_9__356_,data_head_9__355_,data_head_9__354_,data_head_9__353_,
  data_head_9__352_,data_head_9__351_,data_head_9__350_,data_head_9__349_,
  data_head_9__348_,data_head_9__347_,data_head_9__346_,data_head_9__345_,data_head_9__344_,
  data_head_9__343_,data_head_9__342_,data_head_9__341_,data_head_9__340_,
  data_head_9__339_,data_head_9__338_,data_head_9__337_,data_head_9__336_,data_head_9__335_,
  data_head_9__334_,data_head_9__333_,data_head_9__332_,data_head_9__331_,
  data_head_9__330_,data_head_9__329_,data_head_9__328_,data_head_9__327_,data_head_9__326_,
  data_head_9__325_,data_head_9__324_,data_head_9__323_,data_head_9__322_,
  data_head_9__321_,data_head_9__320_,data_head_9__319_,data_head_9__318_,data_head_9__317_,
  data_head_9__316_,data_head_9__315_,data_head_9__314_,data_head_9__313_,
  data_head_9__312_,data_head_9__311_,data_head_9__310_,data_head_9__309_,
  data_head_9__308_,data_head_9__307_,data_head_9__306_,data_head_9__305_,data_head_9__304_,
  data_head_9__303_,data_head_9__302_,data_head_9__301_,data_head_9__300_,
  data_head_9__299_,data_head_9__298_,data_head_9__297_,data_head_9__296_,data_head_9__295_,
  data_head_9__294_,data_head_9__293_,data_head_9__292_,data_head_9__291_,
  data_head_9__290_,data_head_9__289_,data_head_9__288_,data_head_9__287_,data_head_9__286_,
  data_head_9__285_,data_head_9__284_,data_head_9__283_,data_head_9__282_,
  data_head_9__281_,data_head_9__280_,data_head_9__279_,data_head_9__278_,data_head_9__277_,
  data_head_9__276_,data_head_9__275_,data_head_9__274_,data_head_9__273_,
  data_head_9__272_,data_head_9__271_,data_head_9__270_,data_head_9__269_,
  data_head_9__268_,data_head_9__267_,data_head_9__266_,data_head_9__265_,data_head_9__264_,
  data_head_9__263_,data_head_9__262_,data_head_9__261_,data_head_9__260_,
  data_head_9__259_,data_head_9__258_,data_head_9__257_,data_head_9__256_,data_head_9__255_,
  data_head_9__254_,data_head_9__253_,data_head_9__252_,data_head_9__251_,
  data_head_9__250_,data_head_9__249_,data_head_9__248_,data_head_9__247_,data_head_9__246_,
  data_head_9__245_,data_head_9__244_,data_head_9__243_,data_head_9__242_,
  data_head_9__241_,data_head_9__240_,data_head_9__239_,data_head_9__238_,data_head_9__237_,
  data_head_9__236_,data_head_9__235_,data_head_9__234_,data_head_9__233_,
  data_head_9__232_,data_head_9__231_,data_head_9__230_,data_head_9__229_,
  data_head_9__228_,data_head_9__227_,data_head_9__226_,data_head_9__225_,data_head_9__224_,
  data_head_9__223_,data_head_9__222_,data_head_9__221_,data_head_9__220_,
  data_head_9__219_,data_head_9__218_,data_head_9__217_,data_head_9__216_,data_head_9__215_,
  data_head_9__214_,data_head_9__213_,data_head_9__212_,data_head_9__211_,
  data_head_9__210_,data_head_9__209_,data_head_9__208_,data_head_9__207_,data_head_9__206_,
  data_head_9__205_,data_head_9__204_,data_head_9__203_,data_head_9__202_,
  data_head_9__201_,data_head_9__200_,data_head_9__199_,data_head_9__198_,data_head_9__197_,
  data_head_9__196_,data_head_9__195_,data_head_9__194_,data_head_9__193_,
  data_head_9__192_,data_head_9__191_,data_head_9__190_,data_head_9__189_,
  data_head_9__188_,data_head_9__187_,data_head_9__186_,data_head_9__185_,data_head_9__184_,
  data_head_9__183_,data_head_9__182_,data_head_9__181_,data_head_9__180_,
  data_head_9__179_,data_head_9__178_,data_head_9__177_,data_head_9__176_,data_head_9__175_,
  data_head_9__174_,data_head_9__173_,data_head_9__172_,data_head_9__171_,
  data_head_9__170_,data_head_9__169_,data_head_9__168_,data_head_9__167_,data_head_9__166_,
  data_head_9__165_,data_head_9__164_,data_head_9__163_,data_head_9__162_,
  data_head_9__161_,data_head_9__160_,data_head_9__159_,data_head_9__158_,data_head_9__157_,
  data_head_9__156_,data_head_9__155_,data_head_9__154_,data_head_9__153_,
  data_head_9__152_,data_head_9__151_,data_head_9__150_,data_head_9__149_,
  data_head_9__148_,data_head_9__147_,data_head_9__146_,data_head_9__145_,data_head_9__144_,
  data_head_9__143_,data_head_9__142_,data_head_9__141_,data_head_9__140_,
  data_head_9__139_,data_head_9__138_,data_head_9__137_,data_head_9__136_,data_head_9__135_,
  data_head_9__134_,data_head_9__133_,data_head_9__132_,data_head_9__131_,
  data_head_9__130_,data_head_9__129_,data_head_9__128_,data_head_9__127_,data_head_9__126_,
  data_head_9__125_,data_head_9__124_,data_head_9__123_,data_head_9__122_,
  data_head_9__121_,data_head_9__120_,data_head_9__119_,data_head_9__118_,data_head_9__117_,
  data_head_9__116_,data_head_9__115_,data_head_9__114_,data_head_9__113_,
  data_head_9__112_,data_head_9__111_,data_head_9__110_,data_head_9__109_,
  data_head_9__108_,data_head_9__107_,data_head_9__106_,data_head_9__105_,data_head_9__104_,
  data_head_9__103_,data_head_9__102_,data_head_9__101_,data_head_9__100_,
  data_head_9__99_,data_head_9__98_,data_head_9__97_,data_head_9__96_,data_head_9__95_,
  data_head_9__94_,data_head_9__93_,data_head_9__92_,data_head_9__91_,data_head_9__90_,
  data_head_9__89_,data_head_9__88_,data_head_9__87_,data_head_9__86_,data_head_9__85_,
  data_head_9__84_,data_head_9__83_,data_head_9__82_,data_head_9__81_,
  data_head_9__80_,data_head_9__79_,data_head_9__78_,data_head_9__77_,data_head_9__76_,
  data_head_9__75_,data_head_9__74_,data_head_9__73_,data_head_9__72_,data_head_9__71_,
  data_head_9__70_,data_head_9__69_,data_head_9__68_,data_head_9__67_,
  data_head_9__66_,data_head_9__65_,data_head_9__64_,data_head_9__63_,data_head_9__62_,
  data_head_9__61_,data_head_9__60_,data_head_9__59_,data_head_9__58_,data_head_9__57_,
  data_head_9__56_,data_head_9__55_,data_head_9__54_,data_head_9__53_,
  data_head_9__52_,data_head_9__51_,data_head_9__50_,data_head_9__49_,data_head_9__48_,
  data_head_9__47_,data_head_9__46_,data_head_9__45_,data_head_9__44_,data_head_9__43_,
  data_head_9__42_,data_head_9__41_,data_head_9__40_,data_head_9__39_,data_head_9__38_,
  data_head_9__37_,data_head_9__36_,data_head_9__35_,data_head_9__34_,
  data_head_9__33_,data_head_9__32_,data_head_9__31_,data_head_9__30_,data_head_9__29_,
  data_head_9__28_,data_head_9__27_,data_head_9__26_,data_head_9__25_,data_head_9__24_,
  data_head_9__23_,data_head_9__22_,data_head_9__21_,data_head_9__20_,
  data_head_9__19_,data_head_9__18_,data_head_9__17_,data_head_9__16_,data_head_9__15_,
  data_head_9__14_,data_head_9__13_,data_head_9__12_,data_head_9__11_,data_head_9__10_,
  data_head_9__9_,data_head_9__8_,data_head_9__7_,data_head_9__6_,data_head_9__5_,
  data_head_9__4_,data_head_9__3_,data_head_9__2_,data_head_9__1_,data_head_9__0_,
  n_0_net_,valid_head_9__9_,valid_head_9__8_,valid_head_9__7_,valid_head_9__6_,
  valid_head_9__5_,valid_head_9__4_,valid_head_9__3_,valid_head_9__2_,valid_head_9__1_,
  valid_head_9__0_,n_2_net__9_,n_2_net__8_,n_2_net__7_,n_2_net__6_,n_2_net__5_,
  n_2_net__4_,n_2_net__3_,n_2_net__2_,n_2_net__1_,n_2_net__0_,n_3_net__9_,n_3_net__8_,
  n_3_net__7_,n_3_net__6_,n_3_net__5_,n_3_net__4_,n_3_net__3_,n_3_net__2_,
  n_3_net__1_,n_3_net__0_,ready_head_9__9_,ready_head_9__8_,ready_head_9__7_,
  ready_head_9__6_,ready_head_9__5_,ready_head_9__4_,ready_head_9__3_,ready_head_9__2_,
  ready_head_9__1_,ready_head_9__0_,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  n_4_net__1279_,n_4_net__1278_,n_4_net__1277_,n_4_net__1276_,n_4_net__1275_,
  n_4_net__1274_,n_4_net__1273_,n_4_net__1272_,n_4_net__1271_,n_4_net__1270_,n_4_net__1269_,
  n_4_net__1268_,n_4_net__1267_,n_4_net__1266_,n_4_net__1265_,n_4_net__1264_,
  n_4_net__1263_,n_4_net__1262_,n_4_net__1261_,n_4_net__1260_,n_4_net__1259_,
  n_4_net__1258_,n_4_net__1257_,n_4_net__1256_,n_4_net__1255_,n_4_net__1254_,n_4_net__1253_,
  n_4_net__1252_,n_4_net__1251_,n_4_net__1250_,n_4_net__1249_,n_4_net__1248_,
  n_4_net__1247_,n_4_net__1246_,n_4_net__1245_,n_4_net__1244_,n_4_net__1243_,
  n_4_net__1242_,n_4_net__1241_,n_4_net__1240_,n_4_net__1239_,n_4_net__1238_,n_4_net__1237_,
  n_4_net__1236_,n_4_net__1235_,n_4_net__1234_,n_4_net__1233_,n_4_net__1232_,
  n_4_net__1231_,n_4_net__1230_,n_4_net__1229_,n_4_net__1228_,n_4_net__1227_,
  n_4_net__1226_,n_4_net__1225_,n_4_net__1224_,n_4_net__1223_,n_4_net__1222_,n_4_net__1221_,
  n_4_net__1220_,n_4_net__1219_,n_4_net__1218_,n_4_net__1217_,n_4_net__1216_,
  n_4_net__1215_,n_4_net__1214_,n_4_net__1213_,n_4_net__1212_,n_4_net__1211_,
  n_4_net__1210_,n_4_net__1209_,n_4_net__1208_,n_4_net__1207_,n_4_net__1206_,n_4_net__1205_,
  n_4_net__1204_,n_4_net__1203_,n_4_net__1202_,n_4_net__1201_,n_4_net__1200_,
  n_4_net__1199_,n_4_net__1198_,n_4_net__1197_,n_4_net__1196_,n_4_net__1195_,
  n_4_net__1194_,n_4_net__1193_,n_4_net__1192_,n_4_net__1191_,n_4_net__1190_,n_4_net__1189_,
  n_4_net__1188_,n_4_net__1187_,n_4_net__1186_,n_4_net__1185_,n_4_net__1184_,
  n_4_net__1183_,n_4_net__1182_,n_4_net__1181_,n_4_net__1180_,n_4_net__1179_,
  n_4_net__1178_,n_4_net__1177_,n_4_net__1176_,n_4_net__1175_,n_4_net__1174_,n_4_net__1173_,
  n_4_net__1172_,n_4_net__1171_,n_4_net__1170_,n_4_net__1169_,n_4_net__1168_,
  n_4_net__1167_,n_4_net__1166_,n_4_net__1165_,n_4_net__1164_,n_4_net__1163_,
  n_4_net__1162_,n_4_net__1161_,n_4_net__1160_,n_4_net__1159_,n_4_net__1158_,n_4_net__1157_,
  n_4_net__1156_,n_4_net__1155_,n_4_net__1154_,n_4_net__1153_,n_4_net__1152_,
  n_4_net__1151_,n_4_net__1150_,n_4_net__1149_,n_4_net__1148_,n_4_net__1147_,
  n_4_net__1146_,n_4_net__1145_,n_4_net__1144_,n_4_net__1143_,n_4_net__1142_,n_4_net__1141_,
  n_4_net__1140_,n_4_net__1139_,n_4_net__1138_,n_4_net__1137_,n_4_net__1136_,
  n_4_net__1135_,n_4_net__1134_,n_4_net__1133_,n_4_net__1132_,n_4_net__1131_,
  n_4_net__1130_,n_4_net__1129_,n_4_net__1128_,n_4_net__1127_,n_4_net__1126_,n_4_net__1125_,
  n_4_net__1124_,n_4_net__1123_,n_4_net__1122_,n_4_net__1121_,n_4_net__1120_,
  n_4_net__1119_,n_4_net__1118_,n_4_net__1117_,n_4_net__1116_,n_4_net__1115_,
  n_4_net__1114_,n_4_net__1113_,n_4_net__1112_,n_4_net__1111_,n_4_net__1110_,n_4_net__1109_,
  n_4_net__1108_,n_4_net__1107_,n_4_net__1106_,n_4_net__1105_,n_4_net__1104_,
  n_4_net__1103_,n_4_net__1102_,n_4_net__1101_,n_4_net__1100_,n_4_net__1099_,
  n_4_net__1098_,n_4_net__1097_,n_4_net__1096_,n_4_net__1095_,n_4_net__1094_,n_4_net__1093_,
  n_4_net__1092_,n_4_net__1091_,n_4_net__1090_,n_4_net__1089_,n_4_net__1088_,
  n_4_net__1087_,n_4_net__1086_,n_4_net__1085_,n_4_net__1084_,n_4_net__1083_,
  n_4_net__1082_,n_4_net__1081_,n_4_net__1080_,n_4_net__1079_,n_4_net__1078_,n_4_net__1077_,
  n_4_net__1076_,n_4_net__1075_,n_4_net__1074_,n_4_net__1073_,n_4_net__1072_,
  n_4_net__1071_,n_4_net__1070_,n_4_net__1069_,n_4_net__1068_,n_4_net__1067_,
  n_4_net__1066_,n_4_net__1065_,n_4_net__1064_,n_4_net__1063_,n_4_net__1062_,n_4_net__1061_,
  n_4_net__1060_,n_4_net__1059_,n_4_net__1058_,n_4_net__1057_,n_4_net__1056_,
  n_4_net__1055_,n_4_net__1054_,n_4_net__1053_,n_4_net__1052_,n_4_net__1051_,
  n_4_net__1050_,n_4_net__1049_,n_4_net__1048_,n_4_net__1047_,n_4_net__1046_,n_4_net__1045_,
  n_4_net__1044_,n_4_net__1043_,n_4_net__1042_,n_4_net__1041_,n_4_net__1040_,
  n_4_net__1039_,n_4_net__1038_,n_4_net__1037_,n_4_net__1036_,n_4_net__1035_,
  n_4_net__1034_,n_4_net__1033_,n_4_net__1032_,n_4_net__1031_,n_4_net__1030_,n_4_net__1029_,
  n_4_net__1028_,n_4_net__1027_,n_4_net__1026_,n_4_net__1025_,n_4_net__1024_,
  n_4_net__1023_,n_4_net__1022_,n_4_net__1021_,n_4_net__1020_,n_4_net__1019_,
  n_4_net__1018_,n_4_net__1017_,n_4_net__1016_,n_4_net__1015_,n_4_net__1014_,n_4_net__1013_,
  n_4_net__1012_,n_4_net__1011_,n_4_net__1010_,n_4_net__1009_,n_4_net__1008_,
  n_4_net__1007_,n_4_net__1006_,n_4_net__1005_,n_4_net__1004_,n_4_net__1003_,
  n_4_net__1002_,n_4_net__1001_,n_4_net__1000_,n_4_net__999_,n_4_net__998_,n_4_net__997_,
  n_4_net__996_,n_4_net__995_,n_4_net__994_,n_4_net__993_,n_4_net__992_,n_4_net__991_,
  n_4_net__990_,n_4_net__989_,n_4_net__988_,n_4_net__987_,n_4_net__986_,
  n_4_net__985_,n_4_net__984_,n_4_net__983_,n_4_net__982_,n_4_net__981_,n_4_net__980_,
  n_4_net__979_,n_4_net__978_,n_4_net__977_,n_4_net__976_,n_4_net__975_,n_4_net__974_,
  n_4_net__973_,n_4_net__972_,n_4_net__971_,n_4_net__970_,n_4_net__969_,
  n_4_net__968_,n_4_net__967_,n_4_net__966_,n_4_net__965_,n_4_net__964_,n_4_net__963_,
  n_4_net__962_,n_4_net__961_,n_4_net__960_,n_4_net__959_,n_4_net__958_,n_4_net__957_,
  n_4_net__956_,n_4_net__955_,n_4_net__954_,n_4_net__953_,n_4_net__952_,n_4_net__951_,
  n_4_net__950_,n_4_net__949_,n_4_net__948_,n_4_net__947_,n_4_net__946_,
  n_4_net__945_,n_4_net__944_,n_4_net__943_,n_4_net__942_,n_4_net__941_,n_4_net__940_,
  n_4_net__939_,n_4_net__938_,n_4_net__937_,n_4_net__936_,n_4_net__935_,n_4_net__934_,
  n_4_net__933_,n_4_net__932_,n_4_net__931_,n_4_net__930_,n_4_net__929_,
  n_4_net__928_,n_4_net__927_,n_4_net__926_,n_4_net__925_,n_4_net__924_,n_4_net__923_,
  n_4_net__922_,n_4_net__921_,n_4_net__920_,n_4_net__919_,n_4_net__918_,n_4_net__917_,
  n_4_net__916_,n_4_net__915_,n_4_net__914_,n_4_net__913_,n_4_net__912_,n_4_net__911_,
  n_4_net__910_,n_4_net__909_,n_4_net__908_,n_4_net__907_,n_4_net__906_,
  n_4_net__905_,n_4_net__904_,n_4_net__903_,n_4_net__902_,n_4_net__901_,n_4_net__900_,
  n_4_net__899_,n_4_net__898_,n_4_net__897_,n_4_net__896_,n_4_net__895_,n_4_net__894_,
  n_4_net__893_,n_4_net__892_,n_4_net__891_,n_4_net__890_,n_4_net__889_,
  n_4_net__888_,n_4_net__887_,n_4_net__886_,n_4_net__885_,n_4_net__884_,n_4_net__883_,
  n_4_net__882_,n_4_net__881_,n_4_net__880_,n_4_net__879_,n_4_net__878_,n_4_net__877_,
  n_4_net__876_,n_4_net__875_,n_4_net__874_,n_4_net__873_,n_4_net__872_,n_4_net__871_,
  n_4_net__870_,n_4_net__869_,n_4_net__868_,n_4_net__867_,n_4_net__866_,
  n_4_net__865_,n_4_net__864_,n_4_net__863_,n_4_net__862_,n_4_net__861_,n_4_net__860_,
  n_4_net__859_,n_4_net__858_,n_4_net__857_,n_4_net__856_,n_4_net__855_,n_4_net__854_,
  n_4_net__853_,n_4_net__852_,n_4_net__851_,n_4_net__850_,n_4_net__849_,
  n_4_net__848_,n_4_net__847_,n_4_net__846_,n_4_net__845_,n_4_net__844_,n_4_net__843_,
  n_4_net__842_,n_4_net__841_,n_4_net__840_,n_4_net__839_,n_4_net__838_,n_4_net__837_,
  n_4_net__836_,n_4_net__835_,n_4_net__834_,n_4_net__833_,n_4_net__832_,n_4_net__831_,
  n_4_net__830_,n_4_net__829_,n_4_net__828_,n_4_net__827_,n_4_net__826_,
  n_4_net__825_,n_4_net__824_,n_4_net__823_,n_4_net__822_,n_4_net__821_,n_4_net__820_,
  n_4_net__819_,n_4_net__818_,n_4_net__817_,n_4_net__816_,n_4_net__815_,n_4_net__814_,
  n_4_net__813_,n_4_net__812_,n_4_net__811_,n_4_net__810_,n_4_net__809_,
  n_4_net__808_,n_4_net__807_,n_4_net__806_,n_4_net__805_,n_4_net__804_,n_4_net__803_,
  n_4_net__802_,n_4_net__801_,n_4_net__800_,n_4_net__799_,n_4_net__798_,n_4_net__797_,
  n_4_net__796_,n_4_net__795_,n_4_net__794_,n_4_net__793_,n_4_net__792_,n_4_net__791_,
  n_4_net__790_,n_4_net__789_,n_4_net__788_,n_4_net__787_,n_4_net__786_,
  n_4_net__785_,n_4_net__784_,n_4_net__783_,n_4_net__782_,n_4_net__781_,n_4_net__780_,
  n_4_net__779_,n_4_net__778_,n_4_net__777_,n_4_net__776_,n_4_net__775_,n_4_net__774_,
  n_4_net__773_,n_4_net__772_,n_4_net__771_,n_4_net__770_,n_4_net__769_,
  n_4_net__768_,n_4_net__767_,n_4_net__766_,n_4_net__765_,n_4_net__764_,n_4_net__763_,
  n_4_net__762_,n_4_net__761_,n_4_net__760_,n_4_net__759_,n_4_net__758_,n_4_net__757_,
  n_4_net__756_,n_4_net__755_,n_4_net__754_,n_4_net__753_,n_4_net__752_,n_4_net__751_,
  n_4_net__750_,n_4_net__749_,n_4_net__748_,n_4_net__747_,n_4_net__746_,
  n_4_net__745_,n_4_net__744_,n_4_net__743_,n_4_net__742_,n_4_net__741_,n_4_net__740_,
  n_4_net__739_,n_4_net__738_,n_4_net__737_,n_4_net__736_,n_4_net__735_,n_4_net__734_,
  n_4_net__733_,n_4_net__732_,n_4_net__731_,n_4_net__730_,n_4_net__729_,
  n_4_net__728_,n_4_net__727_,n_4_net__726_,n_4_net__725_,n_4_net__724_,n_4_net__723_,
  n_4_net__722_,n_4_net__721_,n_4_net__720_,n_4_net__719_,n_4_net__718_,n_4_net__717_,
  n_4_net__716_,n_4_net__715_,n_4_net__714_,n_4_net__713_,n_4_net__712_,n_4_net__711_,
  n_4_net__710_,n_4_net__709_,n_4_net__708_,n_4_net__707_,n_4_net__706_,
  n_4_net__705_,n_4_net__704_,n_4_net__703_,n_4_net__702_,n_4_net__701_,n_4_net__700_,
  n_4_net__699_,n_4_net__698_,n_4_net__697_,n_4_net__696_,n_4_net__695_,n_4_net__694_,
  n_4_net__693_,n_4_net__692_,n_4_net__691_,n_4_net__690_,n_4_net__689_,
  n_4_net__688_,n_4_net__687_,n_4_net__686_,n_4_net__685_,n_4_net__684_,n_4_net__683_,
  n_4_net__682_,n_4_net__681_,n_4_net__680_,n_4_net__679_,n_4_net__678_,n_4_net__677_,
  n_4_net__676_,n_4_net__675_,n_4_net__674_,n_4_net__673_,n_4_net__672_,n_4_net__671_,
  n_4_net__670_,n_4_net__669_,n_4_net__668_,n_4_net__667_,n_4_net__666_,
  n_4_net__665_,n_4_net__664_,n_4_net__663_,n_4_net__662_,n_4_net__661_,n_4_net__660_,
  n_4_net__659_,n_4_net__658_,n_4_net__657_,n_4_net__656_,n_4_net__655_,n_4_net__654_,
  n_4_net__653_,n_4_net__652_,n_4_net__651_,n_4_net__650_,n_4_net__649_,
  n_4_net__648_,n_4_net__647_,n_4_net__646_,n_4_net__645_,n_4_net__644_,n_4_net__643_,
  n_4_net__642_,n_4_net__641_,n_4_net__640_,n_4_net__639_,n_4_net__638_,n_4_net__637_,
  n_4_net__636_,n_4_net__635_,n_4_net__634_,n_4_net__633_,n_4_net__632_,n_4_net__631_,
  n_4_net__630_,n_4_net__629_,n_4_net__628_,n_4_net__627_,n_4_net__626_,
  n_4_net__625_,n_4_net__624_,n_4_net__623_,n_4_net__622_,n_4_net__621_,n_4_net__620_,
  n_4_net__619_,n_4_net__618_,n_4_net__617_,n_4_net__616_,n_4_net__615_,n_4_net__614_,
  n_4_net__613_,n_4_net__612_,n_4_net__611_,n_4_net__610_,n_4_net__609_,
  n_4_net__608_,n_4_net__607_,n_4_net__606_,n_4_net__605_,n_4_net__604_,n_4_net__603_,
  n_4_net__602_,n_4_net__601_,n_4_net__600_,n_4_net__599_,n_4_net__598_,n_4_net__597_,
  n_4_net__596_,n_4_net__595_,n_4_net__594_,n_4_net__593_,n_4_net__592_,n_4_net__591_,
  n_4_net__590_,n_4_net__589_,n_4_net__588_,n_4_net__587_,n_4_net__586_,
  n_4_net__585_,n_4_net__584_,n_4_net__583_,n_4_net__582_,n_4_net__581_,n_4_net__580_,
  n_4_net__579_,n_4_net__578_,n_4_net__577_,n_4_net__576_,n_4_net__575_,n_4_net__574_,
  n_4_net__573_,n_4_net__572_,n_4_net__571_,n_4_net__570_,n_4_net__569_,
  n_4_net__568_,n_4_net__567_,n_4_net__566_,n_4_net__565_,n_4_net__564_,n_4_net__563_,
  n_4_net__562_,n_4_net__561_,n_4_net__560_,n_4_net__559_,n_4_net__558_,n_4_net__557_,
  n_4_net__556_,n_4_net__555_,n_4_net__554_,n_4_net__553_,n_4_net__552_,n_4_net__551_,
  n_4_net__550_,n_4_net__549_,n_4_net__548_,n_4_net__547_,n_4_net__546_,
  n_4_net__545_,n_4_net__544_,n_4_net__543_,n_4_net__542_,n_4_net__541_,n_4_net__540_,
  n_4_net__539_,n_4_net__538_,n_4_net__537_,n_4_net__536_,n_4_net__535_,n_4_net__534_,
  n_4_net__533_,n_4_net__532_,n_4_net__531_,n_4_net__530_,n_4_net__529_,
  n_4_net__528_,n_4_net__527_,n_4_net__526_,n_4_net__525_,n_4_net__524_,n_4_net__523_,
  n_4_net__522_,n_4_net__521_,n_4_net__520_,n_4_net__519_,n_4_net__518_,n_4_net__517_,
  n_4_net__516_,n_4_net__515_,n_4_net__514_,n_4_net__513_,n_4_net__512_,n_4_net__511_,
  n_4_net__510_,n_4_net__509_,n_4_net__508_,n_4_net__507_,n_4_net__506_,
  n_4_net__505_,n_4_net__504_,n_4_net__503_,n_4_net__502_,n_4_net__501_,n_4_net__500_,
  n_4_net__499_,n_4_net__498_,n_4_net__497_,n_4_net__496_,n_4_net__495_,n_4_net__494_,
  n_4_net__493_,n_4_net__492_,n_4_net__491_,n_4_net__490_,n_4_net__489_,
  n_4_net__488_,n_4_net__487_,n_4_net__486_,n_4_net__485_,n_4_net__484_,n_4_net__483_,
  n_4_net__482_,n_4_net__481_,n_4_net__480_,n_4_net__479_,n_4_net__478_,n_4_net__477_,
  n_4_net__476_,n_4_net__475_,n_4_net__474_,n_4_net__473_,n_4_net__472_,n_4_net__471_,
  n_4_net__470_,n_4_net__469_,n_4_net__468_,n_4_net__467_,n_4_net__466_,
  n_4_net__465_,n_4_net__464_,n_4_net__463_,n_4_net__462_,n_4_net__461_,n_4_net__460_,
  n_4_net__459_,n_4_net__458_,n_4_net__457_,n_4_net__456_,n_4_net__455_,n_4_net__454_,
  n_4_net__453_,n_4_net__452_,n_4_net__451_,n_4_net__450_,n_4_net__449_,
  n_4_net__448_,n_4_net__447_,n_4_net__446_,n_4_net__445_,n_4_net__444_,n_4_net__443_,
  n_4_net__442_,n_4_net__441_,n_4_net__440_,n_4_net__439_,n_4_net__438_,n_4_net__437_,
  n_4_net__436_,n_4_net__435_,n_4_net__434_,n_4_net__433_,n_4_net__432_,n_4_net__431_,
  n_4_net__430_,n_4_net__429_,n_4_net__428_,n_4_net__427_,n_4_net__426_,
  n_4_net__425_,n_4_net__424_,n_4_net__423_,n_4_net__422_,n_4_net__421_,n_4_net__420_,
  n_4_net__419_,n_4_net__418_,n_4_net__417_,n_4_net__416_,n_4_net__415_,n_4_net__414_,
  n_4_net__413_,n_4_net__412_,n_4_net__411_,n_4_net__410_,n_4_net__409_,
  n_4_net__408_,n_4_net__407_,n_4_net__406_,n_4_net__405_,n_4_net__404_,n_4_net__403_,
  n_4_net__402_,n_4_net__401_,n_4_net__400_,n_4_net__399_,n_4_net__398_,n_4_net__397_,
  n_4_net__396_,n_4_net__395_,n_4_net__394_,n_4_net__393_,n_4_net__392_,n_4_net__391_,
  n_4_net__390_,n_4_net__389_,n_4_net__388_,n_4_net__387_,n_4_net__386_,
  n_4_net__385_,n_4_net__384_,n_4_net__383_,n_4_net__382_,n_4_net__381_,n_4_net__380_,
  n_4_net__379_,n_4_net__378_,n_4_net__377_,n_4_net__376_,n_4_net__375_,n_4_net__374_,
  n_4_net__373_,n_4_net__372_,n_4_net__371_,n_4_net__370_,n_4_net__369_,
  n_4_net__368_,n_4_net__367_,n_4_net__366_,n_4_net__365_,n_4_net__364_,n_4_net__363_,
  n_4_net__362_,n_4_net__361_,n_4_net__360_,n_4_net__359_,n_4_net__358_,n_4_net__357_,
  n_4_net__356_,n_4_net__355_,n_4_net__354_,n_4_net__353_,n_4_net__352_,n_4_net__351_,
  n_4_net__350_,n_4_net__349_,n_4_net__348_,n_4_net__347_,n_4_net__346_,
  n_4_net__345_,n_4_net__344_,n_4_net__343_,n_4_net__342_,n_4_net__341_,n_4_net__340_,
  n_4_net__339_,n_4_net__338_,n_4_net__337_,n_4_net__336_,n_4_net__335_,n_4_net__334_,
  n_4_net__333_,n_4_net__332_,n_4_net__331_,n_4_net__330_,n_4_net__329_,
  n_4_net__328_,n_4_net__327_,n_4_net__326_,n_4_net__325_,n_4_net__324_,n_4_net__323_,
  n_4_net__322_,n_4_net__321_,n_4_net__320_,n_4_net__319_,n_4_net__318_,n_4_net__317_,
  n_4_net__316_,n_4_net__315_,n_4_net__314_,n_4_net__313_,n_4_net__312_,n_4_net__311_,
  n_4_net__310_,n_4_net__309_,n_4_net__308_,n_4_net__307_,n_4_net__306_,
  n_4_net__305_,n_4_net__304_,n_4_net__303_,n_4_net__302_,n_4_net__301_,n_4_net__300_,
  n_4_net__299_,n_4_net__298_,n_4_net__297_,n_4_net__296_,n_4_net__295_,n_4_net__294_,
  n_4_net__293_,n_4_net__292_,n_4_net__291_,n_4_net__290_,n_4_net__289_,
  n_4_net__288_,n_4_net__287_,n_4_net__286_,n_4_net__285_,n_4_net__284_,n_4_net__283_,
  n_4_net__282_,n_4_net__281_,n_4_net__280_,n_4_net__279_,n_4_net__278_,n_4_net__277_,
  n_4_net__276_,n_4_net__275_,n_4_net__274_,n_4_net__273_,n_4_net__272_,n_4_net__271_,
  n_4_net__270_,n_4_net__269_,n_4_net__268_,n_4_net__267_,n_4_net__266_,
  n_4_net__265_,n_4_net__264_,n_4_net__263_,n_4_net__262_,n_4_net__261_,n_4_net__260_,
  n_4_net__259_,n_4_net__258_,n_4_net__257_,n_4_net__256_,n_4_net__255_,n_4_net__254_,
  n_4_net__253_,n_4_net__252_,n_4_net__251_,n_4_net__250_,n_4_net__249_,
  n_4_net__248_,n_4_net__247_,n_4_net__246_,n_4_net__245_,n_4_net__244_,n_4_net__243_,
  n_4_net__242_,n_4_net__241_,n_4_net__240_,n_4_net__239_,n_4_net__238_,n_4_net__237_,
  n_4_net__236_,n_4_net__235_,n_4_net__234_,n_4_net__233_,n_4_net__232_,n_4_net__231_,
  n_4_net__230_,n_4_net__229_,n_4_net__228_,n_4_net__227_,n_4_net__226_,
  n_4_net__225_,n_4_net__224_,n_4_net__223_,n_4_net__222_,n_4_net__221_,n_4_net__220_,
  n_4_net__219_,n_4_net__218_,n_4_net__217_,n_4_net__216_,n_4_net__215_,n_4_net__214_,
  n_4_net__213_,n_4_net__212_,n_4_net__211_,n_4_net__210_,n_4_net__209_,
  n_4_net__208_,n_4_net__207_,n_4_net__206_,n_4_net__205_,n_4_net__204_,n_4_net__203_,
  n_4_net__202_,n_4_net__201_,n_4_net__200_,n_4_net__199_,n_4_net__198_,n_4_net__197_,
  n_4_net__196_,n_4_net__195_,n_4_net__194_,n_4_net__193_,n_4_net__192_,n_4_net__191_,
  n_4_net__190_,n_4_net__189_,n_4_net__188_,n_4_net__187_,n_4_net__186_,
  n_4_net__185_,n_4_net__184_,n_4_net__183_,n_4_net__182_,n_4_net__181_,n_4_net__180_,
  n_4_net__179_,n_4_net__178_,n_4_net__177_,n_4_net__176_,n_4_net__175_,n_4_net__174_,
  n_4_net__173_,n_4_net__172_,n_4_net__171_,n_4_net__170_,n_4_net__169_,
  n_4_net__168_,n_4_net__167_,n_4_net__166_,n_4_net__165_,n_4_net__164_,n_4_net__163_,
  n_4_net__162_,n_4_net__161_,n_4_net__160_,n_4_net__159_,n_4_net__158_,n_4_net__157_,
  n_4_net__156_,n_4_net__155_,n_4_net__154_,n_4_net__153_,n_4_net__152_,n_4_net__151_,
  n_4_net__150_,n_4_net__149_,n_4_net__148_,n_4_net__147_,n_4_net__146_,
  n_4_net__145_,n_4_net__144_,n_4_net__143_,n_4_net__142_,n_4_net__141_,n_4_net__140_,
  n_4_net__139_,n_4_net__138_,n_4_net__137_,n_4_net__136_,n_4_net__135_,n_4_net__134_,
  n_4_net__133_,n_4_net__132_,n_4_net__131_,n_4_net__130_,n_4_net__129_,
  n_4_net__128_,n_4_net__127_,n_4_net__126_,n_4_net__125_,n_4_net__124_,n_4_net__123_,
  n_4_net__122_,n_4_net__121_,n_4_net__120_,n_4_net__119_,n_4_net__118_,n_4_net__117_,
  n_4_net__116_,n_4_net__115_,n_4_net__114_,n_4_net__113_,n_4_net__112_,n_4_net__111_,
  n_4_net__110_,n_4_net__109_,n_4_net__108_,n_4_net__107_,n_4_net__106_,
  n_4_net__105_,n_4_net__104_,n_4_net__103_,n_4_net__102_,n_4_net__101_,n_4_net__100_,
  n_4_net__99_,n_4_net__98_,n_4_net__97_,n_4_net__96_,n_4_net__95_,n_4_net__94_,
  n_4_net__93_,n_4_net__92_,n_4_net__91_,n_4_net__90_,n_4_net__89_,n_4_net__88_,
  n_4_net__87_,n_4_net__86_,n_4_net__85_,n_4_net__84_,n_4_net__83_,n_4_net__82_,
  n_4_net__81_,n_4_net__80_,n_4_net__79_,n_4_net__78_,n_4_net__77_,n_4_net__76_,n_4_net__75_,
  n_4_net__74_,n_4_net__73_,n_4_net__72_,n_4_net__71_,n_4_net__70_,n_4_net__69_,
  n_4_net__68_,n_4_net__67_,n_4_net__66_,n_4_net__65_,n_4_net__64_,n_4_net__63_,
  n_4_net__62_,n_4_net__61_,n_4_net__60_,n_4_net__59_,n_4_net__58_,n_4_net__57_,
  n_4_net__56_,n_4_net__55_,n_4_net__54_,n_4_net__53_,n_4_net__52_,n_4_net__51_,
  n_4_net__50_,n_4_net__49_,n_4_net__48_,n_4_net__47_,n_4_net__46_,n_4_net__45_,
  n_4_net__44_,n_4_net__43_,n_4_net__42_,n_4_net__41_,n_4_net__40_,n_4_net__39_,n_4_net__38_,
  n_4_net__37_,n_4_net__36_,n_4_net__35_,n_4_net__34_,n_4_net__33_,n_4_net__32_,
  n_4_net__31_,n_4_net__30_,n_4_net__29_,n_4_net__28_,n_4_net__27_,n_4_net__26_,
  n_4_net__25_,n_4_net__24_,n_4_net__23_,n_4_net__22_,n_4_net__21_,n_4_net__20_,
  n_4_net__19_,n_4_net__18_,n_4_net__17_,n_4_net__16_,n_4_net__15_,n_4_net__14_,
  n_4_net__13_,n_4_net__12_,n_4_net__11_,n_4_net__10_,n_4_net__9_,n_4_net__8_,n_4_net__7_,
  n_4_net__6_,n_4_net__5_,n_4_net__4_,n_4_net__3_,n_4_net__2_,n_4_net__1_,
  n_4_net__0_,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,n_5_net_,N175,N176,N177,
  N178,N179,N180,N181,N182,N183,N184;
  wire [3:0] go_cnt;

  bsg_make_2D_array_width_p128_items_p10
  bm2Da
  (
    .i(data_o_flat),
    .o(data_o)
  );


  bsg_rr_f2f_input_width_p128_num_in_p10_middle_meet_p10
  ic_9__in_chan_bsg_rr_ff_in
  (
    .clk(clk),
    .reset(n_0_net_),
    .valid_i(valid_i),
    .data_i(data_i),
    .data_head_o({ data_head_9__1279_, data_head_9__1278_, data_head_9__1277_, data_head_9__1276_, data_head_9__1275_, data_head_9__1274_, data_head_9__1273_, data_head_9__1272_, data_head_9__1271_, data_head_9__1270_, data_head_9__1269_, data_head_9__1268_, data_head_9__1267_, data_head_9__1266_, data_head_9__1265_, data_head_9__1264_, data_head_9__1263_, data_head_9__1262_, data_head_9__1261_, data_head_9__1260_, data_head_9__1259_, data_head_9__1258_, data_head_9__1257_, data_head_9__1256_, data_head_9__1255_, data_head_9__1254_, data_head_9__1253_, data_head_9__1252_, data_head_9__1251_, data_head_9__1250_, data_head_9__1249_, data_head_9__1248_, data_head_9__1247_, data_head_9__1246_, data_head_9__1245_, data_head_9__1244_, data_head_9__1243_, data_head_9__1242_, data_head_9__1241_, data_head_9__1240_, data_head_9__1239_, data_head_9__1238_, data_head_9__1237_, data_head_9__1236_, data_head_9__1235_, data_head_9__1234_, data_head_9__1233_, data_head_9__1232_, data_head_9__1231_, data_head_9__1230_, data_head_9__1229_, data_head_9__1228_, data_head_9__1227_, data_head_9__1226_, data_head_9__1225_, data_head_9__1224_, data_head_9__1223_, data_head_9__1222_, data_head_9__1221_, data_head_9__1220_, data_head_9__1219_, data_head_9__1218_, data_head_9__1217_, data_head_9__1216_, data_head_9__1215_, data_head_9__1214_, data_head_9__1213_, data_head_9__1212_, data_head_9__1211_, data_head_9__1210_, data_head_9__1209_, data_head_9__1208_, data_head_9__1207_, data_head_9__1206_, data_head_9__1205_, data_head_9__1204_, data_head_9__1203_, data_head_9__1202_, data_head_9__1201_, data_head_9__1200_, data_head_9__1199_, data_head_9__1198_, data_head_9__1197_, data_head_9__1196_, data_head_9__1195_, data_head_9__1194_, data_head_9__1193_, data_head_9__1192_, data_head_9__1191_, data_head_9__1190_, data_head_9__1189_, data_head_9__1188_, data_head_9__1187_, data_head_9__1186_, data_head_9__1185_, data_head_9__1184_, data_head_9__1183_, data_head_9__1182_, data_head_9__1181_, data_head_9__1180_, data_head_9__1179_, data_head_9__1178_, data_head_9__1177_, data_head_9__1176_, data_head_9__1175_, data_head_9__1174_, data_head_9__1173_, data_head_9__1172_, data_head_9__1171_, data_head_9__1170_, data_head_9__1169_, data_head_9__1168_, data_head_9__1167_, data_head_9__1166_, data_head_9__1165_, data_head_9__1164_, data_head_9__1163_, data_head_9__1162_, data_head_9__1161_, data_head_9__1160_, data_head_9__1159_, data_head_9__1158_, data_head_9__1157_, data_head_9__1156_, data_head_9__1155_, data_head_9__1154_, data_head_9__1153_, data_head_9__1152_, data_head_9__1151_, data_head_9__1150_, data_head_9__1149_, data_head_9__1148_, data_head_9__1147_, data_head_9__1146_, data_head_9__1145_, data_head_9__1144_, data_head_9__1143_, data_head_9__1142_, data_head_9__1141_, data_head_9__1140_, data_head_9__1139_, data_head_9__1138_, data_head_9__1137_, data_head_9__1136_, data_head_9__1135_, data_head_9__1134_, data_head_9__1133_, data_head_9__1132_, data_head_9__1131_, data_head_9__1130_, data_head_9__1129_, data_head_9__1128_, data_head_9__1127_, data_head_9__1126_, data_head_9__1125_, data_head_9__1124_, data_head_9__1123_, data_head_9__1122_, data_head_9__1121_, data_head_9__1120_, data_head_9__1119_, data_head_9__1118_, data_head_9__1117_, data_head_9__1116_, data_head_9__1115_, data_head_9__1114_, data_head_9__1113_, data_head_9__1112_, data_head_9__1111_, data_head_9__1110_, data_head_9__1109_, data_head_9__1108_, data_head_9__1107_, data_head_9__1106_, data_head_9__1105_, data_head_9__1104_, data_head_9__1103_, data_head_9__1102_, data_head_9__1101_, data_head_9__1100_, data_head_9__1099_, data_head_9__1098_, data_head_9__1097_, data_head_9__1096_, data_head_9__1095_, data_head_9__1094_, data_head_9__1093_, data_head_9__1092_, data_head_9__1091_, data_head_9__1090_, data_head_9__1089_, data_head_9__1088_, data_head_9__1087_, data_head_9__1086_, data_head_9__1085_, data_head_9__1084_, data_head_9__1083_, data_head_9__1082_, data_head_9__1081_, data_head_9__1080_, data_head_9__1079_, data_head_9__1078_, data_head_9__1077_, data_head_9__1076_, data_head_9__1075_, data_head_9__1074_, data_head_9__1073_, data_head_9__1072_, data_head_9__1071_, data_head_9__1070_, data_head_9__1069_, data_head_9__1068_, data_head_9__1067_, data_head_9__1066_, data_head_9__1065_, data_head_9__1064_, data_head_9__1063_, data_head_9__1062_, data_head_9__1061_, data_head_9__1060_, data_head_9__1059_, data_head_9__1058_, data_head_9__1057_, data_head_9__1056_, data_head_9__1055_, data_head_9__1054_, data_head_9__1053_, data_head_9__1052_, data_head_9__1051_, data_head_9__1050_, data_head_9__1049_, data_head_9__1048_, data_head_9__1047_, data_head_9__1046_, data_head_9__1045_, data_head_9__1044_, data_head_9__1043_, data_head_9__1042_, data_head_9__1041_, data_head_9__1040_, data_head_9__1039_, data_head_9__1038_, data_head_9__1037_, data_head_9__1036_, data_head_9__1035_, data_head_9__1034_, data_head_9__1033_, data_head_9__1032_, data_head_9__1031_, data_head_9__1030_, data_head_9__1029_, data_head_9__1028_, data_head_9__1027_, data_head_9__1026_, data_head_9__1025_, data_head_9__1024_, data_head_9__1023_, data_head_9__1022_, data_head_9__1021_, data_head_9__1020_, data_head_9__1019_, data_head_9__1018_, data_head_9__1017_, data_head_9__1016_, data_head_9__1015_, data_head_9__1014_, data_head_9__1013_, data_head_9__1012_, data_head_9__1011_, data_head_9__1010_, data_head_9__1009_, data_head_9__1008_, data_head_9__1007_, data_head_9__1006_, data_head_9__1005_, data_head_9__1004_, data_head_9__1003_, data_head_9__1002_, data_head_9__1001_, data_head_9__1000_, data_head_9__999_, data_head_9__998_, data_head_9__997_, data_head_9__996_, data_head_9__995_, data_head_9__994_, data_head_9__993_, data_head_9__992_, data_head_9__991_, data_head_9__990_, data_head_9__989_, data_head_9__988_, data_head_9__987_, data_head_9__986_, data_head_9__985_, data_head_9__984_, data_head_9__983_, data_head_9__982_, data_head_9__981_, data_head_9__980_, data_head_9__979_, data_head_9__978_, data_head_9__977_, data_head_9__976_, data_head_9__975_, data_head_9__974_, data_head_9__973_, data_head_9__972_, data_head_9__971_, data_head_9__970_, data_head_9__969_, data_head_9__968_, data_head_9__967_, data_head_9__966_, data_head_9__965_, data_head_9__964_, data_head_9__963_, data_head_9__962_, data_head_9__961_, data_head_9__960_, data_head_9__959_, data_head_9__958_, data_head_9__957_, data_head_9__956_, data_head_9__955_, data_head_9__954_, data_head_9__953_, data_head_9__952_, data_head_9__951_, data_head_9__950_, data_head_9__949_, data_head_9__948_, data_head_9__947_, data_head_9__946_, data_head_9__945_, data_head_9__944_, data_head_9__943_, data_head_9__942_, data_head_9__941_, data_head_9__940_, data_head_9__939_, data_head_9__938_, data_head_9__937_, data_head_9__936_, data_head_9__935_, data_head_9__934_, data_head_9__933_, data_head_9__932_, data_head_9__931_, data_head_9__930_, data_head_9__929_, data_head_9__928_, data_head_9__927_, data_head_9__926_, data_head_9__925_, data_head_9__924_, data_head_9__923_, data_head_9__922_, data_head_9__921_, data_head_9__920_, data_head_9__919_, data_head_9__918_, data_head_9__917_, data_head_9__916_, data_head_9__915_, data_head_9__914_, data_head_9__913_, data_head_9__912_, data_head_9__911_, data_head_9__910_, data_head_9__909_, data_head_9__908_, data_head_9__907_, data_head_9__906_, data_head_9__905_, data_head_9__904_, data_head_9__903_, data_head_9__902_, data_head_9__901_, data_head_9__900_, data_head_9__899_, data_head_9__898_, data_head_9__897_, data_head_9__896_, data_head_9__895_, data_head_9__894_, data_head_9__893_, data_head_9__892_, data_head_9__891_, data_head_9__890_, data_head_9__889_, data_head_9__888_, data_head_9__887_, data_head_9__886_, data_head_9__885_, data_head_9__884_, data_head_9__883_, data_head_9__882_, data_head_9__881_, data_head_9__880_, data_head_9__879_, data_head_9__878_, data_head_9__877_, data_head_9__876_, data_head_9__875_, data_head_9__874_, data_head_9__873_, data_head_9__872_, data_head_9__871_, data_head_9__870_, data_head_9__869_, data_head_9__868_, data_head_9__867_, data_head_9__866_, data_head_9__865_, data_head_9__864_, data_head_9__863_, data_head_9__862_, data_head_9__861_, data_head_9__860_, data_head_9__859_, data_head_9__858_, data_head_9__857_, data_head_9__856_, data_head_9__855_, data_head_9__854_, data_head_9__853_, data_head_9__852_, data_head_9__851_, data_head_9__850_, data_head_9__849_, data_head_9__848_, data_head_9__847_, data_head_9__846_, data_head_9__845_, data_head_9__844_, data_head_9__843_, data_head_9__842_, data_head_9__841_, data_head_9__840_, data_head_9__839_, data_head_9__838_, data_head_9__837_, data_head_9__836_, data_head_9__835_, data_head_9__834_, data_head_9__833_, data_head_9__832_, data_head_9__831_, data_head_9__830_, data_head_9__829_, data_head_9__828_, data_head_9__827_, data_head_9__826_, data_head_9__825_, data_head_9__824_, data_head_9__823_, data_head_9__822_, data_head_9__821_, data_head_9__820_, data_head_9__819_, data_head_9__818_, data_head_9__817_, data_head_9__816_, data_head_9__815_, data_head_9__814_, data_head_9__813_, data_head_9__812_, data_head_9__811_, data_head_9__810_, data_head_9__809_, data_head_9__808_, data_head_9__807_, data_head_9__806_, data_head_9__805_, data_head_9__804_, data_head_9__803_, data_head_9__802_, data_head_9__801_, data_head_9__800_, data_head_9__799_, data_head_9__798_, data_head_9__797_, data_head_9__796_, data_head_9__795_, data_head_9__794_, data_head_9__793_, data_head_9__792_, data_head_9__791_, data_head_9__790_, data_head_9__789_, data_head_9__788_, data_head_9__787_, data_head_9__786_, data_head_9__785_, data_head_9__784_, data_head_9__783_, data_head_9__782_, data_head_9__781_, data_head_9__780_, data_head_9__779_, data_head_9__778_, data_head_9__777_, data_head_9__776_, data_head_9__775_, data_head_9__774_, data_head_9__773_, data_head_9__772_, data_head_9__771_, data_head_9__770_, data_head_9__769_, data_head_9__768_, data_head_9__767_, data_head_9__766_, data_head_9__765_, data_head_9__764_, data_head_9__763_, data_head_9__762_, data_head_9__761_, data_head_9__760_, data_head_9__759_, data_head_9__758_, data_head_9__757_, data_head_9__756_, data_head_9__755_, data_head_9__754_, data_head_9__753_, data_head_9__752_, data_head_9__751_, data_head_9__750_, data_head_9__749_, data_head_9__748_, data_head_9__747_, data_head_9__746_, data_head_9__745_, data_head_9__744_, data_head_9__743_, data_head_9__742_, data_head_9__741_, data_head_9__740_, data_head_9__739_, data_head_9__738_, data_head_9__737_, data_head_9__736_, data_head_9__735_, data_head_9__734_, data_head_9__733_, data_head_9__732_, data_head_9__731_, data_head_9__730_, data_head_9__729_, data_head_9__728_, data_head_9__727_, data_head_9__726_, data_head_9__725_, data_head_9__724_, data_head_9__723_, data_head_9__722_, data_head_9__721_, data_head_9__720_, data_head_9__719_, data_head_9__718_, data_head_9__717_, data_head_9__716_, data_head_9__715_, data_head_9__714_, data_head_9__713_, data_head_9__712_, data_head_9__711_, data_head_9__710_, data_head_9__709_, data_head_9__708_, data_head_9__707_, data_head_9__706_, data_head_9__705_, data_head_9__704_, data_head_9__703_, data_head_9__702_, data_head_9__701_, data_head_9__700_, data_head_9__699_, data_head_9__698_, data_head_9__697_, data_head_9__696_, data_head_9__695_, data_head_9__694_, data_head_9__693_, data_head_9__692_, data_head_9__691_, data_head_9__690_, data_head_9__689_, data_head_9__688_, data_head_9__687_, data_head_9__686_, data_head_9__685_, data_head_9__684_, data_head_9__683_, data_head_9__682_, data_head_9__681_, data_head_9__680_, data_head_9__679_, data_head_9__678_, data_head_9__677_, data_head_9__676_, data_head_9__675_, data_head_9__674_, data_head_9__673_, data_head_9__672_, data_head_9__671_, data_head_9__670_, data_head_9__669_, data_head_9__668_, data_head_9__667_, data_head_9__666_, data_head_9__665_, data_head_9__664_, data_head_9__663_, data_head_9__662_, data_head_9__661_, data_head_9__660_, data_head_9__659_, data_head_9__658_, data_head_9__657_, data_head_9__656_, data_head_9__655_, data_head_9__654_, data_head_9__653_, data_head_9__652_, data_head_9__651_, data_head_9__650_, data_head_9__649_, data_head_9__648_, data_head_9__647_, data_head_9__646_, data_head_9__645_, data_head_9__644_, data_head_9__643_, data_head_9__642_, data_head_9__641_, data_head_9__640_, data_head_9__639_, data_head_9__638_, data_head_9__637_, data_head_9__636_, data_head_9__635_, data_head_9__634_, data_head_9__633_, data_head_9__632_, data_head_9__631_, data_head_9__630_, data_head_9__629_, data_head_9__628_, data_head_9__627_, data_head_9__626_, data_head_9__625_, data_head_9__624_, data_head_9__623_, data_head_9__622_, data_head_9__621_, data_head_9__620_, data_head_9__619_, data_head_9__618_, data_head_9__617_, data_head_9__616_, data_head_9__615_, data_head_9__614_, data_head_9__613_, data_head_9__612_, data_head_9__611_, data_head_9__610_, data_head_9__609_, data_head_9__608_, data_head_9__607_, data_head_9__606_, data_head_9__605_, data_head_9__604_, data_head_9__603_, data_head_9__602_, data_head_9__601_, data_head_9__600_, data_head_9__599_, data_head_9__598_, data_head_9__597_, data_head_9__596_, data_head_9__595_, data_head_9__594_, data_head_9__593_, data_head_9__592_, data_head_9__591_, data_head_9__590_, data_head_9__589_, data_head_9__588_, data_head_9__587_, data_head_9__586_, data_head_9__585_, data_head_9__584_, data_head_9__583_, data_head_9__582_, data_head_9__581_, data_head_9__580_, data_head_9__579_, data_head_9__578_, data_head_9__577_, data_head_9__576_, data_head_9__575_, data_head_9__574_, data_head_9__573_, data_head_9__572_, data_head_9__571_, data_head_9__570_, data_head_9__569_, data_head_9__568_, data_head_9__567_, data_head_9__566_, data_head_9__565_, data_head_9__564_, data_head_9__563_, data_head_9__562_, data_head_9__561_, data_head_9__560_, data_head_9__559_, data_head_9__558_, data_head_9__557_, data_head_9__556_, data_head_9__555_, data_head_9__554_, data_head_9__553_, data_head_9__552_, data_head_9__551_, data_head_9__550_, data_head_9__549_, data_head_9__548_, data_head_9__547_, data_head_9__546_, data_head_9__545_, data_head_9__544_, data_head_9__543_, data_head_9__542_, data_head_9__541_, data_head_9__540_, data_head_9__539_, data_head_9__538_, data_head_9__537_, data_head_9__536_, data_head_9__535_, data_head_9__534_, data_head_9__533_, data_head_9__532_, data_head_9__531_, data_head_9__530_, data_head_9__529_, data_head_9__528_, data_head_9__527_, data_head_9__526_, data_head_9__525_, data_head_9__524_, data_head_9__523_, data_head_9__522_, data_head_9__521_, data_head_9__520_, data_head_9__519_, data_head_9__518_, data_head_9__517_, data_head_9__516_, data_head_9__515_, data_head_9__514_, data_head_9__513_, data_head_9__512_, data_head_9__511_, data_head_9__510_, data_head_9__509_, data_head_9__508_, data_head_9__507_, data_head_9__506_, data_head_9__505_, data_head_9__504_, data_head_9__503_, data_head_9__502_, data_head_9__501_, data_head_9__500_, data_head_9__499_, data_head_9__498_, data_head_9__497_, data_head_9__496_, data_head_9__495_, data_head_9__494_, data_head_9__493_, data_head_9__492_, data_head_9__491_, data_head_9__490_, data_head_9__489_, data_head_9__488_, data_head_9__487_, data_head_9__486_, data_head_9__485_, data_head_9__484_, data_head_9__483_, data_head_9__482_, data_head_9__481_, data_head_9__480_, data_head_9__479_, data_head_9__478_, data_head_9__477_, data_head_9__476_, data_head_9__475_, data_head_9__474_, data_head_9__473_, data_head_9__472_, data_head_9__471_, data_head_9__470_, data_head_9__469_, data_head_9__468_, data_head_9__467_, data_head_9__466_, data_head_9__465_, data_head_9__464_, data_head_9__463_, data_head_9__462_, data_head_9__461_, data_head_9__460_, data_head_9__459_, data_head_9__458_, data_head_9__457_, data_head_9__456_, data_head_9__455_, data_head_9__454_, data_head_9__453_, data_head_9__452_, data_head_9__451_, data_head_9__450_, data_head_9__449_, data_head_9__448_, data_head_9__447_, data_head_9__446_, data_head_9__445_, data_head_9__444_, data_head_9__443_, data_head_9__442_, data_head_9__441_, data_head_9__440_, data_head_9__439_, data_head_9__438_, data_head_9__437_, data_head_9__436_, data_head_9__435_, data_head_9__434_, data_head_9__433_, data_head_9__432_, data_head_9__431_, data_head_9__430_, data_head_9__429_, data_head_9__428_, data_head_9__427_, data_head_9__426_, data_head_9__425_, data_head_9__424_, data_head_9__423_, data_head_9__422_, data_head_9__421_, data_head_9__420_, data_head_9__419_, data_head_9__418_, data_head_9__417_, data_head_9__416_, data_head_9__415_, data_head_9__414_, data_head_9__413_, data_head_9__412_, data_head_9__411_, data_head_9__410_, data_head_9__409_, data_head_9__408_, data_head_9__407_, data_head_9__406_, data_head_9__405_, data_head_9__404_, data_head_9__403_, data_head_9__402_, data_head_9__401_, data_head_9__400_, data_head_9__399_, data_head_9__398_, data_head_9__397_, data_head_9__396_, data_head_9__395_, data_head_9__394_, data_head_9__393_, data_head_9__392_, data_head_9__391_, data_head_9__390_, data_head_9__389_, data_head_9__388_, data_head_9__387_, data_head_9__386_, data_head_9__385_, data_head_9__384_, data_head_9__383_, data_head_9__382_, data_head_9__381_, data_head_9__380_, data_head_9__379_, data_head_9__378_, data_head_9__377_, data_head_9__376_, data_head_9__375_, data_head_9__374_, data_head_9__373_, data_head_9__372_, data_head_9__371_, data_head_9__370_, data_head_9__369_, data_head_9__368_, data_head_9__367_, data_head_9__366_, data_head_9__365_, data_head_9__364_, data_head_9__363_, data_head_9__362_, data_head_9__361_, data_head_9__360_, data_head_9__359_, data_head_9__358_, data_head_9__357_, data_head_9__356_, data_head_9__355_, data_head_9__354_, data_head_9__353_, data_head_9__352_, data_head_9__351_, data_head_9__350_, data_head_9__349_, data_head_9__348_, data_head_9__347_, data_head_9__346_, data_head_9__345_, data_head_9__344_, data_head_9__343_, data_head_9__342_, data_head_9__341_, data_head_9__340_, data_head_9__339_, data_head_9__338_, data_head_9__337_, data_head_9__336_, data_head_9__335_, data_head_9__334_, data_head_9__333_, data_head_9__332_, data_head_9__331_, data_head_9__330_, data_head_9__329_, data_head_9__328_, data_head_9__327_, data_head_9__326_, data_head_9__325_, data_head_9__324_, data_head_9__323_, data_head_9__322_, data_head_9__321_, data_head_9__320_, data_head_9__319_, data_head_9__318_, data_head_9__317_, data_head_9__316_, data_head_9__315_, data_head_9__314_, data_head_9__313_, data_head_9__312_, data_head_9__311_, data_head_9__310_, data_head_9__309_, data_head_9__308_, data_head_9__307_, data_head_9__306_, data_head_9__305_, data_head_9__304_, data_head_9__303_, data_head_9__302_, data_head_9__301_, data_head_9__300_, data_head_9__299_, data_head_9__298_, data_head_9__297_, data_head_9__296_, data_head_9__295_, data_head_9__294_, data_head_9__293_, data_head_9__292_, data_head_9__291_, data_head_9__290_, data_head_9__289_, data_head_9__288_, data_head_9__287_, data_head_9__286_, data_head_9__285_, data_head_9__284_, data_head_9__283_, data_head_9__282_, data_head_9__281_, data_head_9__280_, data_head_9__279_, data_head_9__278_, data_head_9__277_, data_head_9__276_, data_head_9__275_, data_head_9__274_, data_head_9__273_, data_head_9__272_, data_head_9__271_, data_head_9__270_, data_head_9__269_, data_head_9__268_, data_head_9__267_, data_head_9__266_, data_head_9__265_, data_head_9__264_, data_head_9__263_, data_head_9__262_, data_head_9__261_, data_head_9__260_, data_head_9__259_, data_head_9__258_, data_head_9__257_, data_head_9__256_, data_head_9__255_, data_head_9__254_, data_head_9__253_, data_head_9__252_, data_head_9__251_, data_head_9__250_, data_head_9__249_, data_head_9__248_, data_head_9__247_, data_head_9__246_, data_head_9__245_, data_head_9__244_, data_head_9__243_, data_head_9__242_, data_head_9__241_, data_head_9__240_, data_head_9__239_, data_head_9__238_, data_head_9__237_, data_head_9__236_, data_head_9__235_, data_head_9__234_, data_head_9__233_, data_head_9__232_, data_head_9__231_, data_head_9__230_, data_head_9__229_, data_head_9__228_, data_head_9__227_, data_head_9__226_, data_head_9__225_, data_head_9__224_, data_head_9__223_, data_head_9__222_, data_head_9__221_, data_head_9__220_, data_head_9__219_, data_head_9__218_, data_head_9__217_, data_head_9__216_, data_head_9__215_, data_head_9__214_, data_head_9__213_, data_head_9__212_, data_head_9__211_, data_head_9__210_, data_head_9__209_, data_head_9__208_, data_head_9__207_, data_head_9__206_, data_head_9__205_, data_head_9__204_, data_head_9__203_, data_head_9__202_, data_head_9__201_, data_head_9__200_, data_head_9__199_, data_head_9__198_, data_head_9__197_, data_head_9__196_, data_head_9__195_, data_head_9__194_, data_head_9__193_, data_head_9__192_, data_head_9__191_, data_head_9__190_, data_head_9__189_, data_head_9__188_, data_head_9__187_, data_head_9__186_, data_head_9__185_, data_head_9__184_, data_head_9__183_, data_head_9__182_, data_head_9__181_, data_head_9__180_, data_head_9__179_, data_head_9__178_, data_head_9__177_, data_head_9__176_, data_head_9__175_, data_head_9__174_, data_head_9__173_, data_head_9__172_, data_head_9__171_, data_head_9__170_, data_head_9__169_, data_head_9__168_, data_head_9__167_, data_head_9__166_, data_head_9__165_, data_head_9__164_, data_head_9__163_, data_head_9__162_, data_head_9__161_, data_head_9__160_, data_head_9__159_, data_head_9__158_, data_head_9__157_, data_head_9__156_, data_head_9__155_, data_head_9__154_, data_head_9__153_, data_head_9__152_, data_head_9__151_, data_head_9__150_, data_head_9__149_, data_head_9__148_, data_head_9__147_, data_head_9__146_, data_head_9__145_, data_head_9__144_, data_head_9__143_, data_head_9__142_, data_head_9__141_, data_head_9__140_, data_head_9__139_, data_head_9__138_, data_head_9__137_, data_head_9__136_, data_head_9__135_, data_head_9__134_, data_head_9__133_, data_head_9__132_, data_head_9__131_, data_head_9__130_, data_head_9__129_, data_head_9__128_, data_head_9__127_, data_head_9__126_, data_head_9__125_, data_head_9__124_, data_head_9__123_, data_head_9__122_, data_head_9__121_, data_head_9__120_, data_head_9__119_, data_head_9__118_, data_head_9__117_, data_head_9__116_, data_head_9__115_, data_head_9__114_, data_head_9__113_, data_head_9__112_, data_head_9__111_, data_head_9__110_, data_head_9__109_, data_head_9__108_, data_head_9__107_, data_head_9__106_, data_head_9__105_, data_head_9__104_, data_head_9__103_, data_head_9__102_, data_head_9__101_, data_head_9__100_, data_head_9__99_, data_head_9__98_, data_head_9__97_, data_head_9__96_, data_head_9__95_, data_head_9__94_, data_head_9__93_, data_head_9__92_, data_head_9__91_, data_head_9__90_, data_head_9__89_, data_head_9__88_, data_head_9__87_, data_head_9__86_, data_head_9__85_, data_head_9__84_, data_head_9__83_, data_head_9__82_, data_head_9__81_, data_head_9__80_, data_head_9__79_, data_head_9__78_, data_head_9__77_, data_head_9__76_, data_head_9__75_, data_head_9__74_, data_head_9__73_, data_head_9__72_, data_head_9__71_, data_head_9__70_, data_head_9__69_, data_head_9__68_, data_head_9__67_, data_head_9__66_, data_head_9__65_, data_head_9__64_, data_head_9__63_, data_head_9__62_, data_head_9__61_, data_head_9__60_, data_head_9__59_, data_head_9__58_, data_head_9__57_, data_head_9__56_, data_head_9__55_, data_head_9__54_, data_head_9__53_, data_head_9__52_, data_head_9__51_, data_head_9__50_, data_head_9__49_, data_head_9__48_, data_head_9__47_, data_head_9__46_, data_head_9__45_, data_head_9__44_, data_head_9__43_, data_head_9__42_, data_head_9__41_, data_head_9__40_, data_head_9__39_, data_head_9__38_, data_head_9__37_, data_head_9__36_, data_head_9__35_, data_head_9__34_, data_head_9__33_, data_head_9__32_, data_head_9__31_, data_head_9__30_, data_head_9__29_, data_head_9__28_, data_head_9__27_, data_head_9__26_, data_head_9__25_, data_head_9__24_, data_head_9__23_, data_head_9__22_, data_head_9__21_, data_head_9__20_, data_head_9__19_, data_head_9__18_, data_head_9__17_, data_head_9__16_, data_head_9__15_, data_head_9__14_, data_head_9__13_, data_head_9__12_, data_head_9__11_, data_head_9__10_, data_head_9__9_, data_head_9__8_, data_head_9__7_, data_head_9__6_, data_head_9__5_, data_head_9__4_, data_head_9__3_, data_head_9__2_, data_head_9__1_, data_head_9__0_ }),
    .valid_head_o({ valid_head_9__9_, valid_head_9__8_, valid_head_9__7_, valid_head_9__6_, valid_head_9__5_, valid_head_9__4_, valid_head_9__3_, valid_head_9__2_, valid_head_9__1_, valid_head_9__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .yumi_o({ yumi_int_o_9__9_, yumi_int_o_9__8_, yumi_int_o_9__7_, yumi_int_o_9__6_, yumi_int_o_9__5_, yumi_int_o_9__4_, yumi_int_o_9__3_, yumi_int_o_9__2_, yumi_int_o_9__1_, yumi_int_o_9__0_ })
  );


  bsg_rr_f2f_middle_width_p128_middle_meet_p10
  brrf2fm
  (
    .valid_head_i({ n_2_net__9_, n_2_net__8_, n_2_net__7_, n_2_net__6_, n_2_net__5_, n_2_net__4_, n_2_net__3_, n_2_net__2_, n_2_net__1_, n_2_net__0_ }),
    .ready_head_i({ n_3_net__9_, n_3_net__8_, n_3_net__7_, n_3_net__6_, n_3_net__5_, n_3_net__4_, n_3_net__3_, n_3_net__2_, n_3_net__1_, n_3_net__0_ }),
    .go_channels_o(go_channels),
    .go_cnt_o(go_cnt)
  );


  bsg_make_2D_array_width_p128_items_p10
  oc_9__out_chan_bm2Da
  (
    .i({ n_4_net__1279_, n_4_net__1278_, n_4_net__1277_, n_4_net__1276_, n_4_net__1275_, n_4_net__1274_, n_4_net__1273_, n_4_net__1272_, n_4_net__1271_, n_4_net__1270_, n_4_net__1269_, n_4_net__1268_, n_4_net__1267_, n_4_net__1266_, n_4_net__1265_, n_4_net__1264_, n_4_net__1263_, n_4_net__1262_, n_4_net__1261_, n_4_net__1260_, n_4_net__1259_, n_4_net__1258_, n_4_net__1257_, n_4_net__1256_, n_4_net__1255_, n_4_net__1254_, n_4_net__1253_, n_4_net__1252_, n_4_net__1251_, n_4_net__1250_, n_4_net__1249_, n_4_net__1248_, n_4_net__1247_, n_4_net__1246_, n_4_net__1245_, n_4_net__1244_, n_4_net__1243_, n_4_net__1242_, n_4_net__1241_, n_4_net__1240_, n_4_net__1239_, n_4_net__1238_, n_4_net__1237_, n_4_net__1236_, n_4_net__1235_, n_4_net__1234_, n_4_net__1233_, n_4_net__1232_, n_4_net__1231_, n_4_net__1230_, n_4_net__1229_, n_4_net__1228_, n_4_net__1227_, n_4_net__1226_, n_4_net__1225_, n_4_net__1224_, n_4_net__1223_, n_4_net__1222_, n_4_net__1221_, n_4_net__1220_, n_4_net__1219_, n_4_net__1218_, n_4_net__1217_, n_4_net__1216_, n_4_net__1215_, n_4_net__1214_, n_4_net__1213_, n_4_net__1212_, n_4_net__1211_, n_4_net__1210_, n_4_net__1209_, n_4_net__1208_, n_4_net__1207_, n_4_net__1206_, n_4_net__1205_, n_4_net__1204_, n_4_net__1203_, n_4_net__1202_, n_4_net__1201_, n_4_net__1200_, n_4_net__1199_, n_4_net__1198_, n_4_net__1197_, n_4_net__1196_, n_4_net__1195_, n_4_net__1194_, n_4_net__1193_, n_4_net__1192_, n_4_net__1191_, n_4_net__1190_, n_4_net__1189_, n_4_net__1188_, n_4_net__1187_, n_4_net__1186_, n_4_net__1185_, n_4_net__1184_, n_4_net__1183_, n_4_net__1182_, n_4_net__1181_, n_4_net__1180_, n_4_net__1179_, n_4_net__1178_, n_4_net__1177_, n_4_net__1176_, n_4_net__1175_, n_4_net__1174_, n_4_net__1173_, n_4_net__1172_, n_4_net__1171_, n_4_net__1170_, n_4_net__1169_, n_4_net__1168_, n_4_net__1167_, n_4_net__1166_, n_4_net__1165_, n_4_net__1164_, n_4_net__1163_, n_4_net__1162_, n_4_net__1161_, n_4_net__1160_, n_4_net__1159_, n_4_net__1158_, n_4_net__1157_, n_4_net__1156_, n_4_net__1155_, n_4_net__1154_, n_4_net__1153_, n_4_net__1152_, n_4_net__1151_, n_4_net__1150_, n_4_net__1149_, n_4_net__1148_, n_4_net__1147_, n_4_net__1146_, n_4_net__1145_, n_4_net__1144_, n_4_net__1143_, n_4_net__1142_, n_4_net__1141_, n_4_net__1140_, n_4_net__1139_, n_4_net__1138_, n_4_net__1137_, n_4_net__1136_, n_4_net__1135_, n_4_net__1134_, n_4_net__1133_, n_4_net__1132_, n_4_net__1131_, n_4_net__1130_, n_4_net__1129_, n_4_net__1128_, n_4_net__1127_, n_4_net__1126_, n_4_net__1125_, n_4_net__1124_, n_4_net__1123_, n_4_net__1122_, n_4_net__1121_, n_4_net__1120_, n_4_net__1119_, n_4_net__1118_, n_4_net__1117_, n_4_net__1116_, n_4_net__1115_, n_4_net__1114_, n_4_net__1113_, n_4_net__1112_, n_4_net__1111_, n_4_net__1110_, n_4_net__1109_, n_4_net__1108_, n_4_net__1107_, n_4_net__1106_, n_4_net__1105_, n_4_net__1104_, n_4_net__1103_, n_4_net__1102_, n_4_net__1101_, n_4_net__1100_, n_4_net__1099_, n_4_net__1098_, n_4_net__1097_, n_4_net__1096_, n_4_net__1095_, n_4_net__1094_, n_4_net__1093_, n_4_net__1092_, n_4_net__1091_, n_4_net__1090_, n_4_net__1089_, n_4_net__1088_, n_4_net__1087_, n_4_net__1086_, n_4_net__1085_, n_4_net__1084_, n_4_net__1083_, n_4_net__1082_, n_4_net__1081_, n_4_net__1080_, n_4_net__1079_, n_4_net__1078_, n_4_net__1077_, n_4_net__1076_, n_4_net__1075_, n_4_net__1074_, n_4_net__1073_, n_4_net__1072_, n_4_net__1071_, n_4_net__1070_, n_4_net__1069_, n_4_net__1068_, n_4_net__1067_, n_4_net__1066_, n_4_net__1065_, n_4_net__1064_, n_4_net__1063_, n_4_net__1062_, n_4_net__1061_, n_4_net__1060_, n_4_net__1059_, n_4_net__1058_, n_4_net__1057_, n_4_net__1056_, n_4_net__1055_, n_4_net__1054_, n_4_net__1053_, n_4_net__1052_, n_4_net__1051_, n_4_net__1050_, n_4_net__1049_, n_4_net__1048_, n_4_net__1047_, n_4_net__1046_, n_4_net__1045_, n_4_net__1044_, n_4_net__1043_, n_4_net__1042_, n_4_net__1041_, n_4_net__1040_, n_4_net__1039_, n_4_net__1038_, n_4_net__1037_, n_4_net__1036_, n_4_net__1035_, n_4_net__1034_, n_4_net__1033_, n_4_net__1032_, n_4_net__1031_, n_4_net__1030_, n_4_net__1029_, n_4_net__1028_, n_4_net__1027_, n_4_net__1026_, n_4_net__1025_, n_4_net__1024_, n_4_net__1023_, n_4_net__1022_, n_4_net__1021_, n_4_net__1020_, n_4_net__1019_, n_4_net__1018_, n_4_net__1017_, n_4_net__1016_, n_4_net__1015_, n_4_net__1014_, n_4_net__1013_, n_4_net__1012_, n_4_net__1011_, n_4_net__1010_, n_4_net__1009_, n_4_net__1008_, n_4_net__1007_, n_4_net__1006_, n_4_net__1005_, n_4_net__1004_, n_4_net__1003_, n_4_net__1002_, n_4_net__1001_, n_4_net__1000_, n_4_net__999_, n_4_net__998_, n_4_net__997_, n_4_net__996_, n_4_net__995_, n_4_net__994_, n_4_net__993_, n_4_net__992_, n_4_net__991_, n_4_net__990_, n_4_net__989_, n_4_net__988_, n_4_net__987_, n_4_net__986_, n_4_net__985_, n_4_net__984_, n_4_net__983_, n_4_net__982_, n_4_net__981_, n_4_net__980_, n_4_net__979_, n_4_net__978_, n_4_net__977_, n_4_net__976_, n_4_net__975_, n_4_net__974_, n_4_net__973_, n_4_net__972_, n_4_net__971_, n_4_net__970_, n_4_net__969_, n_4_net__968_, n_4_net__967_, n_4_net__966_, n_4_net__965_, n_4_net__964_, n_4_net__963_, n_4_net__962_, n_4_net__961_, n_4_net__960_, n_4_net__959_, n_4_net__958_, n_4_net__957_, n_4_net__956_, n_4_net__955_, n_4_net__954_, n_4_net__953_, n_4_net__952_, n_4_net__951_, n_4_net__950_, n_4_net__949_, n_4_net__948_, n_4_net__947_, n_4_net__946_, n_4_net__945_, n_4_net__944_, n_4_net__943_, n_4_net__942_, n_4_net__941_, n_4_net__940_, n_4_net__939_, n_4_net__938_, n_4_net__937_, n_4_net__936_, n_4_net__935_, n_4_net__934_, n_4_net__933_, n_4_net__932_, n_4_net__931_, n_4_net__930_, n_4_net__929_, n_4_net__928_, n_4_net__927_, n_4_net__926_, n_4_net__925_, n_4_net__924_, n_4_net__923_, n_4_net__922_, n_4_net__921_, n_4_net__920_, n_4_net__919_, n_4_net__918_, n_4_net__917_, n_4_net__916_, n_4_net__915_, n_4_net__914_, n_4_net__913_, n_4_net__912_, n_4_net__911_, n_4_net__910_, n_4_net__909_, n_4_net__908_, n_4_net__907_, n_4_net__906_, n_4_net__905_, n_4_net__904_, n_4_net__903_, n_4_net__902_, n_4_net__901_, n_4_net__900_, n_4_net__899_, n_4_net__898_, n_4_net__897_, n_4_net__896_, n_4_net__895_, n_4_net__894_, n_4_net__893_, n_4_net__892_, n_4_net__891_, n_4_net__890_, n_4_net__889_, n_4_net__888_, n_4_net__887_, n_4_net__886_, n_4_net__885_, n_4_net__884_, n_4_net__883_, n_4_net__882_, n_4_net__881_, n_4_net__880_, n_4_net__879_, n_4_net__878_, n_4_net__877_, n_4_net__876_, n_4_net__875_, n_4_net__874_, n_4_net__873_, n_4_net__872_, n_4_net__871_, n_4_net__870_, n_4_net__869_, n_4_net__868_, n_4_net__867_, n_4_net__866_, n_4_net__865_, n_4_net__864_, n_4_net__863_, n_4_net__862_, n_4_net__861_, n_4_net__860_, n_4_net__859_, n_4_net__858_, n_4_net__857_, n_4_net__856_, n_4_net__855_, n_4_net__854_, n_4_net__853_, n_4_net__852_, n_4_net__851_, n_4_net__850_, n_4_net__849_, n_4_net__848_, n_4_net__847_, n_4_net__846_, n_4_net__845_, n_4_net__844_, n_4_net__843_, n_4_net__842_, n_4_net__841_, n_4_net__840_, n_4_net__839_, n_4_net__838_, n_4_net__837_, n_4_net__836_, n_4_net__835_, n_4_net__834_, n_4_net__833_, n_4_net__832_, n_4_net__831_, n_4_net__830_, n_4_net__829_, n_4_net__828_, n_4_net__827_, n_4_net__826_, n_4_net__825_, n_4_net__824_, n_4_net__823_, n_4_net__822_, n_4_net__821_, n_4_net__820_, n_4_net__819_, n_4_net__818_, n_4_net__817_, n_4_net__816_, n_4_net__815_, n_4_net__814_, n_4_net__813_, n_4_net__812_, n_4_net__811_, n_4_net__810_, n_4_net__809_, n_4_net__808_, n_4_net__807_, n_4_net__806_, n_4_net__805_, n_4_net__804_, n_4_net__803_, n_4_net__802_, n_4_net__801_, n_4_net__800_, n_4_net__799_, n_4_net__798_, n_4_net__797_, n_4_net__796_, n_4_net__795_, n_4_net__794_, n_4_net__793_, n_4_net__792_, n_4_net__791_, n_4_net__790_, n_4_net__789_, n_4_net__788_, n_4_net__787_, n_4_net__786_, n_4_net__785_, n_4_net__784_, n_4_net__783_, n_4_net__782_, n_4_net__781_, n_4_net__780_, n_4_net__779_, n_4_net__778_, n_4_net__777_, n_4_net__776_, n_4_net__775_, n_4_net__774_, n_4_net__773_, n_4_net__772_, n_4_net__771_, n_4_net__770_, n_4_net__769_, n_4_net__768_, n_4_net__767_, n_4_net__766_, n_4_net__765_, n_4_net__764_, n_4_net__763_, n_4_net__762_, n_4_net__761_, n_4_net__760_, n_4_net__759_, n_4_net__758_, n_4_net__757_, n_4_net__756_, n_4_net__755_, n_4_net__754_, n_4_net__753_, n_4_net__752_, n_4_net__751_, n_4_net__750_, n_4_net__749_, n_4_net__748_, n_4_net__747_, n_4_net__746_, n_4_net__745_, n_4_net__744_, n_4_net__743_, n_4_net__742_, n_4_net__741_, n_4_net__740_, n_4_net__739_, n_4_net__738_, n_4_net__737_, n_4_net__736_, n_4_net__735_, n_4_net__734_, n_4_net__733_, n_4_net__732_, n_4_net__731_, n_4_net__730_, n_4_net__729_, n_4_net__728_, n_4_net__727_, n_4_net__726_, n_4_net__725_, n_4_net__724_, n_4_net__723_, n_4_net__722_, n_4_net__721_, n_4_net__720_, n_4_net__719_, n_4_net__718_, n_4_net__717_, n_4_net__716_, n_4_net__715_, n_4_net__714_, n_4_net__713_, n_4_net__712_, n_4_net__711_, n_4_net__710_, n_4_net__709_, n_4_net__708_, n_4_net__707_, n_4_net__706_, n_4_net__705_, n_4_net__704_, n_4_net__703_, n_4_net__702_, n_4_net__701_, n_4_net__700_, n_4_net__699_, n_4_net__698_, n_4_net__697_, n_4_net__696_, n_4_net__695_, n_4_net__694_, n_4_net__693_, n_4_net__692_, n_4_net__691_, n_4_net__690_, n_4_net__689_, n_4_net__688_, n_4_net__687_, n_4_net__686_, n_4_net__685_, n_4_net__684_, n_4_net__683_, n_4_net__682_, n_4_net__681_, n_4_net__680_, n_4_net__679_, n_4_net__678_, n_4_net__677_, n_4_net__676_, n_4_net__675_, n_4_net__674_, n_4_net__673_, n_4_net__672_, n_4_net__671_, n_4_net__670_, n_4_net__669_, n_4_net__668_, n_4_net__667_, n_4_net__666_, n_4_net__665_, n_4_net__664_, n_4_net__663_, n_4_net__662_, n_4_net__661_, n_4_net__660_, n_4_net__659_, n_4_net__658_, n_4_net__657_, n_4_net__656_, n_4_net__655_, n_4_net__654_, n_4_net__653_, n_4_net__652_, n_4_net__651_, n_4_net__650_, n_4_net__649_, n_4_net__648_, n_4_net__647_, n_4_net__646_, n_4_net__645_, n_4_net__644_, n_4_net__643_, n_4_net__642_, n_4_net__641_, n_4_net__640_, n_4_net__639_, n_4_net__638_, n_4_net__637_, n_4_net__636_, n_4_net__635_, n_4_net__634_, n_4_net__633_, n_4_net__632_, n_4_net__631_, n_4_net__630_, n_4_net__629_, n_4_net__628_, n_4_net__627_, n_4_net__626_, n_4_net__625_, n_4_net__624_, n_4_net__623_, n_4_net__622_, n_4_net__621_, n_4_net__620_, n_4_net__619_, n_4_net__618_, n_4_net__617_, n_4_net__616_, n_4_net__615_, n_4_net__614_, n_4_net__613_, n_4_net__612_, n_4_net__611_, n_4_net__610_, n_4_net__609_, n_4_net__608_, n_4_net__607_, n_4_net__606_, n_4_net__605_, n_4_net__604_, n_4_net__603_, n_4_net__602_, n_4_net__601_, n_4_net__600_, n_4_net__599_, n_4_net__598_, n_4_net__597_, n_4_net__596_, n_4_net__595_, n_4_net__594_, n_4_net__593_, n_4_net__592_, n_4_net__591_, n_4_net__590_, n_4_net__589_, n_4_net__588_, n_4_net__587_, n_4_net__586_, n_4_net__585_, n_4_net__584_, n_4_net__583_, n_4_net__582_, n_4_net__581_, n_4_net__580_, n_4_net__579_, n_4_net__578_, n_4_net__577_, n_4_net__576_, n_4_net__575_, n_4_net__574_, n_4_net__573_, n_4_net__572_, n_4_net__571_, n_4_net__570_, n_4_net__569_, n_4_net__568_, n_4_net__567_, n_4_net__566_, n_4_net__565_, n_4_net__564_, n_4_net__563_, n_4_net__562_, n_4_net__561_, n_4_net__560_, n_4_net__559_, n_4_net__558_, n_4_net__557_, n_4_net__556_, n_4_net__555_, n_4_net__554_, n_4_net__553_, n_4_net__552_, n_4_net__551_, n_4_net__550_, n_4_net__549_, n_4_net__548_, n_4_net__547_, n_4_net__546_, n_4_net__545_, n_4_net__544_, n_4_net__543_, n_4_net__542_, n_4_net__541_, n_4_net__540_, n_4_net__539_, n_4_net__538_, n_4_net__537_, n_4_net__536_, n_4_net__535_, n_4_net__534_, n_4_net__533_, n_4_net__532_, n_4_net__531_, n_4_net__530_, n_4_net__529_, n_4_net__528_, n_4_net__527_, n_4_net__526_, n_4_net__525_, n_4_net__524_, n_4_net__523_, n_4_net__522_, n_4_net__521_, n_4_net__520_, n_4_net__519_, n_4_net__518_, n_4_net__517_, n_4_net__516_, n_4_net__515_, n_4_net__514_, n_4_net__513_, n_4_net__512_, n_4_net__511_, n_4_net__510_, n_4_net__509_, n_4_net__508_, n_4_net__507_, n_4_net__506_, n_4_net__505_, n_4_net__504_, n_4_net__503_, n_4_net__502_, n_4_net__501_, n_4_net__500_, n_4_net__499_, n_4_net__498_, n_4_net__497_, n_4_net__496_, n_4_net__495_, n_4_net__494_, n_4_net__493_, n_4_net__492_, n_4_net__491_, n_4_net__490_, n_4_net__489_, n_4_net__488_, n_4_net__487_, n_4_net__486_, n_4_net__485_, n_4_net__484_, n_4_net__483_, n_4_net__482_, n_4_net__481_, n_4_net__480_, n_4_net__479_, n_4_net__478_, n_4_net__477_, n_4_net__476_, n_4_net__475_, n_4_net__474_, n_4_net__473_, n_4_net__472_, n_4_net__471_, n_4_net__470_, n_4_net__469_, n_4_net__468_, n_4_net__467_, n_4_net__466_, n_4_net__465_, n_4_net__464_, n_4_net__463_, n_4_net__462_, n_4_net__461_, n_4_net__460_, n_4_net__459_, n_4_net__458_, n_4_net__457_, n_4_net__456_, n_4_net__455_, n_4_net__454_, n_4_net__453_, n_4_net__452_, n_4_net__451_, n_4_net__450_, n_4_net__449_, n_4_net__448_, n_4_net__447_, n_4_net__446_, n_4_net__445_, n_4_net__444_, n_4_net__443_, n_4_net__442_, n_4_net__441_, n_4_net__440_, n_4_net__439_, n_4_net__438_, n_4_net__437_, n_4_net__436_, n_4_net__435_, n_4_net__434_, n_4_net__433_, n_4_net__432_, n_4_net__431_, n_4_net__430_, n_4_net__429_, n_4_net__428_, n_4_net__427_, n_4_net__426_, n_4_net__425_, n_4_net__424_, n_4_net__423_, n_4_net__422_, n_4_net__421_, n_4_net__420_, n_4_net__419_, n_4_net__418_, n_4_net__417_, n_4_net__416_, n_4_net__415_, n_4_net__414_, n_4_net__413_, n_4_net__412_, n_4_net__411_, n_4_net__410_, n_4_net__409_, n_4_net__408_, n_4_net__407_, n_4_net__406_, n_4_net__405_, n_4_net__404_, n_4_net__403_, n_4_net__402_, n_4_net__401_, n_4_net__400_, n_4_net__399_, n_4_net__398_, n_4_net__397_, n_4_net__396_, n_4_net__395_, n_4_net__394_, n_4_net__393_, n_4_net__392_, n_4_net__391_, n_4_net__390_, n_4_net__389_, n_4_net__388_, n_4_net__387_, n_4_net__386_, n_4_net__385_, n_4_net__384_, n_4_net__383_, n_4_net__382_, n_4_net__381_, n_4_net__380_, n_4_net__379_, n_4_net__378_, n_4_net__377_, n_4_net__376_, n_4_net__375_, n_4_net__374_, n_4_net__373_, n_4_net__372_, n_4_net__371_, n_4_net__370_, n_4_net__369_, n_4_net__368_, n_4_net__367_, n_4_net__366_, n_4_net__365_, n_4_net__364_, n_4_net__363_, n_4_net__362_, n_4_net__361_, n_4_net__360_, n_4_net__359_, n_4_net__358_, n_4_net__357_, n_4_net__356_, n_4_net__355_, n_4_net__354_, n_4_net__353_, n_4_net__352_, n_4_net__351_, n_4_net__350_, n_4_net__349_, n_4_net__348_, n_4_net__347_, n_4_net__346_, n_4_net__345_, n_4_net__344_, n_4_net__343_, n_4_net__342_, n_4_net__341_, n_4_net__340_, n_4_net__339_, n_4_net__338_, n_4_net__337_, n_4_net__336_, n_4_net__335_, n_4_net__334_, n_4_net__333_, n_4_net__332_, n_4_net__331_, n_4_net__330_, n_4_net__329_, n_4_net__328_, n_4_net__327_, n_4_net__326_, n_4_net__325_, n_4_net__324_, n_4_net__323_, n_4_net__322_, n_4_net__321_, n_4_net__320_, n_4_net__319_, n_4_net__318_, n_4_net__317_, n_4_net__316_, n_4_net__315_, n_4_net__314_, n_4_net__313_, n_4_net__312_, n_4_net__311_, n_4_net__310_, n_4_net__309_, n_4_net__308_, n_4_net__307_, n_4_net__306_, n_4_net__305_, n_4_net__304_, n_4_net__303_, n_4_net__302_, n_4_net__301_, n_4_net__300_, n_4_net__299_, n_4_net__298_, n_4_net__297_, n_4_net__296_, n_4_net__295_, n_4_net__294_, n_4_net__293_, n_4_net__292_, n_4_net__291_, n_4_net__290_, n_4_net__289_, n_4_net__288_, n_4_net__287_, n_4_net__286_, n_4_net__285_, n_4_net__284_, n_4_net__283_, n_4_net__282_, n_4_net__281_, n_4_net__280_, n_4_net__279_, n_4_net__278_, n_4_net__277_, n_4_net__276_, n_4_net__275_, n_4_net__274_, n_4_net__273_, n_4_net__272_, n_4_net__271_, n_4_net__270_, n_4_net__269_, n_4_net__268_, n_4_net__267_, n_4_net__266_, n_4_net__265_, n_4_net__264_, n_4_net__263_, n_4_net__262_, n_4_net__261_, n_4_net__260_, n_4_net__259_, n_4_net__258_, n_4_net__257_, n_4_net__256_, n_4_net__255_, n_4_net__254_, n_4_net__253_, n_4_net__252_, n_4_net__251_, n_4_net__250_, n_4_net__249_, n_4_net__248_, n_4_net__247_, n_4_net__246_, n_4_net__245_, n_4_net__244_, n_4_net__243_, n_4_net__242_, n_4_net__241_, n_4_net__240_, n_4_net__239_, n_4_net__238_, n_4_net__237_, n_4_net__236_, n_4_net__235_, n_4_net__234_, n_4_net__233_, n_4_net__232_, n_4_net__231_, n_4_net__230_, n_4_net__229_, n_4_net__228_, n_4_net__227_, n_4_net__226_, n_4_net__225_, n_4_net__224_, n_4_net__223_, n_4_net__222_, n_4_net__221_, n_4_net__220_, n_4_net__219_, n_4_net__218_, n_4_net__217_, n_4_net__216_, n_4_net__215_, n_4_net__214_, n_4_net__213_, n_4_net__212_, n_4_net__211_, n_4_net__210_, n_4_net__209_, n_4_net__208_, n_4_net__207_, n_4_net__206_, n_4_net__205_, n_4_net__204_, n_4_net__203_, n_4_net__202_, n_4_net__201_, n_4_net__200_, n_4_net__199_, n_4_net__198_, n_4_net__197_, n_4_net__196_, n_4_net__195_, n_4_net__194_, n_4_net__193_, n_4_net__192_, n_4_net__191_, n_4_net__190_, n_4_net__189_, n_4_net__188_, n_4_net__187_, n_4_net__186_, n_4_net__185_, n_4_net__184_, n_4_net__183_, n_4_net__182_, n_4_net__181_, n_4_net__180_, n_4_net__179_, n_4_net__178_, n_4_net__177_, n_4_net__176_, n_4_net__175_, n_4_net__174_, n_4_net__173_, n_4_net__172_, n_4_net__171_, n_4_net__170_, n_4_net__169_, n_4_net__168_, n_4_net__167_, n_4_net__166_, n_4_net__165_, n_4_net__164_, n_4_net__163_, n_4_net__162_, n_4_net__161_, n_4_net__160_, n_4_net__159_, n_4_net__158_, n_4_net__157_, n_4_net__156_, n_4_net__155_, n_4_net__154_, n_4_net__153_, n_4_net__152_, n_4_net__151_, n_4_net__150_, n_4_net__149_, n_4_net__148_, n_4_net__147_, n_4_net__146_, n_4_net__145_, n_4_net__144_, n_4_net__143_, n_4_net__142_, n_4_net__141_, n_4_net__140_, n_4_net__139_, n_4_net__138_, n_4_net__137_, n_4_net__136_, n_4_net__135_, n_4_net__134_, n_4_net__133_, n_4_net__132_, n_4_net__131_, n_4_net__130_, n_4_net__129_, n_4_net__128_, n_4_net__127_, n_4_net__126_, n_4_net__125_, n_4_net__124_, n_4_net__123_, n_4_net__122_, n_4_net__121_, n_4_net__120_, n_4_net__119_, n_4_net__118_, n_4_net__117_, n_4_net__116_, n_4_net__115_, n_4_net__114_, n_4_net__113_, n_4_net__112_, n_4_net__111_, n_4_net__110_, n_4_net__109_, n_4_net__108_, n_4_net__107_, n_4_net__106_, n_4_net__105_, n_4_net__104_, n_4_net__103_, n_4_net__102_, n_4_net__101_, n_4_net__100_, n_4_net__99_, n_4_net__98_, n_4_net__97_, n_4_net__96_, n_4_net__95_, n_4_net__94_, n_4_net__93_, n_4_net__92_, n_4_net__91_, n_4_net__90_, n_4_net__89_, n_4_net__88_, n_4_net__87_, n_4_net__86_, n_4_net__85_, n_4_net__84_, n_4_net__83_, n_4_net__82_, n_4_net__81_, n_4_net__80_, n_4_net__79_, n_4_net__78_, n_4_net__77_, n_4_net__76_, n_4_net__75_, n_4_net__74_, n_4_net__73_, n_4_net__72_, n_4_net__71_, n_4_net__70_, n_4_net__69_, n_4_net__68_, n_4_net__67_, n_4_net__66_, n_4_net__65_, n_4_net__64_, n_4_net__63_, n_4_net__62_, n_4_net__61_, n_4_net__60_, n_4_net__59_, n_4_net__58_, n_4_net__57_, n_4_net__56_, n_4_net__55_, n_4_net__54_, n_4_net__53_, n_4_net__52_, n_4_net__51_, n_4_net__50_, n_4_net__49_, n_4_net__48_, n_4_net__47_, n_4_net__46_, n_4_net__45_, n_4_net__44_, n_4_net__43_, n_4_net__42_, n_4_net__41_, n_4_net__40_, n_4_net__39_, n_4_net__38_, n_4_net__37_, n_4_net__36_, n_4_net__35_, n_4_net__34_, n_4_net__33_, n_4_net__32_, n_4_net__31_, n_4_net__30_, n_4_net__29_, n_4_net__28_, n_4_net__27_, n_4_net__26_, n_4_net__25_, n_4_net__24_, n_4_net__23_, n_4_net__22_, n_4_net__21_, n_4_net__20_, n_4_net__19_, n_4_net__18_, n_4_net__17_, n_4_net__16_, n_4_net__15_, n_4_net__14_, n_4_net__13_, n_4_net__12_, n_4_net__11_, n_4_net__10_, n_4_net__9_, n_4_net__8_, n_4_net__7_, n_4_net__6_, n_4_net__5_, n_4_net__4_, n_4_net__3_, n_4_net__2_, n_4_net__1_, n_4_net__0_ }),
    .o(oc_9__out_chan_data_head_array)
  );


  bsg_rr_f2f_output_width_p128_num_out_p10_middle_meet_p10
  oc_9__out_chan_bsg_rr_ff_out
  (
    .clk(clk),
    .reset(n_5_net_),
    .ready_i(ready_i),
    .ready_head_o({ ready_head_9__9_, ready_head_9__8_, ready_head_9__7_, ready_head_9__6_, ready_head_9__5_, ready_head_9__4_, ready_head_9__3_, ready_head_9__2_, ready_head_9__1_, ready_head_9__0_ }),
    .go_channels_i(go_channels),
    .go_cnt_i(go_cnt),
    .data_head_i(oc_9__out_chan_data_head_array),
    .valid_o({ valid_int_o_9__9_, valid_int_o_9__8_, valid_int_o_9__7_, valid_int_o_9__6_, valid_int_o_9__5_, valid_int_o_9__4_, valid_int_o_9__3_, valid_int_o_9__2_, valid_int_o_9__1_, valid_int_o_9__0_ }),
    .data_o({ data_int_o_9__1279_, data_int_o_9__1278_, data_int_o_9__1277_, data_int_o_9__1276_, data_int_o_9__1275_, data_int_o_9__1274_, data_int_o_9__1273_, data_int_o_9__1272_, data_int_o_9__1271_, data_int_o_9__1270_, data_int_o_9__1269_, data_int_o_9__1268_, data_int_o_9__1267_, data_int_o_9__1266_, data_int_o_9__1265_, data_int_o_9__1264_, data_int_o_9__1263_, data_int_o_9__1262_, data_int_o_9__1261_, data_int_o_9__1260_, data_int_o_9__1259_, data_int_o_9__1258_, data_int_o_9__1257_, data_int_o_9__1256_, data_int_o_9__1255_, data_int_o_9__1254_, data_int_o_9__1253_, data_int_o_9__1252_, data_int_o_9__1251_, data_int_o_9__1250_, data_int_o_9__1249_, data_int_o_9__1248_, data_int_o_9__1247_, data_int_o_9__1246_, data_int_o_9__1245_, data_int_o_9__1244_, data_int_o_9__1243_, data_int_o_9__1242_, data_int_o_9__1241_, data_int_o_9__1240_, data_int_o_9__1239_, data_int_o_9__1238_, data_int_o_9__1237_, data_int_o_9__1236_, data_int_o_9__1235_, data_int_o_9__1234_, data_int_o_9__1233_, data_int_o_9__1232_, data_int_o_9__1231_, data_int_o_9__1230_, data_int_o_9__1229_, data_int_o_9__1228_, data_int_o_9__1227_, data_int_o_9__1226_, data_int_o_9__1225_, data_int_o_9__1224_, data_int_o_9__1223_, data_int_o_9__1222_, data_int_o_9__1221_, data_int_o_9__1220_, data_int_o_9__1219_, data_int_o_9__1218_, data_int_o_9__1217_, data_int_o_9__1216_, data_int_o_9__1215_, data_int_o_9__1214_, data_int_o_9__1213_, data_int_o_9__1212_, data_int_o_9__1211_, data_int_o_9__1210_, data_int_o_9__1209_, data_int_o_9__1208_, data_int_o_9__1207_, data_int_o_9__1206_, data_int_o_9__1205_, data_int_o_9__1204_, data_int_o_9__1203_, data_int_o_9__1202_, data_int_o_9__1201_, data_int_o_9__1200_, data_int_o_9__1199_, data_int_o_9__1198_, data_int_o_9__1197_, data_int_o_9__1196_, data_int_o_9__1195_, data_int_o_9__1194_, data_int_o_9__1193_, data_int_o_9__1192_, data_int_o_9__1191_, data_int_o_9__1190_, data_int_o_9__1189_, data_int_o_9__1188_, data_int_o_9__1187_, data_int_o_9__1186_, data_int_o_9__1185_, data_int_o_9__1184_, data_int_o_9__1183_, data_int_o_9__1182_, data_int_o_9__1181_, data_int_o_9__1180_, data_int_o_9__1179_, data_int_o_9__1178_, data_int_o_9__1177_, data_int_o_9__1176_, data_int_o_9__1175_, data_int_o_9__1174_, data_int_o_9__1173_, data_int_o_9__1172_, data_int_o_9__1171_, data_int_o_9__1170_, data_int_o_9__1169_, data_int_o_9__1168_, data_int_o_9__1167_, data_int_o_9__1166_, data_int_o_9__1165_, data_int_o_9__1164_, data_int_o_9__1163_, data_int_o_9__1162_, data_int_o_9__1161_, data_int_o_9__1160_, data_int_o_9__1159_, data_int_o_9__1158_, data_int_o_9__1157_, data_int_o_9__1156_, data_int_o_9__1155_, data_int_o_9__1154_, data_int_o_9__1153_, data_int_o_9__1152_, data_int_o_9__1151_, data_int_o_9__1150_, data_int_o_9__1149_, data_int_o_9__1148_, data_int_o_9__1147_, data_int_o_9__1146_, data_int_o_9__1145_, data_int_o_9__1144_, data_int_o_9__1143_, data_int_o_9__1142_, data_int_o_9__1141_, data_int_o_9__1140_, data_int_o_9__1139_, data_int_o_9__1138_, data_int_o_9__1137_, data_int_o_9__1136_, data_int_o_9__1135_, data_int_o_9__1134_, data_int_o_9__1133_, data_int_o_9__1132_, data_int_o_9__1131_, data_int_o_9__1130_, data_int_o_9__1129_, data_int_o_9__1128_, data_int_o_9__1127_, data_int_o_9__1126_, data_int_o_9__1125_, data_int_o_9__1124_, data_int_o_9__1123_, data_int_o_9__1122_, data_int_o_9__1121_, data_int_o_9__1120_, data_int_o_9__1119_, data_int_o_9__1118_, data_int_o_9__1117_, data_int_o_9__1116_, data_int_o_9__1115_, data_int_o_9__1114_, data_int_o_9__1113_, data_int_o_9__1112_, data_int_o_9__1111_, data_int_o_9__1110_, data_int_o_9__1109_, data_int_o_9__1108_, data_int_o_9__1107_, data_int_o_9__1106_, data_int_o_9__1105_, data_int_o_9__1104_, data_int_o_9__1103_, data_int_o_9__1102_, data_int_o_9__1101_, data_int_o_9__1100_, data_int_o_9__1099_, data_int_o_9__1098_, data_int_o_9__1097_, data_int_o_9__1096_, data_int_o_9__1095_, data_int_o_9__1094_, data_int_o_9__1093_, data_int_o_9__1092_, data_int_o_9__1091_, data_int_o_9__1090_, data_int_o_9__1089_, data_int_o_9__1088_, data_int_o_9__1087_, data_int_o_9__1086_, data_int_o_9__1085_, data_int_o_9__1084_, data_int_o_9__1083_, data_int_o_9__1082_, data_int_o_9__1081_, data_int_o_9__1080_, data_int_o_9__1079_, data_int_o_9__1078_, data_int_o_9__1077_, data_int_o_9__1076_, data_int_o_9__1075_, data_int_o_9__1074_, data_int_o_9__1073_, data_int_o_9__1072_, data_int_o_9__1071_, data_int_o_9__1070_, data_int_o_9__1069_, data_int_o_9__1068_, data_int_o_9__1067_, data_int_o_9__1066_, data_int_o_9__1065_, data_int_o_9__1064_, data_int_o_9__1063_, data_int_o_9__1062_, data_int_o_9__1061_, data_int_o_9__1060_, data_int_o_9__1059_, data_int_o_9__1058_, data_int_o_9__1057_, data_int_o_9__1056_, data_int_o_9__1055_, data_int_o_9__1054_, data_int_o_9__1053_, data_int_o_9__1052_, data_int_o_9__1051_, data_int_o_9__1050_, data_int_o_9__1049_, data_int_o_9__1048_, data_int_o_9__1047_, data_int_o_9__1046_, data_int_o_9__1045_, data_int_o_9__1044_, data_int_o_9__1043_, data_int_o_9__1042_, data_int_o_9__1041_, data_int_o_9__1040_, data_int_o_9__1039_, data_int_o_9__1038_, data_int_o_9__1037_, data_int_o_9__1036_, data_int_o_9__1035_, data_int_o_9__1034_, data_int_o_9__1033_, data_int_o_9__1032_, data_int_o_9__1031_, data_int_o_9__1030_, data_int_o_9__1029_, data_int_o_9__1028_, data_int_o_9__1027_, data_int_o_9__1026_, data_int_o_9__1025_, data_int_o_9__1024_, data_int_o_9__1023_, data_int_o_9__1022_, data_int_o_9__1021_, data_int_o_9__1020_, data_int_o_9__1019_, data_int_o_9__1018_, data_int_o_9__1017_, data_int_o_9__1016_, data_int_o_9__1015_, data_int_o_9__1014_, data_int_o_9__1013_, data_int_o_9__1012_, data_int_o_9__1011_, data_int_o_9__1010_, data_int_o_9__1009_, data_int_o_9__1008_, data_int_o_9__1007_, data_int_o_9__1006_, data_int_o_9__1005_, data_int_o_9__1004_, data_int_o_9__1003_, data_int_o_9__1002_, data_int_o_9__1001_, data_int_o_9__1000_, data_int_o_9__999_, data_int_o_9__998_, data_int_o_9__997_, data_int_o_9__996_, data_int_o_9__995_, data_int_o_9__994_, data_int_o_9__993_, data_int_o_9__992_, data_int_o_9__991_, data_int_o_9__990_, data_int_o_9__989_, data_int_o_9__988_, data_int_o_9__987_, data_int_o_9__986_, data_int_o_9__985_, data_int_o_9__984_, data_int_o_9__983_, data_int_o_9__982_, data_int_o_9__981_, data_int_o_9__980_, data_int_o_9__979_, data_int_o_9__978_, data_int_o_9__977_, data_int_o_9__976_, data_int_o_9__975_, data_int_o_9__974_, data_int_o_9__973_, data_int_o_9__972_, data_int_o_9__971_, data_int_o_9__970_, data_int_o_9__969_, data_int_o_9__968_, data_int_o_9__967_, data_int_o_9__966_, data_int_o_9__965_, data_int_o_9__964_, data_int_o_9__963_, data_int_o_9__962_, data_int_o_9__961_, data_int_o_9__960_, data_int_o_9__959_, data_int_o_9__958_, data_int_o_9__957_, data_int_o_9__956_, data_int_o_9__955_, data_int_o_9__954_, data_int_o_9__953_, data_int_o_9__952_, data_int_o_9__951_, data_int_o_9__950_, data_int_o_9__949_, data_int_o_9__948_, data_int_o_9__947_, data_int_o_9__946_, data_int_o_9__945_, data_int_o_9__944_, data_int_o_9__943_, data_int_o_9__942_, data_int_o_9__941_, data_int_o_9__940_, data_int_o_9__939_, data_int_o_9__938_, data_int_o_9__937_, data_int_o_9__936_, data_int_o_9__935_, data_int_o_9__934_, data_int_o_9__933_, data_int_o_9__932_, data_int_o_9__931_, data_int_o_9__930_, data_int_o_9__929_, data_int_o_9__928_, data_int_o_9__927_, data_int_o_9__926_, data_int_o_9__925_, data_int_o_9__924_, data_int_o_9__923_, data_int_o_9__922_, data_int_o_9__921_, data_int_o_9__920_, data_int_o_9__919_, data_int_o_9__918_, data_int_o_9__917_, data_int_o_9__916_, data_int_o_9__915_, data_int_o_9__914_, data_int_o_9__913_, data_int_o_9__912_, data_int_o_9__911_, data_int_o_9__910_, data_int_o_9__909_, data_int_o_9__908_, data_int_o_9__907_, data_int_o_9__906_, data_int_o_9__905_, data_int_o_9__904_, data_int_o_9__903_, data_int_o_9__902_, data_int_o_9__901_, data_int_o_9__900_, data_int_o_9__899_, data_int_o_9__898_, data_int_o_9__897_, data_int_o_9__896_, data_int_o_9__895_, data_int_o_9__894_, data_int_o_9__893_, data_int_o_9__892_, data_int_o_9__891_, data_int_o_9__890_, data_int_o_9__889_, data_int_o_9__888_, data_int_o_9__887_, data_int_o_9__886_, data_int_o_9__885_, data_int_o_9__884_, data_int_o_9__883_, data_int_o_9__882_, data_int_o_9__881_, data_int_o_9__880_, data_int_o_9__879_, data_int_o_9__878_, data_int_o_9__877_, data_int_o_9__876_, data_int_o_9__875_, data_int_o_9__874_, data_int_o_9__873_, data_int_o_9__872_, data_int_o_9__871_, data_int_o_9__870_, data_int_o_9__869_, data_int_o_9__868_, data_int_o_9__867_, data_int_o_9__866_, data_int_o_9__865_, data_int_o_9__864_, data_int_o_9__863_, data_int_o_9__862_, data_int_o_9__861_, data_int_o_9__860_, data_int_o_9__859_, data_int_o_9__858_, data_int_o_9__857_, data_int_o_9__856_, data_int_o_9__855_, data_int_o_9__854_, data_int_o_9__853_, data_int_o_9__852_, data_int_o_9__851_, data_int_o_9__850_, data_int_o_9__849_, data_int_o_9__848_, data_int_o_9__847_, data_int_o_9__846_, data_int_o_9__845_, data_int_o_9__844_, data_int_o_9__843_, data_int_o_9__842_, data_int_o_9__841_, data_int_o_9__840_, data_int_o_9__839_, data_int_o_9__838_, data_int_o_9__837_, data_int_o_9__836_, data_int_o_9__835_, data_int_o_9__834_, data_int_o_9__833_, data_int_o_9__832_, data_int_o_9__831_, data_int_o_9__830_, data_int_o_9__829_, data_int_o_9__828_, data_int_o_9__827_, data_int_o_9__826_, data_int_o_9__825_, data_int_o_9__824_, data_int_o_9__823_, data_int_o_9__822_, data_int_o_9__821_, data_int_o_9__820_, data_int_o_9__819_, data_int_o_9__818_, data_int_o_9__817_, data_int_o_9__816_, data_int_o_9__815_, data_int_o_9__814_, data_int_o_9__813_, data_int_o_9__812_, data_int_o_9__811_, data_int_o_9__810_, data_int_o_9__809_, data_int_o_9__808_, data_int_o_9__807_, data_int_o_9__806_, data_int_o_9__805_, data_int_o_9__804_, data_int_o_9__803_, data_int_o_9__802_, data_int_o_9__801_, data_int_o_9__800_, data_int_o_9__799_, data_int_o_9__798_, data_int_o_9__797_, data_int_o_9__796_, data_int_o_9__795_, data_int_o_9__794_, data_int_o_9__793_, data_int_o_9__792_, data_int_o_9__791_, data_int_o_9__790_, data_int_o_9__789_, data_int_o_9__788_, data_int_o_9__787_, data_int_o_9__786_, data_int_o_9__785_, data_int_o_9__784_, data_int_o_9__783_, data_int_o_9__782_, data_int_o_9__781_, data_int_o_9__780_, data_int_o_9__779_, data_int_o_9__778_, data_int_o_9__777_, data_int_o_9__776_, data_int_o_9__775_, data_int_o_9__774_, data_int_o_9__773_, data_int_o_9__772_, data_int_o_9__771_, data_int_o_9__770_, data_int_o_9__769_, data_int_o_9__768_, data_int_o_9__767_, data_int_o_9__766_, data_int_o_9__765_, data_int_o_9__764_, data_int_o_9__763_, data_int_o_9__762_, data_int_o_9__761_, data_int_o_9__760_, data_int_o_9__759_, data_int_o_9__758_, data_int_o_9__757_, data_int_o_9__756_, data_int_o_9__755_, data_int_o_9__754_, data_int_o_9__753_, data_int_o_9__752_, data_int_o_9__751_, data_int_o_9__750_, data_int_o_9__749_, data_int_o_9__748_, data_int_o_9__747_, data_int_o_9__746_, data_int_o_9__745_, data_int_o_9__744_, data_int_o_9__743_, data_int_o_9__742_, data_int_o_9__741_, data_int_o_9__740_, data_int_o_9__739_, data_int_o_9__738_, data_int_o_9__737_, data_int_o_9__736_, data_int_o_9__735_, data_int_o_9__734_, data_int_o_9__733_, data_int_o_9__732_, data_int_o_9__731_, data_int_o_9__730_, data_int_o_9__729_, data_int_o_9__728_, data_int_o_9__727_, data_int_o_9__726_, data_int_o_9__725_, data_int_o_9__724_, data_int_o_9__723_, data_int_o_9__722_, data_int_o_9__721_, data_int_o_9__720_, data_int_o_9__719_, data_int_o_9__718_, data_int_o_9__717_, data_int_o_9__716_, data_int_o_9__715_, data_int_o_9__714_, data_int_o_9__713_, data_int_o_9__712_, data_int_o_9__711_, data_int_o_9__710_, data_int_o_9__709_, data_int_o_9__708_, data_int_o_9__707_, data_int_o_9__706_, data_int_o_9__705_, data_int_o_9__704_, data_int_o_9__703_, data_int_o_9__702_, data_int_o_9__701_, data_int_o_9__700_, data_int_o_9__699_, data_int_o_9__698_, data_int_o_9__697_, data_int_o_9__696_, data_int_o_9__695_, data_int_o_9__694_, data_int_o_9__693_, data_int_o_9__692_, data_int_o_9__691_, data_int_o_9__690_, data_int_o_9__689_, data_int_o_9__688_, data_int_o_9__687_, data_int_o_9__686_, data_int_o_9__685_, data_int_o_9__684_, data_int_o_9__683_, data_int_o_9__682_, data_int_o_9__681_, data_int_o_9__680_, data_int_o_9__679_, data_int_o_9__678_, data_int_o_9__677_, data_int_o_9__676_, data_int_o_9__675_, data_int_o_9__674_, data_int_o_9__673_, data_int_o_9__672_, data_int_o_9__671_, data_int_o_9__670_, data_int_o_9__669_, data_int_o_9__668_, data_int_o_9__667_, data_int_o_9__666_, data_int_o_9__665_, data_int_o_9__664_, data_int_o_9__663_, data_int_o_9__662_, data_int_o_9__661_, data_int_o_9__660_, data_int_o_9__659_, data_int_o_9__658_, data_int_o_9__657_, data_int_o_9__656_, data_int_o_9__655_, data_int_o_9__654_, data_int_o_9__653_, data_int_o_9__652_, data_int_o_9__651_, data_int_o_9__650_, data_int_o_9__649_, data_int_o_9__648_, data_int_o_9__647_, data_int_o_9__646_, data_int_o_9__645_, data_int_o_9__644_, data_int_o_9__643_, data_int_o_9__642_, data_int_o_9__641_, data_int_o_9__640_, data_int_o_9__639_, data_int_o_9__638_, data_int_o_9__637_, data_int_o_9__636_, data_int_o_9__635_, data_int_o_9__634_, data_int_o_9__633_, data_int_o_9__632_, data_int_o_9__631_, data_int_o_9__630_, data_int_o_9__629_, data_int_o_9__628_, data_int_o_9__627_, data_int_o_9__626_, data_int_o_9__625_, data_int_o_9__624_, data_int_o_9__623_, data_int_o_9__622_, data_int_o_9__621_, data_int_o_9__620_, data_int_o_9__619_, data_int_o_9__618_, data_int_o_9__617_, data_int_o_9__616_, data_int_o_9__615_, data_int_o_9__614_, data_int_o_9__613_, data_int_o_9__612_, data_int_o_9__611_, data_int_o_9__610_, data_int_o_9__609_, data_int_o_9__608_, data_int_o_9__607_, data_int_o_9__606_, data_int_o_9__605_, data_int_o_9__604_, data_int_o_9__603_, data_int_o_9__602_, data_int_o_9__601_, data_int_o_9__600_, data_int_o_9__599_, data_int_o_9__598_, data_int_o_9__597_, data_int_o_9__596_, data_int_o_9__595_, data_int_o_9__594_, data_int_o_9__593_, data_int_o_9__592_, data_int_o_9__591_, data_int_o_9__590_, data_int_o_9__589_, data_int_o_9__588_, data_int_o_9__587_, data_int_o_9__586_, data_int_o_9__585_, data_int_o_9__584_, data_int_o_9__583_, data_int_o_9__582_, data_int_o_9__581_, data_int_o_9__580_, data_int_o_9__579_, data_int_o_9__578_, data_int_o_9__577_, data_int_o_9__576_, data_int_o_9__575_, data_int_o_9__574_, data_int_o_9__573_, data_int_o_9__572_, data_int_o_9__571_, data_int_o_9__570_, data_int_o_9__569_, data_int_o_9__568_, data_int_o_9__567_, data_int_o_9__566_, data_int_o_9__565_, data_int_o_9__564_, data_int_o_9__563_, data_int_o_9__562_, data_int_o_9__561_, data_int_o_9__560_, data_int_o_9__559_, data_int_o_9__558_, data_int_o_9__557_, data_int_o_9__556_, data_int_o_9__555_, data_int_o_9__554_, data_int_o_9__553_, data_int_o_9__552_, data_int_o_9__551_, data_int_o_9__550_, data_int_o_9__549_, data_int_o_9__548_, data_int_o_9__547_, data_int_o_9__546_, data_int_o_9__545_, data_int_o_9__544_, data_int_o_9__543_, data_int_o_9__542_, data_int_o_9__541_, data_int_o_9__540_, data_int_o_9__539_, data_int_o_9__538_, data_int_o_9__537_, data_int_o_9__536_, data_int_o_9__535_, data_int_o_9__534_, data_int_o_9__533_, data_int_o_9__532_, data_int_o_9__531_, data_int_o_9__530_, data_int_o_9__529_, data_int_o_9__528_, data_int_o_9__527_, data_int_o_9__526_, data_int_o_9__525_, data_int_o_9__524_, data_int_o_9__523_, data_int_o_9__522_, data_int_o_9__521_, data_int_o_9__520_, data_int_o_9__519_, data_int_o_9__518_, data_int_o_9__517_, data_int_o_9__516_, data_int_o_9__515_, data_int_o_9__514_, data_int_o_9__513_, data_int_o_9__512_, data_int_o_9__511_, data_int_o_9__510_, data_int_o_9__509_, data_int_o_9__508_, data_int_o_9__507_, data_int_o_9__506_, data_int_o_9__505_, data_int_o_9__504_, data_int_o_9__503_, data_int_o_9__502_, data_int_o_9__501_, data_int_o_9__500_, data_int_o_9__499_, data_int_o_9__498_, data_int_o_9__497_, data_int_o_9__496_, data_int_o_9__495_, data_int_o_9__494_, data_int_o_9__493_, data_int_o_9__492_, data_int_o_9__491_, data_int_o_9__490_, data_int_o_9__489_, data_int_o_9__488_, data_int_o_9__487_, data_int_o_9__486_, data_int_o_9__485_, data_int_o_9__484_, data_int_o_9__483_, data_int_o_9__482_, data_int_o_9__481_, data_int_o_9__480_, data_int_o_9__479_, data_int_o_9__478_, data_int_o_9__477_, data_int_o_9__476_, data_int_o_9__475_, data_int_o_9__474_, data_int_o_9__473_, data_int_o_9__472_, data_int_o_9__471_, data_int_o_9__470_, data_int_o_9__469_, data_int_o_9__468_, data_int_o_9__467_, data_int_o_9__466_, data_int_o_9__465_, data_int_o_9__464_, data_int_o_9__463_, data_int_o_9__462_, data_int_o_9__461_, data_int_o_9__460_, data_int_o_9__459_, data_int_o_9__458_, data_int_o_9__457_, data_int_o_9__456_, data_int_o_9__455_, data_int_o_9__454_, data_int_o_9__453_, data_int_o_9__452_, data_int_o_9__451_, data_int_o_9__450_, data_int_o_9__449_, data_int_o_9__448_, data_int_o_9__447_, data_int_o_9__446_, data_int_o_9__445_, data_int_o_9__444_, data_int_o_9__443_, data_int_o_9__442_, data_int_o_9__441_, data_int_o_9__440_, data_int_o_9__439_, data_int_o_9__438_, data_int_o_9__437_, data_int_o_9__436_, data_int_o_9__435_, data_int_o_9__434_, data_int_o_9__433_, data_int_o_9__432_, data_int_o_9__431_, data_int_o_9__430_, data_int_o_9__429_, data_int_o_9__428_, data_int_o_9__427_, data_int_o_9__426_, data_int_o_9__425_, data_int_o_9__424_, data_int_o_9__423_, data_int_o_9__422_, data_int_o_9__421_, data_int_o_9__420_, data_int_o_9__419_, data_int_o_9__418_, data_int_o_9__417_, data_int_o_9__416_, data_int_o_9__415_, data_int_o_9__414_, data_int_o_9__413_, data_int_o_9__412_, data_int_o_9__411_, data_int_o_9__410_, data_int_o_9__409_, data_int_o_9__408_, data_int_o_9__407_, data_int_o_9__406_, data_int_o_9__405_, data_int_o_9__404_, data_int_o_9__403_, data_int_o_9__402_, data_int_o_9__401_, data_int_o_9__400_, data_int_o_9__399_, data_int_o_9__398_, data_int_o_9__397_, data_int_o_9__396_, data_int_o_9__395_, data_int_o_9__394_, data_int_o_9__393_, data_int_o_9__392_, data_int_o_9__391_, data_int_o_9__390_, data_int_o_9__389_, data_int_o_9__388_, data_int_o_9__387_, data_int_o_9__386_, data_int_o_9__385_, data_int_o_9__384_, data_int_o_9__383_, data_int_o_9__382_, data_int_o_9__381_, data_int_o_9__380_, data_int_o_9__379_, data_int_o_9__378_, data_int_o_9__377_, data_int_o_9__376_, data_int_o_9__375_, data_int_o_9__374_, data_int_o_9__373_, data_int_o_9__372_, data_int_o_9__371_, data_int_o_9__370_, data_int_o_9__369_, data_int_o_9__368_, data_int_o_9__367_, data_int_o_9__366_, data_int_o_9__365_, data_int_o_9__364_, data_int_o_9__363_, data_int_o_9__362_, data_int_o_9__361_, data_int_o_9__360_, data_int_o_9__359_, data_int_o_9__358_, data_int_o_9__357_, data_int_o_9__356_, data_int_o_9__355_, data_int_o_9__354_, data_int_o_9__353_, data_int_o_9__352_, data_int_o_9__351_, data_int_o_9__350_, data_int_o_9__349_, data_int_o_9__348_, data_int_o_9__347_, data_int_o_9__346_, data_int_o_9__345_, data_int_o_9__344_, data_int_o_9__343_, data_int_o_9__342_, data_int_o_9__341_, data_int_o_9__340_, data_int_o_9__339_, data_int_o_9__338_, data_int_o_9__337_, data_int_o_9__336_, data_int_o_9__335_, data_int_o_9__334_, data_int_o_9__333_, data_int_o_9__332_, data_int_o_9__331_, data_int_o_9__330_, data_int_o_9__329_, data_int_o_9__328_, data_int_o_9__327_, data_int_o_9__326_, data_int_o_9__325_, data_int_o_9__324_, data_int_o_9__323_, data_int_o_9__322_, data_int_o_9__321_, data_int_o_9__320_, data_int_o_9__319_, data_int_o_9__318_, data_int_o_9__317_, data_int_o_9__316_, data_int_o_9__315_, data_int_o_9__314_, data_int_o_9__313_, data_int_o_9__312_, data_int_o_9__311_, data_int_o_9__310_, data_int_o_9__309_, data_int_o_9__308_, data_int_o_9__307_, data_int_o_9__306_, data_int_o_9__305_, data_int_o_9__304_, data_int_o_9__303_, data_int_o_9__302_, data_int_o_9__301_, data_int_o_9__300_, data_int_o_9__299_, data_int_o_9__298_, data_int_o_9__297_, data_int_o_9__296_, data_int_o_9__295_, data_int_o_9__294_, data_int_o_9__293_, data_int_o_9__292_, data_int_o_9__291_, data_int_o_9__290_, data_int_o_9__289_, data_int_o_9__288_, data_int_o_9__287_, data_int_o_9__286_, data_int_o_9__285_, data_int_o_9__284_, data_int_o_9__283_, data_int_o_9__282_, data_int_o_9__281_, data_int_o_9__280_, data_int_o_9__279_, data_int_o_9__278_, data_int_o_9__277_, data_int_o_9__276_, data_int_o_9__275_, data_int_o_9__274_, data_int_o_9__273_, data_int_o_9__272_, data_int_o_9__271_, data_int_o_9__270_, data_int_o_9__269_, data_int_o_9__268_, data_int_o_9__267_, data_int_o_9__266_, data_int_o_9__265_, data_int_o_9__264_, data_int_o_9__263_, data_int_o_9__262_, data_int_o_9__261_, data_int_o_9__260_, data_int_o_9__259_, data_int_o_9__258_, data_int_o_9__257_, data_int_o_9__256_, data_int_o_9__255_, data_int_o_9__254_, data_int_o_9__253_, data_int_o_9__252_, data_int_o_9__251_, data_int_o_9__250_, data_int_o_9__249_, data_int_o_9__248_, data_int_o_9__247_, data_int_o_9__246_, data_int_o_9__245_, data_int_o_9__244_, data_int_o_9__243_, data_int_o_9__242_, data_int_o_9__241_, data_int_o_9__240_, data_int_o_9__239_, data_int_o_9__238_, data_int_o_9__237_, data_int_o_9__236_, data_int_o_9__235_, data_int_o_9__234_, data_int_o_9__233_, data_int_o_9__232_, data_int_o_9__231_, data_int_o_9__230_, data_int_o_9__229_, data_int_o_9__228_, data_int_o_9__227_, data_int_o_9__226_, data_int_o_9__225_, data_int_o_9__224_, data_int_o_9__223_, data_int_o_9__222_, data_int_o_9__221_, data_int_o_9__220_, data_int_o_9__219_, data_int_o_9__218_, data_int_o_9__217_, data_int_o_9__216_, data_int_o_9__215_, data_int_o_9__214_, data_int_o_9__213_, data_int_o_9__212_, data_int_o_9__211_, data_int_o_9__210_, data_int_o_9__209_, data_int_o_9__208_, data_int_o_9__207_, data_int_o_9__206_, data_int_o_9__205_, data_int_o_9__204_, data_int_o_9__203_, data_int_o_9__202_, data_int_o_9__201_, data_int_o_9__200_, data_int_o_9__199_, data_int_o_9__198_, data_int_o_9__197_, data_int_o_9__196_, data_int_o_9__195_, data_int_o_9__194_, data_int_o_9__193_, data_int_o_9__192_, data_int_o_9__191_, data_int_o_9__190_, data_int_o_9__189_, data_int_o_9__188_, data_int_o_9__187_, data_int_o_9__186_, data_int_o_9__185_, data_int_o_9__184_, data_int_o_9__183_, data_int_o_9__182_, data_int_o_9__181_, data_int_o_9__180_, data_int_o_9__179_, data_int_o_9__178_, data_int_o_9__177_, data_int_o_9__176_, data_int_o_9__175_, data_int_o_9__174_, data_int_o_9__173_, data_int_o_9__172_, data_int_o_9__171_, data_int_o_9__170_, data_int_o_9__169_, data_int_o_9__168_, data_int_o_9__167_, data_int_o_9__166_, data_int_o_9__165_, data_int_o_9__164_, data_int_o_9__163_, data_int_o_9__162_, data_int_o_9__161_, data_int_o_9__160_, data_int_o_9__159_, data_int_o_9__158_, data_int_o_9__157_, data_int_o_9__156_, data_int_o_9__155_, data_int_o_9__154_, data_int_o_9__153_, data_int_o_9__152_, data_int_o_9__151_, data_int_o_9__150_, data_int_o_9__149_, data_int_o_9__148_, data_int_o_9__147_, data_int_o_9__146_, data_int_o_9__145_, data_int_o_9__144_, data_int_o_9__143_, data_int_o_9__142_, data_int_o_9__141_, data_int_o_9__140_, data_int_o_9__139_, data_int_o_9__138_, data_int_o_9__137_, data_int_o_9__136_, data_int_o_9__135_, data_int_o_9__134_, data_int_o_9__133_, data_int_o_9__132_, data_int_o_9__131_, data_int_o_9__130_, data_int_o_9__129_, data_int_o_9__128_, data_int_o_9__127_, data_int_o_9__126_, data_int_o_9__125_, data_int_o_9__124_, data_int_o_9__123_, data_int_o_9__122_, data_int_o_9__121_, data_int_o_9__120_, data_int_o_9__119_, data_int_o_9__118_, data_int_o_9__117_, data_int_o_9__116_, data_int_o_9__115_, data_int_o_9__114_, data_int_o_9__113_, data_int_o_9__112_, data_int_o_9__111_, data_int_o_9__110_, data_int_o_9__109_, data_int_o_9__108_, data_int_o_9__107_, data_int_o_9__106_, data_int_o_9__105_, data_int_o_9__104_, data_int_o_9__103_, data_int_o_9__102_, data_int_o_9__101_, data_int_o_9__100_, data_int_o_9__99_, data_int_o_9__98_, data_int_o_9__97_, data_int_o_9__96_, data_int_o_9__95_, data_int_o_9__94_, data_int_o_9__93_, data_int_o_9__92_, data_int_o_9__91_, data_int_o_9__90_, data_int_o_9__89_, data_int_o_9__88_, data_int_o_9__87_, data_int_o_9__86_, data_int_o_9__85_, data_int_o_9__84_, data_int_o_9__83_, data_int_o_9__82_, data_int_o_9__81_, data_int_o_9__80_, data_int_o_9__79_, data_int_o_9__78_, data_int_o_9__77_, data_int_o_9__76_, data_int_o_9__75_, data_int_o_9__74_, data_int_o_9__73_, data_int_o_9__72_, data_int_o_9__71_, data_int_o_9__70_, data_int_o_9__69_, data_int_o_9__68_, data_int_o_9__67_, data_int_o_9__66_, data_int_o_9__65_, data_int_o_9__64_, data_int_o_9__63_, data_int_o_9__62_, data_int_o_9__61_, data_int_o_9__60_, data_int_o_9__59_, data_int_o_9__58_, data_int_o_9__57_, data_int_o_9__56_, data_int_o_9__55_, data_int_o_9__54_, data_int_o_9__53_, data_int_o_9__52_, data_int_o_9__51_, data_int_o_9__50_, data_int_o_9__49_, data_int_o_9__48_, data_int_o_9__47_, data_int_o_9__46_, data_int_o_9__45_, data_int_o_9__44_, data_int_o_9__43_, data_int_o_9__42_, data_int_o_9__41_, data_int_o_9__40_, data_int_o_9__39_, data_int_o_9__38_, data_int_o_9__37_, data_int_o_9__36_, data_int_o_9__35_, data_int_o_9__34_, data_int_o_9__33_, data_int_o_9__32_, data_int_o_9__31_, data_int_o_9__30_, data_int_o_9__29_, data_int_o_9__28_, data_int_o_9__27_, data_int_o_9__26_, data_int_o_9__25_, data_int_o_9__24_, data_int_o_9__23_, data_int_o_9__22_, data_int_o_9__21_, data_int_o_9__20_, data_int_o_9__19_, data_int_o_9__18_, data_int_o_9__17_, data_int_o_9__16_, data_int_o_9__15_, data_int_o_9__14_, data_int_o_9__13_, data_int_o_9__12_, data_int_o_9__11_, data_int_o_9__10_, data_int_o_9__9_, data_int_o_9__8_, data_int_o_9__7_, data_int_o_9__6_, data_int_o_9__5_, data_int_o_9__4_, data_int_o_9__3_, data_int_o_9__2_, data_int_o_9__1_, data_int_o_9__0_ })
  );

  assign N175 = ~in_top_channel_i[3];
  assign N176 = ~in_top_channel_i[0];
  assign N177 = in_top_channel_i[2] | N175;
  assign N178 = in_top_channel_i[1] | N177;
  assign N179 = N176 | N178;
  assign N180 = ~out_top_channel_i[3];
  assign N181 = ~out_top_channel_i[0];
  assign N182 = out_top_channel_i[2] | N180;
  assign N183 = out_top_channel_i[1] | N182;
  assign N184 = N181 | N183;
  assign N125 = N0 & N1 & (N2 & N3);
  assign N0 = ~in_top_channel_i[3];
  assign N1 = ~in_top_channel_i[2];
  assign N2 = ~in_top_channel_i[0];
  assign N3 = ~in_top_channel_i[1];
  assign N126 = in_top_channel_i[3] & N4;
  assign N4 = ~in_top_channel_i[0];
  assign N127 = N5 & N6 & (in_top_channel_i[0] & N7);
  assign N5 = ~in_top_channel_i[3];
  assign N6 = ~in_top_channel_i[2];
  assign N7 = ~in_top_channel_i[1];
  assign N129 = N8 & N9 & in_top_channel_i[1];
  assign N8 = ~in_top_channel_i[2];
  assign N9 = ~in_top_channel_i[0];
  assign N130 = N10 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N10 = ~in_top_channel_i[2];
  assign N131 = in_top_channel_i[2] & N11 & N12;
  assign N11 = ~in_top_channel_i[0];
  assign N12 = ~in_top_channel_i[1];
  assign N132 = in_top_channel_i[2] & in_top_channel_i[0] & N13;
  assign N13 = ~in_top_channel_i[1];
  assign N133 = in_top_channel_i[2] & N14 & in_top_channel_i[1];
  assign N14 = ~in_top_channel_i[0];
  assign N134 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N128 = in_top_channel_i[3] & in_top_channel_i[0];
  assign N135 = N15 & N16 & (N17 & N18);
  assign N15 = ~out_top_channel_i[3];
  assign N16 = ~out_top_channel_i[2];
  assign N17 = ~out_top_channel_i[0];
  assign N18 = ~out_top_channel_i[1];
  assign N136 = out_top_channel_i[3] & N19;
  assign N19 = ~out_top_channel_i[0];
  assign N137 = N20 & N21 & (out_top_channel_i[0] & N22);
  assign N20 = ~out_top_channel_i[3];
  assign N21 = ~out_top_channel_i[2];
  assign N22 = ~out_top_channel_i[1];
  assign N139 = N23 & N24 & out_top_channel_i[1];
  assign N23 = ~out_top_channel_i[2];
  assign N24 = ~out_top_channel_i[0];
  assign N140 = N25 & out_top_channel_i[0] & out_top_channel_i[1];
  assign N25 = ~out_top_channel_i[2];
  assign N141 = out_top_channel_i[2] & N26 & N27;
  assign N26 = ~out_top_channel_i[0];
  assign N27 = ~out_top_channel_i[1];
  assign N142 = out_top_channel_i[2] & out_top_channel_i[0] & N28;
  assign N28 = ~out_top_channel_i[1];
  assign N143 = out_top_channel_i[2] & N29 & out_top_channel_i[1];
  assign N29 = ~out_top_channel_i[0];
  assign N144 = out_top_channel_i[2] & out_top_channel_i[0] & out_top_channel_i[1];
  assign N138 = out_top_channel_i[3] & out_top_channel_i[0];
  assign N145 = N30 & N31 & (N32 & N33);
  assign N30 = ~out_top_channel_i[3];
  assign N31 = ~out_top_channel_i[2];
  assign N32 = ~out_top_channel_i[0];
  assign N33 = ~out_top_channel_i[1];
  assign N146 = out_top_channel_i[3] & N34;
  assign N34 = ~out_top_channel_i[0];
  assign N147 = N35 & N36 & (out_top_channel_i[0] & N37);
  assign N35 = ~out_top_channel_i[3];
  assign N36 = ~out_top_channel_i[2];
  assign N37 = ~out_top_channel_i[1];
  assign N149 = N38 & N39 & out_top_channel_i[1];
  assign N38 = ~out_top_channel_i[2];
  assign N39 = ~out_top_channel_i[0];
  assign N150 = N40 & out_top_channel_i[0] & out_top_channel_i[1];
  assign N40 = ~out_top_channel_i[2];
  assign N151 = out_top_channel_i[2] & N41 & N42;
  assign N41 = ~out_top_channel_i[0];
  assign N42 = ~out_top_channel_i[1];
  assign N152 = out_top_channel_i[2] & out_top_channel_i[0] & N43;
  assign N43 = ~out_top_channel_i[1];
  assign N153 = out_top_channel_i[2] & N44 & out_top_channel_i[1];
  assign N44 = ~out_top_channel_i[0];
  assign N154 = out_top_channel_i[2] & out_top_channel_i[0] & out_top_channel_i[1];
  assign N148 = out_top_channel_i[3] & out_top_channel_i[0];
  assign N155 = N45 & N46 & (N47 & N48);
  assign N45 = ~in_top_channel_i[3];
  assign N46 = ~in_top_channel_i[2];
  assign N47 = ~in_top_channel_i[0];
  assign N48 = ~in_top_channel_i[1];
  assign N156 = in_top_channel_i[3] & N49;
  assign N49 = ~in_top_channel_i[0];
  assign N157 = N50 & N51 & (in_top_channel_i[0] & N52);
  assign N50 = ~in_top_channel_i[3];
  assign N51 = ~in_top_channel_i[2];
  assign N52 = ~in_top_channel_i[1];
  assign N159 = N53 & N54 & in_top_channel_i[1];
  assign N53 = ~in_top_channel_i[2];
  assign N54 = ~in_top_channel_i[0];
  assign N160 = N55 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N55 = ~in_top_channel_i[2];
  assign N161 = in_top_channel_i[2] & N56 & N57;
  assign N56 = ~in_top_channel_i[0];
  assign N57 = ~in_top_channel_i[1];
  assign N162 = in_top_channel_i[2] & in_top_channel_i[0] & N58;
  assign N58 = ~in_top_channel_i[1];
  assign N163 = in_top_channel_i[2] & N59 & in_top_channel_i[1];
  assign N59 = ~in_top_channel_i[0];
  assign N164 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N158 = in_top_channel_i[3] & in_top_channel_i[0];
  assign N165 = N60 & N61 & (N62 & N63);
  assign N60 = ~in_top_channel_i[3];
  assign N61 = ~in_top_channel_i[2];
  assign N62 = ~in_top_channel_i[0];
  assign N63 = ~in_top_channel_i[1];
  assign N166 = in_top_channel_i[3] & N64;
  assign N64 = ~in_top_channel_i[0];
  assign N167 = N65 & N66 & (in_top_channel_i[0] & N67);
  assign N65 = ~in_top_channel_i[3];
  assign N66 = ~in_top_channel_i[2];
  assign N67 = ~in_top_channel_i[1];
  assign N169 = N68 & N69 & in_top_channel_i[1];
  assign N68 = ~in_top_channel_i[2];
  assign N69 = ~in_top_channel_i[0];
  assign N170 = N70 & in_top_channel_i[0] & in_top_channel_i[1];
  assign N70 = ~in_top_channel_i[2];
  assign N171 = in_top_channel_i[2] & N71 & N72;
  assign N71 = ~in_top_channel_i[0];
  assign N72 = ~in_top_channel_i[1];
  assign N172 = in_top_channel_i[2] & in_top_channel_i[0] & N73;
  assign N73 = ~in_top_channel_i[1];
  assign N173 = in_top_channel_i[2] & N74 & in_top_channel_i[1];
  assign N74 = ~in_top_channel_i[0];
  assign N174 = in_top_channel_i[2] & in_top_channel_i[0] & in_top_channel_i[1];
  assign N168 = in_top_channel_i[3] & in_top_channel_i[0];
  assign yumi_o[9] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__9_ : 1'b0;
  assign N75 = N125;
  assign N76 = N127;
  assign N77 = N129;
  assign N78 = N130;
  assign N79 = N131;
  assign N80 = N132;
  assign N81 = N133;
  assign N82 = N134;
  assign N83 = N126;
  assign N84 = N128;
  assign yumi_o[8] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__8_ : 1'b0;
  assign yumi_o[7] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__7_ : 1'b0;
  assign yumi_o[6] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__6_ : 1'b0;
  assign yumi_o[5] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__5_ : 1'b0;
  assign yumi_o[4] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__4_ : 1'b0;
  assign yumi_o[3] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__3_ : 1'b0;
  assign yumi_o[2] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__2_ : 1'b0;
  assign yumi_o[1] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__1_ : 1'b0;
  assign yumi_o[0] = (N75)? 1'b0 : 
                     (N76)? 1'b0 : 
                     (N77)? 1'b0 : 
                     (N78)? 1'b0 : 
                     (N79)? 1'b0 : 
                     (N80)? 1'b0 : 
                     (N81)? 1'b0 : 
                     (N82)? 1'b0 : 
                     (N83)? 1'b0 : 
                     (N84)? yumi_int_o_9__0_ : 1'b0;
  assign valid_o[9] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__9_ : 1'b0;
  assign N85 = N135;
  assign N86 = N137;
  assign N87 = N139;
  assign N88 = N140;
  assign N89 = N141;
  assign N90 = N142;
  assign N91 = N143;
  assign N92 = N144;
  assign N93 = N136;
  assign N94 = N138;
  assign valid_o[8] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__8_ : 1'b0;
  assign valid_o[7] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__7_ : 1'b0;
  assign valid_o[6] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__6_ : 1'b0;
  assign valid_o[5] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__5_ : 1'b0;
  assign valid_o[4] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__4_ : 1'b0;
  assign valid_o[3] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__3_ : 1'b0;
  assign valid_o[2] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__2_ : 1'b0;
  assign valid_o[1] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__1_ : 1'b0;
  assign valid_o[0] = (N85)? 1'b0 : 
                      (N86)? 1'b0 : 
                      (N87)? 1'b0 : 
                      (N88)? 1'b0 : 
                      (N89)? 1'b0 : 
                      (N90)? 1'b0 : 
                      (N91)? 1'b0 : 
                      (N92)? 1'b0 : 
                      (N93)? 1'b0 : 
                      (N94)? valid_int_o_9__0_ : 1'b0;
  assign data_o_flat[1279] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1279_ : 1'b0;
  assign N95 = N145;
  assign N96 = N147;
  assign N97 = N149;
  assign N98 = N150;
  assign N99 = N151;
  assign N100 = N152;
  assign N101 = N153;
  assign N102 = N154;
  assign N103 = N146;
  assign N104 = N148;
  assign data_o_flat[1278] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1278_ : 1'b0;
  assign data_o_flat[1277] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1277_ : 1'b0;
  assign data_o_flat[1276] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1276_ : 1'b0;
  assign data_o_flat[1275] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1275_ : 1'b0;
  assign data_o_flat[1274] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1274_ : 1'b0;
  assign data_o_flat[1273] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1273_ : 1'b0;
  assign data_o_flat[1272] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1272_ : 1'b0;
  assign data_o_flat[1271] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1271_ : 1'b0;
  assign data_o_flat[1270] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1270_ : 1'b0;
  assign data_o_flat[1269] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1269_ : 1'b0;
  assign data_o_flat[1268] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1268_ : 1'b0;
  assign data_o_flat[1267] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1267_ : 1'b0;
  assign data_o_flat[1266] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1266_ : 1'b0;
  assign data_o_flat[1265] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1265_ : 1'b0;
  assign data_o_flat[1264] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1264_ : 1'b0;
  assign data_o_flat[1263] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1263_ : 1'b0;
  assign data_o_flat[1262] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1262_ : 1'b0;
  assign data_o_flat[1261] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1261_ : 1'b0;
  assign data_o_flat[1260] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1260_ : 1'b0;
  assign data_o_flat[1259] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1259_ : 1'b0;
  assign data_o_flat[1258] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1258_ : 1'b0;
  assign data_o_flat[1257] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1257_ : 1'b0;
  assign data_o_flat[1256] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1256_ : 1'b0;
  assign data_o_flat[1255] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1255_ : 1'b0;
  assign data_o_flat[1254] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1254_ : 1'b0;
  assign data_o_flat[1253] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1253_ : 1'b0;
  assign data_o_flat[1252] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1252_ : 1'b0;
  assign data_o_flat[1251] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1251_ : 1'b0;
  assign data_o_flat[1250] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1250_ : 1'b0;
  assign data_o_flat[1249] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1249_ : 1'b0;
  assign data_o_flat[1248] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1248_ : 1'b0;
  assign data_o_flat[1247] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1247_ : 1'b0;
  assign data_o_flat[1246] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1246_ : 1'b0;
  assign data_o_flat[1245] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1245_ : 1'b0;
  assign data_o_flat[1244] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1244_ : 1'b0;
  assign data_o_flat[1243] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1243_ : 1'b0;
  assign data_o_flat[1242] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1242_ : 1'b0;
  assign data_o_flat[1241] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1241_ : 1'b0;
  assign data_o_flat[1240] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1240_ : 1'b0;
  assign data_o_flat[1239] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1239_ : 1'b0;
  assign data_o_flat[1238] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1238_ : 1'b0;
  assign data_o_flat[1237] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1237_ : 1'b0;
  assign data_o_flat[1236] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1236_ : 1'b0;
  assign data_o_flat[1235] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1235_ : 1'b0;
  assign data_o_flat[1234] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1234_ : 1'b0;
  assign data_o_flat[1233] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1233_ : 1'b0;
  assign data_o_flat[1232] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1232_ : 1'b0;
  assign data_o_flat[1231] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1231_ : 1'b0;
  assign data_o_flat[1230] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1230_ : 1'b0;
  assign data_o_flat[1229] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1229_ : 1'b0;
  assign data_o_flat[1228] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1228_ : 1'b0;
  assign data_o_flat[1227] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1227_ : 1'b0;
  assign data_o_flat[1226] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1226_ : 1'b0;
  assign data_o_flat[1225] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1225_ : 1'b0;
  assign data_o_flat[1224] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1224_ : 1'b0;
  assign data_o_flat[1223] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1223_ : 1'b0;
  assign data_o_flat[1222] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1222_ : 1'b0;
  assign data_o_flat[1221] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1221_ : 1'b0;
  assign data_o_flat[1220] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1220_ : 1'b0;
  assign data_o_flat[1219] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1219_ : 1'b0;
  assign data_o_flat[1218] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1218_ : 1'b0;
  assign data_o_flat[1217] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1217_ : 1'b0;
  assign data_o_flat[1216] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1216_ : 1'b0;
  assign data_o_flat[1215] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1215_ : 1'b0;
  assign data_o_flat[1214] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1214_ : 1'b0;
  assign data_o_flat[1213] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1213_ : 1'b0;
  assign data_o_flat[1212] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1212_ : 1'b0;
  assign data_o_flat[1211] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1211_ : 1'b0;
  assign data_o_flat[1210] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1210_ : 1'b0;
  assign data_o_flat[1209] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1209_ : 1'b0;
  assign data_o_flat[1208] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1208_ : 1'b0;
  assign data_o_flat[1207] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1207_ : 1'b0;
  assign data_o_flat[1206] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1206_ : 1'b0;
  assign data_o_flat[1205] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1205_ : 1'b0;
  assign data_o_flat[1204] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1204_ : 1'b0;
  assign data_o_flat[1203] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1203_ : 1'b0;
  assign data_o_flat[1202] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1202_ : 1'b0;
  assign data_o_flat[1201] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1201_ : 1'b0;
  assign data_o_flat[1200] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1200_ : 1'b0;
  assign data_o_flat[1199] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1199_ : 1'b0;
  assign data_o_flat[1198] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1198_ : 1'b0;
  assign data_o_flat[1197] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1197_ : 1'b0;
  assign data_o_flat[1196] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1196_ : 1'b0;
  assign data_o_flat[1195] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1195_ : 1'b0;
  assign data_o_flat[1194] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1194_ : 1'b0;
  assign data_o_flat[1193] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1193_ : 1'b0;
  assign data_o_flat[1192] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1192_ : 1'b0;
  assign data_o_flat[1191] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1191_ : 1'b0;
  assign data_o_flat[1190] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1190_ : 1'b0;
  assign data_o_flat[1189] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1189_ : 1'b0;
  assign data_o_flat[1188] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1188_ : 1'b0;
  assign data_o_flat[1187] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1187_ : 1'b0;
  assign data_o_flat[1186] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1186_ : 1'b0;
  assign data_o_flat[1185] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1185_ : 1'b0;
  assign data_o_flat[1184] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1184_ : 1'b0;
  assign data_o_flat[1183] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1183_ : 1'b0;
  assign data_o_flat[1182] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1182_ : 1'b0;
  assign data_o_flat[1181] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1181_ : 1'b0;
  assign data_o_flat[1180] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1180_ : 1'b0;
  assign data_o_flat[1179] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1179_ : 1'b0;
  assign data_o_flat[1178] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1178_ : 1'b0;
  assign data_o_flat[1177] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1177_ : 1'b0;
  assign data_o_flat[1176] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1176_ : 1'b0;
  assign data_o_flat[1175] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1175_ : 1'b0;
  assign data_o_flat[1174] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1174_ : 1'b0;
  assign data_o_flat[1173] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1173_ : 1'b0;
  assign data_o_flat[1172] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1172_ : 1'b0;
  assign data_o_flat[1171] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1171_ : 1'b0;
  assign data_o_flat[1170] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1170_ : 1'b0;
  assign data_o_flat[1169] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1169_ : 1'b0;
  assign data_o_flat[1168] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1168_ : 1'b0;
  assign data_o_flat[1167] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1167_ : 1'b0;
  assign data_o_flat[1166] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1166_ : 1'b0;
  assign data_o_flat[1165] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1165_ : 1'b0;
  assign data_o_flat[1164] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1164_ : 1'b0;
  assign data_o_flat[1163] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1163_ : 1'b0;
  assign data_o_flat[1162] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1162_ : 1'b0;
  assign data_o_flat[1161] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1161_ : 1'b0;
  assign data_o_flat[1160] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1160_ : 1'b0;
  assign data_o_flat[1159] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1159_ : 1'b0;
  assign data_o_flat[1158] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1158_ : 1'b0;
  assign data_o_flat[1157] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1157_ : 1'b0;
  assign data_o_flat[1156] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1156_ : 1'b0;
  assign data_o_flat[1155] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1155_ : 1'b0;
  assign data_o_flat[1154] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1154_ : 1'b0;
  assign data_o_flat[1153] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1153_ : 1'b0;
  assign data_o_flat[1152] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1152_ : 1'b0;
  assign data_o_flat[1151] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1151_ : 1'b0;
  assign data_o_flat[1150] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1150_ : 1'b0;
  assign data_o_flat[1149] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1149_ : 1'b0;
  assign data_o_flat[1148] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1148_ : 1'b0;
  assign data_o_flat[1147] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1147_ : 1'b0;
  assign data_o_flat[1146] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1146_ : 1'b0;
  assign data_o_flat[1145] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1145_ : 1'b0;
  assign data_o_flat[1144] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1144_ : 1'b0;
  assign data_o_flat[1143] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1143_ : 1'b0;
  assign data_o_flat[1142] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1142_ : 1'b0;
  assign data_o_flat[1141] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1141_ : 1'b0;
  assign data_o_flat[1140] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1140_ : 1'b0;
  assign data_o_flat[1139] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1139_ : 1'b0;
  assign data_o_flat[1138] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1138_ : 1'b0;
  assign data_o_flat[1137] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1137_ : 1'b0;
  assign data_o_flat[1136] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1136_ : 1'b0;
  assign data_o_flat[1135] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1135_ : 1'b0;
  assign data_o_flat[1134] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1134_ : 1'b0;
  assign data_o_flat[1133] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1133_ : 1'b0;
  assign data_o_flat[1132] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1132_ : 1'b0;
  assign data_o_flat[1131] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1131_ : 1'b0;
  assign data_o_flat[1130] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1130_ : 1'b0;
  assign data_o_flat[1129] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1129_ : 1'b0;
  assign data_o_flat[1128] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1128_ : 1'b0;
  assign data_o_flat[1127] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1127_ : 1'b0;
  assign data_o_flat[1126] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1126_ : 1'b0;
  assign data_o_flat[1125] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1125_ : 1'b0;
  assign data_o_flat[1124] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1124_ : 1'b0;
  assign data_o_flat[1123] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1123_ : 1'b0;
  assign data_o_flat[1122] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1122_ : 1'b0;
  assign data_o_flat[1121] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1121_ : 1'b0;
  assign data_o_flat[1120] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1120_ : 1'b0;
  assign data_o_flat[1119] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1119_ : 1'b0;
  assign data_o_flat[1118] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1118_ : 1'b0;
  assign data_o_flat[1117] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1117_ : 1'b0;
  assign data_o_flat[1116] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1116_ : 1'b0;
  assign data_o_flat[1115] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1115_ : 1'b0;
  assign data_o_flat[1114] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1114_ : 1'b0;
  assign data_o_flat[1113] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1113_ : 1'b0;
  assign data_o_flat[1112] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1112_ : 1'b0;
  assign data_o_flat[1111] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1111_ : 1'b0;
  assign data_o_flat[1110] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1110_ : 1'b0;
  assign data_o_flat[1109] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1109_ : 1'b0;
  assign data_o_flat[1108] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1108_ : 1'b0;
  assign data_o_flat[1107] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1107_ : 1'b0;
  assign data_o_flat[1106] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1106_ : 1'b0;
  assign data_o_flat[1105] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1105_ : 1'b0;
  assign data_o_flat[1104] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1104_ : 1'b0;
  assign data_o_flat[1103] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1103_ : 1'b0;
  assign data_o_flat[1102] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1102_ : 1'b0;
  assign data_o_flat[1101] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1101_ : 1'b0;
  assign data_o_flat[1100] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1100_ : 1'b0;
  assign data_o_flat[1099] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1099_ : 1'b0;
  assign data_o_flat[1098] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1098_ : 1'b0;
  assign data_o_flat[1097] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1097_ : 1'b0;
  assign data_o_flat[1096] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1096_ : 1'b0;
  assign data_o_flat[1095] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1095_ : 1'b0;
  assign data_o_flat[1094] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1094_ : 1'b0;
  assign data_o_flat[1093] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1093_ : 1'b0;
  assign data_o_flat[1092] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1092_ : 1'b0;
  assign data_o_flat[1091] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1091_ : 1'b0;
  assign data_o_flat[1090] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1090_ : 1'b0;
  assign data_o_flat[1089] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1089_ : 1'b0;
  assign data_o_flat[1088] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1088_ : 1'b0;
  assign data_o_flat[1087] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1087_ : 1'b0;
  assign data_o_flat[1086] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1086_ : 1'b0;
  assign data_o_flat[1085] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1085_ : 1'b0;
  assign data_o_flat[1084] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1084_ : 1'b0;
  assign data_o_flat[1083] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1083_ : 1'b0;
  assign data_o_flat[1082] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1082_ : 1'b0;
  assign data_o_flat[1081] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1081_ : 1'b0;
  assign data_o_flat[1080] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1080_ : 1'b0;
  assign data_o_flat[1079] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1079_ : 1'b0;
  assign data_o_flat[1078] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1078_ : 1'b0;
  assign data_o_flat[1077] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1077_ : 1'b0;
  assign data_o_flat[1076] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1076_ : 1'b0;
  assign data_o_flat[1075] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1075_ : 1'b0;
  assign data_o_flat[1074] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1074_ : 1'b0;
  assign data_o_flat[1073] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1073_ : 1'b0;
  assign data_o_flat[1072] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1072_ : 1'b0;
  assign data_o_flat[1071] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1071_ : 1'b0;
  assign data_o_flat[1070] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1070_ : 1'b0;
  assign data_o_flat[1069] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1069_ : 1'b0;
  assign data_o_flat[1068] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1068_ : 1'b0;
  assign data_o_flat[1067] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1067_ : 1'b0;
  assign data_o_flat[1066] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1066_ : 1'b0;
  assign data_o_flat[1065] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1065_ : 1'b0;
  assign data_o_flat[1064] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1064_ : 1'b0;
  assign data_o_flat[1063] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1063_ : 1'b0;
  assign data_o_flat[1062] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1062_ : 1'b0;
  assign data_o_flat[1061] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1061_ : 1'b0;
  assign data_o_flat[1060] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1060_ : 1'b0;
  assign data_o_flat[1059] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1059_ : 1'b0;
  assign data_o_flat[1058] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1058_ : 1'b0;
  assign data_o_flat[1057] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1057_ : 1'b0;
  assign data_o_flat[1056] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1056_ : 1'b0;
  assign data_o_flat[1055] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1055_ : 1'b0;
  assign data_o_flat[1054] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1054_ : 1'b0;
  assign data_o_flat[1053] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1053_ : 1'b0;
  assign data_o_flat[1052] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1052_ : 1'b0;
  assign data_o_flat[1051] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1051_ : 1'b0;
  assign data_o_flat[1050] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1050_ : 1'b0;
  assign data_o_flat[1049] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1049_ : 1'b0;
  assign data_o_flat[1048] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1048_ : 1'b0;
  assign data_o_flat[1047] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1047_ : 1'b0;
  assign data_o_flat[1046] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1046_ : 1'b0;
  assign data_o_flat[1045] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1045_ : 1'b0;
  assign data_o_flat[1044] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1044_ : 1'b0;
  assign data_o_flat[1043] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1043_ : 1'b0;
  assign data_o_flat[1042] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1042_ : 1'b0;
  assign data_o_flat[1041] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1041_ : 1'b0;
  assign data_o_flat[1040] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1040_ : 1'b0;
  assign data_o_flat[1039] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1039_ : 1'b0;
  assign data_o_flat[1038] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1038_ : 1'b0;
  assign data_o_flat[1037] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1037_ : 1'b0;
  assign data_o_flat[1036] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1036_ : 1'b0;
  assign data_o_flat[1035] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1035_ : 1'b0;
  assign data_o_flat[1034] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1034_ : 1'b0;
  assign data_o_flat[1033] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1033_ : 1'b0;
  assign data_o_flat[1032] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1032_ : 1'b0;
  assign data_o_flat[1031] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1031_ : 1'b0;
  assign data_o_flat[1030] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1030_ : 1'b0;
  assign data_o_flat[1029] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1029_ : 1'b0;
  assign data_o_flat[1028] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1028_ : 1'b0;
  assign data_o_flat[1027] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1027_ : 1'b0;
  assign data_o_flat[1026] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1026_ : 1'b0;
  assign data_o_flat[1025] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1025_ : 1'b0;
  assign data_o_flat[1024] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1024_ : 1'b0;
  assign data_o_flat[1023] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1023_ : 1'b0;
  assign data_o_flat[1022] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1022_ : 1'b0;
  assign data_o_flat[1021] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1021_ : 1'b0;
  assign data_o_flat[1020] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1020_ : 1'b0;
  assign data_o_flat[1019] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1019_ : 1'b0;
  assign data_o_flat[1018] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1018_ : 1'b0;
  assign data_o_flat[1017] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1017_ : 1'b0;
  assign data_o_flat[1016] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1016_ : 1'b0;
  assign data_o_flat[1015] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1015_ : 1'b0;
  assign data_o_flat[1014] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1014_ : 1'b0;
  assign data_o_flat[1013] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1013_ : 1'b0;
  assign data_o_flat[1012] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1012_ : 1'b0;
  assign data_o_flat[1011] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1011_ : 1'b0;
  assign data_o_flat[1010] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1010_ : 1'b0;
  assign data_o_flat[1009] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1009_ : 1'b0;
  assign data_o_flat[1008] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1008_ : 1'b0;
  assign data_o_flat[1007] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1007_ : 1'b0;
  assign data_o_flat[1006] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1006_ : 1'b0;
  assign data_o_flat[1005] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1005_ : 1'b0;
  assign data_o_flat[1004] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1004_ : 1'b0;
  assign data_o_flat[1003] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1003_ : 1'b0;
  assign data_o_flat[1002] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1002_ : 1'b0;
  assign data_o_flat[1001] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1001_ : 1'b0;
  assign data_o_flat[1000] = (N95)? 1'b0 : 
                             (N96)? 1'b0 : 
                             (N97)? 1'b0 : 
                             (N98)? 1'b0 : 
                             (N99)? 1'b0 : 
                             (N100)? 1'b0 : 
                             (N101)? 1'b0 : 
                             (N102)? 1'b0 : 
                             (N103)? 1'b0 : 
                             (N104)? data_int_o_9__1000_ : 1'b0;
  assign data_o_flat[999] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__999_ : 1'b0;
  assign data_o_flat[998] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__998_ : 1'b0;
  assign data_o_flat[997] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__997_ : 1'b0;
  assign data_o_flat[996] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__996_ : 1'b0;
  assign data_o_flat[995] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__995_ : 1'b0;
  assign data_o_flat[994] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__994_ : 1'b0;
  assign data_o_flat[993] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__993_ : 1'b0;
  assign data_o_flat[992] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__992_ : 1'b0;
  assign data_o_flat[991] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__991_ : 1'b0;
  assign data_o_flat[990] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__990_ : 1'b0;
  assign data_o_flat[989] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__989_ : 1'b0;
  assign data_o_flat[988] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__988_ : 1'b0;
  assign data_o_flat[987] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__987_ : 1'b0;
  assign data_o_flat[986] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__986_ : 1'b0;
  assign data_o_flat[985] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__985_ : 1'b0;
  assign data_o_flat[984] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__984_ : 1'b0;
  assign data_o_flat[983] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__983_ : 1'b0;
  assign data_o_flat[982] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__982_ : 1'b0;
  assign data_o_flat[981] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__981_ : 1'b0;
  assign data_o_flat[980] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__980_ : 1'b0;
  assign data_o_flat[979] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__979_ : 1'b0;
  assign data_o_flat[978] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__978_ : 1'b0;
  assign data_o_flat[977] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__977_ : 1'b0;
  assign data_o_flat[976] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__976_ : 1'b0;
  assign data_o_flat[975] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__975_ : 1'b0;
  assign data_o_flat[974] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__974_ : 1'b0;
  assign data_o_flat[973] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__973_ : 1'b0;
  assign data_o_flat[972] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__972_ : 1'b0;
  assign data_o_flat[971] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__971_ : 1'b0;
  assign data_o_flat[970] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__970_ : 1'b0;
  assign data_o_flat[969] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__969_ : 1'b0;
  assign data_o_flat[968] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__968_ : 1'b0;
  assign data_o_flat[967] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__967_ : 1'b0;
  assign data_o_flat[966] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__966_ : 1'b0;
  assign data_o_flat[965] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__965_ : 1'b0;
  assign data_o_flat[964] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__964_ : 1'b0;
  assign data_o_flat[963] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__963_ : 1'b0;
  assign data_o_flat[962] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__962_ : 1'b0;
  assign data_o_flat[961] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__961_ : 1'b0;
  assign data_o_flat[960] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__960_ : 1'b0;
  assign data_o_flat[959] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__959_ : 1'b0;
  assign data_o_flat[958] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__958_ : 1'b0;
  assign data_o_flat[957] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__957_ : 1'b0;
  assign data_o_flat[956] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__956_ : 1'b0;
  assign data_o_flat[955] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__955_ : 1'b0;
  assign data_o_flat[954] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__954_ : 1'b0;
  assign data_o_flat[953] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__953_ : 1'b0;
  assign data_o_flat[952] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__952_ : 1'b0;
  assign data_o_flat[951] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__951_ : 1'b0;
  assign data_o_flat[950] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__950_ : 1'b0;
  assign data_o_flat[949] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__949_ : 1'b0;
  assign data_o_flat[948] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__948_ : 1'b0;
  assign data_o_flat[947] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__947_ : 1'b0;
  assign data_o_flat[946] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__946_ : 1'b0;
  assign data_o_flat[945] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__945_ : 1'b0;
  assign data_o_flat[944] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__944_ : 1'b0;
  assign data_o_flat[943] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__943_ : 1'b0;
  assign data_o_flat[942] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__942_ : 1'b0;
  assign data_o_flat[941] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__941_ : 1'b0;
  assign data_o_flat[940] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__940_ : 1'b0;
  assign data_o_flat[939] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__939_ : 1'b0;
  assign data_o_flat[938] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__938_ : 1'b0;
  assign data_o_flat[937] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__937_ : 1'b0;
  assign data_o_flat[936] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__936_ : 1'b0;
  assign data_o_flat[935] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__935_ : 1'b0;
  assign data_o_flat[934] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__934_ : 1'b0;
  assign data_o_flat[933] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__933_ : 1'b0;
  assign data_o_flat[932] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__932_ : 1'b0;
  assign data_o_flat[931] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__931_ : 1'b0;
  assign data_o_flat[930] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__930_ : 1'b0;
  assign data_o_flat[929] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__929_ : 1'b0;
  assign data_o_flat[928] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__928_ : 1'b0;
  assign data_o_flat[927] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__927_ : 1'b0;
  assign data_o_flat[926] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__926_ : 1'b0;
  assign data_o_flat[925] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__925_ : 1'b0;
  assign data_o_flat[924] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__924_ : 1'b0;
  assign data_o_flat[923] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__923_ : 1'b0;
  assign data_o_flat[922] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__922_ : 1'b0;
  assign data_o_flat[921] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__921_ : 1'b0;
  assign data_o_flat[920] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__920_ : 1'b0;
  assign data_o_flat[919] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__919_ : 1'b0;
  assign data_o_flat[918] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__918_ : 1'b0;
  assign data_o_flat[917] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__917_ : 1'b0;
  assign data_o_flat[916] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__916_ : 1'b0;
  assign data_o_flat[915] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__915_ : 1'b0;
  assign data_o_flat[914] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__914_ : 1'b0;
  assign data_o_flat[913] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__913_ : 1'b0;
  assign data_o_flat[912] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__912_ : 1'b0;
  assign data_o_flat[911] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__911_ : 1'b0;
  assign data_o_flat[910] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__910_ : 1'b0;
  assign data_o_flat[909] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__909_ : 1'b0;
  assign data_o_flat[908] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__908_ : 1'b0;
  assign data_o_flat[907] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__907_ : 1'b0;
  assign data_o_flat[906] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__906_ : 1'b0;
  assign data_o_flat[905] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__905_ : 1'b0;
  assign data_o_flat[904] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__904_ : 1'b0;
  assign data_o_flat[903] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__903_ : 1'b0;
  assign data_o_flat[902] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__902_ : 1'b0;
  assign data_o_flat[901] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__901_ : 1'b0;
  assign data_o_flat[900] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__900_ : 1'b0;
  assign data_o_flat[899] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__899_ : 1'b0;
  assign data_o_flat[898] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__898_ : 1'b0;
  assign data_o_flat[897] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__897_ : 1'b0;
  assign data_o_flat[896] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__896_ : 1'b0;
  assign data_o_flat[895] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__895_ : 1'b0;
  assign data_o_flat[894] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__894_ : 1'b0;
  assign data_o_flat[893] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__893_ : 1'b0;
  assign data_o_flat[892] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__892_ : 1'b0;
  assign data_o_flat[891] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__891_ : 1'b0;
  assign data_o_flat[890] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__890_ : 1'b0;
  assign data_o_flat[889] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__889_ : 1'b0;
  assign data_o_flat[888] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__888_ : 1'b0;
  assign data_o_flat[887] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__887_ : 1'b0;
  assign data_o_flat[886] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__886_ : 1'b0;
  assign data_o_flat[885] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__885_ : 1'b0;
  assign data_o_flat[884] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__884_ : 1'b0;
  assign data_o_flat[883] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__883_ : 1'b0;
  assign data_o_flat[882] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__882_ : 1'b0;
  assign data_o_flat[881] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__881_ : 1'b0;
  assign data_o_flat[880] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__880_ : 1'b0;
  assign data_o_flat[879] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__879_ : 1'b0;
  assign data_o_flat[878] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__878_ : 1'b0;
  assign data_o_flat[877] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__877_ : 1'b0;
  assign data_o_flat[876] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__876_ : 1'b0;
  assign data_o_flat[875] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__875_ : 1'b0;
  assign data_o_flat[874] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__874_ : 1'b0;
  assign data_o_flat[873] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__873_ : 1'b0;
  assign data_o_flat[872] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__872_ : 1'b0;
  assign data_o_flat[871] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__871_ : 1'b0;
  assign data_o_flat[870] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__870_ : 1'b0;
  assign data_o_flat[869] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__869_ : 1'b0;
  assign data_o_flat[868] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__868_ : 1'b0;
  assign data_o_flat[867] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__867_ : 1'b0;
  assign data_o_flat[866] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__866_ : 1'b0;
  assign data_o_flat[865] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__865_ : 1'b0;
  assign data_o_flat[864] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__864_ : 1'b0;
  assign data_o_flat[863] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__863_ : 1'b0;
  assign data_o_flat[862] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__862_ : 1'b0;
  assign data_o_flat[861] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__861_ : 1'b0;
  assign data_o_flat[860] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__860_ : 1'b0;
  assign data_o_flat[859] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__859_ : 1'b0;
  assign data_o_flat[858] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__858_ : 1'b0;
  assign data_o_flat[857] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__857_ : 1'b0;
  assign data_o_flat[856] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__856_ : 1'b0;
  assign data_o_flat[855] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__855_ : 1'b0;
  assign data_o_flat[854] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__854_ : 1'b0;
  assign data_o_flat[853] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__853_ : 1'b0;
  assign data_o_flat[852] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__852_ : 1'b0;
  assign data_o_flat[851] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__851_ : 1'b0;
  assign data_o_flat[850] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__850_ : 1'b0;
  assign data_o_flat[849] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__849_ : 1'b0;
  assign data_o_flat[848] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__848_ : 1'b0;
  assign data_o_flat[847] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__847_ : 1'b0;
  assign data_o_flat[846] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__846_ : 1'b0;
  assign data_o_flat[845] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__845_ : 1'b0;
  assign data_o_flat[844] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__844_ : 1'b0;
  assign data_o_flat[843] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__843_ : 1'b0;
  assign data_o_flat[842] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__842_ : 1'b0;
  assign data_o_flat[841] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__841_ : 1'b0;
  assign data_o_flat[840] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__840_ : 1'b0;
  assign data_o_flat[839] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__839_ : 1'b0;
  assign data_o_flat[838] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__838_ : 1'b0;
  assign data_o_flat[837] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__837_ : 1'b0;
  assign data_o_flat[836] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__836_ : 1'b0;
  assign data_o_flat[835] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__835_ : 1'b0;
  assign data_o_flat[834] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__834_ : 1'b0;
  assign data_o_flat[833] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__833_ : 1'b0;
  assign data_o_flat[832] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__832_ : 1'b0;
  assign data_o_flat[831] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__831_ : 1'b0;
  assign data_o_flat[830] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__830_ : 1'b0;
  assign data_o_flat[829] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__829_ : 1'b0;
  assign data_o_flat[828] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__828_ : 1'b0;
  assign data_o_flat[827] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__827_ : 1'b0;
  assign data_o_flat[826] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__826_ : 1'b0;
  assign data_o_flat[825] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__825_ : 1'b0;
  assign data_o_flat[824] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__824_ : 1'b0;
  assign data_o_flat[823] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__823_ : 1'b0;
  assign data_o_flat[822] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__822_ : 1'b0;
  assign data_o_flat[821] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__821_ : 1'b0;
  assign data_o_flat[820] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__820_ : 1'b0;
  assign data_o_flat[819] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__819_ : 1'b0;
  assign data_o_flat[818] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__818_ : 1'b0;
  assign data_o_flat[817] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__817_ : 1'b0;
  assign data_o_flat[816] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__816_ : 1'b0;
  assign data_o_flat[815] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__815_ : 1'b0;
  assign data_o_flat[814] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__814_ : 1'b0;
  assign data_o_flat[813] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__813_ : 1'b0;
  assign data_o_flat[812] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__812_ : 1'b0;
  assign data_o_flat[811] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__811_ : 1'b0;
  assign data_o_flat[810] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__810_ : 1'b0;
  assign data_o_flat[809] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__809_ : 1'b0;
  assign data_o_flat[808] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__808_ : 1'b0;
  assign data_o_flat[807] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__807_ : 1'b0;
  assign data_o_flat[806] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__806_ : 1'b0;
  assign data_o_flat[805] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__805_ : 1'b0;
  assign data_o_flat[804] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__804_ : 1'b0;
  assign data_o_flat[803] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__803_ : 1'b0;
  assign data_o_flat[802] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__802_ : 1'b0;
  assign data_o_flat[801] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__801_ : 1'b0;
  assign data_o_flat[800] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__800_ : 1'b0;
  assign data_o_flat[799] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__799_ : 1'b0;
  assign data_o_flat[798] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__798_ : 1'b0;
  assign data_o_flat[797] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__797_ : 1'b0;
  assign data_o_flat[796] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__796_ : 1'b0;
  assign data_o_flat[795] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__795_ : 1'b0;
  assign data_o_flat[794] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__794_ : 1'b0;
  assign data_o_flat[793] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__793_ : 1'b0;
  assign data_o_flat[792] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__792_ : 1'b0;
  assign data_o_flat[791] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__791_ : 1'b0;
  assign data_o_flat[790] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__790_ : 1'b0;
  assign data_o_flat[789] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__789_ : 1'b0;
  assign data_o_flat[788] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__788_ : 1'b0;
  assign data_o_flat[787] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__787_ : 1'b0;
  assign data_o_flat[786] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__786_ : 1'b0;
  assign data_o_flat[785] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__785_ : 1'b0;
  assign data_o_flat[784] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__784_ : 1'b0;
  assign data_o_flat[783] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__783_ : 1'b0;
  assign data_o_flat[782] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__782_ : 1'b0;
  assign data_o_flat[781] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__781_ : 1'b0;
  assign data_o_flat[780] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__780_ : 1'b0;
  assign data_o_flat[779] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__779_ : 1'b0;
  assign data_o_flat[778] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__778_ : 1'b0;
  assign data_o_flat[777] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__777_ : 1'b0;
  assign data_o_flat[776] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__776_ : 1'b0;
  assign data_o_flat[775] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__775_ : 1'b0;
  assign data_o_flat[774] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__774_ : 1'b0;
  assign data_o_flat[773] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__773_ : 1'b0;
  assign data_o_flat[772] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__772_ : 1'b0;
  assign data_o_flat[771] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__771_ : 1'b0;
  assign data_o_flat[770] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__770_ : 1'b0;
  assign data_o_flat[769] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__769_ : 1'b0;
  assign data_o_flat[768] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__768_ : 1'b0;
  assign data_o_flat[767] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__767_ : 1'b0;
  assign data_o_flat[766] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__766_ : 1'b0;
  assign data_o_flat[765] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__765_ : 1'b0;
  assign data_o_flat[764] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__764_ : 1'b0;
  assign data_o_flat[763] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__763_ : 1'b0;
  assign data_o_flat[762] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__762_ : 1'b0;
  assign data_o_flat[761] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__761_ : 1'b0;
  assign data_o_flat[760] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__760_ : 1'b0;
  assign data_o_flat[759] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__759_ : 1'b0;
  assign data_o_flat[758] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__758_ : 1'b0;
  assign data_o_flat[757] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__757_ : 1'b0;
  assign data_o_flat[756] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__756_ : 1'b0;
  assign data_o_flat[755] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__755_ : 1'b0;
  assign data_o_flat[754] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__754_ : 1'b0;
  assign data_o_flat[753] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__753_ : 1'b0;
  assign data_o_flat[752] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__752_ : 1'b0;
  assign data_o_flat[751] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__751_ : 1'b0;
  assign data_o_flat[750] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__750_ : 1'b0;
  assign data_o_flat[749] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__749_ : 1'b0;
  assign data_o_flat[748] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__748_ : 1'b0;
  assign data_o_flat[747] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__747_ : 1'b0;
  assign data_o_flat[746] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__746_ : 1'b0;
  assign data_o_flat[745] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__745_ : 1'b0;
  assign data_o_flat[744] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__744_ : 1'b0;
  assign data_o_flat[743] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__743_ : 1'b0;
  assign data_o_flat[742] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__742_ : 1'b0;
  assign data_o_flat[741] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__741_ : 1'b0;
  assign data_o_flat[740] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__740_ : 1'b0;
  assign data_o_flat[739] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__739_ : 1'b0;
  assign data_o_flat[738] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__738_ : 1'b0;
  assign data_o_flat[737] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__737_ : 1'b0;
  assign data_o_flat[736] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__736_ : 1'b0;
  assign data_o_flat[735] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__735_ : 1'b0;
  assign data_o_flat[734] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__734_ : 1'b0;
  assign data_o_flat[733] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__733_ : 1'b0;
  assign data_o_flat[732] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__732_ : 1'b0;
  assign data_o_flat[731] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__731_ : 1'b0;
  assign data_o_flat[730] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__730_ : 1'b0;
  assign data_o_flat[729] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__729_ : 1'b0;
  assign data_o_flat[728] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__728_ : 1'b0;
  assign data_o_flat[727] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__727_ : 1'b0;
  assign data_o_flat[726] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__726_ : 1'b0;
  assign data_o_flat[725] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__725_ : 1'b0;
  assign data_o_flat[724] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__724_ : 1'b0;
  assign data_o_flat[723] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__723_ : 1'b0;
  assign data_o_flat[722] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__722_ : 1'b0;
  assign data_o_flat[721] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__721_ : 1'b0;
  assign data_o_flat[720] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__720_ : 1'b0;
  assign data_o_flat[719] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__719_ : 1'b0;
  assign data_o_flat[718] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__718_ : 1'b0;
  assign data_o_flat[717] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__717_ : 1'b0;
  assign data_o_flat[716] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__716_ : 1'b0;
  assign data_o_flat[715] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__715_ : 1'b0;
  assign data_o_flat[714] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__714_ : 1'b0;
  assign data_o_flat[713] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__713_ : 1'b0;
  assign data_o_flat[712] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__712_ : 1'b0;
  assign data_o_flat[711] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__711_ : 1'b0;
  assign data_o_flat[710] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__710_ : 1'b0;
  assign data_o_flat[709] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__709_ : 1'b0;
  assign data_o_flat[708] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__708_ : 1'b0;
  assign data_o_flat[707] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__707_ : 1'b0;
  assign data_o_flat[706] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__706_ : 1'b0;
  assign data_o_flat[705] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__705_ : 1'b0;
  assign data_o_flat[704] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__704_ : 1'b0;
  assign data_o_flat[703] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__703_ : 1'b0;
  assign data_o_flat[702] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__702_ : 1'b0;
  assign data_o_flat[701] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__701_ : 1'b0;
  assign data_o_flat[700] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__700_ : 1'b0;
  assign data_o_flat[699] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__699_ : 1'b0;
  assign data_o_flat[698] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__698_ : 1'b0;
  assign data_o_flat[697] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__697_ : 1'b0;
  assign data_o_flat[696] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__696_ : 1'b0;
  assign data_o_flat[695] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__695_ : 1'b0;
  assign data_o_flat[694] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__694_ : 1'b0;
  assign data_o_flat[693] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__693_ : 1'b0;
  assign data_o_flat[692] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__692_ : 1'b0;
  assign data_o_flat[691] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__691_ : 1'b0;
  assign data_o_flat[690] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__690_ : 1'b0;
  assign data_o_flat[689] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__689_ : 1'b0;
  assign data_o_flat[688] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__688_ : 1'b0;
  assign data_o_flat[687] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__687_ : 1'b0;
  assign data_o_flat[686] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__686_ : 1'b0;
  assign data_o_flat[685] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__685_ : 1'b0;
  assign data_o_flat[684] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__684_ : 1'b0;
  assign data_o_flat[683] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__683_ : 1'b0;
  assign data_o_flat[682] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__682_ : 1'b0;
  assign data_o_flat[681] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__681_ : 1'b0;
  assign data_o_flat[680] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__680_ : 1'b0;
  assign data_o_flat[679] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__679_ : 1'b0;
  assign data_o_flat[678] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__678_ : 1'b0;
  assign data_o_flat[677] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__677_ : 1'b0;
  assign data_o_flat[676] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__676_ : 1'b0;
  assign data_o_flat[675] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__675_ : 1'b0;
  assign data_o_flat[674] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__674_ : 1'b0;
  assign data_o_flat[673] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__673_ : 1'b0;
  assign data_o_flat[672] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__672_ : 1'b0;
  assign data_o_flat[671] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__671_ : 1'b0;
  assign data_o_flat[670] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__670_ : 1'b0;
  assign data_o_flat[669] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__669_ : 1'b0;
  assign data_o_flat[668] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__668_ : 1'b0;
  assign data_o_flat[667] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__667_ : 1'b0;
  assign data_o_flat[666] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__666_ : 1'b0;
  assign data_o_flat[665] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__665_ : 1'b0;
  assign data_o_flat[664] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__664_ : 1'b0;
  assign data_o_flat[663] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__663_ : 1'b0;
  assign data_o_flat[662] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__662_ : 1'b0;
  assign data_o_flat[661] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__661_ : 1'b0;
  assign data_o_flat[660] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__660_ : 1'b0;
  assign data_o_flat[659] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__659_ : 1'b0;
  assign data_o_flat[658] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__658_ : 1'b0;
  assign data_o_flat[657] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__657_ : 1'b0;
  assign data_o_flat[656] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__656_ : 1'b0;
  assign data_o_flat[655] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__655_ : 1'b0;
  assign data_o_flat[654] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__654_ : 1'b0;
  assign data_o_flat[653] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__653_ : 1'b0;
  assign data_o_flat[652] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__652_ : 1'b0;
  assign data_o_flat[651] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__651_ : 1'b0;
  assign data_o_flat[650] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__650_ : 1'b0;
  assign data_o_flat[649] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__649_ : 1'b0;
  assign data_o_flat[648] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__648_ : 1'b0;
  assign data_o_flat[647] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__647_ : 1'b0;
  assign data_o_flat[646] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__646_ : 1'b0;
  assign data_o_flat[645] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__645_ : 1'b0;
  assign data_o_flat[644] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__644_ : 1'b0;
  assign data_o_flat[643] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__643_ : 1'b0;
  assign data_o_flat[642] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__642_ : 1'b0;
  assign data_o_flat[641] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__641_ : 1'b0;
  assign data_o_flat[640] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__640_ : 1'b0;
  assign data_o_flat[639] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__639_ : 1'b0;
  assign data_o_flat[638] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__638_ : 1'b0;
  assign data_o_flat[637] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__637_ : 1'b0;
  assign data_o_flat[636] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__636_ : 1'b0;
  assign data_o_flat[635] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__635_ : 1'b0;
  assign data_o_flat[634] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__634_ : 1'b0;
  assign data_o_flat[633] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__633_ : 1'b0;
  assign data_o_flat[632] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__632_ : 1'b0;
  assign data_o_flat[631] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__631_ : 1'b0;
  assign data_o_flat[630] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__630_ : 1'b0;
  assign data_o_flat[629] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__629_ : 1'b0;
  assign data_o_flat[628] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__628_ : 1'b0;
  assign data_o_flat[627] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__627_ : 1'b0;
  assign data_o_flat[626] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__626_ : 1'b0;
  assign data_o_flat[625] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__625_ : 1'b0;
  assign data_o_flat[624] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__624_ : 1'b0;
  assign data_o_flat[623] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__623_ : 1'b0;
  assign data_o_flat[622] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__622_ : 1'b0;
  assign data_o_flat[621] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__621_ : 1'b0;
  assign data_o_flat[620] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__620_ : 1'b0;
  assign data_o_flat[619] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__619_ : 1'b0;
  assign data_o_flat[618] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__618_ : 1'b0;
  assign data_o_flat[617] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__617_ : 1'b0;
  assign data_o_flat[616] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__616_ : 1'b0;
  assign data_o_flat[615] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__615_ : 1'b0;
  assign data_o_flat[614] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__614_ : 1'b0;
  assign data_o_flat[613] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__613_ : 1'b0;
  assign data_o_flat[612] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__612_ : 1'b0;
  assign data_o_flat[611] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__611_ : 1'b0;
  assign data_o_flat[610] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__610_ : 1'b0;
  assign data_o_flat[609] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__609_ : 1'b0;
  assign data_o_flat[608] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__608_ : 1'b0;
  assign data_o_flat[607] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__607_ : 1'b0;
  assign data_o_flat[606] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__606_ : 1'b0;
  assign data_o_flat[605] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__605_ : 1'b0;
  assign data_o_flat[604] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__604_ : 1'b0;
  assign data_o_flat[603] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__603_ : 1'b0;
  assign data_o_flat[602] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__602_ : 1'b0;
  assign data_o_flat[601] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__601_ : 1'b0;
  assign data_o_flat[600] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__600_ : 1'b0;
  assign data_o_flat[599] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__599_ : 1'b0;
  assign data_o_flat[598] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__598_ : 1'b0;
  assign data_o_flat[597] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__597_ : 1'b0;
  assign data_o_flat[596] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__596_ : 1'b0;
  assign data_o_flat[595] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__595_ : 1'b0;
  assign data_o_flat[594] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__594_ : 1'b0;
  assign data_o_flat[593] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__593_ : 1'b0;
  assign data_o_flat[592] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__592_ : 1'b0;
  assign data_o_flat[591] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__591_ : 1'b0;
  assign data_o_flat[590] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__590_ : 1'b0;
  assign data_o_flat[589] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__589_ : 1'b0;
  assign data_o_flat[588] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__588_ : 1'b0;
  assign data_o_flat[587] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__587_ : 1'b0;
  assign data_o_flat[586] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__586_ : 1'b0;
  assign data_o_flat[585] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__585_ : 1'b0;
  assign data_o_flat[584] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__584_ : 1'b0;
  assign data_o_flat[583] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__583_ : 1'b0;
  assign data_o_flat[582] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__582_ : 1'b0;
  assign data_o_flat[581] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__581_ : 1'b0;
  assign data_o_flat[580] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__580_ : 1'b0;
  assign data_o_flat[579] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__579_ : 1'b0;
  assign data_o_flat[578] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__578_ : 1'b0;
  assign data_o_flat[577] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__577_ : 1'b0;
  assign data_o_flat[576] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__576_ : 1'b0;
  assign data_o_flat[575] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__575_ : 1'b0;
  assign data_o_flat[574] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__574_ : 1'b0;
  assign data_o_flat[573] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__573_ : 1'b0;
  assign data_o_flat[572] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__572_ : 1'b0;
  assign data_o_flat[571] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__571_ : 1'b0;
  assign data_o_flat[570] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__570_ : 1'b0;
  assign data_o_flat[569] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__569_ : 1'b0;
  assign data_o_flat[568] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__568_ : 1'b0;
  assign data_o_flat[567] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__567_ : 1'b0;
  assign data_o_flat[566] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__566_ : 1'b0;
  assign data_o_flat[565] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__565_ : 1'b0;
  assign data_o_flat[564] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__564_ : 1'b0;
  assign data_o_flat[563] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__563_ : 1'b0;
  assign data_o_flat[562] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__562_ : 1'b0;
  assign data_o_flat[561] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__561_ : 1'b0;
  assign data_o_flat[560] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__560_ : 1'b0;
  assign data_o_flat[559] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__559_ : 1'b0;
  assign data_o_flat[558] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__558_ : 1'b0;
  assign data_o_flat[557] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__557_ : 1'b0;
  assign data_o_flat[556] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__556_ : 1'b0;
  assign data_o_flat[555] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__555_ : 1'b0;
  assign data_o_flat[554] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__554_ : 1'b0;
  assign data_o_flat[553] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__553_ : 1'b0;
  assign data_o_flat[552] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__552_ : 1'b0;
  assign data_o_flat[551] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__551_ : 1'b0;
  assign data_o_flat[550] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__550_ : 1'b0;
  assign data_o_flat[549] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__549_ : 1'b0;
  assign data_o_flat[548] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__548_ : 1'b0;
  assign data_o_flat[547] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__547_ : 1'b0;
  assign data_o_flat[546] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__546_ : 1'b0;
  assign data_o_flat[545] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__545_ : 1'b0;
  assign data_o_flat[544] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__544_ : 1'b0;
  assign data_o_flat[543] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__543_ : 1'b0;
  assign data_o_flat[542] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__542_ : 1'b0;
  assign data_o_flat[541] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__541_ : 1'b0;
  assign data_o_flat[540] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__540_ : 1'b0;
  assign data_o_flat[539] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__539_ : 1'b0;
  assign data_o_flat[538] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__538_ : 1'b0;
  assign data_o_flat[537] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__537_ : 1'b0;
  assign data_o_flat[536] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__536_ : 1'b0;
  assign data_o_flat[535] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__535_ : 1'b0;
  assign data_o_flat[534] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__534_ : 1'b0;
  assign data_o_flat[533] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__533_ : 1'b0;
  assign data_o_flat[532] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__532_ : 1'b0;
  assign data_o_flat[531] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__531_ : 1'b0;
  assign data_o_flat[530] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__530_ : 1'b0;
  assign data_o_flat[529] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__529_ : 1'b0;
  assign data_o_flat[528] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__528_ : 1'b0;
  assign data_o_flat[527] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__527_ : 1'b0;
  assign data_o_flat[526] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__526_ : 1'b0;
  assign data_o_flat[525] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__525_ : 1'b0;
  assign data_o_flat[524] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__524_ : 1'b0;
  assign data_o_flat[523] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__523_ : 1'b0;
  assign data_o_flat[522] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__522_ : 1'b0;
  assign data_o_flat[521] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__521_ : 1'b0;
  assign data_o_flat[520] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__520_ : 1'b0;
  assign data_o_flat[519] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__519_ : 1'b0;
  assign data_o_flat[518] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__518_ : 1'b0;
  assign data_o_flat[517] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__517_ : 1'b0;
  assign data_o_flat[516] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__516_ : 1'b0;
  assign data_o_flat[515] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__515_ : 1'b0;
  assign data_o_flat[514] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__514_ : 1'b0;
  assign data_o_flat[513] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__513_ : 1'b0;
  assign data_o_flat[512] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__512_ : 1'b0;
  assign data_o_flat[511] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__511_ : 1'b0;
  assign data_o_flat[510] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__510_ : 1'b0;
  assign data_o_flat[509] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__509_ : 1'b0;
  assign data_o_flat[508] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__508_ : 1'b0;
  assign data_o_flat[507] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__507_ : 1'b0;
  assign data_o_flat[506] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__506_ : 1'b0;
  assign data_o_flat[505] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__505_ : 1'b0;
  assign data_o_flat[504] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__504_ : 1'b0;
  assign data_o_flat[503] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__503_ : 1'b0;
  assign data_o_flat[502] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__502_ : 1'b0;
  assign data_o_flat[501] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__501_ : 1'b0;
  assign data_o_flat[500] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__500_ : 1'b0;
  assign data_o_flat[499] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__499_ : 1'b0;
  assign data_o_flat[498] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__498_ : 1'b0;
  assign data_o_flat[497] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__497_ : 1'b0;
  assign data_o_flat[496] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__496_ : 1'b0;
  assign data_o_flat[495] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__495_ : 1'b0;
  assign data_o_flat[494] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__494_ : 1'b0;
  assign data_o_flat[493] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__493_ : 1'b0;
  assign data_o_flat[492] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__492_ : 1'b0;
  assign data_o_flat[491] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__491_ : 1'b0;
  assign data_o_flat[490] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__490_ : 1'b0;
  assign data_o_flat[489] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__489_ : 1'b0;
  assign data_o_flat[488] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__488_ : 1'b0;
  assign data_o_flat[487] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__487_ : 1'b0;
  assign data_o_flat[486] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__486_ : 1'b0;
  assign data_o_flat[485] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__485_ : 1'b0;
  assign data_o_flat[484] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__484_ : 1'b0;
  assign data_o_flat[483] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__483_ : 1'b0;
  assign data_o_flat[482] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__482_ : 1'b0;
  assign data_o_flat[481] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__481_ : 1'b0;
  assign data_o_flat[480] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__480_ : 1'b0;
  assign data_o_flat[479] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__479_ : 1'b0;
  assign data_o_flat[478] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__478_ : 1'b0;
  assign data_o_flat[477] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__477_ : 1'b0;
  assign data_o_flat[476] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__476_ : 1'b0;
  assign data_o_flat[475] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__475_ : 1'b0;
  assign data_o_flat[474] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__474_ : 1'b0;
  assign data_o_flat[473] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__473_ : 1'b0;
  assign data_o_flat[472] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__472_ : 1'b0;
  assign data_o_flat[471] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__471_ : 1'b0;
  assign data_o_flat[470] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__470_ : 1'b0;
  assign data_o_flat[469] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__469_ : 1'b0;
  assign data_o_flat[468] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__468_ : 1'b0;
  assign data_o_flat[467] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__467_ : 1'b0;
  assign data_o_flat[466] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__466_ : 1'b0;
  assign data_o_flat[465] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__465_ : 1'b0;
  assign data_o_flat[464] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__464_ : 1'b0;
  assign data_o_flat[463] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__463_ : 1'b0;
  assign data_o_flat[462] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__462_ : 1'b0;
  assign data_o_flat[461] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__461_ : 1'b0;
  assign data_o_flat[460] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__460_ : 1'b0;
  assign data_o_flat[459] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__459_ : 1'b0;
  assign data_o_flat[458] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__458_ : 1'b0;
  assign data_o_flat[457] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__457_ : 1'b0;
  assign data_o_flat[456] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__456_ : 1'b0;
  assign data_o_flat[455] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__455_ : 1'b0;
  assign data_o_flat[454] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__454_ : 1'b0;
  assign data_o_flat[453] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__453_ : 1'b0;
  assign data_o_flat[452] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__452_ : 1'b0;
  assign data_o_flat[451] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__451_ : 1'b0;
  assign data_o_flat[450] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__450_ : 1'b0;
  assign data_o_flat[449] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__449_ : 1'b0;
  assign data_o_flat[448] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__448_ : 1'b0;
  assign data_o_flat[447] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__447_ : 1'b0;
  assign data_o_flat[446] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__446_ : 1'b0;
  assign data_o_flat[445] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__445_ : 1'b0;
  assign data_o_flat[444] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__444_ : 1'b0;
  assign data_o_flat[443] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__443_ : 1'b0;
  assign data_o_flat[442] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__442_ : 1'b0;
  assign data_o_flat[441] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__441_ : 1'b0;
  assign data_o_flat[440] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__440_ : 1'b0;
  assign data_o_flat[439] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__439_ : 1'b0;
  assign data_o_flat[438] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__438_ : 1'b0;
  assign data_o_flat[437] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__437_ : 1'b0;
  assign data_o_flat[436] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__436_ : 1'b0;
  assign data_o_flat[435] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__435_ : 1'b0;
  assign data_o_flat[434] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__434_ : 1'b0;
  assign data_o_flat[433] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__433_ : 1'b0;
  assign data_o_flat[432] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__432_ : 1'b0;
  assign data_o_flat[431] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__431_ : 1'b0;
  assign data_o_flat[430] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__430_ : 1'b0;
  assign data_o_flat[429] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__429_ : 1'b0;
  assign data_o_flat[428] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__428_ : 1'b0;
  assign data_o_flat[427] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__427_ : 1'b0;
  assign data_o_flat[426] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__426_ : 1'b0;
  assign data_o_flat[425] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__425_ : 1'b0;
  assign data_o_flat[424] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__424_ : 1'b0;
  assign data_o_flat[423] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__423_ : 1'b0;
  assign data_o_flat[422] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__422_ : 1'b0;
  assign data_o_flat[421] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__421_ : 1'b0;
  assign data_o_flat[420] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__420_ : 1'b0;
  assign data_o_flat[419] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__419_ : 1'b0;
  assign data_o_flat[418] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__418_ : 1'b0;
  assign data_o_flat[417] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__417_ : 1'b0;
  assign data_o_flat[416] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__416_ : 1'b0;
  assign data_o_flat[415] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__415_ : 1'b0;
  assign data_o_flat[414] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__414_ : 1'b0;
  assign data_o_flat[413] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__413_ : 1'b0;
  assign data_o_flat[412] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__412_ : 1'b0;
  assign data_o_flat[411] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__411_ : 1'b0;
  assign data_o_flat[410] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__410_ : 1'b0;
  assign data_o_flat[409] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__409_ : 1'b0;
  assign data_o_flat[408] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__408_ : 1'b0;
  assign data_o_flat[407] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__407_ : 1'b0;
  assign data_o_flat[406] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__406_ : 1'b0;
  assign data_o_flat[405] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__405_ : 1'b0;
  assign data_o_flat[404] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__404_ : 1'b0;
  assign data_o_flat[403] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__403_ : 1'b0;
  assign data_o_flat[402] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__402_ : 1'b0;
  assign data_o_flat[401] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__401_ : 1'b0;
  assign data_o_flat[400] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__400_ : 1'b0;
  assign data_o_flat[399] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__399_ : 1'b0;
  assign data_o_flat[398] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__398_ : 1'b0;
  assign data_o_flat[397] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__397_ : 1'b0;
  assign data_o_flat[396] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__396_ : 1'b0;
  assign data_o_flat[395] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__395_ : 1'b0;
  assign data_o_flat[394] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__394_ : 1'b0;
  assign data_o_flat[393] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__393_ : 1'b0;
  assign data_o_flat[392] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__392_ : 1'b0;
  assign data_o_flat[391] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__391_ : 1'b0;
  assign data_o_flat[390] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__390_ : 1'b0;
  assign data_o_flat[389] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__389_ : 1'b0;
  assign data_o_flat[388] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__388_ : 1'b0;
  assign data_o_flat[387] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__387_ : 1'b0;
  assign data_o_flat[386] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__386_ : 1'b0;
  assign data_o_flat[385] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__385_ : 1'b0;
  assign data_o_flat[384] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__384_ : 1'b0;
  assign data_o_flat[383] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__383_ : 1'b0;
  assign data_o_flat[382] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__382_ : 1'b0;
  assign data_o_flat[381] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__381_ : 1'b0;
  assign data_o_flat[380] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__380_ : 1'b0;
  assign data_o_flat[379] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__379_ : 1'b0;
  assign data_o_flat[378] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__378_ : 1'b0;
  assign data_o_flat[377] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__377_ : 1'b0;
  assign data_o_flat[376] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__376_ : 1'b0;
  assign data_o_flat[375] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__375_ : 1'b0;
  assign data_o_flat[374] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__374_ : 1'b0;
  assign data_o_flat[373] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__373_ : 1'b0;
  assign data_o_flat[372] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__372_ : 1'b0;
  assign data_o_flat[371] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__371_ : 1'b0;
  assign data_o_flat[370] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__370_ : 1'b0;
  assign data_o_flat[369] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__369_ : 1'b0;
  assign data_o_flat[368] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__368_ : 1'b0;
  assign data_o_flat[367] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__367_ : 1'b0;
  assign data_o_flat[366] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__366_ : 1'b0;
  assign data_o_flat[365] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__365_ : 1'b0;
  assign data_o_flat[364] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__364_ : 1'b0;
  assign data_o_flat[363] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__363_ : 1'b0;
  assign data_o_flat[362] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__362_ : 1'b0;
  assign data_o_flat[361] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__361_ : 1'b0;
  assign data_o_flat[360] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__360_ : 1'b0;
  assign data_o_flat[359] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__359_ : 1'b0;
  assign data_o_flat[358] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__358_ : 1'b0;
  assign data_o_flat[357] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__357_ : 1'b0;
  assign data_o_flat[356] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__356_ : 1'b0;
  assign data_o_flat[355] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__355_ : 1'b0;
  assign data_o_flat[354] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__354_ : 1'b0;
  assign data_o_flat[353] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__353_ : 1'b0;
  assign data_o_flat[352] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__352_ : 1'b0;
  assign data_o_flat[351] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__351_ : 1'b0;
  assign data_o_flat[350] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__350_ : 1'b0;
  assign data_o_flat[349] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__349_ : 1'b0;
  assign data_o_flat[348] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__348_ : 1'b0;
  assign data_o_flat[347] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__347_ : 1'b0;
  assign data_o_flat[346] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__346_ : 1'b0;
  assign data_o_flat[345] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__345_ : 1'b0;
  assign data_o_flat[344] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__344_ : 1'b0;
  assign data_o_flat[343] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__343_ : 1'b0;
  assign data_o_flat[342] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__342_ : 1'b0;
  assign data_o_flat[341] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__341_ : 1'b0;
  assign data_o_flat[340] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__340_ : 1'b0;
  assign data_o_flat[339] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__339_ : 1'b0;
  assign data_o_flat[338] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__338_ : 1'b0;
  assign data_o_flat[337] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__337_ : 1'b0;
  assign data_o_flat[336] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__336_ : 1'b0;
  assign data_o_flat[335] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__335_ : 1'b0;
  assign data_o_flat[334] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__334_ : 1'b0;
  assign data_o_flat[333] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__333_ : 1'b0;
  assign data_o_flat[332] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__332_ : 1'b0;
  assign data_o_flat[331] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__331_ : 1'b0;
  assign data_o_flat[330] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__330_ : 1'b0;
  assign data_o_flat[329] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__329_ : 1'b0;
  assign data_o_flat[328] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__328_ : 1'b0;
  assign data_o_flat[327] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__327_ : 1'b0;
  assign data_o_flat[326] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__326_ : 1'b0;
  assign data_o_flat[325] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__325_ : 1'b0;
  assign data_o_flat[324] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__324_ : 1'b0;
  assign data_o_flat[323] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__323_ : 1'b0;
  assign data_o_flat[322] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__322_ : 1'b0;
  assign data_o_flat[321] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__321_ : 1'b0;
  assign data_o_flat[320] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__320_ : 1'b0;
  assign data_o_flat[319] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__319_ : 1'b0;
  assign data_o_flat[318] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__318_ : 1'b0;
  assign data_o_flat[317] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__317_ : 1'b0;
  assign data_o_flat[316] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__316_ : 1'b0;
  assign data_o_flat[315] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__315_ : 1'b0;
  assign data_o_flat[314] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__314_ : 1'b0;
  assign data_o_flat[313] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__313_ : 1'b0;
  assign data_o_flat[312] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__312_ : 1'b0;
  assign data_o_flat[311] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__311_ : 1'b0;
  assign data_o_flat[310] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__310_ : 1'b0;
  assign data_o_flat[309] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__309_ : 1'b0;
  assign data_o_flat[308] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__308_ : 1'b0;
  assign data_o_flat[307] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__307_ : 1'b0;
  assign data_o_flat[306] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__306_ : 1'b0;
  assign data_o_flat[305] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__305_ : 1'b0;
  assign data_o_flat[304] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__304_ : 1'b0;
  assign data_o_flat[303] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__303_ : 1'b0;
  assign data_o_flat[302] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__302_ : 1'b0;
  assign data_o_flat[301] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__301_ : 1'b0;
  assign data_o_flat[300] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__300_ : 1'b0;
  assign data_o_flat[299] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__299_ : 1'b0;
  assign data_o_flat[298] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__298_ : 1'b0;
  assign data_o_flat[297] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__297_ : 1'b0;
  assign data_o_flat[296] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__296_ : 1'b0;
  assign data_o_flat[295] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__295_ : 1'b0;
  assign data_o_flat[294] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__294_ : 1'b0;
  assign data_o_flat[293] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__293_ : 1'b0;
  assign data_o_flat[292] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__292_ : 1'b0;
  assign data_o_flat[291] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__291_ : 1'b0;
  assign data_o_flat[290] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__290_ : 1'b0;
  assign data_o_flat[289] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__289_ : 1'b0;
  assign data_o_flat[288] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__288_ : 1'b0;
  assign data_o_flat[287] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__287_ : 1'b0;
  assign data_o_flat[286] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__286_ : 1'b0;
  assign data_o_flat[285] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__285_ : 1'b0;
  assign data_o_flat[284] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__284_ : 1'b0;
  assign data_o_flat[283] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__283_ : 1'b0;
  assign data_o_flat[282] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__282_ : 1'b0;
  assign data_o_flat[281] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__281_ : 1'b0;
  assign data_o_flat[280] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__280_ : 1'b0;
  assign data_o_flat[279] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__279_ : 1'b0;
  assign data_o_flat[278] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__278_ : 1'b0;
  assign data_o_flat[277] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__277_ : 1'b0;
  assign data_o_flat[276] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__276_ : 1'b0;
  assign data_o_flat[275] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__275_ : 1'b0;
  assign data_o_flat[274] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__274_ : 1'b0;
  assign data_o_flat[273] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__273_ : 1'b0;
  assign data_o_flat[272] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__272_ : 1'b0;
  assign data_o_flat[271] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__271_ : 1'b0;
  assign data_o_flat[270] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__270_ : 1'b0;
  assign data_o_flat[269] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__269_ : 1'b0;
  assign data_o_flat[268] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__268_ : 1'b0;
  assign data_o_flat[267] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__267_ : 1'b0;
  assign data_o_flat[266] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__266_ : 1'b0;
  assign data_o_flat[265] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__265_ : 1'b0;
  assign data_o_flat[264] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__264_ : 1'b0;
  assign data_o_flat[263] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__263_ : 1'b0;
  assign data_o_flat[262] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__262_ : 1'b0;
  assign data_o_flat[261] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__261_ : 1'b0;
  assign data_o_flat[260] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__260_ : 1'b0;
  assign data_o_flat[259] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__259_ : 1'b0;
  assign data_o_flat[258] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__258_ : 1'b0;
  assign data_o_flat[257] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__257_ : 1'b0;
  assign data_o_flat[256] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__256_ : 1'b0;
  assign data_o_flat[255] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__255_ : 1'b0;
  assign data_o_flat[254] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__254_ : 1'b0;
  assign data_o_flat[253] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__253_ : 1'b0;
  assign data_o_flat[252] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__252_ : 1'b0;
  assign data_o_flat[251] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__251_ : 1'b0;
  assign data_o_flat[250] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__250_ : 1'b0;
  assign data_o_flat[249] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__249_ : 1'b0;
  assign data_o_flat[248] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__248_ : 1'b0;
  assign data_o_flat[247] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__247_ : 1'b0;
  assign data_o_flat[246] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__246_ : 1'b0;
  assign data_o_flat[245] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__245_ : 1'b0;
  assign data_o_flat[244] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__244_ : 1'b0;
  assign data_o_flat[243] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__243_ : 1'b0;
  assign data_o_flat[242] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__242_ : 1'b0;
  assign data_o_flat[241] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__241_ : 1'b0;
  assign data_o_flat[240] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__240_ : 1'b0;
  assign data_o_flat[239] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__239_ : 1'b0;
  assign data_o_flat[238] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__238_ : 1'b0;
  assign data_o_flat[237] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__237_ : 1'b0;
  assign data_o_flat[236] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__236_ : 1'b0;
  assign data_o_flat[235] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__235_ : 1'b0;
  assign data_o_flat[234] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__234_ : 1'b0;
  assign data_o_flat[233] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__233_ : 1'b0;
  assign data_o_flat[232] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__232_ : 1'b0;
  assign data_o_flat[231] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__231_ : 1'b0;
  assign data_o_flat[230] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__230_ : 1'b0;
  assign data_o_flat[229] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__229_ : 1'b0;
  assign data_o_flat[228] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__228_ : 1'b0;
  assign data_o_flat[227] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__227_ : 1'b0;
  assign data_o_flat[226] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__226_ : 1'b0;
  assign data_o_flat[225] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__225_ : 1'b0;
  assign data_o_flat[224] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__224_ : 1'b0;
  assign data_o_flat[223] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__223_ : 1'b0;
  assign data_o_flat[222] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__222_ : 1'b0;
  assign data_o_flat[221] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__221_ : 1'b0;
  assign data_o_flat[220] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__220_ : 1'b0;
  assign data_o_flat[219] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__219_ : 1'b0;
  assign data_o_flat[218] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__218_ : 1'b0;
  assign data_o_flat[217] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__217_ : 1'b0;
  assign data_o_flat[216] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__216_ : 1'b0;
  assign data_o_flat[215] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__215_ : 1'b0;
  assign data_o_flat[214] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__214_ : 1'b0;
  assign data_o_flat[213] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__213_ : 1'b0;
  assign data_o_flat[212] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__212_ : 1'b0;
  assign data_o_flat[211] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__211_ : 1'b0;
  assign data_o_flat[210] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__210_ : 1'b0;
  assign data_o_flat[209] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__209_ : 1'b0;
  assign data_o_flat[208] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__208_ : 1'b0;
  assign data_o_flat[207] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__207_ : 1'b0;
  assign data_o_flat[206] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__206_ : 1'b0;
  assign data_o_flat[205] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__205_ : 1'b0;
  assign data_o_flat[204] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__204_ : 1'b0;
  assign data_o_flat[203] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__203_ : 1'b0;
  assign data_o_flat[202] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__202_ : 1'b0;
  assign data_o_flat[201] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__201_ : 1'b0;
  assign data_o_flat[200] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__200_ : 1'b0;
  assign data_o_flat[199] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__199_ : 1'b0;
  assign data_o_flat[198] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__198_ : 1'b0;
  assign data_o_flat[197] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__197_ : 1'b0;
  assign data_o_flat[196] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__196_ : 1'b0;
  assign data_o_flat[195] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__195_ : 1'b0;
  assign data_o_flat[194] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__194_ : 1'b0;
  assign data_o_flat[193] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__193_ : 1'b0;
  assign data_o_flat[192] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__192_ : 1'b0;
  assign data_o_flat[191] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__191_ : 1'b0;
  assign data_o_flat[190] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__190_ : 1'b0;
  assign data_o_flat[189] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__189_ : 1'b0;
  assign data_o_flat[188] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__188_ : 1'b0;
  assign data_o_flat[187] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__187_ : 1'b0;
  assign data_o_flat[186] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__186_ : 1'b0;
  assign data_o_flat[185] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__185_ : 1'b0;
  assign data_o_flat[184] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__184_ : 1'b0;
  assign data_o_flat[183] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__183_ : 1'b0;
  assign data_o_flat[182] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__182_ : 1'b0;
  assign data_o_flat[181] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__181_ : 1'b0;
  assign data_o_flat[180] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__180_ : 1'b0;
  assign data_o_flat[179] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__179_ : 1'b0;
  assign data_o_flat[178] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__178_ : 1'b0;
  assign data_o_flat[177] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__177_ : 1'b0;
  assign data_o_flat[176] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__176_ : 1'b0;
  assign data_o_flat[175] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__175_ : 1'b0;
  assign data_o_flat[174] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__174_ : 1'b0;
  assign data_o_flat[173] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__173_ : 1'b0;
  assign data_o_flat[172] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__172_ : 1'b0;
  assign data_o_flat[171] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__171_ : 1'b0;
  assign data_o_flat[170] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__170_ : 1'b0;
  assign data_o_flat[169] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__169_ : 1'b0;
  assign data_o_flat[168] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__168_ : 1'b0;
  assign data_o_flat[167] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__167_ : 1'b0;
  assign data_o_flat[166] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__166_ : 1'b0;
  assign data_o_flat[165] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__165_ : 1'b0;
  assign data_o_flat[164] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__164_ : 1'b0;
  assign data_o_flat[163] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__163_ : 1'b0;
  assign data_o_flat[162] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__162_ : 1'b0;
  assign data_o_flat[161] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__161_ : 1'b0;
  assign data_o_flat[160] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__160_ : 1'b0;
  assign data_o_flat[159] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__159_ : 1'b0;
  assign data_o_flat[158] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__158_ : 1'b0;
  assign data_o_flat[157] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__157_ : 1'b0;
  assign data_o_flat[156] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__156_ : 1'b0;
  assign data_o_flat[155] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__155_ : 1'b0;
  assign data_o_flat[154] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__154_ : 1'b0;
  assign data_o_flat[153] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__153_ : 1'b0;
  assign data_o_flat[152] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__152_ : 1'b0;
  assign data_o_flat[151] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__151_ : 1'b0;
  assign data_o_flat[150] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__150_ : 1'b0;
  assign data_o_flat[149] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__149_ : 1'b0;
  assign data_o_flat[148] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__148_ : 1'b0;
  assign data_o_flat[147] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__147_ : 1'b0;
  assign data_o_flat[146] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__146_ : 1'b0;
  assign data_o_flat[145] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__145_ : 1'b0;
  assign data_o_flat[144] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__144_ : 1'b0;
  assign data_o_flat[143] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__143_ : 1'b0;
  assign data_o_flat[142] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__142_ : 1'b0;
  assign data_o_flat[141] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__141_ : 1'b0;
  assign data_o_flat[140] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__140_ : 1'b0;
  assign data_o_flat[139] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__139_ : 1'b0;
  assign data_o_flat[138] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__138_ : 1'b0;
  assign data_o_flat[137] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__137_ : 1'b0;
  assign data_o_flat[136] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__136_ : 1'b0;
  assign data_o_flat[135] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__135_ : 1'b0;
  assign data_o_flat[134] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__134_ : 1'b0;
  assign data_o_flat[133] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__133_ : 1'b0;
  assign data_o_flat[132] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__132_ : 1'b0;
  assign data_o_flat[131] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__131_ : 1'b0;
  assign data_o_flat[130] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__130_ : 1'b0;
  assign data_o_flat[129] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__129_ : 1'b0;
  assign data_o_flat[128] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__128_ : 1'b0;
  assign data_o_flat[127] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__127_ : 1'b0;
  assign data_o_flat[126] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__126_ : 1'b0;
  assign data_o_flat[125] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__125_ : 1'b0;
  assign data_o_flat[124] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__124_ : 1'b0;
  assign data_o_flat[123] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__123_ : 1'b0;
  assign data_o_flat[122] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__122_ : 1'b0;
  assign data_o_flat[121] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__121_ : 1'b0;
  assign data_o_flat[120] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__120_ : 1'b0;
  assign data_o_flat[119] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__119_ : 1'b0;
  assign data_o_flat[118] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__118_ : 1'b0;
  assign data_o_flat[117] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__117_ : 1'b0;
  assign data_o_flat[116] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__116_ : 1'b0;
  assign data_o_flat[115] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__115_ : 1'b0;
  assign data_o_flat[114] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__114_ : 1'b0;
  assign data_o_flat[113] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__113_ : 1'b0;
  assign data_o_flat[112] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__112_ : 1'b0;
  assign data_o_flat[111] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__111_ : 1'b0;
  assign data_o_flat[110] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__110_ : 1'b0;
  assign data_o_flat[109] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__109_ : 1'b0;
  assign data_o_flat[108] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__108_ : 1'b0;
  assign data_o_flat[107] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__107_ : 1'b0;
  assign data_o_flat[106] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__106_ : 1'b0;
  assign data_o_flat[105] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__105_ : 1'b0;
  assign data_o_flat[104] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__104_ : 1'b0;
  assign data_o_flat[103] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__103_ : 1'b0;
  assign data_o_flat[102] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__102_ : 1'b0;
  assign data_o_flat[101] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__101_ : 1'b0;
  assign data_o_flat[100] = (N95)? 1'b0 : 
                            (N96)? 1'b0 : 
                            (N97)? 1'b0 : 
                            (N98)? 1'b0 : 
                            (N99)? 1'b0 : 
                            (N100)? 1'b0 : 
                            (N101)? 1'b0 : 
                            (N102)? 1'b0 : 
                            (N103)? 1'b0 : 
                            (N104)? data_int_o_9__100_ : 1'b0;
  assign data_o_flat[99] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__99_ : 1'b0;
  assign data_o_flat[98] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__98_ : 1'b0;
  assign data_o_flat[97] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__97_ : 1'b0;
  assign data_o_flat[96] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__96_ : 1'b0;
  assign data_o_flat[95] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__95_ : 1'b0;
  assign data_o_flat[94] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__94_ : 1'b0;
  assign data_o_flat[93] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__93_ : 1'b0;
  assign data_o_flat[92] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__92_ : 1'b0;
  assign data_o_flat[91] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__91_ : 1'b0;
  assign data_o_flat[90] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__90_ : 1'b0;
  assign data_o_flat[89] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__89_ : 1'b0;
  assign data_o_flat[88] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__88_ : 1'b0;
  assign data_o_flat[87] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__87_ : 1'b0;
  assign data_o_flat[86] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__86_ : 1'b0;
  assign data_o_flat[85] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__85_ : 1'b0;
  assign data_o_flat[84] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__84_ : 1'b0;
  assign data_o_flat[83] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__83_ : 1'b0;
  assign data_o_flat[82] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__82_ : 1'b0;
  assign data_o_flat[81] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__81_ : 1'b0;
  assign data_o_flat[80] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__80_ : 1'b0;
  assign data_o_flat[79] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__79_ : 1'b0;
  assign data_o_flat[78] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__78_ : 1'b0;
  assign data_o_flat[77] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__77_ : 1'b0;
  assign data_o_flat[76] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__76_ : 1'b0;
  assign data_o_flat[75] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__75_ : 1'b0;
  assign data_o_flat[74] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__74_ : 1'b0;
  assign data_o_flat[73] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__73_ : 1'b0;
  assign data_o_flat[72] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__72_ : 1'b0;
  assign data_o_flat[71] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__71_ : 1'b0;
  assign data_o_flat[70] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__70_ : 1'b0;
  assign data_o_flat[69] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__69_ : 1'b0;
  assign data_o_flat[68] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__68_ : 1'b0;
  assign data_o_flat[67] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__67_ : 1'b0;
  assign data_o_flat[66] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__66_ : 1'b0;
  assign data_o_flat[65] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__65_ : 1'b0;
  assign data_o_flat[64] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__64_ : 1'b0;
  assign data_o_flat[63] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__63_ : 1'b0;
  assign data_o_flat[62] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__62_ : 1'b0;
  assign data_o_flat[61] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__61_ : 1'b0;
  assign data_o_flat[60] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__60_ : 1'b0;
  assign data_o_flat[59] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__59_ : 1'b0;
  assign data_o_flat[58] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__58_ : 1'b0;
  assign data_o_flat[57] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__57_ : 1'b0;
  assign data_o_flat[56] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__56_ : 1'b0;
  assign data_o_flat[55] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__55_ : 1'b0;
  assign data_o_flat[54] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__54_ : 1'b0;
  assign data_o_flat[53] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__53_ : 1'b0;
  assign data_o_flat[52] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__52_ : 1'b0;
  assign data_o_flat[51] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__51_ : 1'b0;
  assign data_o_flat[50] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__50_ : 1'b0;
  assign data_o_flat[49] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__49_ : 1'b0;
  assign data_o_flat[48] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__48_ : 1'b0;
  assign data_o_flat[47] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__47_ : 1'b0;
  assign data_o_flat[46] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__46_ : 1'b0;
  assign data_o_flat[45] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__45_ : 1'b0;
  assign data_o_flat[44] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__44_ : 1'b0;
  assign data_o_flat[43] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__43_ : 1'b0;
  assign data_o_flat[42] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__42_ : 1'b0;
  assign data_o_flat[41] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__41_ : 1'b0;
  assign data_o_flat[40] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__40_ : 1'b0;
  assign data_o_flat[39] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__39_ : 1'b0;
  assign data_o_flat[38] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__38_ : 1'b0;
  assign data_o_flat[37] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__37_ : 1'b0;
  assign data_o_flat[36] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__36_ : 1'b0;
  assign data_o_flat[35] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__35_ : 1'b0;
  assign data_o_flat[34] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__34_ : 1'b0;
  assign data_o_flat[33] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__33_ : 1'b0;
  assign data_o_flat[32] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__32_ : 1'b0;
  assign data_o_flat[31] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__31_ : 1'b0;
  assign data_o_flat[30] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__30_ : 1'b0;
  assign data_o_flat[29] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__29_ : 1'b0;
  assign data_o_flat[28] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__28_ : 1'b0;
  assign data_o_flat[27] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__27_ : 1'b0;
  assign data_o_flat[26] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__26_ : 1'b0;
  assign data_o_flat[25] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__25_ : 1'b0;
  assign data_o_flat[24] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__24_ : 1'b0;
  assign data_o_flat[23] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__23_ : 1'b0;
  assign data_o_flat[22] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__22_ : 1'b0;
  assign data_o_flat[21] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__21_ : 1'b0;
  assign data_o_flat[20] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__20_ : 1'b0;
  assign data_o_flat[19] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__19_ : 1'b0;
  assign data_o_flat[18] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__18_ : 1'b0;
  assign data_o_flat[17] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__17_ : 1'b0;
  assign data_o_flat[16] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__16_ : 1'b0;
  assign data_o_flat[15] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__15_ : 1'b0;
  assign data_o_flat[14] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__14_ : 1'b0;
  assign data_o_flat[13] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__13_ : 1'b0;
  assign data_o_flat[12] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__12_ : 1'b0;
  assign data_o_flat[11] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__11_ : 1'b0;
  assign data_o_flat[10] = (N95)? 1'b0 : 
                           (N96)? 1'b0 : 
                           (N97)? 1'b0 : 
                           (N98)? 1'b0 : 
                           (N99)? 1'b0 : 
                           (N100)? 1'b0 : 
                           (N101)? 1'b0 : 
                           (N102)? 1'b0 : 
                           (N103)? 1'b0 : 
                           (N104)? data_int_o_9__10_ : 1'b0;
  assign data_o_flat[9] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__9_ : 1'b0;
  assign data_o_flat[8] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__8_ : 1'b0;
  assign data_o_flat[7] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__7_ : 1'b0;
  assign data_o_flat[6] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__6_ : 1'b0;
  assign data_o_flat[5] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__5_ : 1'b0;
  assign data_o_flat[4] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__4_ : 1'b0;
  assign data_o_flat[3] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__3_ : 1'b0;
  assign data_o_flat[2] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__2_ : 1'b0;
  assign data_o_flat[1] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__1_ : 1'b0;
  assign data_o_flat[0] = (N95)? 1'b0 : 
                          (N96)? 1'b0 : 
                          (N97)? 1'b0 : 
                          (N98)? 1'b0 : 
                          (N99)? 1'b0 : 
                          (N100)? 1'b0 : 
                          (N101)? 1'b0 : 
                          (N102)? 1'b0 : 
                          (N103)? 1'b0 : 
                          (N104)? data_int_o_9__0_ : 1'b0;
  assign n_2_net__9_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__9_ : 1'b0;
  assign N105 = N155;
  assign N106 = N157;
  assign N107 = N159;
  assign N108 = N160;
  assign N109 = N161;
  assign N110 = N162;
  assign N111 = N163;
  assign N112 = N164;
  assign N113 = N156;
  assign N114 = N158;
  assign n_2_net__8_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__8_ : 1'b0;
  assign n_2_net__7_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__7_ : 1'b0;
  assign n_2_net__6_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__6_ : 1'b0;
  assign n_2_net__5_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__5_ : 1'b0;
  assign n_2_net__4_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__4_ : 1'b0;
  assign n_2_net__3_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__3_ : 1'b0;
  assign n_2_net__2_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__2_ : 1'b0;
  assign n_2_net__1_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__1_ : 1'b0;
  assign n_2_net__0_ = (N105)? 1'b0 : 
                       (N106)? 1'b0 : 
                       (N107)? 1'b0 : 
                       (N108)? 1'b0 : 
                       (N109)? 1'b0 : 
                       (N110)? 1'b0 : 
                       (N111)? 1'b0 : 
                       (N112)? 1'b0 : 
                       (N113)? 1'b0 : 
                       (N114)? valid_head_9__0_ : 1'b0;
  assign n_3_net__9_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__9_ : 1'b0;
  assign n_3_net__8_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__8_ : 1'b0;
  assign n_3_net__7_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__7_ : 1'b0;
  assign n_3_net__6_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__6_ : 1'b0;
  assign n_3_net__5_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__5_ : 1'b0;
  assign n_3_net__4_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__4_ : 1'b0;
  assign n_3_net__3_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__3_ : 1'b0;
  assign n_3_net__2_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__2_ : 1'b0;
  assign n_3_net__1_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__1_ : 1'b0;
  assign n_3_net__0_ = (N85)? 1'b0 : 
                       (N86)? 1'b0 : 
                       (N87)? 1'b0 : 
                       (N88)? 1'b0 : 
                       (N89)? 1'b0 : 
                       (N90)? 1'b0 : 
                       (N91)? 1'b0 : 
                       (N92)? 1'b0 : 
                       (N93)? 1'b0 : 
                       (N94)? ready_head_9__0_ : 1'b0;
  assign n_4_net__1279_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1279_ : 1'b0;
  assign N115 = N165;
  assign N116 = N167;
  assign N117 = N169;
  assign N118 = N170;
  assign N119 = N171;
  assign N120 = N172;
  assign N121 = N173;
  assign N122 = N174;
  assign N123 = N166;
  assign N124 = N168;
  assign n_4_net__1278_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1278_ : 1'b0;
  assign n_4_net__1277_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1277_ : 1'b0;
  assign n_4_net__1276_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1276_ : 1'b0;
  assign n_4_net__1275_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1275_ : 1'b0;
  assign n_4_net__1274_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1274_ : 1'b0;
  assign n_4_net__1273_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1273_ : 1'b0;
  assign n_4_net__1272_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1272_ : 1'b0;
  assign n_4_net__1271_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1271_ : 1'b0;
  assign n_4_net__1270_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1270_ : 1'b0;
  assign n_4_net__1269_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1269_ : 1'b0;
  assign n_4_net__1268_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1268_ : 1'b0;
  assign n_4_net__1267_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1267_ : 1'b0;
  assign n_4_net__1266_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1266_ : 1'b0;
  assign n_4_net__1265_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1265_ : 1'b0;
  assign n_4_net__1264_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1264_ : 1'b0;
  assign n_4_net__1263_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1263_ : 1'b0;
  assign n_4_net__1262_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1262_ : 1'b0;
  assign n_4_net__1261_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1261_ : 1'b0;
  assign n_4_net__1260_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1260_ : 1'b0;
  assign n_4_net__1259_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1259_ : 1'b0;
  assign n_4_net__1258_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1258_ : 1'b0;
  assign n_4_net__1257_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1257_ : 1'b0;
  assign n_4_net__1256_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1256_ : 1'b0;
  assign n_4_net__1255_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1255_ : 1'b0;
  assign n_4_net__1254_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1254_ : 1'b0;
  assign n_4_net__1253_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1253_ : 1'b0;
  assign n_4_net__1252_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1252_ : 1'b0;
  assign n_4_net__1251_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1251_ : 1'b0;
  assign n_4_net__1250_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1250_ : 1'b0;
  assign n_4_net__1249_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1249_ : 1'b0;
  assign n_4_net__1248_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1248_ : 1'b0;
  assign n_4_net__1247_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1247_ : 1'b0;
  assign n_4_net__1246_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1246_ : 1'b0;
  assign n_4_net__1245_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1245_ : 1'b0;
  assign n_4_net__1244_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1244_ : 1'b0;
  assign n_4_net__1243_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1243_ : 1'b0;
  assign n_4_net__1242_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1242_ : 1'b0;
  assign n_4_net__1241_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1241_ : 1'b0;
  assign n_4_net__1240_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1240_ : 1'b0;
  assign n_4_net__1239_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1239_ : 1'b0;
  assign n_4_net__1238_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1238_ : 1'b0;
  assign n_4_net__1237_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1237_ : 1'b0;
  assign n_4_net__1236_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1236_ : 1'b0;
  assign n_4_net__1235_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1235_ : 1'b0;
  assign n_4_net__1234_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1234_ : 1'b0;
  assign n_4_net__1233_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1233_ : 1'b0;
  assign n_4_net__1232_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1232_ : 1'b0;
  assign n_4_net__1231_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1231_ : 1'b0;
  assign n_4_net__1230_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1230_ : 1'b0;
  assign n_4_net__1229_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1229_ : 1'b0;
  assign n_4_net__1228_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1228_ : 1'b0;
  assign n_4_net__1227_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1227_ : 1'b0;
  assign n_4_net__1226_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1226_ : 1'b0;
  assign n_4_net__1225_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1225_ : 1'b0;
  assign n_4_net__1224_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1224_ : 1'b0;
  assign n_4_net__1223_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1223_ : 1'b0;
  assign n_4_net__1222_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1222_ : 1'b0;
  assign n_4_net__1221_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1221_ : 1'b0;
  assign n_4_net__1220_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1220_ : 1'b0;
  assign n_4_net__1219_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1219_ : 1'b0;
  assign n_4_net__1218_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1218_ : 1'b0;
  assign n_4_net__1217_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1217_ : 1'b0;
  assign n_4_net__1216_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1216_ : 1'b0;
  assign n_4_net__1215_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1215_ : 1'b0;
  assign n_4_net__1214_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1214_ : 1'b0;
  assign n_4_net__1213_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1213_ : 1'b0;
  assign n_4_net__1212_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1212_ : 1'b0;
  assign n_4_net__1211_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1211_ : 1'b0;
  assign n_4_net__1210_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1210_ : 1'b0;
  assign n_4_net__1209_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1209_ : 1'b0;
  assign n_4_net__1208_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1208_ : 1'b0;
  assign n_4_net__1207_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1207_ : 1'b0;
  assign n_4_net__1206_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1206_ : 1'b0;
  assign n_4_net__1205_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1205_ : 1'b0;
  assign n_4_net__1204_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1204_ : 1'b0;
  assign n_4_net__1203_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1203_ : 1'b0;
  assign n_4_net__1202_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1202_ : 1'b0;
  assign n_4_net__1201_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1201_ : 1'b0;
  assign n_4_net__1200_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1200_ : 1'b0;
  assign n_4_net__1199_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1199_ : 1'b0;
  assign n_4_net__1198_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1198_ : 1'b0;
  assign n_4_net__1197_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1197_ : 1'b0;
  assign n_4_net__1196_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1196_ : 1'b0;
  assign n_4_net__1195_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1195_ : 1'b0;
  assign n_4_net__1194_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1194_ : 1'b0;
  assign n_4_net__1193_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1193_ : 1'b0;
  assign n_4_net__1192_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1192_ : 1'b0;
  assign n_4_net__1191_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1191_ : 1'b0;
  assign n_4_net__1190_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1190_ : 1'b0;
  assign n_4_net__1189_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1189_ : 1'b0;
  assign n_4_net__1188_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1188_ : 1'b0;
  assign n_4_net__1187_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1187_ : 1'b0;
  assign n_4_net__1186_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1186_ : 1'b0;
  assign n_4_net__1185_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1185_ : 1'b0;
  assign n_4_net__1184_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1184_ : 1'b0;
  assign n_4_net__1183_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1183_ : 1'b0;
  assign n_4_net__1182_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1182_ : 1'b0;
  assign n_4_net__1181_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1181_ : 1'b0;
  assign n_4_net__1180_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1180_ : 1'b0;
  assign n_4_net__1179_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1179_ : 1'b0;
  assign n_4_net__1178_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1178_ : 1'b0;
  assign n_4_net__1177_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1177_ : 1'b0;
  assign n_4_net__1176_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1176_ : 1'b0;
  assign n_4_net__1175_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1175_ : 1'b0;
  assign n_4_net__1174_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1174_ : 1'b0;
  assign n_4_net__1173_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1173_ : 1'b0;
  assign n_4_net__1172_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1172_ : 1'b0;
  assign n_4_net__1171_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1171_ : 1'b0;
  assign n_4_net__1170_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1170_ : 1'b0;
  assign n_4_net__1169_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1169_ : 1'b0;
  assign n_4_net__1168_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1168_ : 1'b0;
  assign n_4_net__1167_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1167_ : 1'b0;
  assign n_4_net__1166_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1166_ : 1'b0;
  assign n_4_net__1165_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1165_ : 1'b0;
  assign n_4_net__1164_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1164_ : 1'b0;
  assign n_4_net__1163_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1163_ : 1'b0;
  assign n_4_net__1162_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1162_ : 1'b0;
  assign n_4_net__1161_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1161_ : 1'b0;
  assign n_4_net__1160_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1160_ : 1'b0;
  assign n_4_net__1159_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1159_ : 1'b0;
  assign n_4_net__1158_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1158_ : 1'b0;
  assign n_4_net__1157_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1157_ : 1'b0;
  assign n_4_net__1156_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1156_ : 1'b0;
  assign n_4_net__1155_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1155_ : 1'b0;
  assign n_4_net__1154_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1154_ : 1'b0;
  assign n_4_net__1153_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1153_ : 1'b0;
  assign n_4_net__1152_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1152_ : 1'b0;
  assign n_4_net__1151_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1151_ : 1'b0;
  assign n_4_net__1150_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1150_ : 1'b0;
  assign n_4_net__1149_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1149_ : 1'b0;
  assign n_4_net__1148_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1148_ : 1'b0;
  assign n_4_net__1147_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1147_ : 1'b0;
  assign n_4_net__1146_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1146_ : 1'b0;
  assign n_4_net__1145_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1145_ : 1'b0;
  assign n_4_net__1144_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1144_ : 1'b0;
  assign n_4_net__1143_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1143_ : 1'b0;
  assign n_4_net__1142_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1142_ : 1'b0;
  assign n_4_net__1141_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1141_ : 1'b0;
  assign n_4_net__1140_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1140_ : 1'b0;
  assign n_4_net__1139_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1139_ : 1'b0;
  assign n_4_net__1138_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1138_ : 1'b0;
  assign n_4_net__1137_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1137_ : 1'b0;
  assign n_4_net__1136_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1136_ : 1'b0;
  assign n_4_net__1135_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1135_ : 1'b0;
  assign n_4_net__1134_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1134_ : 1'b0;
  assign n_4_net__1133_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1133_ : 1'b0;
  assign n_4_net__1132_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1132_ : 1'b0;
  assign n_4_net__1131_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1131_ : 1'b0;
  assign n_4_net__1130_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1130_ : 1'b0;
  assign n_4_net__1129_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1129_ : 1'b0;
  assign n_4_net__1128_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1128_ : 1'b0;
  assign n_4_net__1127_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1127_ : 1'b0;
  assign n_4_net__1126_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1126_ : 1'b0;
  assign n_4_net__1125_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1125_ : 1'b0;
  assign n_4_net__1124_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1124_ : 1'b0;
  assign n_4_net__1123_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1123_ : 1'b0;
  assign n_4_net__1122_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1122_ : 1'b0;
  assign n_4_net__1121_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1121_ : 1'b0;
  assign n_4_net__1120_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1120_ : 1'b0;
  assign n_4_net__1119_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1119_ : 1'b0;
  assign n_4_net__1118_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1118_ : 1'b0;
  assign n_4_net__1117_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1117_ : 1'b0;
  assign n_4_net__1116_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1116_ : 1'b0;
  assign n_4_net__1115_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1115_ : 1'b0;
  assign n_4_net__1114_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1114_ : 1'b0;
  assign n_4_net__1113_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1113_ : 1'b0;
  assign n_4_net__1112_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1112_ : 1'b0;
  assign n_4_net__1111_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1111_ : 1'b0;
  assign n_4_net__1110_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1110_ : 1'b0;
  assign n_4_net__1109_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1109_ : 1'b0;
  assign n_4_net__1108_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1108_ : 1'b0;
  assign n_4_net__1107_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1107_ : 1'b0;
  assign n_4_net__1106_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1106_ : 1'b0;
  assign n_4_net__1105_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1105_ : 1'b0;
  assign n_4_net__1104_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1104_ : 1'b0;
  assign n_4_net__1103_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1103_ : 1'b0;
  assign n_4_net__1102_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1102_ : 1'b0;
  assign n_4_net__1101_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1101_ : 1'b0;
  assign n_4_net__1100_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1100_ : 1'b0;
  assign n_4_net__1099_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1099_ : 1'b0;
  assign n_4_net__1098_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1098_ : 1'b0;
  assign n_4_net__1097_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1097_ : 1'b0;
  assign n_4_net__1096_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1096_ : 1'b0;
  assign n_4_net__1095_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1095_ : 1'b0;
  assign n_4_net__1094_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1094_ : 1'b0;
  assign n_4_net__1093_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1093_ : 1'b0;
  assign n_4_net__1092_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1092_ : 1'b0;
  assign n_4_net__1091_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1091_ : 1'b0;
  assign n_4_net__1090_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1090_ : 1'b0;
  assign n_4_net__1089_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1089_ : 1'b0;
  assign n_4_net__1088_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1088_ : 1'b0;
  assign n_4_net__1087_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1087_ : 1'b0;
  assign n_4_net__1086_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1086_ : 1'b0;
  assign n_4_net__1085_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1085_ : 1'b0;
  assign n_4_net__1084_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1084_ : 1'b0;
  assign n_4_net__1083_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1083_ : 1'b0;
  assign n_4_net__1082_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1082_ : 1'b0;
  assign n_4_net__1081_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1081_ : 1'b0;
  assign n_4_net__1080_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1080_ : 1'b0;
  assign n_4_net__1079_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1079_ : 1'b0;
  assign n_4_net__1078_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1078_ : 1'b0;
  assign n_4_net__1077_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1077_ : 1'b0;
  assign n_4_net__1076_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1076_ : 1'b0;
  assign n_4_net__1075_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1075_ : 1'b0;
  assign n_4_net__1074_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1074_ : 1'b0;
  assign n_4_net__1073_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1073_ : 1'b0;
  assign n_4_net__1072_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1072_ : 1'b0;
  assign n_4_net__1071_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1071_ : 1'b0;
  assign n_4_net__1070_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1070_ : 1'b0;
  assign n_4_net__1069_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1069_ : 1'b0;
  assign n_4_net__1068_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1068_ : 1'b0;
  assign n_4_net__1067_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1067_ : 1'b0;
  assign n_4_net__1066_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1066_ : 1'b0;
  assign n_4_net__1065_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1065_ : 1'b0;
  assign n_4_net__1064_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1064_ : 1'b0;
  assign n_4_net__1063_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1063_ : 1'b0;
  assign n_4_net__1062_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1062_ : 1'b0;
  assign n_4_net__1061_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1061_ : 1'b0;
  assign n_4_net__1060_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1060_ : 1'b0;
  assign n_4_net__1059_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1059_ : 1'b0;
  assign n_4_net__1058_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1058_ : 1'b0;
  assign n_4_net__1057_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1057_ : 1'b0;
  assign n_4_net__1056_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1056_ : 1'b0;
  assign n_4_net__1055_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1055_ : 1'b0;
  assign n_4_net__1054_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1054_ : 1'b0;
  assign n_4_net__1053_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1053_ : 1'b0;
  assign n_4_net__1052_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1052_ : 1'b0;
  assign n_4_net__1051_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1051_ : 1'b0;
  assign n_4_net__1050_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1050_ : 1'b0;
  assign n_4_net__1049_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1049_ : 1'b0;
  assign n_4_net__1048_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1048_ : 1'b0;
  assign n_4_net__1047_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1047_ : 1'b0;
  assign n_4_net__1046_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1046_ : 1'b0;
  assign n_4_net__1045_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1045_ : 1'b0;
  assign n_4_net__1044_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1044_ : 1'b0;
  assign n_4_net__1043_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1043_ : 1'b0;
  assign n_4_net__1042_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1042_ : 1'b0;
  assign n_4_net__1041_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1041_ : 1'b0;
  assign n_4_net__1040_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1040_ : 1'b0;
  assign n_4_net__1039_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1039_ : 1'b0;
  assign n_4_net__1038_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1038_ : 1'b0;
  assign n_4_net__1037_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1037_ : 1'b0;
  assign n_4_net__1036_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1036_ : 1'b0;
  assign n_4_net__1035_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1035_ : 1'b0;
  assign n_4_net__1034_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1034_ : 1'b0;
  assign n_4_net__1033_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1033_ : 1'b0;
  assign n_4_net__1032_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1032_ : 1'b0;
  assign n_4_net__1031_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1031_ : 1'b0;
  assign n_4_net__1030_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1030_ : 1'b0;
  assign n_4_net__1029_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1029_ : 1'b0;
  assign n_4_net__1028_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1028_ : 1'b0;
  assign n_4_net__1027_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1027_ : 1'b0;
  assign n_4_net__1026_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1026_ : 1'b0;
  assign n_4_net__1025_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1025_ : 1'b0;
  assign n_4_net__1024_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1024_ : 1'b0;
  assign n_4_net__1023_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1023_ : 1'b0;
  assign n_4_net__1022_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1022_ : 1'b0;
  assign n_4_net__1021_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1021_ : 1'b0;
  assign n_4_net__1020_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1020_ : 1'b0;
  assign n_4_net__1019_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1019_ : 1'b0;
  assign n_4_net__1018_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1018_ : 1'b0;
  assign n_4_net__1017_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1017_ : 1'b0;
  assign n_4_net__1016_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1016_ : 1'b0;
  assign n_4_net__1015_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1015_ : 1'b0;
  assign n_4_net__1014_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1014_ : 1'b0;
  assign n_4_net__1013_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1013_ : 1'b0;
  assign n_4_net__1012_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1012_ : 1'b0;
  assign n_4_net__1011_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1011_ : 1'b0;
  assign n_4_net__1010_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1010_ : 1'b0;
  assign n_4_net__1009_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1009_ : 1'b0;
  assign n_4_net__1008_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1008_ : 1'b0;
  assign n_4_net__1007_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1007_ : 1'b0;
  assign n_4_net__1006_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1006_ : 1'b0;
  assign n_4_net__1005_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1005_ : 1'b0;
  assign n_4_net__1004_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1004_ : 1'b0;
  assign n_4_net__1003_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1003_ : 1'b0;
  assign n_4_net__1002_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1002_ : 1'b0;
  assign n_4_net__1001_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1001_ : 1'b0;
  assign n_4_net__1000_ = (N115)? 1'b0 : 
                          (N116)? 1'b0 : 
                          (N117)? 1'b0 : 
                          (N118)? 1'b0 : 
                          (N119)? 1'b0 : 
                          (N120)? 1'b0 : 
                          (N121)? 1'b0 : 
                          (N122)? 1'b0 : 
                          (N123)? 1'b0 : 
                          (N124)? data_head_9__1000_ : 1'b0;
  assign n_4_net__999_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__999_ : 1'b0;
  assign n_4_net__998_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__998_ : 1'b0;
  assign n_4_net__997_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__997_ : 1'b0;
  assign n_4_net__996_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__996_ : 1'b0;
  assign n_4_net__995_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__995_ : 1'b0;
  assign n_4_net__994_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__994_ : 1'b0;
  assign n_4_net__993_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__993_ : 1'b0;
  assign n_4_net__992_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__992_ : 1'b0;
  assign n_4_net__991_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__991_ : 1'b0;
  assign n_4_net__990_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__990_ : 1'b0;
  assign n_4_net__989_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__989_ : 1'b0;
  assign n_4_net__988_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__988_ : 1'b0;
  assign n_4_net__987_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__987_ : 1'b0;
  assign n_4_net__986_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__986_ : 1'b0;
  assign n_4_net__985_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__985_ : 1'b0;
  assign n_4_net__984_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__984_ : 1'b0;
  assign n_4_net__983_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__983_ : 1'b0;
  assign n_4_net__982_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__982_ : 1'b0;
  assign n_4_net__981_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__981_ : 1'b0;
  assign n_4_net__980_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__980_ : 1'b0;
  assign n_4_net__979_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__979_ : 1'b0;
  assign n_4_net__978_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__978_ : 1'b0;
  assign n_4_net__977_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__977_ : 1'b0;
  assign n_4_net__976_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__976_ : 1'b0;
  assign n_4_net__975_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__975_ : 1'b0;
  assign n_4_net__974_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__974_ : 1'b0;
  assign n_4_net__973_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__973_ : 1'b0;
  assign n_4_net__972_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__972_ : 1'b0;
  assign n_4_net__971_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__971_ : 1'b0;
  assign n_4_net__970_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__970_ : 1'b0;
  assign n_4_net__969_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__969_ : 1'b0;
  assign n_4_net__968_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__968_ : 1'b0;
  assign n_4_net__967_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__967_ : 1'b0;
  assign n_4_net__966_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__966_ : 1'b0;
  assign n_4_net__965_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__965_ : 1'b0;
  assign n_4_net__964_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__964_ : 1'b0;
  assign n_4_net__963_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__963_ : 1'b0;
  assign n_4_net__962_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__962_ : 1'b0;
  assign n_4_net__961_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__961_ : 1'b0;
  assign n_4_net__960_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__960_ : 1'b0;
  assign n_4_net__959_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__959_ : 1'b0;
  assign n_4_net__958_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__958_ : 1'b0;
  assign n_4_net__957_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__957_ : 1'b0;
  assign n_4_net__956_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__956_ : 1'b0;
  assign n_4_net__955_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__955_ : 1'b0;
  assign n_4_net__954_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__954_ : 1'b0;
  assign n_4_net__953_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__953_ : 1'b0;
  assign n_4_net__952_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__952_ : 1'b0;
  assign n_4_net__951_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__951_ : 1'b0;
  assign n_4_net__950_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__950_ : 1'b0;
  assign n_4_net__949_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__949_ : 1'b0;
  assign n_4_net__948_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__948_ : 1'b0;
  assign n_4_net__947_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__947_ : 1'b0;
  assign n_4_net__946_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__946_ : 1'b0;
  assign n_4_net__945_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__945_ : 1'b0;
  assign n_4_net__944_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__944_ : 1'b0;
  assign n_4_net__943_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__943_ : 1'b0;
  assign n_4_net__942_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__942_ : 1'b0;
  assign n_4_net__941_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__941_ : 1'b0;
  assign n_4_net__940_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__940_ : 1'b0;
  assign n_4_net__939_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__939_ : 1'b0;
  assign n_4_net__938_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__938_ : 1'b0;
  assign n_4_net__937_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__937_ : 1'b0;
  assign n_4_net__936_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__936_ : 1'b0;
  assign n_4_net__935_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__935_ : 1'b0;
  assign n_4_net__934_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__934_ : 1'b0;
  assign n_4_net__933_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__933_ : 1'b0;
  assign n_4_net__932_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__932_ : 1'b0;
  assign n_4_net__931_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__931_ : 1'b0;
  assign n_4_net__930_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__930_ : 1'b0;
  assign n_4_net__929_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__929_ : 1'b0;
  assign n_4_net__928_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__928_ : 1'b0;
  assign n_4_net__927_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__927_ : 1'b0;
  assign n_4_net__926_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__926_ : 1'b0;
  assign n_4_net__925_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__925_ : 1'b0;
  assign n_4_net__924_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__924_ : 1'b0;
  assign n_4_net__923_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__923_ : 1'b0;
  assign n_4_net__922_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__922_ : 1'b0;
  assign n_4_net__921_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__921_ : 1'b0;
  assign n_4_net__920_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__920_ : 1'b0;
  assign n_4_net__919_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__919_ : 1'b0;
  assign n_4_net__918_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__918_ : 1'b0;
  assign n_4_net__917_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__917_ : 1'b0;
  assign n_4_net__916_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__916_ : 1'b0;
  assign n_4_net__915_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__915_ : 1'b0;
  assign n_4_net__914_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__914_ : 1'b0;
  assign n_4_net__913_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__913_ : 1'b0;
  assign n_4_net__912_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__912_ : 1'b0;
  assign n_4_net__911_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__911_ : 1'b0;
  assign n_4_net__910_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__910_ : 1'b0;
  assign n_4_net__909_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__909_ : 1'b0;
  assign n_4_net__908_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__908_ : 1'b0;
  assign n_4_net__907_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__907_ : 1'b0;
  assign n_4_net__906_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__906_ : 1'b0;
  assign n_4_net__905_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__905_ : 1'b0;
  assign n_4_net__904_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__904_ : 1'b0;
  assign n_4_net__903_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__903_ : 1'b0;
  assign n_4_net__902_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__902_ : 1'b0;
  assign n_4_net__901_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__901_ : 1'b0;
  assign n_4_net__900_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__900_ : 1'b0;
  assign n_4_net__899_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__899_ : 1'b0;
  assign n_4_net__898_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__898_ : 1'b0;
  assign n_4_net__897_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__897_ : 1'b0;
  assign n_4_net__896_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__896_ : 1'b0;
  assign n_4_net__895_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__895_ : 1'b0;
  assign n_4_net__894_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__894_ : 1'b0;
  assign n_4_net__893_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__893_ : 1'b0;
  assign n_4_net__892_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__892_ : 1'b0;
  assign n_4_net__891_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__891_ : 1'b0;
  assign n_4_net__890_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__890_ : 1'b0;
  assign n_4_net__889_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__889_ : 1'b0;
  assign n_4_net__888_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__888_ : 1'b0;
  assign n_4_net__887_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__887_ : 1'b0;
  assign n_4_net__886_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__886_ : 1'b0;
  assign n_4_net__885_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__885_ : 1'b0;
  assign n_4_net__884_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__884_ : 1'b0;
  assign n_4_net__883_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__883_ : 1'b0;
  assign n_4_net__882_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__882_ : 1'b0;
  assign n_4_net__881_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__881_ : 1'b0;
  assign n_4_net__880_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__880_ : 1'b0;
  assign n_4_net__879_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__879_ : 1'b0;
  assign n_4_net__878_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__878_ : 1'b0;
  assign n_4_net__877_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__877_ : 1'b0;
  assign n_4_net__876_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__876_ : 1'b0;
  assign n_4_net__875_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__875_ : 1'b0;
  assign n_4_net__874_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__874_ : 1'b0;
  assign n_4_net__873_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__873_ : 1'b0;
  assign n_4_net__872_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__872_ : 1'b0;
  assign n_4_net__871_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__871_ : 1'b0;
  assign n_4_net__870_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__870_ : 1'b0;
  assign n_4_net__869_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__869_ : 1'b0;
  assign n_4_net__868_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__868_ : 1'b0;
  assign n_4_net__867_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__867_ : 1'b0;
  assign n_4_net__866_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__866_ : 1'b0;
  assign n_4_net__865_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__865_ : 1'b0;
  assign n_4_net__864_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__864_ : 1'b0;
  assign n_4_net__863_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__863_ : 1'b0;
  assign n_4_net__862_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__862_ : 1'b0;
  assign n_4_net__861_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__861_ : 1'b0;
  assign n_4_net__860_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__860_ : 1'b0;
  assign n_4_net__859_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__859_ : 1'b0;
  assign n_4_net__858_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__858_ : 1'b0;
  assign n_4_net__857_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__857_ : 1'b0;
  assign n_4_net__856_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__856_ : 1'b0;
  assign n_4_net__855_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__855_ : 1'b0;
  assign n_4_net__854_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__854_ : 1'b0;
  assign n_4_net__853_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__853_ : 1'b0;
  assign n_4_net__852_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__852_ : 1'b0;
  assign n_4_net__851_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__851_ : 1'b0;
  assign n_4_net__850_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__850_ : 1'b0;
  assign n_4_net__849_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__849_ : 1'b0;
  assign n_4_net__848_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__848_ : 1'b0;
  assign n_4_net__847_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__847_ : 1'b0;
  assign n_4_net__846_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__846_ : 1'b0;
  assign n_4_net__845_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__845_ : 1'b0;
  assign n_4_net__844_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__844_ : 1'b0;
  assign n_4_net__843_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__843_ : 1'b0;
  assign n_4_net__842_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__842_ : 1'b0;
  assign n_4_net__841_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__841_ : 1'b0;
  assign n_4_net__840_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__840_ : 1'b0;
  assign n_4_net__839_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__839_ : 1'b0;
  assign n_4_net__838_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__838_ : 1'b0;
  assign n_4_net__837_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__837_ : 1'b0;
  assign n_4_net__836_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__836_ : 1'b0;
  assign n_4_net__835_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__835_ : 1'b0;
  assign n_4_net__834_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__834_ : 1'b0;
  assign n_4_net__833_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__833_ : 1'b0;
  assign n_4_net__832_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__832_ : 1'b0;
  assign n_4_net__831_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__831_ : 1'b0;
  assign n_4_net__830_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__830_ : 1'b0;
  assign n_4_net__829_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__829_ : 1'b0;
  assign n_4_net__828_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__828_ : 1'b0;
  assign n_4_net__827_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__827_ : 1'b0;
  assign n_4_net__826_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__826_ : 1'b0;
  assign n_4_net__825_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__825_ : 1'b0;
  assign n_4_net__824_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__824_ : 1'b0;
  assign n_4_net__823_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__823_ : 1'b0;
  assign n_4_net__822_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__822_ : 1'b0;
  assign n_4_net__821_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__821_ : 1'b0;
  assign n_4_net__820_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__820_ : 1'b0;
  assign n_4_net__819_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__819_ : 1'b0;
  assign n_4_net__818_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__818_ : 1'b0;
  assign n_4_net__817_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__817_ : 1'b0;
  assign n_4_net__816_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__816_ : 1'b0;
  assign n_4_net__815_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__815_ : 1'b0;
  assign n_4_net__814_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__814_ : 1'b0;
  assign n_4_net__813_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__813_ : 1'b0;
  assign n_4_net__812_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__812_ : 1'b0;
  assign n_4_net__811_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__811_ : 1'b0;
  assign n_4_net__810_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__810_ : 1'b0;
  assign n_4_net__809_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__809_ : 1'b0;
  assign n_4_net__808_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__808_ : 1'b0;
  assign n_4_net__807_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__807_ : 1'b0;
  assign n_4_net__806_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__806_ : 1'b0;
  assign n_4_net__805_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__805_ : 1'b0;
  assign n_4_net__804_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__804_ : 1'b0;
  assign n_4_net__803_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__803_ : 1'b0;
  assign n_4_net__802_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__802_ : 1'b0;
  assign n_4_net__801_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__801_ : 1'b0;
  assign n_4_net__800_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__800_ : 1'b0;
  assign n_4_net__799_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__799_ : 1'b0;
  assign n_4_net__798_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__798_ : 1'b0;
  assign n_4_net__797_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__797_ : 1'b0;
  assign n_4_net__796_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__796_ : 1'b0;
  assign n_4_net__795_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__795_ : 1'b0;
  assign n_4_net__794_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__794_ : 1'b0;
  assign n_4_net__793_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__793_ : 1'b0;
  assign n_4_net__792_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__792_ : 1'b0;
  assign n_4_net__791_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__791_ : 1'b0;
  assign n_4_net__790_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__790_ : 1'b0;
  assign n_4_net__789_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__789_ : 1'b0;
  assign n_4_net__788_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__788_ : 1'b0;
  assign n_4_net__787_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__787_ : 1'b0;
  assign n_4_net__786_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__786_ : 1'b0;
  assign n_4_net__785_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__785_ : 1'b0;
  assign n_4_net__784_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__784_ : 1'b0;
  assign n_4_net__783_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__783_ : 1'b0;
  assign n_4_net__782_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__782_ : 1'b0;
  assign n_4_net__781_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__781_ : 1'b0;
  assign n_4_net__780_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__780_ : 1'b0;
  assign n_4_net__779_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__779_ : 1'b0;
  assign n_4_net__778_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__778_ : 1'b0;
  assign n_4_net__777_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__777_ : 1'b0;
  assign n_4_net__776_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__776_ : 1'b0;
  assign n_4_net__775_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__775_ : 1'b0;
  assign n_4_net__774_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__774_ : 1'b0;
  assign n_4_net__773_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__773_ : 1'b0;
  assign n_4_net__772_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__772_ : 1'b0;
  assign n_4_net__771_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__771_ : 1'b0;
  assign n_4_net__770_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__770_ : 1'b0;
  assign n_4_net__769_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__769_ : 1'b0;
  assign n_4_net__768_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__768_ : 1'b0;
  assign n_4_net__767_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__767_ : 1'b0;
  assign n_4_net__766_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__766_ : 1'b0;
  assign n_4_net__765_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__765_ : 1'b0;
  assign n_4_net__764_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__764_ : 1'b0;
  assign n_4_net__763_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__763_ : 1'b0;
  assign n_4_net__762_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__762_ : 1'b0;
  assign n_4_net__761_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__761_ : 1'b0;
  assign n_4_net__760_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__760_ : 1'b0;
  assign n_4_net__759_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__759_ : 1'b0;
  assign n_4_net__758_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__758_ : 1'b0;
  assign n_4_net__757_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__757_ : 1'b0;
  assign n_4_net__756_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__756_ : 1'b0;
  assign n_4_net__755_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__755_ : 1'b0;
  assign n_4_net__754_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__754_ : 1'b0;
  assign n_4_net__753_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__753_ : 1'b0;
  assign n_4_net__752_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__752_ : 1'b0;
  assign n_4_net__751_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__751_ : 1'b0;
  assign n_4_net__750_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__750_ : 1'b0;
  assign n_4_net__749_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__749_ : 1'b0;
  assign n_4_net__748_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__748_ : 1'b0;
  assign n_4_net__747_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__747_ : 1'b0;
  assign n_4_net__746_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__746_ : 1'b0;
  assign n_4_net__745_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__745_ : 1'b0;
  assign n_4_net__744_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__744_ : 1'b0;
  assign n_4_net__743_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__743_ : 1'b0;
  assign n_4_net__742_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__742_ : 1'b0;
  assign n_4_net__741_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__741_ : 1'b0;
  assign n_4_net__740_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__740_ : 1'b0;
  assign n_4_net__739_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__739_ : 1'b0;
  assign n_4_net__738_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__738_ : 1'b0;
  assign n_4_net__737_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__737_ : 1'b0;
  assign n_4_net__736_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__736_ : 1'b0;
  assign n_4_net__735_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__735_ : 1'b0;
  assign n_4_net__734_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__734_ : 1'b0;
  assign n_4_net__733_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__733_ : 1'b0;
  assign n_4_net__732_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__732_ : 1'b0;
  assign n_4_net__731_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__731_ : 1'b0;
  assign n_4_net__730_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__730_ : 1'b0;
  assign n_4_net__729_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__729_ : 1'b0;
  assign n_4_net__728_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__728_ : 1'b0;
  assign n_4_net__727_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__727_ : 1'b0;
  assign n_4_net__726_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__726_ : 1'b0;
  assign n_4_net__725_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__725_ : 1'b0;
  assign n_4_net__724_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__724_ : 1'b0;
  assign n_4_net__723_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__723_ : 1'b0;
  assign n_4_net__722_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__722_ : 1'b0;
  assign n_4_net__721_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__721_ : 1'b0;
  assign n_4_net__720_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__720_ : 1'b0;
  assign n_4_net__719_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__719_ : 1'b0;
  assign n_4_net__718_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__718_ : 1'b0;
  assign n_4_net__717_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__717_ : 1'b0;
  assign n_4_net__716_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__716_ : 1'b0;
  assign n_4_net__715_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__715_ : 1'b0;
  assign n_4_net__714_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__714_ : 1'b0;
  assign n_4_net__713_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__713_ : 1'b0;
  assign n_4_net__712_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__712_ : 1'b0;
  assign n_4_net__711_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__711_ : 1'b0;
  assign n_4_net__710_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__710_ : 1'b0;
  assign n_4_net__709_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__709_ : 1'b0;
  assign n_4_net__708_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__708_ : 1'b0;
  assign n_4_net__707_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__707_ : 1'b0;
  assign n_4_net__706_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__706_ : 1'b0;
  assign n_4_net__705_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__705_ : 1'b0;
  assign n_4_net__704_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__704_ : 1'b0;
  assign n_4_net__703_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__703_ : 1'b0;
  assign n_4_net__702_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__702_ : 1'b0;
  assign n_4_net__701_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__701_ : 1'b0;
  assign n_4_net__700_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__700_ : 1'b0;
  assign n_4_net__699_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__699_ : 1'b0;
  assign n_4_net__698_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__698_ : 1'b0;
  assign n_4_net__697_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__697_ : 1'b0;
  assign n_4_net__696_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__696_ : 1'b0;
  assign n_4_net__695_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__695_ : 1'b0;
  assign n_4_net__694_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__694_ : 1'b0;
  assign n_4_net__693_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__693_ : 1'b0;
  assign n_4_net__692_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__692_ : 1'b0;
  assign n_4_net__691_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__691_ : 1'b0;
  assign n_4_net__690_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__690_ : 1'b0;
  assign n_4_net__689_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__689_ : 1'b0;
  assign n_4_net__688_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__688_ : 1'b0;
  assign n_4_net__687_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__687_ : 1'b0;
  assign n_4_net__686_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__686_ : 1'b0;
  assign n_4_net__685_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__685_ : 1'b0;
  assign n_4_net__684_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__684_ : 1'b0;
  assign n_4_net__683_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__683_ : 1'b0;
  assign n_4_net__682_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__682_ : 1'b0;
  assign n_4_net__681_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__681_ : 1'b0;
  assign n_4_net__680_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__680_ : 1'b0;
  assign n_4_net__679_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__679_ : 1'b0;
  assign n_4_net__678_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__678_ : 1'b0;
  assign n_4_net__677_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__677_ : 1'b0;
  assign n_4_net__676_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__676_ : 1'b0;
  assign n_4_net__675_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__675_ : 1'b0;
  assign n_4_net__674_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__674_ : 1'b0;
  assign n_4_net__673_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__673_ : 1'b0;
  assign n_4_net__672_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__672_ : 1'b0;
  assign n_4_net__671_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__671_ : 1'b0;
  assign n_4_net__670_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__670_ : 1'b0;
  assign n_4_net__669_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__669_ : 1'b0;
  assign n_4_net__668_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__668_ : 1'b0;
  assign n_4_net__667_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__667_ : 1'b0;
  assign n_4_net__666_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__666_ : 1'b0;
  assign n_4_net__665_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__665_ : 1'b0;
  assign n_4_net__664_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__664_ : 1'b0;
  assign n_4_net__663_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__663_ : 1'b0;
  assign n_4_net__662_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__662_ : 1'b0;
  assign n_4_net__661_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__661_ : 1'b0;
  assign n_4_net__660_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__660_ : 1'b0;
  assign n_4_net__659_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__659_ : 1'b0;
  assign n_4_net__658_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__658_ : 1'b0;
  assign n_4_net__657_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__657_ : 1'b0;
  assign n_4_net__656_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__656_ : 1'b0;
  assign n_4_net__655_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__655_ : 1'b0;
  assign n_4_net__654_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__654_ : 1'b0;
  assign n_4_net__653_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__653_ : 1'b0;
  assign n_4_net__652_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__652_ : 1'b0;
  assign n_4_net__651_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__651_ : 1'b0;
  assign n_4_net__650_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__650_ : 1'b0;
  assign n_4_net__649_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__649_ : 1'b0;
  assign n_4_net__648_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__648_ : 1'b0;
  assign n_4_net__647_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__647_ : 1'b0;
  assign n_4_net__646_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__646_ : 1'b0;
  assign n_4_net__645_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__645_ : 1'b0;
  assign n_4_net__644_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__644_ : 1'b0;
  assign n_4_net__643_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__643_ : 1'b0;
  assign n_4_net__642_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__642_ : 1'b0;
  assign n_4_net__641_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__641_ : 1'b0;
  assign n_4_net__640_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__640_ : 1'b0;
  assign n_4_net__639_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__639_ : 1'b0;
  assign n_4_net__638_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__638_ : 1'b0;
  assign n_4_net__637_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__637_ : 1'b0;
  assign n_4_net__636_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__636_ : 1'b0;
  assign n_4_net__635_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__635_ : 1'b0;
  assign n_4_net__634_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__634_ : 1'b0;
  assign n_4_net__633_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__633_ : 1'b0;
  assign n_4_net__632_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__632_ : 1'b0;
  assign n_4_net__631_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__631_ : 1'b0;
  assign n_4_net__630_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__630_ : 1'b0;
  assign n_4_net__629_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__629_ : 1'b0;
  assign n_4_net__628_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__628_ : 1'b0;
  assign n_4_net__627_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__627_ : 1'b0;
  assign n_4_net__626_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__626_ : 1'b0;
  assign n_4_net__625_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__625_ : 1'b0;
  assign n_4_net__624_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__624_ : 1'b0;
  assign n_4_net__623_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__623_ : 1'b0;
  assign n_4_net__622_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__622_ : 1'b0;
  assign n_4_net__621_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__621_ : 1'b0;
  assign n_4_net__620_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__620_ : 1'b0;
  assign n_4_net__619_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__619_ : 1'b0;
  assign n_4_net__618_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__618_ : 1'b0;
  assign n_4_net__617_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__617_ : 1'b0;
  assign n_4_net__616_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__616_ : 1'b0;
  assign n_4_net__615_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__615_ : 1'b0;
  assign n_4_net__614_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__614_ : 1'b0;
  assign n_4_net__613_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__613_ : 1'b0;
  assign n_4_net__612_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__612_ : 1'b0;
  assign n_4_net__611_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__611_ : 1'b0;
  assign n_4_net__610_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__610_ : 1'b0;
  assign n_4_net__609_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__609_ : 1'b0;
  assign n_4_net__608_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__608_ : 1'b0;
  assign n_4_net__607_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__607_ : 1'b0;
  assign n_4_net__606_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__606_ : 1'b0;
  assign n_4_net__605_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__605_ : 1'b0;
  assign n_4_net__604_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__604_ : 1'b0;
  assign n_4_net__603_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__603_ : 1'b0;
  assign n_4_net__602_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__602_ : 1'b0;
  assign n_4_net__601_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__601_ : 1'b0;
  assign n_4_net__600_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__600_ : 1'b0;
  assign n_4_net__599_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__599_ : 1'b0;
  assign n_4_net__598_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__598_ : 1'b0;
  assign n_4_net__597_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__597_ : 1'b0;
  assign n_4_net__596_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__596_ : 1'b0;
  assign n_4_net__595_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__595_ : 1'b0;
  assign n_4_net__594_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__594_ : 1'b0;
  assign n_4_net__593_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__593_ : 1'b0;
  assign n_4_net__592_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__592_ : 1'b0;
  assign n_4_net__591_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__591_ : 1'b0;
  assign n_4_net__590_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__590_ : 1'b0;
  assign n_4_net__589_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__589_ : 1'b0;
  assign n_4_net__588_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__588_ : 1'b0;
  assign n_4_net__587_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__587_ : 1'b0;
  assign n_4_net__586_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__586_ : 1'b0;
  assign n_4_net__585_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__585_ : 1'b0;
  assign n_4_net__584_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__584_ : 1'b0;
  assign n_4_net__583_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__583_ : 1'b0;
  assign n_4_net__582_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__582_ : 1'b0;
  assign n_4_net__581_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__581_ : 1'b0;
  assign n_4_net__580_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__580_ : 1'b0;
  assign n_4_net__579_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__579_ : 1'b0;
  assign n_4_net__578_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__578_ : 1'b0;
  assign n_4_net__577_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__577_ : 1'b0;
  assign n_4_net__576_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__576_ : 1'b0;
  assign n_4_net__575_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__575_ : 1'b0;
  assign n_4_net__574_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__574_ : 1'b0;
  assign n_4_net__573_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__573_ : 1'b0;
  assign n_4_net__572_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__572_ : 1'b0;
  assign n_4_net__571_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__571_ : 1'b0;
  assign n_4_net__570_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__570_ : 1'b0;
  assign n_4_net__569_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__569_ : 1'b0;
  assign n_4_net__568_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__568_ : 1'b0;
  assign n_4_net__567_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__567_ : 1'b0;
  assign n_4_net__566_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__566_ : 1'b0;
  assign n_4_net__565_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__565_ : 1'b0;
  assign n_4_net__564_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__564_ : 1'b0;
  assign n_4_net__563_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__563_ : 1'b0;
  assign n_4_net__562_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__562_ : 1'b0;
  assign n_4_net__561_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__561_ : 1'b0;
  assign n_4_net__560_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__560_ : 1'b0;
  assign n_4_net__559_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__559_ : 1'b0;
  assign n_4_net__558_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__558_ : 1'b0;
  assign n_4_net__557_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__557_ : 1'b0;
  assign n_4_net__556_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__556_ : 1'b0;
  assign n_4_net__555_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__555_ : 1'b0;
  assign n_4_net__554_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__554_ : 1'b0;
  assign n_4_net__553_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__553_ : 1'b0;
  assign n_4_net__552_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__552_ : 1'b0;
  assign n_4_net__551_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__551_ : 1'b0;
  assign n_4_net__550_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__550_ : 1'b0;
  assign n_4_net__549_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__549_ : 1'b0;
  assign n_4_net__548_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__548_ : 1'b0;
  assign n_4_net__547_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__547_ : 1'b0;
  assign n_4_net__546_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__546_ : 1'b0;
  assign n_4_net__545_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__545_ : 1'b0;
  assign n_4_net__544_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__544_ : 1'b0;
  assign n_4_net__543_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__543_ : 1'b0;
  assign n_4_net__542_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__542_ : 1'b0;
  assign n_4_net__541_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__541_ : 1'b0;
  assign n_4_net__540_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__540_ : 1'b0;
  assign n_4_net__539_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__539_ : 1'b0;
  assign n_4_net__538_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__538_ : 1'b0;
  assign n_4_net__537_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__537_ : 1'b0;
  assign n_4_net__536_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__536_ : 1'b0;
  assign n_4_net__535_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__535_ : 1'b0;
  assign n_4_net__534_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__534_ : 1'b0;
  assign n_4_net__533_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__533_ : 1'b0;
  assign n_4_net__532_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__532_ : 1'b0;
  assign n_4_net__531_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__531_ : 1'b0;
  assign n_4_net__530_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__530_ : 1'b0;
  assign n_4_net__529_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__529_ : 1'b0;
  assign n_4_net__528_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__528_ : 1'b0;
  assign n_4_net__527_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__527_ : 1'b0;
  assign n_4_net__526_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__526_ : 1'b0;
  assign n_4_net__525_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__525_ : 1'b0;
  assign n_4_net__524_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__524_ : 1'b0;
  assign n_4_net__523_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__523_ : 1'b0;
  assign n_4_net__522_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__522_ : 1'b0;
  assign n_4_net__521_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__521_ : 1'b0;
  assign n_4_net__520_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__520_ : 1'b0;
  assign n_4_net__519_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__519_ : 1'b0;
  assign n_4_net__518_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__518_ : 1'b0;
  assign n_4_net__517_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__517_ : 1'b0;
  assign n_4_net__516_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__516_ : 1'b0;
  assign n_4_net__515_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__515_ : 1'b0;
  assign n_4_net__514_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__514_ : 1'b0;
  assign n_4_net__513_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__513_ : 1'b0;
  assign n_4_net__512_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__512_ : 1'b0;
  assign n_4_net__511_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__511_ : 1'b0;
  assign n_4_net__510_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__510_ : 1'b0;
  assign n_4_net__509_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__509_ : 1'b0;
  assign n_4_net__508_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__508_ : 1'b0;
  assign n_4_net__507_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__507_ : 1'b0;
  assign n_4_net__506_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__506_ : 1'b0;
  assign n_4_net__505_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__505_ : 1'b0;
  assign n_4_net__504_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__504_ : 1'b0;
  assign n_4_net__503_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__503_ : 1'b0;
  assign n_4_net__502_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__502_ : 1'b0;
  assign n_4_net__501_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__501_ : 1'b0;
  assign n_4_net__500_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__500_ : 1'b0;
  assign n_4_net__499_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__499_ : 1'b0;
  assign n_4_net__498_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__498_ : 1'b0;
  assign n_4_net__497_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__497_ : 1'b0;
  assign n_4_net__496_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__496_ : 1'b0;
  assign n_4_net__495_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__495_ : 1'b0;
  assign n_4_net__494_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__494_ : 1'b0;
  assign n_4_net__493_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__493_ : 1'b0;
  assign n_4_net__492_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__492_ : 1'b0;
  assign n_4_net__491_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__491_ : 1'b0;
  assign n_4_net__490_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__490_ : 1'b0;
  assign n_4_net__489_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__489_ : 1'b0;
  assign n_4_net__488_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__488_ : 1'b0;
  assign n_4_net__487_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__487_ : 1'b0;
  assign n_4_net__486_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__486_ : 1'b0;
  assign n_4_net__485_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__485_ : 1'b0;
  assign n_4_net__484_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__484_ : 1'b0;
  assign n_4_net__483_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__483_ : 1'b0;
  assign n_4_net__482_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__482_ : 1'b0;
  assign n_4_net__481_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__481_ : 1'b0;
  assign n_4_net__480_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__480_ : 1'b0;
  assign n_4_net__479_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__479_ : 1'b0;
  assign n_4_net__478_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__478_ : 1'b0;
  assign n_4_net__477_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__477_ : 1'b0;
  assign n_4_net__476_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__476_ : 1'b0;
  assign n_4_net__475_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__475_ : 1'b0;
  assign n_4_net__474_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__474_ : 1'b0;
  assign n_4_net__473_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__473_ : 1'b0;
  assign n_4_net__472_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__472_ : 1'b0;
  assign n_4_net__471_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__471_ : 1'b0;
  assign n_4_net__470_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__470_ : 1'b0;
  assign n_4_net__469_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__469_ : 1'b0;
  assign n_4_net__468_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__468_ : 1'b0;
  assign n_4_net__467_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__467_ : 1'b0;
  assign n_4_net__466_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__466_ : 1'b0;
  assign n_4_net__465_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__465_ : 1'b0;
  assign n_4_net__464_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__464_ : 1'b0;
  assign n_4_net__463_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__463_ : 1'b0;
  assign n_4_net__462_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__462_ : 1'b0;
  assign n_4_net__461_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__461_ : 1'b0;
  assign n_4_net__460_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__460_ : 1'b0;
  assign n_4_net__459_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__459_ : 1'b0;
  assign n_4_net__458_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__458_ : 1'b0;
  assign n_4_net__457_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__457_ : 1'b0;
  assign n_4_net__456_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__456_ : 1'b0;
  assign n_4_net__455_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__455_ : 1'b0;
  assign n_4_net__454_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__454_ : 1'b0;
  assign n_4_net__453_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__453_ : 1'b0;
  assign n_4_net__452_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__452_ : 1'b0;
  assign n_4_net__451_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__451_ : 1'b0;
  assign n_4_net__450_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__450_ : 1'b0;
  assign n_4_net__449_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__449_ : 1'b0;
  assign n_4_net__448_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__448_ : 1'b0;
  assign n_4_net__447_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__447_ : 1'b0;
  assign n_4_net__446_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__446_ : 1'b0;
  assign n_4_net__445_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__445_ : 1'b0;
  assign n_4_net__444_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__444_ : 1'b0;
  assign n_4_net__443_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__443_ : 1'b0;
  assign n_4_net__442_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__442_ : 1'b0;
  assign n_4_net__441_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__441_ : 1'b0;
  assign n_4_net__440_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__440_ : 1'b0;
  assign n_4_net__439_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__439_ : 1'b0;
  assign n_4_net__438_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__438_ : 1'b0;
  assign n_4_net__437_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__437_ : 1'b0;
  assign n_4_net__436_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__436_ : 1'b0;
  assign n_4_net__435_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__435_ : 1'b0;
  assign n_4_net__434_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__434_ : 1'b0;
  assign n_4_net__433_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__433_ : 1'b0;
  assign n_4_net__432_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__432_ : 1'b0;
  assign n_4_net__431_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__431_ : 1'b0;
  assign n_4_net__430_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__430_ : 1'b0;
  assign n_4_net__429_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__429_ : 1'b0;
  assign n_4_net__428_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__428_ : 1'b0;
  assign n_4_net__427_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__427_ : 1'b0;
  assign n_4_net__426_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__426_ : 1'b0;
  assign n_4_net__425_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__425_ : 1'b0;
  assign n_4_net__424_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__424_ : 1'b0;
  assign n_4_net__423_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__423_ : 1'b0;
  assign n_4_net__422_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__422_ : 1'b0;
  assign n_4_net__421_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__421_ : 1'b0;
  assign n_4_net__420_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__420_ : 1'b0;
  assign n_4_net__419_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__419_ : 1'b0;
  assign n_4_net__418_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__418_ : 1'b0;
  assign n_4_net__417_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__417_ : 1'b0;
  assign n_4_net__416_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__416_ : 1'b0;
  assign n_4_net__415_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__415_ : 1'b0;
  assign n_4_net__414_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__414_ : 1'b0;
  assign n_4_net__413_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__413_ : 1'b0;
  assign n_4_net__412_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__412_ : 1'b0;
  assign n_4_net__411_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__411_ : 1'b0;
  assign n_4_net__410_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__410_ : 1'b0;
  assign n_4_net__409_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__409_ : 1'b0;
  assign n_4_net__408_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__408_ : 1'b0;
  assign n_4_net__407_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__407_ : 1'b0;
  assign n_4_net__406_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__406_ : 1'b0;
  assign n_4_net__405_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__405_ : 1'b0;
  assign n_4_net__404_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__404_ : 1'b0;
  assign n_4_net__403_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__403_ : 1'b0;
  assign n_4_net__402_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__402_ : 1'b0;
  assign n_4_net__401_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__401_ : 1'b0;
  assign n_4_net__400_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__400_ : 1'b0;
  assign n_4_net__399_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__399_ : 1'b0;
  assign n_4_net__398_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__398_ : 1'b0;
  assign n_4_net__397_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__397_ : 1'b0;
  assign n_4_net__396_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__396_ : 1'b0;
  assign n_4_net__395_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__395_ : 1'b0;
  assign n_4_net__394_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__394_ : 1'b0;
  assign n_4_net__393_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__393_ : 1'b0;
  assign n_4_net__392_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__392_ : 1'b0;
  assign n_4_net__391_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__391_ : 1'b0;
  assign n_4_net__390_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__390_ : 1'b0;
  assign n_4_net__389_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__389_ : 1'b0;
  assign n_4_net__388_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__388_ : 1'b0;
  assign n_4_net__387_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__387_ : 1'b0;
  assign n_4_net__386_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__386_ : 1'b0;
  assign n_4_net__385_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__385_ : 1'b0;
  assign n_4_net__384_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__384_ : 1'b0;
  assign n_4_net__383_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__383_ : 1'b0;
  assign n_4_net__382_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__382_ : 1'b0;
  assign n_4_net__381_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__381_ : 1'b0;
  assign n_4_net__380_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__380_ : 1'b0;
  assign n_4_net__379_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__379_ : 1'b0;
  assign n_4_net__378_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__378_ : 1'b0;
  assign n_4_net__377_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__377_ : 1'b0;
  assign n_4_net__376_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__376_ : 1'b0;
  assign n_4_net__375_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__375_ : 1'b0;
  assign n_4_net__374_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__374_ : 1'b0;
  assign n_4_net__373_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__373_ : 1'b0;
  assign n_4_net__372_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__372_ : 1'b0;
  assign n_4_net__371_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__371_ : 1'b0;
  assign n_4_net__370_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__370_ : 1'b0;
  assign n_4_net__369_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__369_ : 1'b0;
  assign n_4_net__368_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__368_ : 1'b0;
  assign n_4_net__367_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__367_ : 1'b0;
  assign n_4_net__366_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__366_ : 1'b0;
  assign n_4_net__365_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__365_ : 1'b0;
  assign n_4_net__364_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__364_ : 1'b0;
  assign n_4_net__363_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__363_ : 1'b0;
  assign n_4_net__362_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__362_ : 1'b0;
  assign n_4_net__361_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__361_ : 1'b0;
  assign n_4_net__360_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__360_ : 1'b0;
  assign n_4_net__359_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__359_ : 1'b0;
  assign n_4_net__358_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__358_ : 1'b0;
  assign n_4_net__357_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__357_ : 1'b0;
  assign n_4_net__356_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__356_ : 1'b0;
  assign n_4_net__355_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__355_ : 1'b0;
  assign n_4_net__354_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__354_ : 1'b0;
  assign n_4_net__353_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__353_ : 1'b0;
  assign n_4_net__352_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__352_ : 1'b0;
  assign n_4_net__351_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__351_ : 1'b0;
  assign n_4_net__350_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__350_ : 1'b0;
  assign n_4_net__349_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__349_ : 1'b0;
  assign n_4_net__348_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__348_ : 1'b0;
  assign n_4_net__347_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__347_ : 1'b0;
  assign n_4_net__346_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__346_ : 1'b0;
  assign n_4_net__345_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__345_ : 1'b0;
  assign n_4_net__344_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__344_ : 1'b0;
  assign n_4_net__343_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__343_ : 1'b0;
  assign n_4_net__342_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__342_ : 1'b0;
  assign n_4_net__341_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__341_ : 1'b0;
  assign n_4_net__340_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__340_ : 1'b0;
  assign n_4_net__339_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__339_ : 1'b0;
  assign n_4_net__338_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__338_ : 1'b0;
  assign n_4_net__337_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__337_ : 1'b0;
  assign n_4_net__336_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__336_ : 1'b0;
  assign n_4_net__335_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__335_ : 1'b0;
  assign n_4_net__334_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__334_ : 1'b0;
  assign n_4_net__333_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__333_ : 1'b0;
  assign n_4_net__332_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__332_ : 1'b0;
  assign n_4_net__331_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__331_ : 1'b0;
  assign n_4_net__330_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__330_ : 1'b0;
  assign n_4_net__329_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__329_ : 1'b0;
  assign n_4_net__328_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__328_ : 1'b0;
  assign n_4_net__327_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__327_ : 1'b0;
  assign n_4_net__326_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__326_ : 1'b0;
  assign n_4_net__325_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__325_ : 1'b0;
  assign n_4_net__324_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__324_ : 1'b0;
  assign n_4_net__323_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__323_ : 1'b0;
  assign n_4_net__322_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__322_ : 1'b0;
  assign n_4_net__321_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__321_ : 1'b0;
  assign n_4_net__320_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__320_ : 1'b0;
  assign n_4_net__319_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__319_ : 1'b0;
  assign n_4_net__318_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__318_ : 1'b0;
  assign n_4_net__317_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__317_ : 1'b0;
  assign n_4_net__316_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__316_ : 1'b0;
  assign n_4_net__315_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__315_ : 1'b0;
  assign n_4_net__314_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__314_ : 1'b0;
  assign n_4_net__313_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__313_ : 1'b0;
  assign n_4_net__312_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__312_ : 1'b0;
  assign n_4_net__311_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__311_ : 1'b0;
  assign n_4_net__310_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__310_ : 1'b0;
  assign n_4_net__309_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__309_ : 1'b0;
  assign n_4_net__308_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__308_ : 1'b0;
  assign n_4_net__307_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__307_ : 1'b0;
  assign n_4_net__306_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__306_ : 1'b0;
  assign n_4_net__305_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__305_ : 1'b0;
  assign n_4_net__304_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__304_ : 1'b0;
  assign n_4_net__303_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__303_ : 1'b0;
  assign n_4_net__302_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__302_ : 1'b0;
  assign n_4_net__301_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__301_ : 1'b0;
  assign n_4_net__300_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__300_ : 1'b0;
  assign n_4_net__299_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__299_ : 1'b0;
  assign n_4_net__298_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__298_ : 1'b0;
  assign n_4_net__297_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__297_ : 1'b0;
  assign n_4_net__296_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__296_ : 1'b0;
  assign n_4_net__295_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__295_ : 1'b0;
  assign n_4_net__294_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__294_ : 1'b0;
  assign n_4_net__293_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__293_ : 1'b0;
  assign n_4_net__292_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__292_ : 1'b0;
  assign n_4_net__291_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__291_ : 1'b0;
  assign n_4_net__290_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__290_ : 1'b0;
  assign n_4_net__289_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__289_ : 1'b0;
  assign n_4_net__288_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__288_ : 1'b0;
  assign n_4_net__287_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__287_ : 1'b0;
  assign n_4_net__286_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__286_ : 1'b0;
  assign n_4_net__285_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__285_ : 1'b0;
  assign n_4_net__284_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__284_ : 1'b0;
  assign n_4_net__283_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__283_ : 1'b0;
  assign n_4_net__282_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__282_ : 1'b0;
  assign n_4_net__281_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__281_ : 1'b0;
  assign n_4_net__280_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__280_ : 1'b0;
  assign n_4_net__279_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__279_ : 1'b0;
  assign n_4_net__278_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__278_ : 1'b0;
  assign n_4_net__277_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__277_ : 1'b0;
  assign n_4_net__276_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__276_ : 1'b0;
  assign n_4_net__275_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__275_ : 1'b0;
  assign n_4_net__274_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__274_ : 1'b0;
  assign n_4_net__273_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__273_ : 1'b0;
  assign n_4_net__272_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__272_ : 1'b0;
  assign n_4_net__271_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__271_ : 1'b0;
  assign n_4_net__270_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__270_ : 1'b0;
  assign n_4_net__269_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__269_ : 1'b0;
  assign n_4_net__268_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__268_ : 1'b0;
  assign n_4_net__267_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__267_ : 1'b0;
  assign n_4_net__266_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__266_ : 1'b0;
  assign n_4_net__265_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__265_ : 1'b0;
  assign n_4_net__264_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__264_ : 1'b0;
  assign n_4_net__263_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__263_ : 1'b0;
  assign n_4_net__262_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__262_ : 1'b0;
  assign n_4_net__261_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__261_ : 1'b0;
  assign n_4_net__260_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__260_ : 1'b0;
  assign n_4_net__259_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__259_ : 1'b0;
  assign n_4_net__258_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__258_ : 1'b0;
  assign n_4_net__257_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__257_ : 1'b0;
  assign n_4_net__256_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__256_ : 1'b0;
  assign n_4_net__255_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__255_ : 1'b0;
  assign n_4_net__254_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__254_ : 1'b0;
  assign n_4_net__253_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__253_ : 1'b0;
  assign n_4_net__252_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__252_ : 1'b0;
  assign n_4_net__251_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__251_ : 1'b0;
  assign n_4_net__250_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__250_ : 1'b0;
  assign n_4_net__249_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__249_ : 1'b0;
  assign n_4_net__248_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__248_ : 1'b0;
  assign n_4_net__247_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__247_ : 1'b0;
  assign n_4_net__246_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__246_ : 1'b0;
  assign n_4_net__245_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__245_ : 1'b0;
  assign n_4_net__244_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__244_ : 1'b0;
  assign n_4_net__243_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__243_ : 1'b0;
  assign n_4_net__242_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__242_ : 1'b0;
  assign n_4_net__241_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__241_ : 1'b0;
  assign n_4_net__240_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__240_ : 1'b0;
  assign n_4_net__239_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__239_ : 1'b0;
  assign n_4_net__238_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__238_ : 1'b0;
  assign n_4_net__237_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__237_ : 1'b0;
  assign n_4_net__236_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__236_ : 1'b0;
  assign n_4_net__235_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__235_ : 1'b0;
  assign n_4_net__234_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__234_ : 1'b0;
  assign n_4_net__233_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__233_ : 1'b0;
  assign n_4_net__232_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__232_ : 1'b0;
  assign n_4_net__231_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__231_ : 1'b0;
  assign n_4_net__230_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__230_ : 1'b0;
  assign n_4_net__229_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__229_ : 1'b0;
  assign n_4_net__228_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__228_ : 1'b0;
  assign n_4_net__227_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__227_ : 1'b0;
  assign n_4_net__226_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__226_ : 1'b0;
  assign n_4_net__225_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__225_ : 1'b0;
  assign n_4_net__224_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__224_ : 1'b0;
  assign n_4_net__223_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__223_ : 1'b0;
  assign n_4_net__222_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__222_ : 1'b0;
  assign n_4_net__221_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__221_ : 1'b0;
  assign n_4_net__220_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__220_ : 1'b0;
  assign n_4_net__219_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__219_ : 1'b0;
  assign n_4_net__218_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__218_ : 1'b0;
  assign n_4_net__217_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__217_ : 1'b0;
  assign n_4_net__216_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__216_ : 1'b0;
  assign n_4_net__215_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__215_ : 1'b0;
  assign n_4_net__214_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__214_ : 1'b0;
  assign n_4_net__213_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__213_ : 1'b0;
  assign n_4_net__212_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__212_ : 1'b0;
  assign n_4_net__211_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__211_ : 1'b0;
  assign n_4_net__210_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__210_ : 1'b0;
  assign n_4_net__209_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__209_ : 1'b0;
  assign n_4_net__208_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__208_ : 1'b0;
  assign n_4_net__207_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__207_ : 1'b0;
  assign n_4_net__206_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__206_ : 1'b0;
  assign n_4_net__205_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__205_ : 1'b0;
  assign n_4_net__204_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__204_ : 1'b0;
  assign n_4_net__203_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__203_ : 1'b0;
  assign n_4_net__202_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__202_ : 1'b0;
  assign n_4_net__201_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__201_ : 1'b0;
  assign n_4_net__200_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__200_ : 1'b0;
  assign n_4_net__199_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__199_ : 1'b0;
  assign n_4_net__198_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__198_ : 1'b0;
  assign n_4_net__197_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__197_ : 1'b0;
  assign n_4_net__196_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__196_ : 1'b0;
  assign n_4_net__195_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__195_ : 1'b0;
  assign n_4_net__194_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__194_ : 1'b0;
  assign n_4_net__193_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__193_ : 1'b0;
  assign n_4_net__192_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__192_ : 1'b0;
  assign n_4_net__191_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__191_ : 1'b0;
  assign n_4_net__190_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__190_ : 1'b0;
  assign n_4_net__189_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__189_ : 1'b0;
  assign n_4_net__188_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__188_ : 1'b0;
  assign n_4_net__187_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__187_ : 1'b0;
  assign n_4_net__186_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__186_ : 1'b0;
  assign n_4_net__185_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__185_ : 1'b0;
  assign n_4_net__184_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__184_ : 1'b0;
  assign n_4_net__183_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__183_ : 1'b0;
  assign n_4_net__182_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__182_ : 1'b0;
  assign n_4_net__181_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__181_ : 1'b0;
  assign n_4_net__180_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__180_ : 1'b0;
  assign n_4_net__179_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__179_ : 1'b0;
  assign n_4_net__178_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__178_ : 1'b0;
  assign n_4_net__177_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__177_ : 1'b0;
  assign n_4_net__176_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__176_ : 1'b0;
  assign n_4_net__175_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__175_ : 1'b0;
  assign n_4_net__174_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__174_ : 1'b0;
  assign n_4_net__173_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__173_ : 1'b0;
  assign n_4_net__172_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__172_ : 1'b0;
  assign n_4_net__171_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__171_ : 1'b0;
  assign n_4_net__170_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__170_ : 1'b0;
  assign n_4_net__169_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__169_ : 1'b0;
  assign n_4_net__168_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__168_ : 1'b0;
  assign n_4_net__167_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__167_ : 1'b0;
  assign n_4_net__166_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__166_ : 1'b0;
  assign n_4_net__165_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__165_ : 1'b0;
  assign n_4_net__164_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__164_ : 1'b0;
  assign n_4_net__163_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__163_ : 1'b0;
  assign n_4_net__162_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__162_ : 1'b0;
  assign n_4_net__161_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__161_ : 1'b0;
  assign n_4_net__160_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__160_ : 1'b0;
  assign n_4_net__159_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__159_ : 1'b0;
  assign n_4_net__158_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__158_ : 1'b0;
  assign n_4_net__157_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__157_ : 1'b0;
  assign n_4_net__156_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__156_ : 1'b0;
  assign n_4_net__155_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__155_ : 1'b0;
  assign n_4_net__154_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__154_ : 1'b0;
  assign n_4_net__153_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__153_ : 1'b0;
  assign n_4_net__152_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__152_ : 1'b0;
  assign n_4_net__151_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__151_ : 1'b0;
  assign n_4_net__150_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__150_ : 1'b0;
  assign n_4_net__149_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__149_ : 1'b0;
  assign n_4_net__148_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__148_ : 1'b0;
  assign n_4_net__147_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__147_ : 1'b0;
  assign n_4_net__146_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__146_ : 1'b0;
  assign n_4_net__145_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__145_ : 1'b0;
  assign n_4_net__144_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__144_ : 1'b0;
  assign n_4_net__143_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__143_ : 1'b0;
  assign n_4_net__142_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__142_ : 1'b0;
  assign n_4_net__141_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__141_ : 1'b0;
  assign n_4_net__140_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__140_ : 1'b0;
  assign n_4_net__139_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__139_ : 1'b0;
  assign n_4_net__138_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__138_ : 1'b0;
  assign n_4_net__137_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__137_ : 1'b0;
  assign n_4_net__136_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__136_ : 1'b0;
  assign n_4_net__135_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__135_ : 1'b0;
  assign n_4_net__134_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__134_ : 1'b0;
  assign n_4_net__133_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__133_ : 1'b0;
  assign n_4_net__132_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__132_ : 1'b0;
  assign n_4_net__131_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__131_ : 1'b0;
  assign n_4_net__130_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__130_ : 1'b0;
  assign n_4_net__129_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__129_ : 1'b0;
  assign n_4_net__128_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__128_ : 1'b0;
  assign n_4_net__127_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__127_ : 1'b0;
  assign n_4_net__126_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__126_ : 1'b0;
  assign n_4_net__125_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__125_ : 1'b0;
  assign n_4_net__124_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__124_ : 1'b0;
  assign n_4_net__123_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__123_ : 1'b0;
  assign n_4_net__122_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__122_ : 1'b0;
  assign n_4_net__121_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__121_ : 1'b0;
  assign n_4_net__120_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__120_ : 1'b0;
  assign n_4_net__119_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__119_ : 1'b0;
  assign n_4_net__118_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__118_ : 1'b0;
  assign n_4_net__117_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__117_ : 1'b0;
  assign n_4_net__116_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__116_ : 1'b0;
  assign n_4_net__115_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__115_ : 1'b0;
  assign n_4_net__114_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__114_ : 1'b0;
  assign n_4_net__113_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__113_ : 1'b0;
  assign n_4_net__112_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__112_ : 1'b0;
  assign n_4_net__111_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__111_ : 1'b0;
  assign n_4_net__110_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__110_ : 1'b0;
  assign n_4_net__109_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__109_ : 1'b0;
  assign n_4_net__108_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__108_ : 1'b0;
  assign n_4_net__107_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__107_ : 1'b0;
  assign n_4_net__106_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__106_ : 1'b0;
  assign n_4_net__105_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__105_ : 1'b0;
  assign n_4_net__104_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__104_ : 1'b0;
  assign n_4_net__103_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__103_ : 1'b0;
  assign n_4_net__102_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__102_ : 1'b0;
  assign n_4_net__101_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__101_ : 1'b0;
  assign n_4_net__100_ = (N115)? 1'b0 : 
                         (N116)? 1'b0 : 
                         (N117)? 1'b0 : 
                         (N118)? 1'b0 : 
                         (N119)? 1'b0 : 
                         (N120)? 1'b0 : 
                         (N121)? 1'b0 : 
                         (N122)? 1'b0 : 
                         (N123)? 1'b0 : 
                         (N124)? data_head_9__100_ : 1'b0;
  assign n_4_net__99_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__99_ : 1'b0;
  assign n_4_net__98_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__98_ : 1'b0;
  assign n_4_net__97_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__97_ : 1'b0;
  assign n_4_net__96_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__96_ : 1'b0;
  assign n_4_net__95_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__95_ : 1'b0;
  assign n_4_net__94_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__94_ : 1'b0;
  assign n_4_net__93_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__93_ : 1'b0;
  assign n_4_net__92_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__92_ : 1'b0;
  assign n_4_net__91_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__91_ : 1'b0;
  assign n_4_net__90_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__90_ : 1'b0;
  assign n_4_net__89_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__89_ : 1'b0;
  assign n_4_net__88_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__88_ : 1'b0;
  assign n_4_net__87_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__87_ : 1'b0;
  assign n_4_net__86_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__86_ : 1'b0;
  assign n_4_net__85_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__85_ : 1'b0;
  assign n_4_net__84_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__84_ : 1'b0;
  assign n_4_net__83_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__83_ : 1'b0;
  assign n_4_net__82_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__82_ : 1'b0;
  assign n_4_net__81_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__81_ : 1'b0;
  assign n_4_net__80_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__80_ : 1'b0;
  assign n_4_net__79_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__79_ : 1'b0;
  assign n_4_net__78_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__78_ : 1'b0;
  assign n_4_net__77_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__77_ : 1'b0;
  assign n_4_net__76_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__76_ : 1'b0;
  assign n_4_net__75_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__75_ : 1'b0;
  assign n_4_net__74_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__74_ : 1'b0;
  assign n_4_net__73_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__73_ : 1'b0;
  assign n_4_net__72_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__72_ : 1'b0;
  assign n_4_net__71_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__71_ : 1'b0;
  assign n_4_net__70_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__70_ : 1'b0;
  assign n_4_net__69_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__69_ : 1'b0;
  assign n_4_net__68_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__68_ : 1'b0;
  assign n_4_net__67_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__67_ : 1'b0;
  assign n_4_net__66_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__66_ : 1'b0;
  assign n_4_net__65_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__65_ : 1'b0;
  assign n_4_net__64_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__64_ : 1'b0;
  assign n_4_net__63_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__63_ : 1'b0;
  assign n_4_net__62_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__62_ : 1'b0;
  assign n_4_net__61_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__61_ : 1'b0;
  assign n_4_net__60_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__60_ : 1'b0;
  assign n_4_net__59_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__59_ : 1'b0;
  assign n_4_net__58_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__58_ : 1'b0;
  assign n_4_net__57_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__57_ : 1'b0;
  assign n_4_net__56_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__56_ : 1'b0;
  assign n_4_net__55_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__55_ : 1'b0;
  assign n_4_net__54_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__54_ : 1'b0;
  assign n_4_net__53_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__53_ : 1'b0;
  assign n_4_net__52_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__52_ : 1'b0;
  assign n_4_net__51_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__51_ : 1'b0;
  assign n_4_net__50_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__50_ : 1'b0;
  assign n_4_net__49_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__49_ : 1'b0;
  assign n_4_net__48_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__48_ : 1'b0;
  assign n_4_net__47_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__47_ : 1'b0;
  assign n_4_net__46_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__46_ : 1'b0;
  assign n_4_net__45_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__45_ : 1'b0;
  assign n_4_net__44_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__44_ : 1'b0;
  assign n_4_net__43_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__43_ : 1'b0;
  assign n_4_net__42_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__42_ : 1'b0;
  assign n_4_net__41_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__41_ : 1'b0;
  assign n_4_net__40_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__40_ : 1'b0;
  assign n_4_net__39_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__39_ : 1'b0;
  assign n_4_net__38_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__38_ : 1'b0;
  assign n_4_net__37_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__37_ : 1'b0;
  assign n_4_net__36_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__36_ : 1'b0;
  assign n_4_net__35_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__35_ : 1'b0;
  assign n_4_net__34_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__34_ : 1'b0;
  assign n_4_net__33_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__33_ : 1'b0;
  assign n_4_net__32_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__32_ : 1'b0;
  assign n_4_net__31_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__31_ : 1'b0;
  assign n_4_net__30_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__30_ : 1'b0;
  assign n_4_net__29_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__29_ : 1'b0;
  assign n_4_net__28_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__28_ : 1'b0;
  assign n_4_net__27_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__27_ : 1'b0;
  assign n_4_net__26_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__26_ : 1'b0;
  assign n_4_net__25_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__25_ : 1'b0;
  assign n_4_net__24_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__24_ : 1'b0;
  assign n_4_net__23_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__23_ : 1'b0;
  assign n_4_net__22_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__22_ : 1'b0;
  assign n_4_net__21_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__21_ : 1'b0;
  assign n_4_net__20_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__20_ : 1'b0;
  assign n_4_net__19_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__19_ : 1'b0;
  assign n_4_net__18_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__18_ : 1'b0;
  assign n_4_net__17_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__17_ : 1'b0;
  assign n_4_net__16_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__16_ : 1'b0;
  assign n_4_net__15_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__15_ : 1'b0;
  assign n_4_net__14_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__14_ : 1'b0;
  assign n_4_net__13_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__13_ : 1'b0;
  assign n_4_net__12_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__12_ : 1'b0;
  assign n_4_net__11_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__11_ : 1'b0;
  assign n_4_net__10_ = (N115)? 1'b0 : 
                        (N116)? 1'b0 : 
                        (N117)? 1'b0 : 
                        (N118)? 1'b0 : 
                        (N119)? 1'b0 : 
                        (N120)? 1'b0 : 
                        (N121)? 1'b0 : 
                        (N122)? 1'b0 : 
                        (N123)? 1'b0 : 
                        (N124)? data_head_9__10_ : 1'b0;
  assign n_4_net__9_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__9_ : 1'b0;
  assign n_4_net__8_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__8_ : 1'b0;
  assign n_4_net__7_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__7_ : 1'b0;
  assign n_4_net__6_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__6_ : 1'b0;
  assign n_4_net__5_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__5_ : 1'b0;
  assign n_4_net__4_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__4_ : 1'b0;
  assign n_4_net__3_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__3_ : 1'b0;
  assign n_4_net__2_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__2_ : 1'b0;
  assign n_4_net__1_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__1_ : 1'b0;
  assign n_4_net__0_ = (N115)? 1'b0 : 
                       (N116)? 1'b0 : 
                       (N117)? 1'b0 : 
                       (N118)? 1'b0 : 
                       (N119)? 1'b0 : 
                       (N120)? 1'b0 : 
                       (N121)? 1'b0 : 
                       (N122)? 1'b0 : 
                       (N123)? 1'b0 : 
                       (N124)? data_head_9__0_ : 1'b0;
  assign n_0_net_ = reset | N179;
  assign n_5_net_ = reset | N184;

endmodule



module bsg_assembler_out
(
  clk,
  reset,
  calibration_done_i,
  valid_i,
  data_i,
  ready_o,
  in_top_channel_i,
  out_top_channel_i,
  valid_o,
  data_o,
  ready_i
);

  input [1279:0] data_i;
  input [3:0] in_top_channel_i;
  input [3:0] out_top_channel_i;
  output [9:0] valid_o;
  output [1279:0] data_o;
  input [9:0] ready_i;
  input clk;
  input reset;
  input calibration_done_i;
  input valid_i;
  output ready_o;
  wire [9:0] valid_o,fifo_not_full_vec,fifo_valid_vec,fifo_deq_vec;
  wire [1279:0] data_o,fifo_data_vec;
  wire ready_o,n_0_net_,n_1_net_,n_2_net_,n_3_net_,n_4_net_,n_5_net_,n_6_net_,n_7_net_,
  n_8_net_,n_9_net_,N0,N1,N2,N3,N4,N5,N6,N7,N8;

  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_0__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[0]),
    .data_i(data_i[127:0]),
    .v_i(n_0_net_),
    .v_o(fifo_valid_vec[0]),
    .data_o(fifo_data_vec[127:0]),
    .yumi_i(fifo_deq_vec[0])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_1__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[1]),
    .data_i(data_i[255:128]),
    .v_i(n_1_net_),
    .v_o(fifo_valid_vec[1]),
    .data_o(fifo_data_vec[255:128]),
    .yumi_i(fifo_deq_vec[1])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_2__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[2]),
    .data_i(data_i[383:256]),
    .v_i(n_2_net_),
    .v_o(fifo_valid_vec[2]),
    .data_o(fifo_data_vec[383:256]),
    .yumi_i(fifo_deq_vec[2])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_3__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[3]),
    .data_i(data_i[511:384]),
    .v_i(n_3_net_),
    .v_o(fifo_valid_vec[3]),
    .data_o(fifo_data_vec[511:384]),
    .yumi_i(fifo_deq_vec[3])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_4__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[4]),
    .data_i(data_i[639:512]),
    .v_i(n_4_net_),
    .v_o(fifo_valid_vec[4]),
    .data_o(fifo_data_vec[639:512]),
    .yumi_i(fifo_deq_vec[4])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_5__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[5]),
    .data_i(data_i[767:640]),
    .v_i(n_5_net_),
    .v_o(fifo_valid_vec[5]),
    .data_o(fifo_data_vec[767:640]),
    .yumi_i(fifo_deq_vec[5])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_6__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[6]),
    .data_i(data_i[895:768]),
    .v_i(n_6_net_),
    .v_o(fifo_valid_vec[6]),
    .data_o(fifo_data_vec[895:768]),
    .yumi_i(fifo_deq_vec[6])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_7__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[7]),
    .data_i(data_i[1023:896]),
    .v_i(n_7_net_),
    .v_o(fifo_valid_vec[7]),
    .data_o(fifo_data_vec[1023:896]),
    .yumi_i(fifo_deq_vec[7])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_8__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[8]),
    .data_i(data_i[1151:1024]),
    .v_i(n_8_net_),
    .v_o(fifo_valid_vec[8]),
    .data_o(fifo_data_vec[1151:1024]),
    .yumi_i(fifo_deq_vec[8])
  );


  bsg_two_fifo_width_p128_ready_THEN_valid_p1
  fifos_9__ring_packet_fifo
  (
    .clk_i(clk),
    .reset_i(reset),
    .ready_o(fifo_not_full_vec[9]),
    .data_i(data_i[1279:1152]),
    .v_i(n_9_net_),
    .v_o(fifo_valid_vec[9]),
    .data_o(fifo_data_vec[1279:1152]),
    .yumi_i(fifo_deq_vec[9])
  );


  bsg_round_robin_fifo_to_fifo_width_p128_num_in_p10_num_out_p10_out_channel_count_mask_p512
  rr_fifo_to_fifo
  (
    .clk(clk),
    .reset(reset),
    .valid_i(fifo_valid_vec),
    .data_i(fifo_data_vec),
    .yumi_o(fifo_deq_vec),
    .in_top_channel_i(in_top_channel_i),
    .out_top_channel_i(out_top_channel_i),
    .valid_o(valid_o),
    .data_o(data_o),
    .ready_i(ready_i)
  );

  assign ready_o = N8 & calibration_done_i;
  assign N8 = N7 & fifo_not_full_vec[0];
  assign N7 = N6 & fifo_not_full_vec[1];
  assign N6 = N5 & fifo_not_full_vec[2];
  assign N5 = N4 & fifo_not_full_vec[3];
  assign N4 = N3 & fifo_not_full_vec[4];
  assign N3 = N2 & fifo_not_full_vec[5];
  assign N2 = N1 & fifo_not_full_vec[6];
  assign N1 = N0 & fifo_not_full_vec[7];
  assign N0 = fifo_not_full_vec[9] & fifo_not_full_vec[8];
  assign n_0_net_ = valid_i & ready_o;
  assign n_1_net_ = valid_i & ready_o;
  assign n_2_net_ = valid_i & ready_o;
  assign n_3_net_ = valid_i & ready_o;
  assign n_4_net_ = valid_i & ready_o;
  assign n_5_net_ = valid_i & ready_o;
  assign n_6_net_ = valid_i & ready_o;
  assign n_7_net_ = valid_i & ready_o;
  assign n_8_net_ = valid_i & ready_o;
  assign n_9_net_ = valid_i & ready_o;

endmodule

