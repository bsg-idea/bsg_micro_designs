

module top
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;

  bsg_fifo_1r1w_narrowed
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .v_o(v_o)
  );


endmodule



module bsg_circular_ptr_slots_p50_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [5:0] o;
  output [5:0] n_o;
  input clk;
  input reset_i;
  wire [5:0] o,n_o,ptr_nowrap;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9;
  wire [6:0] ptr_wrap;
  reg o_5_sv2v_reg,o_4_sv2v_reg,o_3_sv2v_reg,o_2_sv2v_reg,o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[5] = o_5_sv2v_reg;
  assign o[4] = o_4_sv2v_reg;
  assign o[3] = o_3_sv2v_reg;
  assign o[2] = o_2_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign ptr_nowrap = o + add_i[0];
  assign { N8, N7, N6, N5, N4, N3, N2 } = o - { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 };
  assign ptr_wrap = { N8, N7, N6, N5, N4, N3, N2 } + add_i[0];
  assign n_o = (N0)? ptr_wrap[5:0] : 
               (N1)? ptr_nowrap : 1'b0;
  assign N0 = N9;
  assign N1 = ptr_wrap[6];
  assign N9 = ~ptr_wrap[6];

  always @(posedge clk) begin
    if(reset_i) begin
      o_5_sv2v_reg <= 1'b0;
      o_4_sv2v_reg <= 1'b0;
      o_3_sv2v_reg <= 1'b0;
      o_2_sv2v_reg <= 1'b0;
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_5_sv2v_reg <= n_o[5];
      o_4_sv2v_reg <= n_o[4];
      o_3_sv2v_reg <= n_o[3];
      o_2_sv2v_reg <= n_o[2];
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p50
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [5:0] wptr_r_o;
  output [5:0] rptr_r_o;
  output [5:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [5:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,N0,N1,N2,enq_r,deq_r,N3,equal_ptrs,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,
  sv2v_dc_4,sv2v_dc_5,sv2v_dc_6;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p50_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p50_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N3 = (N0)? 1'b1 : 
              (N2)? 1'b0 : 1'b0;
  assign N0 = N1;
  assign N1 = enq_i | deq_i;
  assign N2 = ~N1;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N3) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p50_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [31:0] w_data_i;
  input [5:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448;
  wire [1599:0] mem;
  reg mem_1599_sv2v_reg,mem_1598_sv2v_reg,mem_1597_sv2v_reg,mem_1596_sv2v_reg,
  mem_1595_sv2v_reg,mem_1594_sv2v_reg,mem_1593_sv2v_reg,mem_1592_sv2v_reg,
  mem_1591_sv2v_reg,mem_1590_sv2v_reg,mem_1589_sv2v_reg,mem_1588_sv2v_reg,mem_1587_sv2v_reg,
  mem_1586_sv2v_reg,mem_1585_sv2v_reg,mem_1584_sv2v_reg,mem_1583_sv2v_reg,
  mem_1582_sv2v_reg,mem_1581_sv2v_reg,mem_1580_sv2v_reg,mem_1579_sv2v_reg,mem_1578_sv2v_reg,
  mem_1577_sv2v_reg,mem_1576_sv2v_reg,mem_1575_sv2v_reg,mem_1574_sv2v_reg,
  mem_1573_sv2v_reg,mem_1572_sv2v_reg,mem_1571_sv2v_reg,mem_1570_sv2v_reg,mem_1569_sv2v_reg,
  mem_1568_sv2v_reg,mem_1567_sv2v_reg,mem_1566_sv2v_reg,mem_1565_sv2v_reg,
  mem_1564_sv2v_reg,mem_1563_sv2v_reg,mem_1562_sv2v_reg,mem_1561_sv2v_reg,mem_1560_sv2v_reg,
  mem_1559_sv2v_reg,mem_1558_sv2v_reg,mem_1557_sv2v_reg,mem_1556_sv2v_reg,
  mem_1555_sv2v_reg,mem_1554_sv2v_reg,mem_1553_sv2v_reg,mem_1552_sv2v_reg,
  mem_1551_sv2v_reg,mem_1550_sv2v_reg,mem_1549_sv2v_reg,mem_1548_sv2v_reg,mem_1547_sv2v_reg,
  mem_1546_sv2v_reg,mem_1545_sv2v_reg,mem_1544_sv2v_reg,mem_1543_sv2v_reg,
  mem_1542_sv2v_reg,mem_1541_sv2v_reg,mem_1540_sv2v_reg,mem_1539_sv2v_reg,mem_1538_sv2v_reg,
  mem_1537_sv2v_reg,mem_1536_sv2v_reg,mem_1535_sv2v_reg,mem_1534_sv2v_reg,
  mem_1533_sv2v_reg,mem_1532_sv2v_reg,mem_1531_sv2v_reg,mem_1530_sv2v_reg,mem_1529_sv2v_reg,
  mem_1528_sv2v_reg,mem_1527_sv2v_reg,mem_1526_sv2v_reg,mem_1525_sv2v_reg,
  mem_1524_sv2v_reg,mem_1523_sv2v_reg,mem_1522_sv2v_reg,mem_1521_sv2v_reg,mem_1520_sv2v_reg,
  mem_1519_sv2v_reg,mem_1518_sv2v_reg,mem_1517_sv2v_reg,mem_1516_sv2v_reg,
  mem_1515_sv2v_reg,mem_1514_sv2v_reg,mem_1513_sv2v_reg,mem_1512_sv2v_reg,
  mem_1511_sv2v_reg,mem_1510_sv2v_reg,mem_1509_sv2v_reg,mem_1508_sv2v_reg,mem_1507_sv2v_reg,
  mem_1506_sv2v_reg,mem_1505_sv2v_reg,mem_1504_sv2v_reg,mem_1503_sv2v_reg,
  mem_1502_sv2v_reg,mem_1501_sv2v_reg,mem_1500_sv2v_reg,mem_1499_sv2v_reg,mem_1498_sv2v_reg,
  mem_1497_sv2v_reg,mem_1496_sv2v_reg,mem_1495_sv2v_reg,mem_1494_sv2v_reg,
  mem_1493_sv2v_reg,mem_1492_sv2v_reg,mem_1491_sv2v_reg,mem_1490_sv2v_reg,mem_1489_sv2v_reg,
  mem_1488_sv2v_reg,mem_1487_sv2v_reg,mem_1486_sv2v_reg,mem_1485_sv2v_reg,
  mem_1484_sv2v_reg,mem_1483_sv2v_reg,mem_1482_sv2v_reg,mem_1481_sv2v_reg,mem_1480_sv2v_reg,
  mem_1479_sv2v_reg,mem_1478_sv2v_reg,mem_1477_sv2v_reg,mem_1476_sv2v_reg,
  mem_1475_sv2v_reg,mem_1474_sv2v_reg,mem_1473_sv2v_reg,mem_1472_sv2v_reg,
  mem_1471_sv2v_reg,mem_1470_sv2v_reg,mem_1469_sv2v_reg,mem_1468_sv2v_reg,mem_1467_sv2v_reg,
  mem_1466_sv2v_reg,mem_1465_sv2v_reg,mem_1464_sv2v_reg,mem_1463_sv2v_reg,
  mem_1462_sv2v_reg,mem_1461_sv2v_reg,mem_1460_sv2v_reg,mem_1459_sv2v_reg,mem_1458_sv2v_reg,
  mem_1457_sv2v_reg,mem_1456_sv2v_reg,mem_1455_sv2v_reg,mem_1454_sv2v_reg,
  mem_1453_sv2v_reg,mem_1452_sv2v_reg,mem_1451_sv2v_reg,mem_1450_sv2v_reg,mem_1449_sv2v_reg,
  mem_1448_sv2v_reg,mem_1447_sv2v_reg,mem_1446_sv2v_reg,mem_1445_sv2v_reg,
  mem_1444_sv2v_reg,mem_1443_sv2v_reg,mem_1442_sv2v_reg,mem_1441_sv2v_reg,mem_1440_sv2v_reg,
  mem_1439_sv2v_reg,mem_1438_sv2v_reg,mem_1437_sv2v_reg,mem_1436_sv2v_reg,
  mem_1435_sv2v_reg,mem_1434_sv2v_reg,mem_1433_sv2v_reg,mem_1432_sv2v_reg,
  mem_1431_sv2v_reg,mem_1430_sv2v_reg,mem_1429_sv2v_reg,mem_1428_sv2v_reg,mem_1427_sv2v_reg,
  mem_1426_sv2v_reg,mem_1425_sv2v_reg,mem_1424_sv2v_reg,mem_1423_sv2v_reg,
  mem_1422_sv2v_reg,mem_1421_sv2v_reg,mem_1420_sv2v_reg,mem_1419_sv2v_reg,mem_1418_sv2v_reg,
  mem_1417_sv2v_reg,mem_1416_sv2v_reg,mem_1415_sv2v_reg,mem_1414_sv2v_reg,
  mem_1413_sv2v_reg,mem_1412_sv2v_reg,mem_1411_sv2v_reg,mem_1410_sv2v_reg,mem_1409_sv2v_reg,
  mem_1408_sv2v_reg,mem_1407_sv2v_reg,mem_1406_sv2v_reg,mem_1405_sv2v_reg,
  mem_1404_sv2v_reg,mem_1403_sv2v_reg,mem_1402_sv2v_reg,mem_1401_sv2v_reg,mem_1400_sv2v_reg,
  mem_1399_sv2v_reg,mem_1398_sv2v_reg,mem_1397_sv2v_reg,mem_1396_sv2v_reg,
  mem_1395_sv2v_reg,mem_1394_sv2v_reg,mem_1393_sv2v_reg,mem_1392_sv2v_reg,
  mem_1391_sv2v_reg,mem_1390_sv2v_reg,mem_1389_sv2v_reg,mem_1388_sv2v_reg,mem_1387_sv2v_reg,
  mem_1386_sv2v_reg,mem_1385_sv2v_reg,mem_1384_sv2v_reg,mem_1383_sv2v_reg,
  mem_1382_sv2v_reg,mem_1381_sv2v_reg,mem_1380_sv2v_reg,mem_1379_sv2v_reg,mem_1378_sv2v_reg,
  mem_1377_sv2v_reg,mem_1376_sv2v_reg,mem_1375_sv2v_reg,mem_1374_sv2v_reg,
  mem_1373_sv2v_reg,mem_1372_sv2v_reg,mem_1371_sv2v_reg,mem_1370_sv2v_reg,mem_1369_sv2v_reg,
  mem_1368_sv2v_reg,mem_1367_sv2v_reg,mem_1366_sv2v_reg,mem_1365_sv2v_reg,
  mem_1364_sv2v_reg,mem_1363_sv2v_reg,mem_1362_sv2v_reg,mem_1361_sv2v_reg,mem_1360_sv2v_reg,
  mem_1359_sv2v_reg,mem_1358_sv2v_reg,mem_1357_sv2v_reg,mem_1356_sv2v_reg,
  mem_1355_sv2v_reg,mem_1354_sv2v_reg,mem_1353_sv2v_reg,mem_1352_sv2v_reg,
  mem_1351_sv2v_reg,mem_1350_sv2v_reg,mem_1349_sv2v_reg,mem_1348_sv2v_reg,mem_1347_sv2v_reg,
  mem_1346_sv2v_reg,mem_1345_sv2v_reg,mem_1344_sv2v_reg,mem_1343_sv2v_reg,
  mem_1342_sv2v_reg,mem_1341_sv2v_reg,mem_1340_sv2v_reg,mem_1339_sv2v_reg,mem_1338_sv2v_reg,
  mem_1337_sv2v_reg,mem_1336_sv2v_reg,mem_1335_sv2v_reg,mem_1334_sv2v_reg,
  mem_1333_sv2v_reg,mem_1332_sv2v_reg,mem_1331_sv2v_reg,mem_1330_sv2v_reg,mem_1329_sv2v_reg,
  mem_1328_sv2v_reg,mem_1327_sv2v_reg,mem_1326_sv2v_reg,mem_1325_sv2v_reg,
  mem_1324_sv2v_reg,mem_1323_sv2v_reg,mem_1322_sv2v_reg,mem_1321_sv2v_reg,mem_1320_sv2v_reg,
  mem_1319_sv2v_reg,mem_1318_sv2v_reg,mem_1317_sv2v_reg,mem_1316_sv2v_reg,
  mem_1315_sv2v_reg,mem_1314_sv2v_reg,mem_1313_sv2v_reg,mem_1312_sv2v_reg,
  mem_1311_sv2v_reg,mem_1310_sv2v_reg,mem_1309_sv2v_reg,mem_1308_sv2v_reg,mem_1307_sv2v_reg,
  mem_1306_sv2v_reg,mem_1305_sv2v_reg,mem_1304_sv2v_reg,mem_1303_sv2v_reg,
  mem_1302_sv2v_reg,mem_1301_sv2v_reg,mem_1300_sv2v_reg,mem_1299_sv2v_reg,mem_1298_sv2v_reg,
  mem_1297_sv2v_reg,mem_1296_sv2v_reg,mem_1295_sv2v_reg,mem_1294_sv2v_reg,
  mem_1293_sv2v_reg,mem_1292_sv2v_reg,mem_1291_sv2v_reg,mem_1290_sv2v_reg,mem_1289_sv2v_reg,
  mem_1288_sv2v_reg,mem_1287_sv2v_reg,mem_1286_sv2v_reg,mem_1285_sv2v_reg,
  mem_1284_sv2v_reg,mem_1283_sv2v_reg,mem_1282_sv2v_reg,mem_1281_sv2v_reg,mem_1280_sv2v_reg,
  mem_1279_sv2v_reg,mem_1278_sv2v_reg,mem_1277_sv2v_reg,mem_1276_sv2v_reg,
  mem_1275_sv2v_reg,mem_1274_sv2v_reg,mem_1273_sv2v_reg,mem_1272_sv2v_reg,
  mem_1271_sv2v_reg,mem_1270_sv2v_reg,mem_1269_sv2v_reg,mem_1268_sv2v_reg,mem_1267_sv2v_reg,
  mem_1266_sv2v_reg,mem_1265_sv2v_reg,mem_1264_sv2v_reg,mem_1263_sv2v_reg,
  mem_1262_sv2v_reg,mem_1261_sv2v_reg,mem_1260_sv2v_reg,mem_1259_sv2v_reg,mem_1258_sv2v_reg,
  mem_1257_sv2v_reg,mem_1256_sv2v_reg,mem_1255_sv2v_reg,mem_1254_sv2v_reg,
  mem_1253_sv2v_reg,mem_1252_sv2v_reg,mem_1251_sv2v_reg,mem_1250_sv2v_reg,mem_1249_sv2v_reg,
  mem_1248_sv2v_reg,mem_1247_sv2v_reg,mem_1246_sv2v_reg,mem_1245_sv2v_reg,
  mem_1244_sv2v_reg,mem_1243_sv2v_reg,mem_1242_sv2v_reg,mem_1241_sv2v_reg,mem_1240_sv2v_reg,
  mem_1239_sv2v_reg,mem_1238_sv2v_reg,mem_1237_sv2v_reg,mem_1236_sv2v_reg,
  mem_1235_sv2v_reg,mem_1234_sv2v_reg,mem_1233_sv2v_reg,mem_1232_sv2v_reg,
  mem_1231_sv2v_reg,mem_1230_sv2v_reg,mem_1229_sv2v_reg,mem_1228_sv2v_reg,mem_1227_sv2v_reg,
  mem_1226_sv2v_reg,mem_1225_sv2v_reg,mem_1224_sv2v_reg,mem_1223_sv2v_reg,
  mem_1222_sv2v_reg,mem_1221_sv2v_reg,mem_1220_sv2v_reg,mem_1219_sv2v_reg,mem_1218_sv2v_reg,
  mem_1217_sv2v_reg,mem_1216_sv2v_reg,mem_1215_sv2v_reg,mem_1214_sv2v_reg,
  mem_1213_sv2v_reg,mem_1212_sv2v_reg,mem_1211_sv2v_reg,mem_1210_sv2v_reg,mem_1209_sv2v_reg,
  mem_1208_sv2v_reg,mem_1207_sv2v_reg,mem_1206_sv2v_reg,mem_1205_sv2v_reg,
  mem_1204_sv2v_reg,mem_1203_sv2v_reg,mem_1202_sv2v_reg,mem_1201_sv2v_reg,mem_1200_sv2v_reg,
  mem_1199_sv2v_reg,mem_1198_sv2v_reg,mem_1197_sv2v_reg,mem_1196_sv2v_reg,
  mem_1195_sv2v_reg,mem_1194_sv2v_reg,mem_1193_sv2v_reg,mem_1192_sv2v_reg,
  mem_1191_sv2v_reg,mem_1190_sv2v_reg,mem_1189_sv2v_reg,mem_1188_sv2v_reg,mem_1187_sv2v_reg,
  mem_1186_sv2v_reg,mem_1185_sv2v_reg,mem_1184_sv2v_reg,mem_1183_sv2v_reg,
  mem_1182_sv2v_reg,mem_1181_sv2v_reg,mem_1180_sv2v_reg,mem_1179_sv2v_reg,mem_1178_sv2v_reg,
  mem_1177_sv2v_reg,mem_1176_sv2v_reg,mem_1175_sv2v_reg,mem_1174_sv2v_reg,
  mem_1173_sv2v_reg,mem_1172_sv2v_reg,mem_1171_sv2v_reg,mem_1170_sv2v_reg,mem_1169_sv2v_reg,
  mem_1168_sv2v_reg,mem_1167_sv2v_reg,mem_1166_sv2v_reg,mem_1165_sv2v_reg,
  mem_1164_sv2v_reg,mem_1163_sv2v_reg,mem_1162_sv2v_reg,mem_1161_sv2v_reg,mem_1160_sv2v_reg,
  mem_1159_sv2v_reg,mem_1158_sv2v_reg,mem_1157_sv2v_reg,mem_1156_sv2v_reg,
  mem_1155_sv2v_reg,mem_1154_sv2v_reg,mem_1153_sv2v_reg,mem_1152_sv2v_reg,
  mem_1151_sv2v_reg,mem_1150_sv2v_reg,mem_1149_sv2v_reg,mem_1148_sv2v_reg,mem_1147_sv2v_reg,
  mem_1146_sv2v_reg,mem_1145_sv2v_reg,mem_1144_sv2v_reg,mem_1143_sv2v_reg,
  mem_1142_sv2v_reg,mem_1141_sv2v_reg,mem_1140_sv2v_reg,mem_1139_sv2v_reg,mem_1138_sv2v_reg,
  mem_1137_sv2v_reg,mem_1136_sv2v_reg,mem_1135_sv2v_reg,mem_1134_sv2v_reg,
  mem_1133_sv2v_reg,mem_1132_sv2v_reg,mem_1131_sv2v_reg,mem_1130_sv2v_reg,mem_1129_sv2v_reg,
  mem_1128_sv2v_reg,mem_1127_sv2v_reg,mem_1126_sv2v_reg,mem_1125_sv2v_reg,
  mem_1124_sv2v_reg,mem_1123_sv2v_reg,mem_1122_sv2v_reg,mem_1121_sv2v_reg,mem_1120_sv2v_reg,
  mem_1119_sv2v_reg,mem_1118_sv2v_reg,mem_1117_sv2v_reg,mem_1116_sv2v_reg,
  mem_1115_sv2v_reg,mem_1114_sv2v_reg,mem_1113_sv2v_reg,mem_1112_sv2v_reg,
  mem_1111_sv2v_reg,mem_1110_sv2v_reg,mem_1109_sv2v_reg,mem_1108_sv2v_reg,mem_1107_sv2v_reg,
  mem_1106_sv2v_reg,mem_1105_sv2v_reg,mem_1104_sv2v_reg,mem_1103_sv2v_reg,
  mem_1102_sv2v_reg,mem_1101_sv2v_reg,mem_1100_sv2v_reg,mem_1099_sv2v_reg,mem_1098_sv2v_reg,
  mem_1097_sv2v_reg,mem_1096_sv2v_reg,mem_1095_sv2v_reg,mem_1094_sv2v_reg,
  mem_1093_sv2v_reg,mem_1092_sv2v_reg,mem_1091_sv2v_reg,mem_1090_sv2v_reg,mem_1089_sv2v_reg,
  mem_1088_sv2v_reg,mem_1087_sv2v_reg,mem_1086_sv2v_reg,mem_1085_sv2v_reg,
  mem_1084_sv2v_reg,mem_1083_sv2v_reg,mem_1082_sv2v_reg,mem_1081_sv2v_reg,mem_1080_sv2v_reg,
  mem_1079_sv2v_reg,mem_1078_sv2v_reg,mem_1077_sv2v_reg,mem_1076_sv2v_reg,
  mem_1075_sv2v_reg,mem_1074_sv2v_reg,mem_1073_sv2v_reg,mem_1072_sv2v_reg,
  mem_1071_sv2v_reg,mem_1070_sv2v_reg,mem_1069_sv2v_reg,mem_1068_sv2v_reg,mem_1067_sv2v_reg,
  mem_1066_sv2v_reg,mem_1065_sv2v_reg,mem_1064_sv2v_reg,mem_1063_sv2v_reg,
  mem_1062_sv2v_reg,mem_1061_sv2v_reg,mem_1060_sv2v_reg,mem_1059_sv2v_reg,mem_1058_sv2v_reg,
  mem_1057_sv2v_reg,mem_1056_sv2v_reg,mem_1055_sv2v_reg,mem_1054_sv2v_reg,
  mem_1053_sv2v_reg,mem_1052_sv2v_reg,mem_1051_sv2v_reg,mem_1050_sv2v_reg,mem_1049_sv2v_reg,
  mem_1048_sv2v_reg,mem_1047_sv2v_reg,mem_1046_sv2v_reg,mem_1045_sv2v_reg,
  mem_1044_sv2v_reg,mem_1043_sv2v_reg,mem_1042_sv2v_reg,mem_1041_sv2v_reg,mem_1040_sv2v_reg,
  mem_1039_sv2v_reg,mem_1038_sv2v_reg,mem_1037_sv2v_reg,mem_1036_sv2v_reg,
  mem_1035_sv2v_reg,mem_1034_sv2v_reg,mem_1033_sv2v_reg,mem_1032_sv2v_reg,
  mem_1031_sv2v_reg,mem_1030_sv2v_reg,mem_1029_sv2v_reg,mem_1028_sv2v_reg,mem_1027_sv2v_reg,
  mem_1026_sv2v_reg,mem_1025_sv2v_reg,mem_1024_sv2v_reg,mem_1023_sv2v_reg,
  mem_1022_sv2v_reg,mem_1021_sv2v_reg,mem_1020_sv2v_reg,mem_1019_sv2v_reg,mem_1018_sv2v_reg,
  mem_1017_sv2v_reg,mem_1016_sv2v_reg,mem_1015_sv2v_reg,mem_1014_sv2v_reg,
  mem_1013_sv2v_reg,mem_1012_sv2v_reg,mem_1011_sv2v_reg,mem_1010_sv2v_reg,mem_1009_sv2v_reg,
  mem_1008_sv2v_reg,mem_1007_sv2v_reg,mem_1006_sv2v_reg,mem_1005_sv2v_reg,
  mem_1004_sv2v_reg,mem_1003_sv2v_reg,mem_1002_sv2v_reg,mem_1001_sv2v_reg,mem_1000_sv2v_reg,
  mem_999_sv2v_reg,mem_998_sv2v_reg,mem_997_sv2v_reg,mem_996_sv2v_reg,
  mem_995_sv2v_reg,mem_994_sv2v_reg,mem_993_sv2v_reg,mem_992_sv2v_reg,mem_991_sv2v_reg,
  mem_990_sv2v_reg,mem_989_sv2v_reg,mem_988_sv2v_reg,mem_987_sv2v_reg,mem_986_sv2v_reg,
  mem_985_sv2v_reg,mem_984_sv2v_reg,mem_983_sv2v_reg,mem_982_sv2v_reg,
  mem_981_sv2v_reg,mem_980_sv2v_reg,mem_979_sv2v_reg,mem_978_sv2v_reg,mem_977_sv2v_reg,
  mem_976_sv2v_reg,mem_975_sv2v_reg,mem_974_sv2v_reg,mem_973_sv2v_reg,mem_972_sv2v_reg,
  mem_971_sv2v_reg,mem_970_sv2v_reg,mem_969_sv2v_reg,mem_968_sv2v_reg,
  mem_967_sv2v_reg,mem_966_sv2v_reg,mem_965_sv2v_reg,mem_964_sv2v_reg,mem_963_sv2v_reg,
  mem_962_sv2v_reg,mem_961_sv2v_reg,mem_960_sv2v_reg,mem_959_sv2v_reg,mem_958_sv2v_reg,
  mem_957_sv2v_reg,mem_956_sv2v_reg,mem_955_sv2v_reg,mem_954_sv2v_reg,mem_953_sv2v_reg,
  mem_952_sv2v_reg,mem_951_sv2v_reg,mem_950_sv2v_reg,mem_949_sv2v_reg,
  mem_948_sv2v_reg,mem_947_sv2v_reg,mem_946_sv2v_reg,mem_945_sv2v_reg,mem_944_sv2v_reg,
  mem_943_sv2v_reg,mem_942_sv2v_reg,mem_941_sv2v_reg,mem_940_sv2v_reg,mem_939_sv2v_reg,
  mem_938_sv2v_reg,mem_937_sv2v_reg,mem_936_sv2v_reg,mem_935_sv2v_reg,
  mem_934_sv2v_reg,mem_933_sv2v_reg,mem_932_sv2v_reg,mem_931_sv2v_reg,mem_930_sv2v_reg,
  mem_929_sv2v_reg,mem_928_sv2v_reg,mem_927_sv2v_reg,mem_926_sv2v_reg,mem_925_sv2v_reg,
  mem_924_sv2v_reg,mem_923_sv2v_reg,mem_922_sv2v_reg,mem_921_sv2v_reg,mem_920_sv2v_reg,
  mem_919_sv2v_reg,mem_918_sv2v_reg,mem_917_sv2v_reg,mem_916_sv2v_reg,
  mem_915_sv2v_reg,mem_914_sv2v_reg,mem_913_sv2v_reg,mem_912_sv2v_reg,mem_911_sv2v_reg,
  mem_910_sv2v_reg,mem_909_sv2v_reg,mem_908_sv2v_reg,mem_907_sv2v_reg,mem_906_sv2v_reg,
  mem_905_sv2v_reg,mem_904_sv2v_reg,mem_903_sv2v_reg,mem_902_sv2v_reg,
  mem_901_sv2v_reg,mem_900_sv2v_reg,mem_899_sv2v_reg,mem_898_sv2v_reg,mem_897_sv2v_reg,
  mem_896_sv2v_reg,mem_895_sv2v_reg,mem_894_sv2v_reg,mem_893_sv2v_reg,mem_892_sv2v_reg,
  mem_891_sv2v_reg,mem_890_sv2v_reg,mem_889_sv2v_reg,mem_888_sv2v_reg,
  mem_887_sv2v_reg,mem_886_sv2v_reg,mem_885_sv2v_reg,mem_884_sv2v_reg,mem_883_sv2v_reg,
  mem_882_sv2v_reg,mem_881_sv2v_reg,mem_880_sv2v_reg,mem_879_sv2v_reg,mem_878_sv2v_reg,
  mem_877_sv2v_reg,mem_876_sv2v_reg,mem_875_sv2v_reg,mem_874_sv2v_reg,mem_873_sv2v_reg,
  mem_872_sv2v_reg,mem_871_sv2v_reg,mem_870_sv2v_reg,mem_869_sv2v_reg,
  mem_868_sv2v_reg,mem_867_sv2v_reg,mem_866_sv2v_reg,mem_865_sv2v_reg,mem_864_sv2v_reg,
  mem_863_sv2v_reg,mem_862_sv2v_reg,mem_861_sv2v_reg,mem_860_sv2v_reg,mem_859_sv2v_reg,
  mem_858_sv2v_reg,mem_857_sv2v_reg,mem_856_sv2v_reg,mem_855_sv2v_reg,
  mem_854_sv2v_reg,mem_853_sv2v_reg,mem_852_sv2v_reg,mem_851_sv2v_reg,mem_850_sv2v_reg,
  mem_849_sv2v_reg,mem_848_sv2v_reg,mem_847_sv2v_reg,mem_846_sv2v_reg,mem_845_sv2v_reg,
  mem_844_sv2v_reg,mem_843_sv2v_reg,mem_842_sv2v_reg,mem_841_sv2v_reg,mem_840_sv2v_reg,
  mem_839_sv2v_reg,mem_838_sv2v_reg,mem_837_sv2v_reg,mem_836_sv2v_reg,
  mem_835_sv2v_reg,mem_834_sv2v_reg,mem_833_sv2v_reg,mem_832_sv2v_reg,mem_831_sv2v_reg,
  mem_830_sv2v_reg,mem_829_sv2v_reg,mem_828_sv2v_reg,mem_827_sv2v_reg,mem_826_sv2v_reg,
  mem_825_sv2v_reg,mem_824_sv2v_reg,mem_823_sv2v_reg,mem_822_sv2v_reg,
  mem_821_sv2v_reg,mem_820_sv2v_reg,mem_819_sv2v_reg,mem_818_sv2v_reg,mem_817_sv2v_reg,
  mem_816_sv2v_reg,mem_815_sv2v_reg,mem_814_sv2v_reg,mem_813_sv2v_reg,mem_812_sv2v_reg,
  mem_811_sv2v_reg,mem_810_sv2v_reg,mem_809_sv2v_reg,mem_808_sv2v_reg,
  mem_807_sv2v_reg,mem_806_sv2v_reg,mem_805_sv2v_reg,mem_804_sv2v_reg,mem_803_sv2v_reg,
  mem_802_sv2v_reg,mem_801_sv2v_reg,mem_800_sv2v_reg,mem_799_sv2v_reg,mem_798_sv2v_reg,
  mem_797_sv2v_reg,mem_796_sv2v_reg,mem_795_sv2v_reg,mem_794_sv2v_reg,mem_793_sv2v_reg,
  mem_792_sv2v_reg,mem_791_sv2v_reg,mem_790_sv2v_reg,mem_789_sv2v_reg,
  mem_788_sv2v_reg,mem_787_sv2v_reg,mem_786_sv2v_reg,mem_785_sv2v_reg,mem_784_sv2v_reg,
  mem_783_sv2v_reg,mem_782_sv2v_reg,mem_781_sv2v_reg,mem_780_sv2v_reg,mem_779_sv2v_reg,
  mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,mem_775_sv2v_reg,
  mem_774_sv2v_reg,mem_773_sv2v_reg,mem_772_sv2v_reg,mem_771_sv2v_reg,mem_770_sv2v_reg,
  mem_769_sv2v_reg,mem_768_sv2v_reg,mem_767_sv2v_reg,mem_766_sv2v_reg,mem_765_sv2v_reg,
  mem_764_sv2v_reg,mem_763_sv2v_reg,mem_762_sv2v_reg,mem_761_sv2v_reg,mem_760_sv2v_reg,
  mem_759_sv2v_reg,mem_758_sv2v_reg,mem_757_sv2v_reg,mem_756_sv2v_reg,
  mem_755_sv2v_reg,mem_754_sv2v_reg,mem_753_sv2v_reg,mem_752_sv2v_reg,mem_751_sv2v_reg,
  mem_750_sv2v_reg,mem_749_sv2v_reg,mem_748_sv2v_reg,mem_747_sv2v_reg,mem_746_sv2v_reg,
  mem_745_sv2v_reg,mem_744_sv2v_reg,mem_743_sv2v_reg,mem_742_sv2v_reg,
  mem_741_sv2v_reg,mem_740_sv2v_reg,mem_739_sv2v_reg,mem_738_sv2v_reg,mem_737_sv2v_reg,
  mem_736_sv2v_reg,mem_735_sv2v_reg,mem_734_sv2v_reg,mem_733_sv2v_reg,mem_732_sv2v_reg,
  mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,mem_728_sv2v_reg,
  mem_727_sv2v_reg,mem_726_sv2v_reg,mem_725_sv2v_reg,mem_724_sv2v_reg,mem_723_sv2v_reg,
  mem_722_sv2v_reg,mem_721_sv2v_reg,mem_720_sv2v_reg,mem_719_sv2v_reg,mem_718_sv2v_reg,
  mem_717_sv2v_reg,mem_716_sv2v_reg,mem_715_sv2v_reg,mem_714_sv2v_reg,mem_713_sv2v_reg,
  mem_712_sv2v_reg,mem_711_sv2v_reg,mem_710_sv2v_reg,mem_709_sv2v_reg,
  mem_708_sv2v_reg,mem_707_sv2v_reg,mem_706_sv2v_reg,mem_705_sv2v_reg,mem_704_sv2v_reg,
  mem_703_sv2v_reg,mem_702_sv2v_reg,mem_701_sv2v_reg,mem_700_sv2v_reg,mem_699_sv2v_reg,
  mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,mem_695_sv2v_reg,
  mem_694_sv2v_reg,mem_693_sv2v_reg,mem_692_sv2v_reg,mem_691_sv2v_reg,mem_690_sv2v_reg,
  mem_689_sv2v_reg,mem_688_sv2v_reg,mem_687_sv2v_reg,mem_686_sv2v_reg,mem_685_sv2v_reg,
  mem_684_sv2v_reg,mem_683_sv2v_reg,mem_682_sv2v_reg,mem_681_sv2v_reg,mem_680_sv2v_reg,
  mem_679_sv2v_reg,mem_678_sv2v_reg,mem_677_sv2v_reg,mem_676_sv2v_reg,
  mem_675_sv2v_reg,mem_674_sv2v_reg,mem_673_sv2v_reg,mem_672_sv2v_reg,mem_671_sv2v_reg,
  mem_670_sv2v_reg,mem_669_sv2v_reg,mem_668_sv2v_reg,mem_667_sv2v_reg,mem_666_sv2v_reg,
  mem_665_sv2v_reg,mem_664_sv2v_reg,mem_663_sv2v_reg,mem_662_sv2v_reg,
  mem_661_sv2v_reg,mem_660_sv2v_reg,mem_659_sv2v_reg,mem_658_sv2v_reg,mem_657_sv2v_reg,
  mem_656_sv2v_reg,mem_655_sv2v_reg,mem_654_sv2v_reg,mem_653_sv2v_reg,mem_652_sv2v_reg,
  mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,mem_648_sv2v_reg,
  mem_647_sv2v_reg,mem_646_sv2v_reg,mem_645_sv2v_reg,mem_644_sv2v_reg,mem_643_sv2v_reg,
  mem_642_sv2v_reg,mem_641_sv2v_reg,mem_640_sv2v_reg,mem_639_sv2v_reg,mem_638_sv2v_reg,
  mem_637_sv2v_reg,mem_636_sv2v_reg,mem_635_sv2v_reg,mem_634_sv2v_reg,mem_633_sv2v_reg,
  mem_632_sv2v_reg,mem_631_sv2v_reg,mem_630_sv2v_reg,mem_629_sv2v_reg,
  mem_628_sv2v_reg,mem_627_sv2v_reg,mem_626_sv2v_reg,mem_625_sv2v_reg,mem_624_sv2v_reg,
  mem_623_sv2v_reg,mem_622_sv2v_reg,mem_621_sv2v_reg,mem_620_sv2v_reg,mem_619_sv2v_reg,
  mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,mem_615_sv2v_reg,
  mem_614_sv2v_reg,mem_613_sv2v_reg,mem_612_sv2v_reg,mem_611_sv2v_reg,mem_610_sv2v_reg,
  mem_609_sv2v_reg,mem_608_sv2v_reg,mem_607_sv2v_reg,mem_606_sv2v_reg,mem_605_sv2v_reg,
  mem_604_sv2v_reg,mem_603_sv2v_reg,mem_602_sv2v_reg,mem_601_sv2v_reg,mem_600_sv2v_reg,
  mem_599_sv2v_reg,mem_598_sv2v_reg,mem_597_sv2v_reg,mem_596_sv2v_reg,
  mem_595_sv2v_reg,mem_594_sv2v_reg,mem_593_sv2v_reg,mem_592_sv2v_reg,mem_591_sv2v_reg,
  mem_590_sv2v_reg,mem_589_sv2v_reg,mem_588_sv2v_reg,mem_587_sv2v_reg,mem_586_sv2v_reg,
  mem_585_sv2v_reg,mem_584_sv2v_reg,mem_583_sv2v_reg,mem_582_sv2v_reg,
  mem_581_sv2v_reg,mem_580_sv2v_reg,mem_579_sv2v_reg,mem_578_sv2v_reg,mem_577_sv2v_reg,
  mem_576_sv2v_reg,mem_575_sv2v_reg,mem_574_sv2v_reg,mem_573_sv2v_reg,mem_572_sv2v_reg,
  mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,mem_568_sv2v_reg,
  mem_567_sv2v_reg,mem_566_sv2v_reg,mem_565_sv2v_reg,mem_564_sv2v_reg,mem_563_sv2v_reg,
  mem_562_sv2v_reg,mem_561_sv2v_reg,mem_560_sv2v_reg,mem_559_sv2v_reg,mem_558_sv2v_reg,
  mem_557_sv2v_reg,mem_556_sv2v_reg,mem_555_sv2v_reg,mem_554_sv2v_reg,mem_553_sv2v_reg,
  mem_552_sv2v_reg,mem_551_sv2v_reg,mem_550_sv2v_reg,mem_549_sv2v_reg,
  mem_548_sv2v_reg,mem_547_sv2v_reg,mem_546_sv2v_reg,mem_545_sv2v_reg,mem_544_sv2v_reg,
  mem_543_sv2v_reg,mem_542_sv2v_reg,mem_541_sv2v_reg,mem_540_sv2v_reg,mem_539_sv2v_reg,
  mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,mem_535_sv2v_reg,
  mem_534_sv2v_reg,mem_533_sv2v_reg,mem_532_sv2v_reg,mem_531_sv2v_reg,mem_530_sv2v_reg,
  mem_529_sv2v_reg,mem_528_sv2v_reg,mem_527_sv2v_reg,mem_526_sv2v_reg,mem_525_sv2v_reg,
  mem_524_sv2v_reg,mem_523_sv2v_reg,mem_522_sv2v_reg,mem_521_sv2v_reg,mem_520_sv2v_reg,
  mem_519_sv2v_reg,mem_518_sv2v_reg,mem_517_sv2v_reg,mem_516_sv2v_reg,
  mem_515_sv2v_reg,mem_514_sv2v_reg,mem_513_sv2v_reg,mem_512_sv2v_reg,mem_511_sv2v_reg,
  mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,mem_507_sv2v_reg,mem_506_sv2v_reg,
  mem_505_sv2v_reg,mem_504_sv2v_reg,mem_503_sv2v_reg,mem_502_sv2v_reg,
  mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,mem_497_sv2v_reg,
  mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,mem_493_sv2v_reg,mem_492_sv2v_reg,
  mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,mem_488_sv2v_reg,
  mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,mem_483_sv2v_reg,
  mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,mem_479_sv2v_reg,mem_478_sv2v_reg,
  mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,mem_474_sv2v_reg,mem_473_sv2v_reg,
  mem_472_sv2v_reg,mem_471_sv2v_reg,mem_470_sv2v_reg,mem_469_sv2v_reg,
  mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,mem_464_sv2v_reg,
  mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,mem_460_sv2v_reg,mem_459_sv2v_reg,
  mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,mem_455_sv2v_reg,
  mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,mem_450_sv2v_reg,
  mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,mem_446_sv2v_reg,mem_445_sv2v_reg,
  mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,mem_441_sv2v_reg,mem_440_sv2v_reg,
  mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,mem_436_sv2v_reg,
  mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,mem_431_sv2v_reg,
  mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,mem_427_sv2v_reg,mem_426_sv2v_reg,
  mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,mem_422_sv2v_reg,
  mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,mem_417_sv2v_reg,
  mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,mem_413_sv2v_reg,mem_412_sv2v_reg,
  mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,mem_408_sv2v_reg,
  mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,mem_403_sv2v_reg,
  mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,mem_399_sv2v_reg,mem_398_sv2v_reg,
  mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,mem_394_sv2v_reg,mem_393_sv2v_reg,
  mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,mem_389_sv2v_reg,
  mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,mem_384_sv2v_reg,
  mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,mem_380_sv2v_reg,mem_379_sv2v_reg,
  mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,mem_375_sv2v_reg,
  mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,mem_370_sv2v_reg,
  mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,mem_366_sv2v_reg,mem_365_sv2v_reg,
  mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,mem_361_sv2v_reg,mem_360_sv2v_reg,
  mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,mem_356_sv2v_reg,
  mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,mem_351_sv2v_reg,
  mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,mem_347_sv2v_reg,mem_346_sv2v_reg,
  mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,mem_342_sv2v_reg,
  mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,mem_337_sv2v_reg,
  mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,mem_333_sv2v_reg,mem_332_sv2v_reg,
  mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,mem_328_sv2v_reg,
  mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,mem_323_sv2v_reg,
  mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,mem_319_sv2v_reg,mem_318_sv2v_reg,
  mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,mem_314_sv2v_reg,mem_313_sv2v_reg,
  mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,mem_309_sv2v_reg,
  mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,mem_304_sv2v_reg,
  mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,mem_300_sv2v_reg,mem_299_sv2v_reg,
  mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,mem_295_sv2v_reg,
  mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,mem_290_sv2v_reg,
  mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,mem_286_sv2v_reg,mem_285_sv2v_reg,
  mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,mem_281_sv2v_reg,mem_280_sv2v_reg,
  mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,mem_276_sv2v_reg,
  mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,mem_271_sv2v_reg,
  mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,mem_267_sv2v_reg,mem_266_sv2v_reg,
  mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,mem_262_sv2v_reg,
  mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,mem_257_sv2v_reg,
  mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,
  mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,
  mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,
  mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,
  mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,mem_233_sv2v_reg,
  mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,mem_229_sv2v_reg,
  mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,
  mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,mem_219_sv2v_reg,
  mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,mem_215_sv2v_reg,
  mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,
  mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,
  mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,mem_200_sv2v_reg,
  mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,mem_196_sv2v_reg,
  mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,
  mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,mem_186_sv2v_reg,
  mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,mem_182_sv2v_reg,
  mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,
  mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,
  mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,
  mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,
  mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,
  mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,mem_153_sv2v_reg,
  mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,mem_149_sv2v_reg,
  mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,
  mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,mem_139_sv2v_reg,
  mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,mem_135_sv2v_reg,
  mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,
  mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,
  mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,mem_120_sv2v_reg,
  mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,mem_116_sv2v_reg,
  mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,
  mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,mem_106_sv2v_reg,
  mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,mem_102_sv2v_reg,
  mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,
  mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,
  mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,
  mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,
  mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,
  mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,
  mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,
  mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,
  mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,
  mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,
  mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,
  mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,
  mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,
  mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,
  mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,
  mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,
  mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,
  mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,
  mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,
  mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,
  mem_0_sv2v_reg;
  assign mem[1599] = mem_1599_sv2v_reg;
  assign mem[1598] = mem_1598_sv2v_reg;
  assign mem[1597] = mem_1597_sv2v_reg;
  assign mem[1596] = mem_1596_sv2v_reg;
  assign mem[1595] = mem_1595_sv2v_reg;
  assign mem[1594] = mem_1594_sv2v_reg;
  assign mem[1593] = mem_1593_sv2v_reg;
  assign mem[1592] = mem_1592_sv2v_reg;
  assign mem[1591] = mem_1591_sv2v_reg;
  assign mem[1590] = mem_1590_sv2v_reg;
  assign mem[1589] = mem_1589_sv2v_reg;
  assign mem[1588] = mem_1588_sv2v_reg;
  assign mem[1587] = mem_1587_sv2v_reg;
  assign mem[1586] = mem_1586_sv2v_reg;
  assign mem[1585] = mem_1585_sv2v_reg;
  assign mem[1584] = mem_1584_sv2v_reg;
  assign mem[1583] = mem_1583_sv2v_reg;
  assign mem[1582] = mem_1582_sv2v_reg;
  assign mem[1581] = mem_1581_sv2v_reg;
  assign mem[1580] = mem_1580_sv2v_reg;
  assign mem[1579] = mem_1579_sv2v_reg;
  assign mem[1578] = mem_1578_sv2v_reg;
  assign mem[1577] = mem_1577_sv2v_reg;
  assign mem[1576] = mem_1576_sv2v_reg;
  assign mem[1575] = mem_1575_sv2v_reg;
  assign mem[1574] = mem_1574_sv2v_reg;
  assign mem[1573] = mem_1573_sv2v_reg;
  assign mem[1572] = mem_1572_sv2v_reg;
  assign mem[1571] = mem_1571_sv2v_reg;
  assign mem[1570] = mem_1570_sv2v_reg;
  assign mem[1569] = mem_1569_sv2v_reg;
  assign mem[1568] = mem_1568_sv2v_reg;
  assign mem[1567] = mem_1567_sv2v_reg;
  assign mem[1566] = mem_1566_sv2v_reg;
  assign mem[1565] = mem_1565_sv2v_reg;
  assign mem[1564] = mem_1564_sv2v_reg;
  assign mem[1563] = mem_1563_sv2v_reg;
  assign mem[1562] = mem_1562_sv2v_reg;
  assign mem[1561] = mem_1561_sv2v_reg;
  assign mem[1560] = mem_1560_sv2v_reg;
  assign mem[1559] = mem_1559_sv2v_reg;
  assign mem[1558] = mem_1558_sv2v_reg;
  assign mem[1557] = mem_1557_sv2v_reg;
  assign mem[1556] = mem_1556_sv2v_reg;
  assign mem[1555] = mem_1555_sv2v_reg;
  assign mem[1554] = mem_1554_sv2v_reg;
  assign mem[1553] = mem_1553_sv2v_reg;
  assign mem[1552] = mem_1552_sv2v_reg;
  assign mem[1551] = mem_1551_sv2v_reg;
  assign mem[1550] = mem_1550_sv2v_reg;
  assign mem[1549] = mem_1549_sv2v_reg;
  assign mem[1548] = mem_1548_sv2v_reg;
  assign mem[1547] = mem_1547_sv2v_reg;
  assign mem[1546] = mem_1546_sv2v_reg;
  assign mem[1545] = mem_1545_sv2v_reg;
  assign mem[1544] = mem_1544_sv2v_reg;
  assign mem[1543] = mem_1543_sv2v_reg;
  assign mem[1542] = mem_1542_sv2v_reg;
  assign mem[1541] = mem_1541_sv2v_reg;
  assign mem[1540] = mem_1540_sv2v_reg;
  assign mem[1539] = mem_1539_sv2v_reg;
  assign mem[1538] = mem_1538_sv2v_reg;
  assign mem[1537] = mem_1537_sv2v_reg;
  assign mem[1536] = mem_1536_sv2v_reg;
  assign mem[1535] = mem_1535_sv2v_reg;
  assign mem[1534] = mem_1534_sv2v_reg;
  assign mem[1533] = mem_1533_sv2v_reg;
  assign mem[1532] = mem_1532_sv2v_reg;
  assign mem[1531] = mem_1531_sv2v_reg;
  assign mem[1530] = mem_1530_sv2v_reg;
  assign mem[1529] = mem_1529_sv2v_reg;
  assign mem[1528] = mem_1528_sv2v_reg;
  assign mem[1527] = mem_1527_sv2v_reg;
  assign mem[1526] = mem_1526_sv2v_reg;
  assign mem[1525] = mem_1525_sv2v_reg;
  assign mem[1524] = mem_1524_sv2v_reg;
  assign mem[1523] = mem_1523_sv2v_reg;
  assign mem[1522] = mem_1522_sv2v_reg;
  assign mem[1521] = mem_1521_sv2v_reg;
  assign mem[1520] = mem_1520_sv2v_reg;
  assign mem[1519] = mem_1519_sv2v_reg;
  assign mem[1518] = mem_1518_sv2v_reg;
  assign mem[1517] = mem_1517_sv2v_reg;
  assign mem[1516] = mem_1516_sv2v_reg;
  assign mem[1515] = mem_1515_sv2v_reg;
  assign mem[1514] = mem_1514_sv2v_reg;
  assign mem[1513] = mem_1513_sv2v_reg;
  assign mem[1512] = mem_1512_sv2v_reg;
  assign mem[1511] = mem_1511_sv2v_reg;
  assign mem[1510] = mem_1510_sv2v_reg;
  assign mem[1509] = mem_1509_sv2v_reg;
  assign mem[1508] = mem_1508_sv2v_reg;
  assign mem[1507] = mem_1507_sv2v_reg;
  assign mem[1506] = mem_1506_sv2v_reg;
  assign mem[1505] = mem_1505_sv2v_reg;
  assign mem[1504] = mem_1504_sv2v_reg;
  assign mem[1503] = mem_1503_sv2v_reg;
  assign mem[1502] = mem_1502_sv2v_reg;
  assign mem[1501] = mem_1501_sv2v_reg;
  assign mem[1500] = mem_1500_sv2v_reg;
  assign mem[1499] = mem_1499_sv2v_reg;
  assign mem[1498] = mem_1498_sv2v_reg;
  assign mem[1497] = mem_1497_sv2v_reg;
  assign mem[1496] = mem_1496_sv2v_reg;
  assign mem[1495] = mem_1495_sv2v_reg;
  assign mem[1494] = mem_1494_sv2v_reg;
  assign mem[1493] = mem_1493_sv2v_reg;
  assign mem[1492] = mem_1492_sv2v_reg;
  assign mem[1491] = mem_1491_sv2v_reg;
  assign mem[1490] = mem_1490_sv2v_reg;
  assign mem[1489] = mem_1489_sv2v_reg;
  assign mem[1488] = mem_1488_sv2v_reg;
  assign mem[1487] = mem_1487_sv2v_reg;
  assign mem[1486] = mem_1486_sv2v_reg;
  assign mem[1485] = mem_1485_sv2v_reg;
  assign mem[1484] = mem_1484_sv2v_reg;
  assign mem[1483] = mem_1483_sv2v_reg;
  assign mem[1482] = mem_1482_sv2v_reg;
  assign mem[1481] = mem_1481_sv2v_reg;
  assign mem[1480] = mem_1480_sv2v_reg;
  assign mem[1479] = mem_1479_sv2v_reg;
  assign mem[1478] = mem_1478_sv2v_reg;
  assign mem[1477] = mem_1477_sv2v_reg;
  assign mem[1476] = mem_1476_sv2v_reg;
  assign mem[1475] = mem_1475_sv2v_reg;
  assign mem[1474] = mem_1474_sv2v_reg;
  assign mem[1473] = mem_1473_sv2v_reg;
  assign mem[1472] = mem_1472_sv2v_reg;
  assign mem[1471] = mem_1471_sv2v_reg;
  assign mem[1470] = mem_1470_sv2v_reg;
  assign mem[1469] = mem_1469_sv2v_reg;
  assign mem[1468] = mem_1468_sv2v_reg;
  assign mem[1467] = mem_1467_sv2v_reg;
  assign mem[1466] = mem_1466_sv2v_reg;
  assign mem[1465] = mem_1465_sv2v_reg;
  assign mem[1464] = mem_1464_sv2v_reg;
  assign mem[1463] = mem_1463_sv2v_reg;
  assign mem[1462] = mem_1462_sv2v_reg;
  assign mem[1461] = mem_1461_sv2v_reg;
  assign mem[1460] = mem_1460_sv2v_reg;
  assign mem[1459] = mem_1459_sv2v_reg;
  assign mem[1458] = mem_1458_sv2v_reg;
  assign mem[1457] = mem_1457_sv2v_reg;
  assign mem[1456] = mem_1456_sv2v_reg;
  assign mem[1455] = mem_1455_sv2v_reg;
  assign mem[1454] = mem_1454_sv2v_reg;
  assign mem[1453] = mem_1453_sv2v_reg;
  assign mem[1452] = mem_1452_sv2v_reg;
  assign mem[1451] = mem_1451_sv2v_reg;
  assign mem[1450] = mem_1450_sv2v_reg;
  assign mem[1449] = mem_1449_sv2v_reg;
  assign mem[1448] = mem_1448_sv2v_reg;
  assign mem[1447] = mem_1447_sv2v_reg;
  assign mem[1446] = mem_1446_sv2v_reg;
  assign mem[1445] = mem_1445_sv2v_reg;
  assign mem[1444] = mem_1444_sv2v_reg;
  assign mem[1443] = mem_1443_sv2v_reg;
  assign mem[1442] = mem_1442_sv2v_reg;
  assign mem[1441] = mem_1441_sv2v_reg;
  assign mem[1440] = mem_1440_sv2v_reg;
  assign mem[1439] = mem_1439_sv2v_reg;
  assign mem[1438] = mem_1438_sv2v_reg;
  assign mem[1437] = mem_1437_sv2v_reg;
  assign mem[1436] = mem_1436_sv2v_reg;
  assign mem[1435] = mem_1435_sv2v_reg;
  assign mem[1434] = mem_1434_sv2v_reg;
  assign mem[1433] = mem_1433_sv2v_reg;
  assign mem[1432] = mem_1432_sv2v_reg;
  assign mem[1431] = mem_1431_sv2v_reg;
  assign mem[1430] = mem_1430_sv2v_reg;
  assign mem[1429] = mem_1429_sv2v_reg;
  assign mem[1428] = mem_1428_sv2v_reg;
  assign mem[1427] = mem_1427_sv2v_reg;
  assign mem[1426] = mem_1426_sv2v_reg;
  assign mem[1425] = mem_1425_sv2v_reg;
  assign mem[1424] = mem_1424_sv2v_reg;
  assign mem[1423] = mem_1423_sv2v_reg;
  assign mem[1422] = mem_1422_sv2v_reg;
  assign mem[1421] = mem_1421_sv2v_reg;
  assign mem[1420] = mem_1420_sv2v_reg;
  assign mem[1419] = mem_1419_sv2v_reg;
  assign mem[1418] = mem_1418_sv2v_reg;
  assign mem[1417] = mem_1417_sv2v_reg;
  assign mem[1416] = mem_1416_sv2v_reg;
  assign mem[1415] = mem_1415_sv2v_reg;
  assign mem[1414] = mem_1414_sv2v_reg;
  assign mem[1413] = mem_1413_sv2v_reg;
  assign mem[1412] = mem_1412_sv2v_reg;
  assign mem[1411] = mem_1411_sv2v_reg;
  assign mem[1410] = mem_1410_sv2v_reg;
  assign mem[1409] = mem_1409_sv2v_reg;
  assign mem[1408] = mem_1408_sv2v_reg;
  assign mem[1407] = mem_1407_sv2v_reg;
  assign mem[1406] = mem_1406_sv2v_reg;
  assign mem[1405] = mem_1405_sv2v_reg;
  assign mem[1404] = mem_1404_sv2v_reg;
  assign mem[1403] = mem_1403_sv2v_reg;
  assign mem[1402] = mem_1402_sv2v_reg;
  assign mem[1401] = mem_1401_sv2v_reg;
  assign mem[1400] = mem_1400_sv2v_reg;
  assign mem[1399] = mem_1399_sv2v_reg;
  assign mem[1398] = mem_1398_sv2v_reg;
  assign mem[1397] = mem_1397_sv2v_reg;
  assign mem[1396] = mem_1396_sv2v_reg;
  assign mem[1395] = mem_1395_sv2v_reg;
  assign mem[1394] = mem_1394_sv2v_reg;
  assign mem[1393] = mem_1393_sv2v_reg;
  assign mem[1392] = mem_1392_sv2v_reg;
  assign mem[1391] = mem_1391_sv2v_reg;
  assign mem[1390] = mem_1390_sv2v_reg;
  assign mem[1389] = mem_1389_sv2v_reg;
  assign mem[1388] = mem_1388_sv2v_reg;
  assign mem[1387] = mem_1387_sv2v_reg;
  assign mem[1386] = mem_1386_sv2v_reg;
  assign mem[1385] = mem_1385_sv2v_reg;
  assign mem[1384] = mem_1384_sv2v_reg;
  assign mem[1383] = mem_1383_sv2v_reg;
  assign mem[1382] = mem_1382_sv2v_reg;
  assign mem[1381] = mem_1381_sv2v_reg;
  assign mem[1380] = mem_1380_sv2v_reg;
  assign mem[1379] = mem_1379_sv2v_reg;
  assign mem[1378] = mem_1378_sv2v_reg;
  assign mem[1377] = mem_1377_sv2v_reg;
  assign mem[1376] = mem_1376_sv2v_reg;
  assign mem[1375] = mem_1375_sv2v_reg;
  assign mem[1374] = mem_1374_sv2v_reg;
  assign mem[1373] = mem_1373_sv2v_reg;
  assign mem[1372] = mem_1372_sv2v_reg;
  assign mem[1371] = mem_1371_sv2v_reg;
  assign mem[1370] = mem_1370_sv2v_reg;
  assign mem[1369] = mem_1369_sv2v_reg;
  assign mem[1368] = mem_1368_sv2v_reg;
  assign mem[1367] = mem_1367_sv2v_reg;
  assign mem[1366] = mem_1366_sv2v_reg;
  assign mem[1365] = mem_1365_sv2v_reg;
  assign mem[1364] = mem_1364_sv2v_reg;
  assign mem[1363] = mem_1363_sv2v_reg;
  assign mem[1362] = mem_1362_sv2v_reg;
  assign mem[1361] = mem_1361_sv2v_reg;
  assign mem[1360] = mem_1360_sv2v_reg;
  assign mem[1359] = mem_1359_sv2v_reg;
  assign mem[1358] = mem_1358_sv2v_reg;
  assign mem[1357] = mem_1357_sv2v_reg;
  assign mem[1356] = mem_1356_sv2v_reg;
  assign mem[1355] = mem_1355_sv2v_reg;
  assign mem[1354] = mem_1354_sv2v_reg;
  assign mem[1353] = mem_1353_sv2v_reg;
  assign mem[1352] = mem_1352_sv2v_reg;
  assign mem[1351] = mem_1351_sv2v_reg;
  assign mem[1350] = mem_1350_sv2v_reg;
  assign mem[1349] = mem_1349_sv2v_reg;
  assign mem[1348] = mem_1348_sv2v_reg;
  assign mem[1347] = mem_1347_sv2v_reg;
  assign mem[1346] = mem_1346_sv2v_reg;
  assign mem[1345] = mem_1345_sv2v_reg;
  assign mem[1344] = mem_1344_sv2v_reg;
  assign mem[1343] = mem_1343_sv2v_reg;
  assign mem[1342] = mem_1342_sv2v_reg;
  assign mem[1341] = mem_1341_sv2v_reg;
  assign mem[1340] = mem_1340_sv2v_reg;
  assign mem[1339] = mem_1339_sv2v_reg;
  assign mem[1338] = mem_1338_sv2v_reg;
  assign mem[1337] = mem_1337_sv2v_reg;
  assign mem[1336] = mem_1336_sv2v_reg;
  assign mem[1335] = mem_1335_sv2v_reg;
  assign mem[1334] = mem_1334_sv2v_reg;
  assign mem[1333] = mem_1333_sv2v_reg;
  assign mem[1332] = mem_1332_sv2v_reg;
  assign mem[1331] = mem_1331_sv2v_reg;
  assign mem[1330] = mem_1330_sv2v_reg;
  assign mem[1329] = mem_1329_sv2v_reg;
  assign mem[1328] = mem_1328_sv2v_reg;
  assign mem[1327] = mem_1327_sv2v_reg;
  assign mem[1326] = mem_1326_sv2v_reg;
  assign mem[1325] = mem_1325_sv2v_reg;
  assign mem[1324] = mem_1324_sv2v_reg;
  assign mem[1323] = mem_1323_sv2v_reg;
  assign mem[1322] = mem_1322_sv2v_reg;
  assign mem[1321] = mem_1321_sv2v_reg;
  assign mem[1320] = mem_1320_sv2v_reg;
  assign mem[1319] = mem_1319_sv2v_reg;
  assign mem[1318] = mem_1318_sv2v_reg;
  assign mem[1317] = mem_1317_sv2v_reg;
  assign mem[1316] = mem_1316_sv2v_reg;
  assign mem[1315] = mem_1315_sv2v_reg;
  assign mem[1314] = mem_1314_sv2v_reg;
  assign mem[1313] = mem_1313_sv2v_reg;
  assign mem[1312] = mem_1312_sv2v_reg;
  assign mem[1311] = mem_1311_sv2v_reg;
  assign mem[1310] = mem_1310_sv2v_reg;
  assign mem[1309] = mem_1309_sv2v_reg;
  assign mem[1308] = mem_1308_sv2v_reg;
  assign mem[1307] = mem_1307_sv2v_reg;
  assign mem[1306] = mem_1306_sv2v_reg;
  assign mem[1305] = mem_1305_sv2v_reg;
  assign mem[1304] = mem_1304_sv2v_reg;
  assign mem[1303] = mem_1303_sv2v_reg;
  assign mem[1302] = mem_1302_sv2v_reg;
  assign mem[1301] = mem_1301_sv2v_reg;
  assign mem[1300] = mem_1300_sv2v_reg;
  assign mem[1299] = mem_1299_sv2v_reg;
  assign mem[1298] = mem_1298_sv2v_reg;
  assign mem[1297] = mem_1297_sv2v_reg;
  assign mem[1296] = mem_1296_sv2v_reg;
  assign mem[1295] = mem_1295_sv2v_reg;
  assign mem[1294] = mem_1294_sv2v_reg;
  assign mem[1293] = mem_1293_sv2v_reg;
  assign mem[1292] = mem_1292_sv2v_reg;
  assign mem[1291] = mem_1291_sv2v_reg;
  assign mem[1290] = mem_1290_sv2v_reg;
  assign mem[1289] = mem_1289_sv2v_reg;
  assign mem[1288] = mem_1288_sv2v_reg;
  assign mem[1287] = mem_1287_sv2v_reg;
  assign mem[1286] = mem_1286_sv2v_reg;
  assign mem[1285] = mem_1285_sv2v_reg;
  assign mem[1284] = mem_1284_sv2v_reg;
  assign mem[1283] = mem_1283_sv2v_reg;
  assign mem[1282] = mem_1282_sv2v_reg;
  assign mem[1281] = mem_1281_sv2v_reg;
  assign mem[1280] = mem_1280_sv2v_reg;
  assign mem[1279] = mem_1279_sv2v_reg;
  assign mem[1278] = mem_1278_sv2v_reg;
  assign mem[1277] = mem_1277_sv2v_reg;
  assign mem[1276] = mem_1276_sv2v_reg;
  assign mem[1275] = mem_1275_sv2v_reg;
  assign mem[1274] = mem_1274_sv2v_reg;
  assign mem[1273] = mem_1273_sv2v_reg;
  assign mem[1272] = mem_1272_sv2v_reg;
  assign mem[1271] = mem_1271_sv2v_reg;
  assign mem[1270] = mem_1270_sv2v_reg;
  assign mem[1269] = mem_1269_sv2v_reg;
  assign mem[1268] = mem_1268_sv2v_reg;
  assign mem[1267] = mem_1267_sv2v_reg;
  assign mem[1266] = mem_1266_sv2v_reg;
  assign mem[1265] = mem_1265_sv2v_reg;
  assign mem[1264] = mem_1264_sv2v_reg;
  assign mem[1263] = mem_1263_sv2v_reg;
  assign mem[1262] = mem_1262_sv2v_reg;
  assign mem[1261] = mem_1261_sv2v_reg;
  assign mem[1260] = mem_1260_sv2v_reg;
  assign mem[1259] = mem_1259_sv2v_reg;
  assign mem[1258] = mem_1258_sv2v_reg;
  assign mem[1257] = mem_1257_sv2v_reg;
  assign mem[1256] = mem_1256_sv2v_reg;
  assign mem[1255] = mem_1255_sv2v_reg;
  assign mem[1254] = mem_1254_sv2v_reg;
  assign mem[1253] = mem_1253_sv2v_reg;
  assign mem[1252] = mem_1252_sv2v_reg;
  assign mem[1251] = mem_1251_sv2v_reg;
  assign mem[1250] = mem_1250_sv2v_reg;
  assign mem[1249] = mem_1249_sv2v_reg;
  assign mem[1248] = mem_1248_sv2v_reg;
  assign mem[1247] = mem_1247_sv2v_reg;
  assign mem[1246] = mem_1246_sv2v_reg;
  assign mem[1245] = mem_1245_sv2v_reg;
  assign mem[1244] = mem_1244_sv2v_reg;
  assign mem[1243] = mem_1243_sv2v_reg;
  assign mem[1242] = mem_1242_sv2v_reg;
  assign mem[1241] = mem_1241_sv2v_reg;
  assign mem[1240] = mem_1240_sv2v_reg;
  assign mem[1239] = mem_1239_sv2v_reg;
  assign mem[1238] = mem_1238_sv2v_reg;
  assign mem[1237] = mem_1237_sv2v_reg;
  assign mem[1236] = mem_1236_sv2v_reg;
  assign mem[1235] = mem_1235_sv2v_reg;
  assign mem[1234] = mem_1234_sv2v_reg;
  assign mem[1233] = mem_1233_sv2v_reg;
  assign mem[1232] = mem_1232_sv2v_reg;
  assign mem[1231] = mem_1231_sv2v_reg;
  assign mem[1230] = mem_1230_sv2v_reg;
  assign mem[1229] = mem_1229_sv2v_reg;
  assign mem[1228] = mem_1228_sv2v_reg;
  assign mem[1227] = mem_1227_sv2v_reg;
  assign mem[1226] = mem_1226_sv2v_reg;
  assign mem[1225] = mem_1225_sv2v_reg;
  assign mem[1224] = mem_1224_sv2v_reg;
  assign mem[1223] = mem_1223_sv2v_reg;
  assign mem[1222] = mem_1222_sv2v_reg;
  assign mem[1221] = mem_1221_sv2v_reg;
  assign mem[1220] = mem_1220_sv2v_reg;
  assign mem[1219] = mem_1219_sv2v_reg;
  assign mem[1218] = mem_1218_sv2v_reg;
  assign mem[1217] = mem_1217_sv2v_reg;
  assign mem[1216] = mem_1216_sv2v_reg;
  assign mem[1215] = mem_1215_sv2v_reg;
  assign mem[1214] = mem_1214_sv2v_reg;
  assign mem[1213] = mem_1213_sv2v_reg;
  assign mem[1212] = mem_1212_sv2v_reg;
  assign mem[1211] = mem_1211_sv2v_reg;
  assign mem[1210] = mem_1210_sv2v_reg;
  assign mem[1209] = mem_1209_sv2v_reg;
  assign mem[1208] = mem_1208_sv2v_reg;
  assign mem[1207] = mem_1207_sv2v_reg;
  assign mem[1206] = mem_1206_sv2v_reg;
  assign mem[1205] = mem_1205_sv2v_reg;
  assign mem[1204] = mem_1204_sv2v_reg;
  assign mem[1203] = mem_1203_sv2v_reg;
  assign mem[1202] = mem_1202_sv2v_reg;
  assign mem[1201] = mem_1201_sv2v_reg;
  assign mem[1200] = mem_1200_sv2v_reg;
  assign mem[1199] = mem_1199_sv2v_reg;
  assign mem[1198] = mem_1198_sv2v_reg;
  assign mem[1197] = mem_1197_sv2v_reg;
  assign mem[1196] = mem_1196_sv2v_reg;
  assign mem[1195] = mem_1195_sv2v_reg;
  assign mem[1194] = mem_1194_sv2v_reg;
  assign mem[1193] = mem_1193_sv2v_reg;
  assign mem[1192] = mem_1192_sv2v_reg;
  assign mem[1191] = mem_1191_sv2v_reg;
  assign mem[1190] = mem_1190_sv2v_reg;
  assign mem[1189] = mem_1189_sv2v_reg;
  assign mem[1188] = mem_1188_sv2v_reg;
  assign mem[1187] = mem_1187_sv2v_reg;
  assign mem[1186] = mem_1186_sv2v_reg;
  assign mem[1185] = mem_1185_sv2v_reg;
  assign mem[1184] = mem_1184_sv2v_reg;
  assign mem[1183] = mem_1183_sv2v_reg;
  assign mem[1182] = mem_1182_sv2v_reg;
  assign mem[1181] = mem_1181_sv2v_reg;
  assign mem[1180] = mem_1180_sv2v_reg;
  assign mem[1179] = mem_1179_sv2v_reg;
  assign mem[1178] = mem_1178_sv2v_reg;
  assign mem[1177] = mem_1177_sv2v_reg;
  assign mem[1176] = mem_1176_sv2v_reg;
  assign mem[1175] = mem_1175_sv2v_reg;
  assign mem[1174] = mem_1174_sv2v_reg;
  assign mem[1173] = mem_1173_sv2v_reg;
  assign mem[1172] = mem_1172_sv2v_reg;
  assign mem[1171] = mem_1171_sv2v_reg;
  assign mem[1170] = mem_1170_sv2v_reg;
  assign mem[1169] = mem_1169_sv2v_reg;
  assign mem[1168] = mem_1168_sv2v_reg;
  assign mem[1167] = mem_1167_sv2v_reg;
  assign mem[1166] = mem_1166_sv2v_reg;
  assign mem[1165] = mem_1165_sv2v_reg;
  assign mem[1164] = mem_1164_sv2v_reg;
  assign mem[1163] = mem_1163_sv2v_reg;
  assign mem[1162] = mem_1162_sv2v_reg;
  assign mem[1161] = mem_1161_sv2v_reg;
  assign mem[1160] = mem_1160_sv2v_reg;
  assign mem[1159] = mem_1159_sv2v_reg;
  assign mem[1158] = mem_1158_sv2v_reg;
  assign mem[1157] = mem_1157_sv2v_reg;
  assign mem[1156] = mem_1156_sv2v_reg;
  assign mem[1155] = mem_1155_sv2v_reg;
  assign mem[1154] = mem_1154_sv2v_reg;
  assign mem[1153] = mem_1153_sv2v_reg;
  assign mem[1152] = mem_1152_sv2v_reg;
  assign mem[1151] = mem_1151_sv2v_reg;
  assign mem[1150] = mem_1150_sv2v_reg;
  assign mem[1149] = mem_1149_sv2v_reg;
  assign mem[1148] = mem_1148_sv2v_reg;
  assign mem[1147] = mem_1147_sv2v_reg;
  assign mem[1146] = mem_1146_sv2v_reg;
  assign mem[1145] = mem_1145_sv2v_reg;
  assign mem[1144] = mem_1144_sv2v_reg;
  assign mem[1143] = mem_1143_sv2v_reg;
  assign mem[1142] = mem_1142_sv2v_reg;
  assign mem[1141] = mem_1141_sv2v_reg;
  assign mem[1140] = mem_1140_sv2v_reg;
  assign mem[1139] = mem_1139_sv2v_reg;
  assign mem[1138] = mem_1138_sv2v_reg;
  assign mem[1137] = mem_1137_sv2v_reg;
  assign mem[1136] = mem_1136_sv2v_reg;
  assign mem[1135] = mem_1135_sv2v_reg;
  assign mem[1134] = mem_1134_sv2v_reg;
  assign mem[1133] = mem_1133_sv2v_reg;
  assign mem[1132] = mem_1132_sv2v_reg;
  assign mem[1131] = mem_1131_sv2v_reg;
  assign mem[1130] = mem_1130_sv2v_reg;
  assign mem[1129] = mem_1129_sv2v_reg;
  assign mem[1128] = mem_1128_sv2v_reg;
  assign mem[1127] = mem_1127_sv2v_reg;
  assign mem[1126] = mem_1126_sv2v_reg;
  assign mem[1125] = mem_1125_sv2v_reg;
  assign mem[1124] = mem_1124_sv2v_reg;
  assign mem[1123] = mem_1123_sv2v_reg;
  assign mem[1122] = mem_1122_sv2v_reg;
  assign mem[1121] = mem_1121_sv2v_reg;
  assign mem[1120] = mem_1120_sv2v_reg;
  assign mem[1119] = mem_1119_sv2v_reg;
  assign mem[1118] = mem_1118_sv2v_reg;
  assign mem[1117] = mem_1117_sv2v_reg;
  assign mem[1116] = mem_1116_sv2v_reg;
  assign mem[1115] = mem_1115_sv2v_reg;
  assign mem[1114] = mem_1114_sv2v_reg;
  assign mem[1113] = mem_1113_sv2v_reg;
  assign mem[1112] = mem_1112_sv2v_reg;
  assign mem[1111] = mem_1111_sv2v_reg;
  assign mem[1110] = mem_1110_sv2v_reg;
  assign mem[1109] = mem_1109_sv2v_reg;
  assign mem[1108] = mem_1108_sv2v_reg;
  assign mem[1107] = mem_1107_sv2v_reg;
  assign mem[1106] = mem_1106_sv2v_reg;
  assign mem[1105] = mem_1105_sv2v_reg;
  assign mem[1104] = mem_1104_sv2v_reg;
  assign mem[1103] = mem_1103_sv2v_reg;
  assign mem[1102] = mem_1102_sv2v_reg;
  assign mem[1101] = mem_1101_sv2v_reg;
  assign mem[1100] = mem_1100_sv2v_reg;
  assign mem[1099] = mem_1099_sv2v_reg;
  assign mem[1098] = mem_1098_sv2v_reg;
  assign mem[1097] = mem_1097_sv2v_reg;
  assign mem[1096] = mem_1096_sv2v_reg;
  assign mem[1095] = mem_1095_sv2v_reg;
  assign mem[1094] = mem_1094_sv2v_reg;
  assign mem[1093] = mem_1093_sv2v_reg;
  assign mem[1092] = mem_1092_sv2v_reg;
  assign mem[1091] = mem_1091_sv2v_reg;
  assign mem[1090] = mem_1090_sv2v_reg;
  assign mem[1089] = mem_1089_sv2v_reg;
  assign mem[1088] = mem_1088_sv2v_reg;
  assign mem[1087] = mem_1087_sv2v_reg;
  assign mem[1086] = mem_1086_sv2v_reg;
  assign mem[1085] = mem_1085_sv2v_reg;
  assign mem[1084] = mem_1084_sv2v_reg;
  assign mem[1083] = mem_1083_sv2v_reg;
  assign mem[1082] = mem_1082_sv2v_reg;
  assign mem[1081] = mem_1081_sv2v_reg;
  assign mem[1080] = mem_1080_sv2v_reg;
  assign mem[1079] = mem_1079_sv2v_reg;
  assign mem[1078] = mem_1078_sv2v_reg;
  assign mem[1077] = mem_1077_sv2v_reg;
  assign mem[1076] = mem_1076_sv2v_reg;
  assign mem[1075] = mem_1075_sv2v_reg;
  assign mem[1074] = mem_1074_sv2v_reg;
  assign mem[1073] = mem_1073_sv2v_reg;
  assign mem[1072] = mem_1072_sv2v_reg;
  assign mem[1071] = mem_1071_sv2v_reg;
  assign mem[1070] = mem_1070_sv2v_reg;
  assign mem[1069] = mem_1069_sv2v_reg;
  assign mem[1068] = mem_1068_sv2v_reg;
  assign mem[1067] = mem_1067_sv2v_reg;
  assign mem[1066] = mem_1066_sv2v_reg;
  assign mem[1065] = mem_1065_sv2v_reg;
  assign mem[1064] = mem_1064_sv2v_reg;
  assign mem[1063] = mem_1063_sv2v_reg;
  assign mem[1062] = mem_1062_sv2v_reg;
  assign mem[1061] = mem_1061_sv2v_reg;
  assign mem[1060] = mem_1060_sv2v_reg;
  assign mem[1059] = mem_1059_sv2v_reg;
  assign mem[1058] = mem_1058_sv2v_reg;
  assign mem[1057] = mem_1057_sv2v_reg;
  assign mem[1056] = mem_1056_sv2v_reg;
  assign mem[1055] = mem_1055_sv2v_reg;
  assign mem[1054] = mem_1054_sv2v_reg;
  assign mem[1053] = mem_1053_sv2v_reg;
  assign mem[1052] = mem_1052_sv2v_reg;
  assign mem[1051] = mem_1051_sv2v_reg;
  assign mem[1050] = mem_1050_sv2v_reg;
  assign mem[1049] = mem_1049_sv2v_reg;
  assign mem[1048] = mem_1048_sv2v_reg;
  assign mem[1047] = mem_1047_sv2v_reg;
  assign mem[1046] = mem_1046_sv2v_reg;
  assign mem[1045] = mem_1045_sv2v_reg;
  assign mem[1044] = mem_1044_sv2v_reg;
  assign mem[1043] = mem_1043_sv2v_reg;
  assign mem[1042] = mem_1042_sv2v_reg;
  assign mem[1041] = mem_1041_sv2v_reg;
  assign mem[1040] = mem_1040_sv2v_reg;
  assign mem[1039] = mem_1039_sv2v_reg;
  assign mem[1038] = mem_1038_sv2v_reg;
  assign mem[1037] = mem_1037_sv2v_reg;
  assign mem[1036] = mem_1036_sv2v_reg;
  assign mem[1035] = mem_1035_sv2v_reg;
  assign mem[1034] = mem_1034_sv2v_reg;
  assign mem[1033] = mem_1033_sv2v_reg;
  assign mem[1032] = mem_1032_sv2v_reg;
  assign mem[1031] = mem_1031_sv2v_reg;
  assign mem[1030] = mem_1030_sv2v_reg;
  assign mem[1029] = mem_1029_sv2v_reg;
  assign mem[1028] = mem_1028_sv2v_reg;
  assign mem[1027] = mem_1027_sv2v_reg;
  assign mem[1026] = mem_1026_sv2v_reg;
  assign mem[1025] = mem_1025_sv2v_reg;
  assign mem[1024] = mem_1024_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign N424 = ~w_addr_i[5];
  assign N425 = w_addr_i[3] & w_addr_i[4];
  assign N426 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N427 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N428 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N429 = w_addr_i[5] & N426;
  assign N430 = w_addr_i[5] & N427;
  assign N431 = w_addr_i[5] & N428;
  assign N432 = N424 & N425;
  assign N433 = N424 & N426;
  assign N434 = N424 & N427;
  assign N435 = N424 & N428;
  assign N436 = ~w_addr_i[2];
  assign N437 = w_addr_i[0] & w_addr_i[1];
  assign N438 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N439 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N440 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N441 = w_addr_i[2] & N437;
  assign N442 = w_addr_i[2] & N438;
  assign N443 = w_addr_i[2] & N439;
  assign N444 = w_addr_i[2] & N440;
  assign N445 = N436 & N437;
  assign N446 = N436 & N438;
  assign N447 = N436 & N439;
  assign N448 = N436 & N440;
  assign N373 = N429 & N447;
  assign N372 = N429 & N448;
  assign N371 = N430 & N441;
  assign N370 = N430 & N442;
  assign N369 = N430 & N443;
  assign N368 = N430 & N444;
  assign N367 = N430 & N445;
  assign N366 = N430 & N446;
  assign N365 = N430 & N447;
  assign N364 = N430 & N448;
  assign N363 = N431 & N441;
  assign N362 = N431 & N442;
  assign N361 = N431 & N443;
  assign N360 = N431 & N444;
  assign N359 = N431 & N445;
  assign N358 = N431 & N446;
  assign N357 = N431 & N447;
  assign N356 = N431 & N448;
  assign N355 = N432 & N441;
  assign N354 = N432 & N442;
  assign N353 = N432 & N443;
  assign N352 = N432 & N444;
  assign N351 = N432 & N445;
  assign N350 = N432 & N446;
  assign N349 = N432 & N447;
  assign N348 = N432 & N448;
  assign N347 = N433 & N441;
  assign N346 = N433 & N442;
  assign N345 = N433 & N443;
  assign N344 = N433 & N444;
  assign N343 = N433 & N445;
  assign N342 = N433 & N446;
  assign N341 = N433 & N447;
  assign N340 = N433 & N448;
  assign N339 = N434 & N441;
  assign N338 = N434 & N442;
  assign N337 = N434 & N443;
  assign N336 = N434 & N444;
  assign N335 = N434 & N445;
  assign N334 = N434 & N446;
  assign N333 = N434 & N447;
  assign N332 = N434 & N448;
  assign N331 = N435 & N441;
  assign N330 = N435 & N442;
  assign N329 = N435 & N443;
  assign N328 = N435 & N444;
  assign N327 = N435 & N445;
  assign N326 = N435 & N446;
  assign N325 = N435 & N447;
  assign N324 = N435 & N448;
  assign N8 = N12 & N13;
  assign N9 = N8 & N14;
  assign N10 = N9 & N15;
  assign N11 = N10 & N16;
  assign N273 = N11 & N17;
  assign N12 = ~r_addr_i[5];
  assign N13 = ~r_addr_i[4];
  assign N14 = ~r_addr_i[3];
  assign N15 = ~r_addr_i[2];
  assign N16 = ~r_addr_i[0];
  assign N17 = ~r_addr_i[1];
  assign N18 = r_addr_i[5] & N22;
  assign N19 = N18 & N23;
  assign N20 = N19 & N24;
  assign N21 = N20 & N25;
  assign N274 = N21 & N26;
  assign N22 = ~r_addr_i[4];
  assign N23 = ~r_addr_i[3];
  assign N24 = ~r_addr_i[2];
  assign N25 = ~r_addr_i[0];
  assign N26 = ~r_addr_i[1];
  assign N27 = N31 & N32;
  assign N28 = N27 & N33;
  assign N29 = N28 & N34;
  assign N30 = N29 & r_addr_i[0];
  assign N275 = N30 & N35;
  assign N31 = ~r_addr_i[5];
  assign N32 = ~r_addr_i[4];
  assign N33 = ~r_addr_i[3];
  assign N34 = ~r_addr_i[2];
  assign N35 = ~r_addr_i[1];
  assign N36 = N40 & N41;
  assign N37 = N36 & N42;
  assign N38 = N37 & N43;
  assign N39 = N38 & N44;
  assign N277 = N39 & r_addr_i[1];
  assign N40 = ~r_addr_i[5];
  assign N41 = ~r_addr_i[4];
  assign N42 = ~r_addr_i[3];
  assign N43 = ~r_addr_i[2];
  assign N44 = ~r_addr_i[0];
  assign N45 = N49 & N50;
  assign N46 = N45 & N51;
  assign N47 = N46 & N52;
  assign N48 = N47 & r_addr_i[0];
  assign N279 = N48 & r_addr_i[1];
  assign N49 = ~r_addr_i[5];
  assign N50 = ~r_addr_i[4];
  assign N51 = ~r_addr_i[3];
  assign N52 = ~r_addr_i[2];
  assign N53 = N57 & N58;
  assign N54 = N53 & N59;
  assign N55 = N54 & r_addr_i[2];
  assign N56 = N55 & N60;
  assign N281 = N56 & N61;
  assign N57 = ~r_addr_i[5];
  assign N58 = ~r_addr_i[4];
  assign N59 = ~r_addr_i[3];
  assign N60 = ~r_addr_i[0];
  assign N61 = ~r_addr_i[1];
  assign N62 = N66 & N67;
  assign N63 = N62 & N68;
  assign N64 = N63 & r_addr_i[2];
  assign N65 = N64 & r_addr_i[0];
  assign N283 = N65 & N69;
  assign N66 = ~r_addr_i[5];
  assign N67 = ~r_addr_i[4];
  assign N68 = ~r_addr_i[3];
  assign N69 = ~r_addr_i[1];
  assign N70 = N74 & N75;
  assign N71 = N70 & N76;
  assign N72 = N71 & r_addr_i[2];
  assign N73 = N72 & N77;
  assign N285 = N73 & r_addr_i[1];
  assign N74 = ~r_addr_i[5];
  assign N75 = ~r_addr_i[4];
  assign N76 = ~r_addr_i[3];
  assign N77 = ~r_addr_i[0];
  assign N78 = N82 & N83;
  assign N79 = N78 & N84;
  assign N80 = N79 & r_addr_i[2];
  assign N81 = N80 & r_addr_i[0];
  assign N287 = N81 & r_addr_i[1];
  assign N82 = ~r_addr_i[5];
  assign N83 = ~r_addr_i[4];
  assign N84 = ~r_addr_i[3];
  assign N85 = N89 & N90;
  assign N86 = N85 & r_addr_i[3];
  assign N87 = N86 & N91;
  assign N88 = N87 & N92;
  assign N289 = N88 & N93;
  assign N89 = ~r_addr_i[5];
  assign N90 = ~r_addr_i[4];
  assign N91 = ~r_addr_i[2];
  assign N92 = ~r_addr_i[0];
  assign N93 = ~r_addr_i[1];
  assign N94 = N98 & N99;
  assign N95 = N94 & r_addr_i[3];
  assign N96 = N95 & N100;
  assign N97 = N96 & r_addr_i[0];
  assign N291 = N97 & N101;
  assign N98 = ~r_addr_i[5];
  assign N99 = ~r_addr_i[4];
  assign N100 = ~r_addr_i[2];
  assign N101 = ~r_addr_i[1];
  assign N102 = N106 & N107;
  assign N103 = N102 & r_addr_i[3];
  assign N104 = N103 & N108;
  assign N105 = N104 & N109;
  assign N293 = N105 & r_addr_i[1];
  assign N106 = ~r_addr_i[5];
  assign N107 = ~r_addr_i[4];
  assign N108 = ~r_addr_i[2];
  assign N109 = ~r_addr_i[0];
  assign N110 = N114 & N115;
  assign N111 = N110 & r_addr_i[3];
  assign N112 = N111 & N116;
  assign N113 = N112 & r_addr_i[0];
  assign N295 = N113 & r_addr_i[1];
  assign N114 = ~r_addr_i[5];
  assign N115 = ~r_addr_i[4];
  assign N116 = ~r_addr_i[2];
  assign N117 = N121 & N122;
  assign N118 = N117 & r_addr_i[3];
  assign N119 = N118 & r_addr_i[2];
  assign N120 = N119 & N123;
  assign N297 = N120 & N124;
  assign N121 = ~r_addr_i[5];
  assign N122 = ~r_addr_i[4];
  assign N123 = ~r_addr_i[0];
  assign N124 = ~r_addr_i[1];
  assign N125 = N129 & N130;
  assign N126 = N125 & r_addr_i[3];
  assign N127 = N126 & r_addr_i[2];
  assign N128 = N127 & r_addr_i[0];
  assign N299 = N128 & N131;
  assign N129 = ~r_addr_i[5];
  assign N130 = ~r_addr_i[4];
  assign N131 = ~r_addr_i[1];
  assign N132 = N136 & N137;
  assign N133 = N132 & r_addr_i[3];
  assign N134 = N133 & r_addr_i[2];
  assign N135 = N134 & N138;
  assign N301 = N135 & r_addr_i[1];
  assign N136 = ~r_addr_i[5];
  assign N137 = ~r_addr_i[4];
  assign N138 = ~r_addr_i[0];
  assign N139 = N143 & N144;
  assign N140 = N139 & r_addr_i[3];
  assign N141 = N140 & r_addr_i[2];
  assign N142 = N141 & r_addr_i[0];
  assign N303 = N142 & r_addr_i[1];
  assign N143 = ~r_addr_i[5];
  assign N144 = ~r_addr_i[4];
  assign N145 = N149 & r_addr_i[4];
  assign N146 = N145 & N150;
  assign N147 = N146 & N151;
  assign N148 = N147 & N152;
  assign N305 = N148 & N153;
  assign N149 = ~r_addr_i[5];
  assign N150 = ~r_addr_i[3];
  assign N151 = ~r_addr_i[2];
  assign N152 = ~r_addr_i[0];
  assign N153 = ~r_addr_i[1];
  assign N154 = N158 & r_addr_i[4];
  assign N155 = N154 & N159;
  assign N156 = N155 & N160;
  assign N157 = N156 & r_addr_i[0];
  assign N307 = N157 & N161;
  assign N158 = ~r_addr_i[5];
  assign N159 = ~r_addr_i[3];
  assign N160 = ~r_addr_i[2];
  assign N161 = ~r_addr_i[1];
  assign N309 = r_addr_i[4] & N162 & (N163 & N164) & r_addr_i[1];
  assign N162 = ~r_addr_i[3];
  assign N163 = ~r_addr_i[2];
  assign N164 = ~r_addr_i[0];
  assign N310 = r_addr_i[4] & N165 & (N166 & r_addr_i[0]) & r_addr_i[1];
  assign N165 = ~r_addr_i[3];
  assign N166 = ~r_addr_i[2];
  assign N311 = r_addr_i[4] & N167 & (r_addr_i[2] & N168) & N169;
  assign N167 = ~r_addr_i[3];
  assign N168 = ~r_addr_i[0];
  assign N169 = ~r_addr_i[1];
  assign N312 = r_addr_i[4] & N170 & (r_addr_i[2] & r_addr_i[0]) & N171;
  assign N170 = ~r_addr_i[3];
  assign N171 = ~r_addr_i[1];
  assign N313 = r_addr_i[4] & N172 & (r_addr_i[2] & N173) & r_addr_i[1];
  assign N172 = ~r_addr_i[3];
  assign N173 = ~r_addr_i[0];
  assign N314 = r_addr_i[4] & N174 & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N174 = ~r_addr_i[3];
  assign N315 = r_addr_i[4] & r_addr_i[3] & (N175 & N176) & N177;
  assign N175 = ~r_addr_i[2];
  assign N176 = ~r_addr_i[0];
  assign N177 = ~r_addr_i[1];
  assign N316 = r_addr_i[4] & r_addr_i[3] & (N178 & r_addr_i[0]) & N179;
  assign N178 = ~r_addr_i[2];
  assign N179 = ~r_addr_i[1];
  assign N317 = r_addr_i[4] & r_addr_i[3] & (N180 & N181) & r_addr_i[1];
  assign N180 = ~r_addr_i[2];
  assign N181 = ~r_addr_i[0];
  assign N318 = r_addr_i[4] & r_addr_i[3] & (N182 & r_addr_i[0]) & r_addr_i[1];
  assign N182 = ~r_addr_i[2];
  assign N319 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & N183) & N184;
  assign N183 = ~r_addr_i[0];
  assign N184 = ~r_addr_i[1];
  assign N320 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & N185;
  assign N185 = ~r_addr_i[1];
  assign N321 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & N186) & r_addr_i[1];
  assign N186 = ~r_addr_i[0];
  assign N322 = r_addr_i[4] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N187 = r_addr_i[5] & N191;
  assign N188 = N187 & N192;
  assign N189 = N188 & N193;
  assign N190 = N189 & r_addr_i[0];
  assign N276 = N190 & N194;
  assign N191 = ~r_addr_i[4];
  assign N192 = ~r_addr_i[3];
  assign N193 = ~r_addr_i[2];
  assign N194 = ~r_addr_i[1];
  assign N278 = r_addr_i[5] & N195 & (N196 & N197) & r_addr_i[1];
  assign N195 = ~r_addr_i[3];
  assign N196 = ~r_addr_i[2];
  assign N197 = ~r_addr_i[0];
  assign N280 = r_addr_i[5] & N198 & (N199 & r_addr_i[0]) & r_addr_i[1];
  assign N198 = ~r_addr_i[3];
  assign N199 = ~r_addr_i[2];
  assign N282 = r_addr_i[5] & N200 & (r_addr_i[2] & N201) & N202;
  assign N200 = ~r_addr_i[3];
  assign N201 = ~r_addr_i[0];
  assign N202 = ~r_addr_i[1];
  assign N284 = r_addr_i[5] & N203 & (r_addr_i[2] & r_addr_i[0]) & N204;
  assign N203 = ~r_addr_i[3];
  assign N204 = ~r_addr_i[1];
  assign N286 = r_addr_i[5] & N205 & (r_addr_i[2] & N206) & r_addr_i[1];
  assign N205 = ~r_addr_i[3];
  assign N206 = ~r_addr_i[0];
  assign N288 = r_addr_i[5] & N207 & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N207 = ~r_addr_i[3];
  assign N290 = r_addr_i[5] & r_addr_i[3] & (N208 & N209) & N210;
  assign N208 = ~r_addr_i[2];
  assign N209 = ~r_addr_i[0];
  assign N210 = ~r_addr_i[1];
  assign N292 = r_addr_i[5] & r_addr_i[3] & (N211 & r_addr_i[0]) & N212;
  assign N211 = ~r_addr_i[2];
  assign N212 = ~r_addr_i[1];
  assign N294 = r_addr_i[5] & r_addr_i[3] & (N213 & N214) & r_addr_i[1];
  assign N213 = ~r_addr_i[2];
  assign N214 = ~r_addr_i[0];
  assign N296 = r_addr_i[5] & r_addr_i[3] & (N215 & r_addr_i[0]) & r_addr_i[1];
  assign N215 = ~r_addr_i[2];
  assign N298 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & N216) & N217;
  assign N216 = ~r_addr_i[0];
  assign N217 = ~r_addr_i[1];
  assign N300 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & N218;
  assign N218 = ~r_addr_i[1];
  assign N302 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & N219) & r_addr_i[1];
  assign N219 = ~r_addr_i[0];
  assign N304 = r_addr_i[5] & r_addr_i[3] & (r_addr_i[2] & r_addr_i[0]) & r_addr_i[1];
  assign N306 = r_addr_i[5] & r_addr_i[4] & N220;
  assign N220 = ~r_addr_i[0];
  assign N308 = r_addr_i[5] & r_addr_i[4] & r_addr_i[0];
  assign { N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374 } = (N221)? { N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324 } : 
                                                                                                                                                                                                                                                                                                                          (N222)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N221 = w_v_i;
  assign N222 = N323;
  assign r_data_o[31] = (N223)? mem[31] : 
                        (N224)? mem[63] : 
                        (N225)? mem[95] : 
                        (N226)? mem[127] : 
                        (N227)? mem[159] : 
                        (N228)? mem[191] : 
                        (N229)? mem[223] : 
                        (N230)? mem[255] : 
                        (N231)? mem[287] : 
                        (N232)? mem[319] : 
                        (N233)? mem[351] : 
                        (N234)? mem[383] : 
                        (N235)? mem[415] : 
                        (N236)? mem[447] : 
                        (N237)? mem[479] : 
                        (N238)? mem[511] : 
                        (N239)? mem[543] : 
                        (N240)? mem[575] : 
                        (N241)? mem[607] : 
                        (N242)? mem[639] : 
                        (N243)? mem[671] : 
                        (N244)? mem[703] : 
                        (N245)? mem[735] : 
                        (N246)? mem[767] : 
                        (N247)? mem[799] : 
                        (N248)? mem[831] : 
                        (N249)? mem[863] : 
                        (N250)? mem[895] : 
                        (N251)? mem[927] : 
                        (N252)? mem[959] : 
                        (N253)? mem[991] : 
                        (N254)? mem[1023] : 
                        (N255)? mem[1055] : 
                        (N256)? mem[1087] : 
                        (N257)? mem[1119] : 
                        (N258)? mem[1151] : 
                        (N259)? mem[1183] : 
                        (N260)? mem[1215] : 
                        (N261)? mem[1247] : 
                        (N262)? mem[1279] : 
                        (N263)? mem[1311] : 
                        (N264)? mem[1343] : 
                        (N265)? mem[1375] : 
                        (N266)? mem[1407] : 
                        (N267)? mem[1439] : 
                        (N268)? mem[1471] : 
                        (N269)? mem[1503] : 
                        (N270)? mem[1535] : 
                        (N271)? mem[1567] : 
                        (N272)? mem[1599] : 1'b0;
  assign N223 = N273;
  assign N224 = N275;
  assign N225 = N277;
  assign N226 = N279;
  assign N227 = N281;
  assign N228 = N283;
  assign N229 = N285;
  assign N230 = N287;
  assign N231 = N289;
  assign N232 = N291;
  assign N233 = N293;
  assign N234 = N295;
  assign N235 = N297;
  assign N236 = N299;
  assign N237 = N301;
  assign N238 = N303;
  assign N239 = N305;
  assign N240 = N307;
  assign N241 = N309;
  assign N242 = N310;
  assign N243 = N311;
  assign N244 = N312;
  assign N245 = N313;
  assign N246 = N314;
  assign N247 = N315;
  assign N248 = N316;
  assign N249 = N317;
  assign N250 = N318;
  assign N251 = N319;
  assign N252 = N320;
  assign N253 = N321;
  assign N254 = N322;
  assign N255 = N274;
  assign N256 = N276;
  assign N257 = N278;
  assign N258 = N280;
  assign N259 = N282;
  assign N260 = N284;
  assign N261 = N286;
  assign N262 = N288;
  assign N263 = N290;
  assign N264 = N292;
  assign N265 = N294;
  assign N266 = N296;
  assign N267 = N298;
  assign N268 = N300;
  assign N269 = N302;
  assign N270 = N304;
  assign N271 = N306;
  assign N272 = N308;
  assign r_data_o[30] = (N223)? mem[30] : 
                        (N224)? mem[62] : 
                        (N225)? mem[94] : 
                        (N226)? mem[126] : 
                        (N227)? mem[158] : 
                        (N228)? mem[190] : 
                        (N229)? mem[222] : 
                        (N230)? mem[254] : 
                        (N231)? mem[286] : 
                        (N232)? mem[318] : 
                        (N233)? mem[350] : 
                        (N234)? mem[382] : 
                        (N235)? mem[414] : 
                        (N236)? mem[446] : 
                        (N237)? mem[478] : 
                        (N238)? mem[510] : 
                        (N239)? mem[542] : 
                        (N240)? mem[574] : 
                        (N241)? mem[606] : 
                        (N242)? mem[638] : 
                        (N243)? mem[670] : 
                        (N244)? mem[702] : 
                        (N245)? mem[734] : 
                        (N246)? mem[766] : 
                        (N247)? mem[798] : 
                        (N248)? mem[830] : 
                        (N249)? mem[862] : 
                        (N250)? mem[894] : 
                        (N251)? mem[926] : 
                        (N252)? mem[958] : 
                        (N253)? mem[990] : 
                        (N254)? mem[1022] : 
                        (N255)? mem[1054] : 
                        (N256)? mem[1086] : 
                        (N257)? mem[1118] : 
                        (N258)? mem[1150] : 
                        (N259)? mem[1182] : 
                        (N260)? mem[1214] : 
                        (N261)? mem[1246] : 
                        (N262)? mem[1278] : 
                        (N263)? mem[1310] : 
                        (N264)? mem[1342] : 
                        (N265)? mem[1374] : 
                        (N266)? mem[1406] : 
                        (N267)? mem[1438] : 
                        (N268)? mem[1470] : 
                        (N269)? mem[1502] : 
                        (N270)? mem[1534] : 
                        (N271)? mem[1566] : 
                        (N272)? mem[1598] : 1'b0;
  assign r_data_o[29] = (N223)? mem[29] : 
                        (N224)? mem[61] : 
                        (N225)? mem[93] : 
                        (N226)? mem[125] : 
                        (N227)? mem[157] : 
                        (N228)? mem[189] : 
                        (N229)? mem[221] : 
                        (N230)? mem[253] : 
                        (N231)? mem[285] : 
                        (N232)? mem[317] : 
                        (N233)? mem[349] : 
                        (N234)? mem[381] : 
                        (N235)? mem[413] : 
                        (N236)? mem[445] : 
                        (N237)? mem[477] : 
                        (N238)? mem[509] : 
                        (N239)? mem[541] : 
                        (N240)? mem[573] : 
                        (N241)? mem[605] : 
                        (N242)? mem[637] : 
                        (N243)? mem[669] : 
                        (N244)? mem[701] : 
                        (N245)? mem[733] : 
                        (N246)? mem[765] : 
                        (N247)? mem[797] : 
                        (N248)? mem[829] : 
                        (N249)? mem[861] : 
                        (N250)? mem[893] : 
                        (N251)? mem[925] : 
                        (N252)? mem[957] : 
                        (N253)? mem[989] : 
                        (N254)? mem[1021] : 
                        (N255)? mem[1053] : 
                        (N256)? mem[1085] : 
                        (N257)? mem[1117] : 
                        (N258)? mem[1149] : 
                        (N259)? mem[1181] : 
                        (N260)? mem[1213] : 
                        (N261)? mem[1245] : 
                        (N262)? mem[1277] : 
                        (N263)? mem[1309] : 
                        (N264)? mem[1341] : 
                        (N265)? mem[1373] : 
                        (N266)? mem[1405] : 
                        (N267)? mem[1437] : 
                        (N268)? mem[1469] : 
                        (N269)? mem[1501] : 
                        (N270)? mem[1533] : 
                        (N271)? mem[1565] : 
                        (N272)? mem[1597] : 1'b0;
  assign r_data_o[28] = (N223)? mem[28] : 
                        (N224)? mem[60] : 
                        (N225)? mem[92] : 
                        (N226)? mem[124] : 
                        (N227)? mem[156] : 
                        (N228)? mem[188] : 
                        (N229)? mem[220] : 
                        (N230)? mem[252] : 
                        (N231)? mem[284] : 
                        (N232)? mem[316] : 
                        (N233)? mem[348] : 
                        (N234)? mem[380] : 
                        (N235)? mem[412] : 
                        (N236)? mem[444] : 
                        (N237)? mem[476] : 
                        (N238)? mem[508] : 
                        (N239)? mem[540] : 
                        (N240)? mem[572] : 
                        (N241)? mem[604] : 
                        (N242)? mem[636] : 
                        (N243)? mem[668] : 
                        (N244)? mem[700] : 
                        (N245)? mem[732] : 
                        (N246)? mem[764] : 
                        (N247)? mem[796] : 
                        (N248)? mem[828] : 
                        (N249)? mem[860] : 
                        (N250)? mem[892] : 
                        (N251)? mem[924] : 
                        (N252)? mem[956] : 
                        (N253)? mem[988] : 
                        (N254)? mem[1020] : 
                        (N255)? mem[1052] : 
                        (N256)? mem[1084] : 
                        (N257)? mem[1116] : 
                        (N258)? mem[1148] : 
                        (N259)? mem[1180] : 
                        (N260)? mem[1212] : 
                        (N261)? mem[1244] : 
                        (N262)? mem[1276] : 
                        (N263)? mem[1308] : 
                        (N264)? mem[1340] : 
                        (N265)? mem[1372] : 
                        (N266)? mem[1404] : 
                        (N267)? mem[1436] : 
                        (N268)? mem[1468] : 
                        (N269)? mem[1500] : 
                        (N270)? mem[1532] : 
                        (N271)? mem[1564] : 
                        (N272)? mem[1596] : 1'b0;
  assign r_data_o[27] = (N223)? mem[27] : 
                        (N224)? mem[59] : 
                        (N225)? mem[91] : 
                        (N226)? mem[123] : 
                        (N227)? mem[155] : 
                        (N228)? mem[187] : 
                        (N229)? mem[219] : 
                        (N230)? mem[251] : 
                        (N231)? mem[283] : 
                        (N232)? mem[315] : 
                        (N233)? mem[347] : 
                        (N234)? mem[379] : 
                        (N235)? mem[411] : 
                        (N236)? mem[443] : 
                        (N237)? mem[475] : 
                        (N238)? mem[507] : 
                        (N239)? mem[539] : 
                        (N240)? mem[571] : 
                        (N241)? mem[603] : 
                        (N242)? mem[635] : 
                        (N243)? mem[667] : 
                        (N244)? mem[699] : 
                        (N245)? mem[731] : 
                        (N246)? mem[763] : 
                        (N247)? mem[795] : 
                        (N248)? mem[827] : 
                        (N249)? mem[859] : 
                        (N250)? mem[891] : 
                        (N251)? mem[923] : 
                        (N252)? mem[955] : 
                        (N253)? mem[987] : 
                        (N254)? mem[1019] : 
                        (N255)? mem[1051] : 
                        (N256)? mem[1083] : 
                        (N257)? mem[1115] : 
                        (N258)? mem[1147] : 
                        (N259)? mem[1179] : 
                        (N260)? mem[1211] : 
                        (N261)? mem[1243] : 
                        (N262)? mem[1275] : 
                        (N263)? mem[1307] : 
                        (N264)? mem[1339] : 
                        (N265)? mem[1371] : 
                        (N266)? mem[1403] : 
                        (N267)? mem[1435] : 
                        (N268)? mem[1467] : 
                        (N269)? mem[1499] : 
                        (N270)? mem[1531] : 
                        (N271)? mem[1563] : 
                        (N272)? mem[1595] : 1'b0;
  assign r_data_o[26] = (N223)? mem[26] : 
                        (N224)? mem[58] : 
                        (N225)? mem[90] : 
                        (N226)? mem[122] : 
                        (N227)? mem[154] : 
                        (N228)? mem[186] : 
                        (N229)? mem[218] : 
                        (N230)? mem[250] : 
                        (N231)? mem[282] : 
                        (N232)? mem[314] : 
                        (N233)? mem[346] : 
                        (N234)? mem[378] : 
                        (N235)? mem[410] : 
                        (N236)? mem[442] : 
                        (N237)? mem[474] : 
                        (N238)? mem[506] : 
                        (N239)? mem[538] : 
                        (N240)? mem[570] : 
                        (N241)? mem[602] : 
                        (N242)? mem[634] : 
                        (N243)? mem[666] : 
                        (N244)? mem[698] : 
                        (N245)? mem[730] : 
                        (N246)? mem[762] : 
                        (N247)? mem[794] : 
                        (N248)? mem[826] : 
                        (N249)? mem[858] : 
                        (N250)? mem[890] : 
                        (N251)? mem[922] : 
                        (N252)? mem[954] : 
                        (N253)? mem[986] : 
                        (N254)? mem[1018] : 
                        (N255)? mem[1050] : 
                        (N256)? mem[1082] : 
                        (N257)? mem[1114] : 
                        (N258)? mem[1146] : 
                        (N259)? mem[1178] : 
                        (N260)? mem[1210] : 
                        (N261)? mem[1242] : 
                        (N262)? mem[1274] : 
                        (N263)? mem[1306] : 
                        (N264)? mem[1338] : 
                        (N265)? mem[1370] : 
                        (N266)? mem[1402] : 
                        (N267)? mem[1434] : 
                        (N268)? mem[1466] : 
                        (N269)? mem[1498] : 
                        (N270)? mem[1530] : 
                        (N271)? mem[1562] : 
                        (N272)? mem[1594] : 1'b0;
  assign r_data_o[25] = (N223)? mem[25] : 
                        (N224)? mem[57] : 
                        (N225)? mem[89] : 
                        (N226)? mem[121] : 
                        (N227)? mem[153] : 
                        (N228)? mem[185] : 
                        (N229)? mem[217] : 
                        (N230)? mem[249] : 
                        (N231)? mem[281] : 
                        (N232)? mem[313] : 
                        (N233)? mem[345] : 
                        (N234)? mem[377] : 
                        (N235)? mem[409] : 
                        (N236)? mem[441] : 
                        (N237)? mem[473] : 
                        (N238)? mem[505] : 
                        (N239)? mem[537] : 
                        (N240)? mem[569] : 
                        (N241)? mem[601] : 
                        (N242)? mem[633] : 
                        (N243)? mem[665] : 
                        (N244)? mem[697] : 
                        (N245)? mem[729] : 
                        (N246)? mem[761] : 
                        (N247)? mem[793] : 
                        (N248)? mem[825] : 
                        (N249)? mem[857] : 
                        (N250)? mem[889] : 
                        (N251)? mem[921] : 
                        (N252)? mem[953] : 
                        (N253)? mem[985] : 
                        (N254)? mem[1017] : 
                        (N255)? mem[1049] : 
                        (N256)? mem[1081] : 
                        (N257)? mem[1113] : 
                        (N258)? mem[1145] : 
                        (N259)? mem[1177] : 
                        (N260)? mem[1209] : 
                        (N261)? mem[1241] : 
                        (N262)? mem[1273] : 
                        (N263)? mem[1305] : 
                        (N264)? mem[1337] : 
                        (N265)? mem[1369] : 
                        (N266)? mem[1401] : 
                        (N267)? mem[1433] : 
                        (N268)? mem[1465] : 
                        (N269)? mem[1497] : 
                        (N270)? mem[1529] : 
                        (N271)? mem[1561] : 
                        (N272)? mem[1593] : 1'b0;
  assign r_data_o[24] = (N223)? mem[24] : 
                        (N224)? mem[56] : 
                        (N225)? mem[88] : 
                        (N226)? mem[120] : 
                        (N227)? mem[152] : 
                        (N228)? mem[184] : 
                        (N229)? mem[216] : 
                        (N230)? mem[248] : 
                        (N231)? mem[280] : 
                        (N232)? mem[312] : 
                        (N233)? mem[344] : 
                        (N234)? mem[376] : 
                        (N235)? mem[408] : 
                        (N236)? mem[440] : 
                        (N237)? mem[472] : 
                        (N238)? mem[504] : 
                        (N239)? mem[536] : 
                        (N240)? mem[568] : 
                        (N241)? mem[600] : 
                        (N242)? mem[632] : 
                        (N243)? mem[664] : 
                        (N244)? mem[696] : 
                        (N245)? mem[728] : 
                        (N246)? mem[760] : 
                        (N247)? mem[792] : 
                        (N248)? mem[824] : 
                        (N249)? mem[856] : 
                        (N250)? mem[888] : 
                        (N251)? mem[920] : 
                        (N252)? mem[952] : 
                        (N253)? mem[984] : 
                        (N254)? mem[1016] : 
                        (N255)? mem[1048] : 
                        (N256)? mem[1080] : 
                        (N257)? mem[1112] : 
                        (N258)? mem[1144] : 
                        (N259)? mem[1176] : 
                        (N260)? mem[1208] : 
                        (N261)? mem[1240] : 
                        (N262)? mem[1272] : 
                        (N263)? mem[1304] : 
                        (N264)? mem[1336] : 
                        (N265)? mem[1368] : 
                        (N266)? mem[1400] : 
                        (N267)? mem[1432] : 
                        (N268)? mem[1464] : 
                        (N269)? mem[1496] : 
                        (N270)? mem[1528] : 
                        (N271)? mem[1560] : 
                        (N272)? mem[1592] : 1'b0;
  assign r_data_o[23] = (N223)? mem[23] : 
                        (N224)? mem[55] : 
                        (N225)? mem[87] : 
                        (N226)? mem[119] : 
                        (N227)? mem[151] : 
                        (N228)? mem[183] : 
                        (N229)? mem[215] : 
                        (N230)? mem[247] : 
                        (N231)? mem[279] : 
                        (N232)? mem[311] : 
                        (N233)? mem[343] : 
                        (N234)? mem[375] : 
                        (N235)? mem[407] : 
                        (N236)? mem[439] : 
                        (N237)? mem[471] : 
                        (N238)? mem[503] : 
                        (N239)? mem[535] : 
                        (N240)? mem[567] : 
                        (N241)? mem[599] : 
                        (N242)? mem[631] : 
                        (N243)? mem[663] : 
                        (N244)? mem[695] : 
                        (N245)? mem[727] : 
                        (N246)? mem[759] : 
                        (N247)? mem[791] : 
                        (N248)? mem[823] : 
                        (N249)? mem[855] : 
                        (N250)? mem[887] : 
                        (N251)? mem[919] : 
                        (N252)? mem[951] : 
                        (N253)? mem[983] : 
                        (N254)? mem[1015] : 
                        (N255)? mem[1047] : 
                        (N256)? mem[1079] : 
                        (N257)? mem[1111] : 
                        (N258)? mem[1143] : 
                        (N259)? mem[1175] : 
                        (N260)? mem[1207] : 
                        (N261)? mem[1239] : 
                        (N262)? mem[1271] : 
                        (N263)? mem[1303] : 
                        (N264)? mem[1335] : 
                        (N265)? mem[1367] : 
                        (N266)? mem[1399] : 
                        (N267)? mem[1431] : 
                        (N268)? mem[1463] : 
                        (N269)? mem[1495] : 
                        (N270)? mem[1527] : 
                        (N271)? mem[1559] : 
                        (N272)? mem[1591] : 1'b0;
  assign r_data_o[22] = (N223)? mem[22] : 
                        (N224)? mem[54] : 
                        (N225)? mem[86] : 
                        (N226)? mem[118] : 
                        (N227)? mem[150] : 
                        (N228)? mem[182] : 
                        (N229)? mem[214] : 
                        (N230)? mem[246] : 
                        (N231)? mem[278] : 
                        (N232)? mem[310] : 
                        (N233)? mem[342] : 
                        (N234)? mem[374] : 
                        (N235)? mem[406] : 
                        (N236)? mem[438] : 
                        (N237)? mem[470] : 
                        (N238)? mem[502] : 
                        (N239)? mem[534] : 
                        (N240)? mem[566] : 
                        (N241)? mem[598] : 
                        (N242)? mem[630] : 
                        (N243)? mem[662] : 
                        (N244)? mem[694] : 
                        (N245)? mem[726] : 
                        (N246)? mem[758] : 
                        (N247)? mem[790] : 
                        (N248)? mem[822] : 
                        (N249)? mem[854] : 
                        (N250)? mem[886] : 
                        (N251)? mem[918] : 
                        (N252)? mem[950] : 
                        (N253)? mem[982] : 
                        (N254)? mem[1014] : 
                        (N255)? mem[1046] : 
                        (N256)? mem[1078] : 
                        (N257)? mem[1110] : 
                        (N258)? mem[1142] : 
                        (N259)? mem[1174] : 
                        (N260)? mem[1206] : 
                        (N261)? mem[1238] : 
                        (N262)? mem[1270] : 
                        (N263)? mem[1302] : 
                        (N264)? mem[1334] : 
                        (N265)? mem[1366] : 
                        (N266)? mem[1398] : 
                        (N267)? mem[1430] : 
                        (N268)? mem[1462] : 
                        (N269)? mem[1494] : 
                        (N270)? mem[1526] : 
                        (N271)? mem[1558] : 
                        (N272)? mem[1590] : 1'b0;
  assign r_data_o[21] = (N223)? mem[21] : 
                        (N224)? mem[53] : 
                        (N225)? mem[85] : 
                        (N226)? mem[117] : 
                        (N227)? mem[149] : 
                        (N228)? mem[181] : 
                        (N229)? mem[213] : 
                        (N230)? mem[245] : 
                        (N231)? mem[277] : 
                        (N232)? mem[309] : 
                        (N233)? mem[341] : 
                        (N234)? mem[373] : 
                        (N235)? mem[405] : 
                        (N236)? mem[437] : 
                        (N237)? mem[469] : 
                        (N238)? mem[501] : 
                        (N239)? mem[533] : 
                        (N240)? mem[565] : 
                        (N241)? mem[597] : 
                        (N242)? mem[629] : 
                        (N243)? mem[661] : 
                        (N244)? mem[693] : 
                        (N245)? mem[725] : 
                        (N246)? mem[757] : 
                        (N247)? mem[789] : 
                        (N248)? mem[821] : 
                        (N249)? mem[853] : 
                        (N250)? mem[885] : 
                        (N251)? mem[917] : 
                        (N252)? mem[949] : 
                        (N253)? mem[981] : 
                        (N254)? mem[1013] : 
                        (N255)? mem[1045] : 
                        (N256)? mem[1077] : 
                        (N257)? mem[1109] : 
                        (N258)? mem[1141] : 
                        (N259)? mem[1173] : 
                        (N260)? mem[1205] : 
                        (N261)? mem[1237] : 
                        (N262)? mem[1269] : 
                        (N263)? mem[1301] : 
                        (N264)? mem[1333] : 
                        (N265)? mem[1365] : 
                        (N266)? mem[1397] : 
                        (N267)? mem[1429] : 
                        (N268)? mem[1461] : 
                        (N269)? mem[1493] : 
                        (N270)? mem[1525] : 
                        (N271)? mem[1557] : 
                        (N272)? mem[1589] : 1'b0;
  assign r_data_o[20] = (N223)? mem[20] : 
                        (N224)? mem[52] : 
                        (N225)? mem[84] : 
                        (N226)? mem[116] : 
                        (N227)? mem[148] : 
                        (N228)? mem[180] : 
                        (N229)? mem[212] : 
                        (N230)? mem[244] : 
                        (N231)? mem[276] : 
                        (N232)? mem[308] : 
                        (N233)? mem[340] : 
                        (N234)? mem[372] : 
                        (N235)? mem[404] : 
                        (N236)? mem[436] : 
                        (N237)? mem[468] : 
                        (N238)? mem[500] : 
                        (N239)? mem[532] : 
                        (N240)? mem[564] : 
                        (N241)? mem[596] : 
                        (N242)? mem[628] : 
                        (N243)? mem[660] : 
                        (N244)? mem[692] : 
                        (N245)? mem[724] : 
                        (N246)? mem[756] : 
                        (N247)? mem[788] : 
                        (N248)? mem[820] : 
                        (N249)? mem[852] : 
                        (N250)? mem[884] : 
                        (N251)? mem[916] : 
                        (N252)? mem[948] : 
                        (N253)? mem[980] : 
                        (N254)? mem[1012] : 
                        (N255)? mem[1044] : 
                        (N256)? mem[1076] : 
                        (N257)? mem[1108] : 
                        (N258)? mem[1140] : 
                        (N259)? mem[1172] : 
                        (N260)? mem[1204] : 
                        (N261)? mem[1236] : 
                        (N262)? mem[1268] : 
                        (N263)? mem[1300] : 
                        (N264)? mem[1332] : 
                        (N265)? mem[1364] : 
                        (N266)? mem[1396] : 
                        (N267)? mem[1428] : 
                        (N268)? mem[1460] : 
                        (N269)? mem[1492] : 
                        (N270)? mem[1524] : 
                        (N271)? mem[1556] : 
                        (N272)? mem[1588] : 1'b0;
  assign r_data_o[19] = (N223)? mem[19] : 
                        (N224)? mem[51] : 
                        (N225)? mem[83] : 
                        (N226)? mem[115] : 
                        (N227)? mem[147] : 
                        (N228)? mem[179] : 
                        (N229)? mem[211] : 
                        (N230)? mem[243] : 
                        (N231)? mem[275] : 
                        (N232)? mem[307] : 
                        (N233)? mem[339] : 
                        (N234)? mem[371] : 
                        (N235)? mem[403] : 
                        (N236)? mem[435] : 
                        (N237)? mem[467] : 
                        (N238)? mem[499] : 
                        (N239)? mem[531] : 
                        (N240)? mem[563] : 
                        (N241)? mem[595] : 
                        (N242)? mem[627] : 
                        (N243)? mem[659] : 
                        (N244)? mem[691] : 
                        (N245)? mem[723] : 
                        (N246)? mem[755] : 
                        (N247)? mem[787] : 
                        (N248)? mem[819] : 
                        (N249)? mem[851] : 
                        (N250)? mem[883] : 
                        (N251)? mem[915] : 
                        (N252)? mem[947] : 
                        (N253)? mem[979] : 
                        (N254)? mem[1011] : 
                        (N255)? mem[1043] : 
                        (N256)? mem[1075] : 
                        (N257)? mem[1107] : 
                        (N258)? mem[1139] : 
                        (N259)? mem[1171] : 
                        (N260)? mem[1203] : 
                        (N261)? mem[1235] : 
                        (N262)? mem[1267] : 
                        (N263)? mem[1299] : 
                        (N264)? mem[1331] : 
                        (N265)? mem[1363] : 
                        (N266)? mem[1395] : 
                        (N267)? mem[1427] : 
                        (N268)? mem[1459] : 
                        (N269)? mem[1491] : 
                        (N270)? mem[1523] : 
                        (N271)? mem[1555] : 
                        (N272)? mem[1587] : 1'b0;
  assign r_data_o[18] = (N223)? mem[18] : 
                        (N224)? mem[50] : 
                        (N225)? mem[82] : 
                        (N226)? mem[114] : 
                        (N227)? mem[146] : 
                        (N228)? mem[178] : 
                        (N229)? mem[210] : 
                        (N230)? mem[242] : 
                        (N231)? mem[274] : 
                        (N232)? mem[306] : 
                        (N233)? mem[338] : 
                        (N234)? mem[370] : 
                        (N235)? mem[402] : 
                        (N236)? mem[434] : 
                        (N237)? mem[466] : 
                        (N238)? mem[498] : 
                        (N239)? mem[530] : 
                        (N240)? mem[562] : 
                        (N241)? mem[594] : 
                        (N242)? mem[626] : 
                        (N243)? mem[658] : 
                        (N244)? mem[690] : 
                        (N245)? mem[722] : 
                        (N246)? mem[754] : 
                        (N247)? mem[786] : 
                        (N248)? mem[818] : 
                        (N249)? mem[850] : 
                        (N250)? mem[882] : 
                        (N251)? mem[914] : 
                        (N252)? mem[946] : 
                        (N253)? mem[978] : 
                        (N254)? mem[1010] : 
                        (N255)? mem[1042] : 
                        (N256)? mem[1074] : 
                        (N257)? mem[1106] : 
                        (N258)? mem[1138] : 
                        (N259)? mem[1170] : 
                        (N260)? mem[1202] : 
                        (N261)? mem[1234] : 
                        (N262)? mem[1266] : 
                        (N263)? mem[1298] : 
                        (N264)? mem[1330] : 
                        (N265)? mem[1362] : 
                        (N266)? mem[1394] : 
                        (N267)? mem[1426] : 
                        (N268)? mem[1458] : 
                        (N269)? mem[1490] : 
                        (N270)? mem[1522] : 
                        (N271)? mem[1554] : 
                        (N272)? mem[1586] : 1'b0;
  assign r_data_o[17] = (N223)? mem[17] : 
                        (N224)? mem[49] : 
                        (N225)? mem[81] : 
                        (N226)? mem[113] : 
                        (N227)? mem[145] : 
                        (N228)? mem[177] : 
                        (N229)? mem[209] : 
                        (N230)? mem[241] : 
                        (N231)? mem[273] : 
                        (N232)? mem[305] : 
                        (N233)? mem[337] : 
                        (N234)? mem[369] : 
                        (N235)? mem[401] : 
                        (N236)? mem[433] : 
                        (N237)? mem[465] : 
                        (N238)? mem[497] : 
                        (N239)? mem[529] : 
                        (N240)? mem[561] : 
                        (N241)? mem[593] : 
                        (N242)? mem[625] : 
                        (N243)? mem[657] : 
                        (N244)? mem[689] : 
                        (N245)? mem[721] : 
                        (N246)? mem[753] : 
                        (N247)? mem[785] : 
                        (N248)? mem[817] : 
                        (N249)? mem[849] : 
                        (N250)? mem[881] : 
                        (N251)? mem[913] : 
                        (N252)? mem[945] : 
                        (N253)? mem[977] : 
                        (N254)? mem[1009] : 
                        (N255)? mem[1041] : 
                        (N256)? mem[1073] : 
                        (N257)? mem[1105] : 
                        (N258)? mem[1137] : 
                        (N259)? mem[1169] : 
                        (N260)? mem[1201] : 
                        (N261)? mem[1233] : 
                        (N262)? mem[1265] : 
                        (N263)? mem[1297] : 
                        (N264)? mem[1329] : 
                        (N265)? mem[1361] : 
                        (N266)? mem[1393] : 
                        (N267)? mem[1425] : 
                        (N268)? mem[1457] : 
                        (N269)? mem[1489] : 
                        (N270)? mem[1521] : 
                        (N271)? mem[1553] : 
                        (N272)? mem[1585] : 1'b0;
  assign r_data_o[16] = (N223)? mem[16] : 
                        (N224)? mem[48] : 
                        (N225)? mem[80] : 
                        (N226)? mem[112] : 
                        (N227)? mem[144] : 
                        (N228)? mem[176] : 
                        (N229)? mem[208] : 
                        (N230)? mem[240] : 
                        (N231)? mem[272] : 
                        (N232)? mem[304] : 
                        (N233)? mem[336] : 
                        (N234)? mem[368] : 
                        (N235)? mem[400] : 
                        (N236)? mem[432] : 
                        (N237)? mem[464] : 
                        (N238)? mem[496] : 
                        (N239)? mem[528] : 
                        (N240)? mem[560] : 
                        (N241)? mem[592] : 
                        (N242)? mem[624] : 
                        (N243)? mem[656] : 
                        (N244)? mem[688] : 
                        (N245)? mem[720] : 
                        (N246)? mem[752] : 
                        (N247)? mem[784] : 
                        (N248)? mem[816] : 
                        (N249)? mem[848] : 
                        (N250)? mem[880] : 
                        (N251)? mem[912] : 
                        (N252)? mem[944] : 
                        (N253)? mem[976] : 
                        (N254)? mem[1008] : 
                        (N255)? mem[1040] : 
                        (N256)? mem[1072] : 
                        (N257)? mem[1104] : 
                        (N258)? mem[1136] : 
                        (N259)? mem[1168] : 
                        (N260)? mem[1200] : 
                        (N261)? mem[1232] : 
                        (N262)? mem[1264] : 
                        (N263)? mem[1296] : 
                        (N264)? mem[1328] : 
                        (N265)? mem[1360] : 
                        (N266)? mem[1392] : 
                        (N267)? mem[1424] : 
                        (N268)? mem[1456] : 
                        (N269)? mem[1488] : 
                        (N270)? mem[1520] : 
                        (N271)? mem[1552] : 
                        (N272)? mem[1584] : 1'b0;
  assign r_data_o[15] = (N223)? mem[15] : 
                        (N224)? mem[47] : 
                        (N225)? mem[79] : 
                        (N226)? mem[111] : 
                        (N227)? mem[143] : 
                        (N228)? mem[175] : 
                        (N229)? mem[207] : 
                        (N230)? mem[239] : 
                        (N231)? mem[271] : 
                        (N232)? mem[303] : 
                        (N233)? mem[335] : 
                        (N234)? mem[367] : 
                        (N235)? mem[399] : 
                        (N236)? mem[431] : 
                        (N237)? mem[463] : 
                        (N238)? mem[495] : 
                        (N239)? mem[527] : 
                        (N240)? mem[559] : 
                        (N241)? mem[591] : 
                        (N242)? mem[623] : 
                        (N243)? mem[655] : 
                        (N244)? mem[687] : 
                        (N245)? mem[719] : 
                        (N246)? mem[751] : 
                        (N247)? mem[783] : 
                        (N248)? mem[815] : 
                        (N249)? mem[847] : 
                        (N250)? mem[879] : 
                        (N251)? mem[911] : 
                        (N252)? mem[943] : 
                        (N253)? mem[975] : 
                        (N254)? mem[1007] : 
                        (N255)? mem[1039] : 
                        (N256)? mem[1071] : 
                        (N257)? mem[1103] : 
                        (N258)? mem[1135] : 
                        (N259)? mem[1167] : 
                        (N260)? mem[1199] : 
                        (N261)? mem[1231] : 
                        (N262)? mem[1263] : 
                        (N263)? mem[1295] : 
                        (N264)? mem[1327] : 
                        (N265)? mem[1359] : 
                        (N266)? mem[1391] : 
                        (N267)? mem[1423] : 
                        (N268)? mem[1455] : 
                        (N269)? mem[1487] : 
                        (N270)? mem[1519] : 
                        (N271)? mem[1551] : 
                        (N272)? mem[1583] : 1'b0;
  assign r_data_o[14] = (N223)? mem[14] : 
                        (N224)? mem[46] : 
                        (N225)? mem[78] : 
                        (N226)? mem[110] : 
                        (N227)? mem[142] : 
                        (N228)? mem[174] : 
                        (N229)? mem[206] : 
                        (N230)? mem[238] : 
                        (N231)? mem[270] : 
                        (N232)? mem[302] : 
                        (N233)? mem[334] : 
                        (N234)? mem[366] : 
                        (N235)? mem[398] : 
                        (N236)? mem[430] : 
                        (N237)? mem[462] : 
                        (N238)? mem[494] : 
                        (N239)? mem[526] : 
                        (N240)? mem[558] : 
                        (N241)? mem[590] : 
                        (N242)? mem[622] : 
                        (N243)? mem[654] : 
                        (N244)? mem[686] : 
                        (N245)? mem[718] : 
                        (N246)? mem[750] : 
                        (N247)? mem[782] : 
                        (N248)? mem[814] : 
                        (N249)? mem[846] : 
                        (N250)? mem[878] : 
                        (N251)? mem[910] : 
                        (N252)? mem[942] : 
                        (N253)? mem[974] : 
                        (N254)? mem[1006] : 
                        (N255)? mem[1038] : 
                        (N256)? mem[1070] : 
                        (N257)? mem[1102] : 
                        (N258)? mem[1134] : 
                        (N259)? mem[1166] : 
                        (N260)? mem[1198] : 
                        (N261)? mem[1230] : 
                        (N262)? mem[1262] : 
                        (N263)? mem[1294] : 
                        (N264)? mem[1326] : 
                        (N265)? mem[1358] : 
                        (N266)? mem[1390] : 
                        (N267)? mem[1422] : 
                        (N268)? mem[1454] : 
                        (N269)? mem[1486] : 
                        (N270)? mem[1518] : 
                        (N271)? mem[1550] : 
                        (N272)? mem[1582] : 1'b0;
  assign r_data_o[13] = (N223)? mem[13] : 
                        (N224)? mem[45] : 
                        (N225)? mem[77] : 
                        (N226)? mem[109] : 
                        (N227)? mem[141] : 
                        (N228)? mem[173] : 
                        (N229)? mem[205] : 
                        (N230)? mem[237] : 
                        (N231)? mem[269] : 
                        (N232)? mem[301] : 
                        (N233)? mem[333] : 
                        (N234)? mem[365] : 
                        (N235)? mem[397] : 
                        (N236)? mem[429] : 
                        (N237)? mem[461] : 
                        (N238)? mem[493] : 
                        (N239)? mem[525] : 
                        (N240)? mem[557] : 
                        (N241)? mem[589] : 
                        (N242)? mem[621] : 
                        (N243)? mem[653] : 
                        (N244)? mem[685] : 
                        (N245)? mem[717] : 
                        (N246)? mem[749] : 
                        (N247)? mem[781] : 
                        (N248)? mem[813] : 
                        (N249)? mem[845] : 
                        (N250)? mem[877] : 
                        (N251)? mem[909] : 
                        (N252)? mem[941] : 
                        (N253)? mem[973] : 
                        (N254)? mem[1005] : 
                        (N255)? mem[1037] : 
                        (N256)? mem[1069] : 
                        (N257)? mem[1101] : 
                        (N258)? mem[1133] : 
                        (N259)? mem[1165] : 
                        (N260)? mem[1197] : 
                        (N261)? mem[1229] : 
                        (N262)? mem[1261] : 
                        (N263)? mem[1293] : 
                        (N264)? mem[1325] : 
                        (N265)? mem[1357] : 
                        (N266)? mem[1389] : 
                        (N267)? mem[1421] : 
                        (N268)? mem[1453] : 
                        (N269)? mem[1485] : 
                        (N270)? mem[1517] : 
                        (N271)? mem[1549] : 
                        (N272)? mem[1581] : 1'b0;
  assign r_data_o[12] = (N223)? mem[12] : 
                        (N224)? mem[44] : 
                        (N225)? mem[76] : 
                        (N226)? mem[108] : 
                        (N227)? mem[140] : 
                        (N228)? mem[172] : 
                        (N229)? mem[204] : 
                        (N230)? mem[236] : 
                        (N231)? mem[268] : 
                        (N232)? mem[300] : 
                        (N233)? mem[332] : 
                        (N234)? mem[364] : 
                        (N235)? mem[396] : 
                        (N236)? mem[428] : 
                        (N237)? mem[460] : 
                        (N238)? mem[492] : 
                        (N239)? mem[524] : 
                        (N240)? mem[556] : 
                        (N241)? mem[588] : 
                        (N242)? mem[620] : 
                        (N243)? mem[652] : 
                        (N244)? mem[684] : 
                        (N245)? mem[716] : 
                        (N246)? mem[748] : 
                        (N247)? mem[780] : 
                        (N248)? mem[812] : 
                        (N249)? mem[844] : 
                        (N250)? mem[876] : 
                        (N251)? mem[908] : 
                        (N252)? mem[940] : 
                        (N253)? mem[972] : 
                        (N254)? mem[1004] : 
                        (N255)? mem[1036] : 
                        (N256)? mem[1068] : 
                        (N257)? mem[1100] : 
                        (N258)? mem[1132] : 
                        (N259)? mem[1164] : 
                        (N260)? mem[1196] : 
                        (N261)? mem[1228] : 
                        (N262)? mem[1260] : 
                        (N263)? mem[1292] : 
                        (N264)? mem[1324] : 
                        (N265)? mem[1356] : 
                        (N266)? mem[1388] : 
                        (N267)? mem[1420] : 
                        (N268)? mem[1452] : 
                        (N269)? mem[1484] : 
                        (N270)? mem[1516] : 
                        (N271)? mem[1548] : 
                        (N272)? mem[1580] : 1'b0;
  assign r_data_o[11] = (N223)? mem[11] : 
                        (N224)? mem[43] : 
                        (N225)? mem[75] : 
                        (N226)? mem[107] : 
                        (N227)? mem[139] : 
                        (N228)? mem[171] : 
                        (N229)? mem[203] : 
                        (N230)? mem[235] : 
                        (N231)? mem[267] : 
                        (N232)? mem[299] : 
                        (N233)? mem[331] : 
                        (N234)? mem[363] : 
                        (N235)? mem[395] : 
                        (N236)? mem[427] : 
                        (N237)? mem[459] : 
                        (N238)? mem[491] : 
                        (N239)? mem[523] : 
                        (N240)? mem[555] : 
                        (N241)? mem[587] : 
                        (N242)? mem[619] : 
                        (N243)? mem[651] : 
                        (N244)? mem[683] : 
                        (N245)? mem[715] : 
                        (N246)? mem[747] : 
                        (N247)? mem[779] : 
                        (N248)? mem[811] : 
                        (N249)? mem[843] : 
                        (N250)? mem[875] : 
                        (N251)? mem[907] : 
                        (N252)? mem[939] : 
                        (N253)? mem[971] : 
                        (N254)? mem[1003] : 
                        (N255)? mem[1035] : 
                        (N256)? mem[1067] : 
                        (N257)? mem[1099] : 
                        (N258)? mem[1131] : 
                        (N259)? mem[1163] : 
                        (N260)? mem[1195] : 
                        (N261)? mem[1227] : 
                        (N262)? mem[1259] : 
                        (N263)? mem[1291] : 
                        (N264)? mem[1323] : 
                        (N265)? mem[1355] : 
                        (N266)? mem[1387] : 
                        (N267)? mem[1419] : 
                        (N268)? mem[1451] : 
                        (N269)? mem[1483] : 
                        (N270)? mem[1515] : 
                        (N271)? mem[1547] : 
                        (N272)? mem[1579] : 1'b0;
  assign r_data_o[10] = (N223)? mem[10] : 
                        (N224)? mem[42] : 
                        (N225)? mem[74] : 
                        (N226)? mem[106] : 
                        (N227)? mem[138] : 
                        (N228)? mem[170] : 
                        (N229)? mem[202] : 
                        (N230)? mem[234] : 
                        (N231)? mem[266] : 
                        (N232)? mem[298] : 
                        (N233)? mem[330] : 
                        (N234)? mem[362] : 
                        (N235)? mem[394] : 
                        (N236)? mem[426] : 
                        (N237)? mem[458] : 
                        (N238)? mem[490] : 
                        (N239)? mem[522] : 
                        (N240)? mem[554] : 
                        (N241)? mem[586] : 
                        (N242)? mem[618] : 
                        (N243)? mem[650] : 
                        (N244)? mem[682] : 
                        (N245)? mem[714] : 
                        (N246)? mem[746] : 
                        (N247)? mem[778] : 
                        (N248)? mem[810] : 
                        (N249)? mem[842] : 
                        (N250)? mem[874] : 
                        (N251)? mem[906] : 
                        (N252)? mem[938] : 
                        (N253)? mem[970] : 
                        (N254)? mem[1002] : 
                        (N255)? mem[1034] : 
                        (N256)? mem[1066] : 
                        (N257)? mem[1098] : 
                        (N258)? mem[1130] : 
                        (N259)? mem[1162] : 
                        (N260)? mem[1194] : 
                        (N261)? mem[1226] : 
                        (N262)? mem[1258] : 
                        (N263)? mem[1290] : 
                        (N264)? mem[1322] : 
                        (N265)? mem[1354] : 
                        (N266)? mem[1386] : 
                        (N267)? mem[1418] : 
                        (N268)? mem[1450] : 
                        (N269)? mem[1482] : 
                        (N270)? mem[1514] : 
                        (N271)? mem[1546] : 
                        (N272)? mem[1578] : 1'b0;
  assign r_data_o[9] = (N223)? mem[9] : 
                       (N224)? mem[41] : 
                       (N225)? mem[73] : 
                       (N226)? mem[105] : 
                       (N227)? mem[137] : 
                       (N228)? mem[169] : 
                       (N229)? mem[201] : 
                       (N230)? mem[233] : 
                       (N231)? mem[265] : 
                       (N232)? mem[297] : 
                       (N233)? mem[329] : 
                       (N234)? mem[361] : 
                       (N235)? mem[393] : 
                       (N236)? mem[425] : 
                       (N237)? mem[457] : 
                       (N238)? mem[489] : 
                       (N239)? mem[521] : 
                       (N240)? mem[553] : 
                       (N241)? mem[585] : 
                       (N242)? mem[617] : 
                       (N243)? mem[649] : 
                       (N244)? mem[681] : 
                       (N245)? mem[713] : 
                       (N246)? mem[745] : 
                       (N247)? mem[777] : 
                       (N248)? mem[809] : 
                       (N249)? mem[841] : 
                       (N250)? mem[873] : 
                       (N251)? mem[905] : 
                       (N252)? mem[937] : 
                       (N253)? mem[969] : 
                       (N254)? mem[1001] : 
                       (N255)? mem[1033] : 
                       (N256)? mem[1065] : 
                       (N257)? mem[1097] : 
                       (N258)? mem[1129] : 
                       (N259)? mem[1161] : 
                       (N260)? mem[1193] : 
                       (N261)? mem[1225] : 
                       (N262)? mem[1257] : 
                       (N263)? mem[1289] : 
                       (N264)? mem[1321] : 
                       (N265)? mem[1353] : 
                       (N266)? mem[1385] : 
                       (N267)? mem[1417] : 
                       (N268)? mem[1449] : 
                       (N269)? mem[1481] : 
                       (N270)? mem[1513] : 
                       (N271)? mem[1545] : 
                       (N272)? mem[1577] : 1'b0;
  assign r_data_o[8] = (N223)? mem[8] : 
                       (N224)? mem[40] : 
                       (N225)? mem[72] : 
                       (N226)? mem[104] : 
                       (N227)? mem[136] : 
                       (N228)? mem[168] : 
                       (N229)? mem[200] : 
                       (N230)? mem[232] : 
                       (N231)? mem[264] : 
                       (N232)? mem[296] : 
                       (N233)? mem[328] : 
                       (N234)? mem[360] : 
                       (N235)? mem[392] : 
                       (N236)? mem[424] : 
                       (N237)? mem[456] : 
                       (N238)? mem[488] : 
                       (N239)? mem[520] : 
                       (N240)? mem[552] : 
                       (N241)? mem[584] : 
                       (N242)? mem[616] : 
                       (N243)? mem[648] : 
                       (N244)? mem[680] : 
                       (N245)? mem[712] : 
                       (N246)? mem[744] : 
                       (N247)? mem[776] : 
                       (N248)? mem[808] : 
                       (N249)? mem[840] : 
                       (N250)? mem[872] : 
                       (N251)? mem[904] : 
                       (N252)? mem[936] : 
                       (N253)? mem[968] : 
                       (N254)? mem[1000] : 
                       (N255)? mem[1032] : 
                       (N256)? mem[1064] : 
                       (N257)? mem[1096] : 
                       (N258)? mem[1128] : 
                       (N259)? mem[1160] : 
                       (N260)? mem[1192] : 
                       (N261)? mem[1224] : 
                       (N262)? mem[1256] : 
                       (N263)? mem[1288] : 
                       (N264)? mem[1320] : 
                       (N265)? mem[1352] : 
                       (N266)? mem[1384] : 
                       (N267)? mem[1416] : 
                       (N268)? mem[1448] : 
                       (N269)? mem[1480] : 
                       (N270)? mem[1512] : 
                       (N271)? mem[1544] : 
                       (N272)? mem[1576] : 1'b0;
  assign r_data_o[7] = (N223)? mem[7] : 
                       (N224)? mem[39] : 
                       (N225)? mem[71] : 
                       (N226)? mem[103] : 
                       (N227)? mem[135] : 
                       (N228)? mem[167] : 
                       (N229)? mem[199] : 
                       (N230)? mem[231] : 
                       (N231)? mem[263] : 
                       (N232)? mem[295] : 
                       (N233)? mem[327] : 
                       (N234)? mem[359] : 
                       (N235)? mem[391] : 
                       (N236)? mem[423] : 
                       (N237)? mem[455] : 
                       (N238)? mem[487] : 
                       (N239)? mem[519] : 
                       (N240)? mem[551] : 
                       (N241)? mem[583] : 
                       (N242)? mem[615] : 
                       (N243)? mem[647] : 
                       (N244)? mem[679] : 
                       (N245)? mem[711] : 
                       (N246)? mem[743] : 
                       (N247)? mem[775] : 
                       (N248)? mem[807] : 
                       (N249)? mem[839] : 
                       (N250)? mem[871] : 
                       (N251)? mem[903] : 
                       (N252)? mem[935] : 
                       (N253)? mem[967] : 
                       (N254)? mem[999] : 
                       (N255)? mem[1031] : 
                       (N256)? mem[1063] : 
                       (N257)? mem[1095] : 
                       (N258)? mem[1127] : 
                       (N259)? mem[1159] : 
                       (N260)? mem[1191] : 
                       (N261)? mem[1223] : 
                       (N262)? mem[1255] : 
                       (N263)? mem[1287] : 
                       (N264)? mem[1319] : 
                       (N265)? mem[1351] : 
                       (N266)? mem[1383] : 
                       (N267)? mem[1415] : 
                       (N268)? mem[1447] : 
                       (N269)? mem[1479] : 
                       (N270)? mem[1511] : 
                       (N271)? mem[1543] : 
                       (N272)? mem[1575] : 1'b0;
  assign r_data_o[6] = (N223)? mem[6] : 
                       (N224)? mem[38] : 
                       (N225)? mem[70] : 
                       (N226)? mem[102] : 
                       (N227)? mem[134] : 
                       (N228)? mem[166] : 
                       (N229)? mem[198] : 
                       (N230)? mem[230] : 
                       (N231)? mem[262] : 
                       (N232)? mem[294] : 
                       (N233)? mem[326] : 
                       (N234)? mem[358] : 
                       (N235)? mem[390] : 
                       (N236)? mem[422] : 
                       (N237)? mem[454] : 
                       (N238)? mem[486] : 
                       (N239)? mem[518] : 
                       (N240)? mem[550] : 
                       (N241)? mem[582] : 
                       (N242)? mem[614] : 
                       (N243)? mem[646] : 
                       (N244)? mem[678] : 
                       (N245)? mem[710] : 
                       (N246)? mem[742] : 
                       (N247)? mem[774] : 
                       (N248)? mem[806] : 
                       (N249)? mem[838] : 
                       (N250)? mem[870] : 
                       (N251)? mem[902] : 
                       (N252)? mem[934] : 
                       (N253)? mem[966] : 
                       (N254)? mem[998] : 
                       (N255)? mem[1030] : 
                       (N256)? mem[1062] : 
                       (N257)? mem[1094] : 
                       (N258)? mem[1126] : 
                       (N259)? mem[1158] : 
                       (N260)? mem[1190] : 
                       (N261)? mem[1222] : 
                       (N262)? mem[1254] : 
                       (N263)? mem[1286] : 
                       (N264)? mem[1318] : 
                       (N265)? mem[1350] : 
                       (N266)? mem[1382] : 
                       (N267)? mem[1414] : 
                       (N268)? mem[1446] : 
                       (N269)? mem[1478] : 
                       (N270)? mem[1510] : 
                       (N271)? mem[1542] : 
                       (N272)? mem[1574] : 1'b0;
  assign r_data_o[5] = (N223)? mem[5] : 
                       (N224)? mem[37] : 
                       (N225)? mem[69] : 
                       (N226)? mem[101] : 
                       (N227)? mem[133] : 
                       (N228)? mem[165] : 
                       (N229)? mem[197] : 
                       (N230)? mem[229] : 
                       (N231)? mem[261] : 
                       (N232)? mem[293] : 
                       (N233)? mem[325] : 
                       (N234)? mem[357] : 
                       (N235)? mem[389] : 
                       (N236)? mem[421] : 
                       (N237)? mem[453] : 
                       (N238)? mem[485] : 
                       (N239)? mem[517] : 
                       (N240)? mem[549] : 
                       (N241)? mem[581] : 
                       (N242)? mem[613] : 
                       (N243)? mem[645] : 
                       (N244)? mem[677] : 
                       (N245)? mem[709] : 
                       (N246)? mem[741] : 
                       (N247)? mem[773] : 
                       (N248)? mem[805] : 
                       (N249)? mem[837] : 
                       (N250)? mem[869] : 
                       (N251)? mem[901] : 
                       (N252)? mem[933] : 
                       (N253)? mem[965] : 
                       (N254)? mem[997] : 
                       (N255)? mem[1029] : 
                       (N256)? mem[1061] : 
                       (N257)? mem[1093] : 
                       (N258)? mem[1125] : 
                       (N259)? mem[1157] : 
                       (N260)? mem[1189] : 
                       (N261)? mem[1221] : 
                       (N262)? mem[1253] : 
                       (N263)? mem[1285] : 
                       (N264)? mem[1317] : 
                       (N265)? mem[1349] : 
                       (N266)? mem[1381] : 
                       (N267)? mem[1413] : 
                       (N268)? mem[1445] : 
                       (N269)? mem[1477] : 
                       (N270)? mem[1509] : 
                       (N271)? mem[1541] : 
                       (N272)? mem[1573] : 1'b0;
  assign r_data_o[4] = (N223)? mem[4] : 
                       (N224)? mem[36] : 
                       (N225)? mem[68] : 
                       (N226)? mem[100] : 
                       (N227)? mem[132] : 
                       (N228)? mem[164] : 
                       (N229)? mem[196] : 
                       (N230)? mem[228] : 
                       (N231)? mem[260] : 
                       (N232)? mem[292] : 
                       (N233)? mem[324] : 
                       (N234)? mem[356] : 
                       (N235)? mem[388] : 
                       (N236)? mem[420] : 
                       (N237)? mem[452] : 
                       (N238)? mem[484] : 
                       (N239)? mem[516] : 
                       (N240)? mem[548] : 
                       (N241)? mem[580] : 
                       (N242)? mem[612] : 
                       (N243)? mem[644] : 
                       (N244)? mem[676] : 
                       (N245)? mem[708] : 
                       (N246)? mem[740] : 
                       (N247)? mem[772] : 
                       (N248)? mem[804] : 
                       (N249)? mem[836] : 
                       (N250)? mem[868] : 
                       (N251)? mem[900] : 
                       (N252)? mem[932] : 
                       (N253)? mem[964] : 
                       (N254)? mem[996] : 
                       (N255)? mem[1028] : 
                       (N256)? mem[1060] : 
                       (N257)? mem[1092] : 
                       (N258)? mem[1124] : 
                       (N259)? mem[1156] : 
                       (N260)? mem[1188] : 
                       (N261)? mem[1220] : 
                       (N262)? mem[1252] : 
                       (N263)? mem[1284] : 
                       (N264)? mem[1316] : 
                       (N265)? mem[1348] : 
                       (N266)? mem[1380] : 
                       (N267)? mem[1412] : 
                       (N268)? mem[1444] : 
                       (N269)? mem[1476] : 
                       (N270)? mem[1508] : 
                       (N271)? mem[1540] : 
                       (N272)? mem[1572] : 1'b0;
  assign r_data_o[3] = (N223)? mem[3] : 
                       (N224)? mem[35] : 
                       (N225)? mem[67] : 
                       (N226)? mem[99] : 
                       (N227)? mem[131] : 
                       (N228)? mem[163] : 
                       (N229)? mem[195] : 
                       (N230)? mem[227] : 
                       (N231)? mem[259] : 
                       (N232)? mem[291] : 
                       (N233)? mem[323] : 
                       (N234)? mem[355] : 
                       (N235)? mem[387] : 
                       (N236)? mem[419] : 
                       (N237)? mem[451] : 
                       (N238)? mem[483] : 
                       (N239)? mem[515] : 
                       (N240)? mem[547] : 
                       (N241)? mem[579] : 
                       (N242)? mem[611] : 
                       (N243)? mem[643] : 
                       (N244)? mem[675] : 
                       (N245)? mem[707] : 
                       (N246)? mem[739] : 
                       (N247)? mem[771] : 
                       (N248)? mem[803] : 
                       (N249)? mem[835] : 
                       (N250)? mem[867] : 
                       (N251)? mem[899] : 
                       (N252)? mem[931] : 
                       (N253)? mem[963] : 
                       (N254)? mem[995] : 
                       (N255)? mem[1027] : 
                       (N256)? mem[1059] : 
                       (N257)? mem[1091] : 
                       (N258)? mem[1123] : 
                       (N259)? mem[1155] : 
                       (N260)? mem[1187] : 
                       (N261)? mem[1219] : 
                       (N262)? mem[1251] : 
                       (N263)? mem[1283] : 
                       (N264)? mem[1315] : 
                       (N265)? mem[1347] : 
                       (N266)? mem[1379] : 
                       (N267)? mem[1411] : 
                       (N268)? mem[1443] : 
                       (N269)? mem[1475] : 
                       (N270)? mem[1507] : 
                       (N271)? mem[1539] : 
                       (N272)? mem[1571] : 1'b0;
  assign r_data_o[2] = (N223)? mem[2] : 
                       (N224)? mem[34] : 
                       (N225)? mem[66] : 
                       (N226)? mem[98] : 
                       (N227)? mem[130] : 
                       (N228)? mem[162] : 
                       (N229)? mem[194] : 
                       (N230)? mem[226] : 
                       (N231)? mem[258] : 
                       (N232)? mem[290] : 
                       (N233)? mem[322] : 
                       (N234)? mem[354] : 
                       (N235)? mem[386] : 
                       (N236)? mem[418] : 
                       (N237)? mem[450] : 
                       (N238)? mem[482] : 
                       (N239)? mem[514] : 
                       (N240)? mem[546] : 
                       (N241)? mem[578] : 
                       (N242)? mem[610] : 
                       (N243)? mem[642] : 
                       (N244)? mem[674] : 
                       (N245)? mem[706] : 
                       (N246)? mem[738] : 
                       (N247)? mem[770] : 
                       (N248)? mem[802] : 
                       (N249)? mem[834] : 
                       (N250)? mem[866] : 
                       (N251)? mem[898] : 
                       (N252)? mem[930] : 
                       (N253)? mem[962] : 
                       (N254)? mem[994] : 
                       (N255)? mem[1026] : 
                       (N256)? mem[1058] : 
                       (N257)? mem[1090] : 
                       (N258)? mem[1122] : 
                       (N259)? mem[1154] : 
                       (N260)? mem[1186] : 
                       (N261)? mem[1218] : 
                       (N262)? mem[1250] : 
                       (N263)? mem[1282] : 
                       (N264)? mem[1314] : 
                       (N265)? mem[1346] : 
                       (N266)? mem[1378] : 
                       (N267)? mem[1410] : 
                       (N268)? mem[1442] : 
                       (N269)? mem[1474] : 
                       (N270)? mem[1506] : 
                       (N271)? mem[1538] : 
                       (N272)? mem[1570] : 1'b0;
  assign r_data_o[1] = (N223)? mem[1] : 
                       (N224)? mem[33] : 
                       (N225)? mem[65] : 
                       (N226)? mem[97] : 
                       (N227)? mem[129] : 
                       (N228)? mem[161] : 
                       (N229)? mem[193] : 
                       (N230)? mem[225] : 
                       (N231)? mem[257] : 
                       (N232)? mem[289] : 
                       (N233)? mem[321] : 
                       (N234)? mem[353] : 
                       (N235)? mem[385] : 
                       (N236)? mem[417] : 
                       (N237)? mem[449] : 
                       (N238)? mem[481] : 
                       (N239)? mem[513] : 
                       (N240)? mem[545] : 
                       (N241)? mem[577] : 
                       (N242)? mem[609] : 
                       (N243)? mem[641] : 
                       (N244)? mem[673] : 
                       (N245)? mem[705] : 
                       (N246)? mem[737] : 
                       (N247)? mem[769] : 
                       (N248)? mem[801] : 
                       (N249)? mem[833] : 
                       (N250)? mem[865] : 
                       (N251)? mem[897] : 
                       (N252)? mem[929] : 
                       (N253)? mem[961] : 
                       (N254)? mem[993] : 
                       (N255)? mem[1025] : 
                       (N256)? mem[1057] : 
                       (N257)? mem[1089] : 
                       (N258)? mem[1121] : 
                       (N259)? mem[1153] : 
                       (N260)? mem[1185] : 
                       (N261)? mem[1217] : 
                       (N262)? mem[1249] : 
                       (N263)? mem[1281] : 
                       (N264)? mem[1313] : 
                       (N265)? mem[1345] : 
                       (N266)? mem[1377] : 
                       (N267)? mem[1409] : 
                       (N268)? mem[1441] : 
                       (N269)? mem[1473] : 
                       (N270)? mem[1505] : 
                       (N271)? mem[1537] : 
                       (N272)? mem[1569] : 1'b0;
  assign r_data_o[0] = (N223)? mem[0] : 
                       (N224)? mem[32] : 
                       (N225)? mem[64] : 
                       (N226)? mem[96] : 
                       (N227)? mem[128] : 
                       (N228)? mem[160] : 
                       (N229)? mem[192] : 
                       (N230)? mem[224] : 
                       (N231)? mem[256] : 
                       (N232)? mem[288] : 
                       (N233)? mem[320] : 
                       (N234)? mem[352] : 
                       (N235)? mem[384] : 
                       (N236)? mem[416] : 
                       (N237)? mem[448] : 
                       (N238)? mem[480] : 
                       (N239)? mem[512] : 
                       (N240)? mem[544] : 
                       (N241)? mem[576] : 
                       (N242)? mem[608] : 
                       (N243)? mem[640] : 
                       (N244)? mem[672] : 
                       (N245)? mem[704] : 
                       (N246)? mem[736] : 
                       (N247)? mem[768] : 
                       (N248)? mem[800] : 
                       (N249)? mem[832] : 
                       (N250)? mem[864] : 
                       (N251)? mem[896] : 
                       (N252)? mem[928] : 
                       (N253)? mem[960] : 
                       (N254)? mem[992] : 
                       (N255)? mem[1024] : 
                       (N256)? mem[1056] : 
                       (N257)? mem[1088] : 
                       (N258)? mem[1120] : 
                       (N259)? mem[1152] : 
                       (N260)? mem[1184] : 
                       (N261)? mem[1216] : 
                       (N262)? mem[1248] : 
                       (N263)? mem[1280] : 
                       (N264)? mem[1312] : 
                       (N265)? mem[1344] : 
                       (N266)? mem[1376] : 
                       (N267)? mem[1408] : 
                       (N268)? mem[1440] : 
                       (N269)? mem[1472] : 
                       (N270)? mem[1504] : 
                       (N271)? mem[1536] : 
                       (N272)? mem[1568] : 1'b0;
  assign N323 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N423) begin
      mem_1599_sv2v_reg <= w_data_i[31];
      mem_1598_sv2v_reg <= w_data_i[30];
      mem_1597_sv2v_reg <= w_data_i[29];
      mem_1596_sv2v_reg <= w_data_i[28];
      mem_1595_sv2v_reg <= w_data_i[27];
      mem_1594_sv2v_reg <= w_data_i[26];
      mem_1593_sv2v_reg <= w_data_i[25];
      mem_1592_sv2v_reg <= w_data_i[24];
      mem_1591_sv2v_reg <= w_data_i[23];
      mem_1590_sv2v_reg <= w_data_i[22];
      mem_1589_sv2v_reg <= w_data_i[21];
      mem_1588_sv2v_reg <= w_data_i[20];
      mem_1587_sv2v_reg <= w_data_i[19];
      mem_1586_sv2v_reg <= w_data_i[18];
      mem_1585_sv2v_reg <= w_data_i[17];
      mem_1584_sv2v_reg <= w_data_i[16];
      mem_1583_sv2v_reg <= w_data_i[15];
      mem_1582_sv2v_reg <= w_data_i[14];
      mem_1581_sv2v_reg <= w_data_i[13];
      mem_1580_sv2v_reg <= w_data_i[12];
      mem_1579_sv2v_reg <= w_data_i[11];
      mem_1578_sv2v_reg <= w_data_i[10];
      mem_1577_sv2v_reg <= w_data_i[9];
      mem_1576_sv2v_reg <= w_data_i[8];
      mem_1575_sv2v_reg <= w_data_i[7];
      mem_1574_sv2v_reg <= w_data_i[6];
      mem_1573_sv2v_reg <= w_data_i[5];
      mem_1572_sv2v_reg <= w_data_i[4];
      mem_1571_sv2v_reg <= w_data_i[3];
      mem_1570_sv2v_reg <= w_data_i[2];
      mem_1569_sv2v_reg <= w_data_i[1];
      mem_1568_sv2v_reg <= w_data_i[0];
    end 
    if(N422) begin
      mem_1567_sv2v_reg <= w_data_i[31];
      mem_1566_sv2v_reg <= w_data_i[30];
      mem_1565_sv2v_reg <= w_data_i[29];
      mem_1564_sv2v_reg <= w_data_i[28];
      mem_1563_sv2v_reg <= w_data_i[27];
      mem_1562_sv2v_reg <= w_data_i[26];
      mem_1561_sv2v_reg <= w_data_i[25];
      mem_1560_sv2v_reg <= w_data_i[24];
      mem_1559_sv2v_reg <= w_data_i[23];
      mem_1558_sv2v_reg <= w_data_i[22];
      mem_1557_sv2v_reg <= w_data_i[21];
      mem_1556_sv2v_reg <= w_data_i[20];
      mem_1555_sv2v_reg <= w_data_i[19];
      mem_1554_sv2v_reg <= w_data_i[18];
      mem_1553_sv2v_reg <= w_data_i[17];
      mem_1552_sv2v_reg <= w_data_i[16];
      mem_1551_sv2v_reg <= w_data_i[15];
      mem_1550_sv2v_reg <= w_data_i[14];
      mem_1549_sv2v_reg <= w_data_i[13];
      mem_1548_sv2v_reg <= w_data_i[12];
      mem_1547_sv2v_reg <= w_data_i[11];
      mem_1546_sv2v_reg <= w_data_i[10];
      mem_1545_sv2v_reg <= w_data_i[9];
      mem_1544_sv2v_reg <= w_data_i[8];
      mem_1543_sv2v_reg <= w_data_i[7];
      mem_1542_sv2v_reg <= w_data_i[6];
      mem_1541_sv2v_reg <= w_data_i[5];
      mem_1540_sv2v_reg <= w_data_i[4];
      mem_1539_sv2v_reg <= w_data_i[3];
      mem_1538_sv2v_reg <= w_data_i[2];
      mem_1537_sv2v_reg <= w_data_i[1];
      mem_1536_sv2v_reg <= w_data_i[0];
    end 
    if(N421) begin
      mem_1535_sv2v_reg <= w_data_i[31];
      mem_1534_sv2v_reg <= w_data_i[30];
      mem_1533_sv2v_reg <= w_data_i[29];
      mem_1532_sv2v_reg <= w_data_i[28];
      mem_1531_sv2v_reg <= w_data_i[27];
      mem_1530_sv2v_reg <= w_data_i[26];
      mem_1529_sv2v_reg <= w_data_i[25];
      mem_1528_sv2v_reg <= w_data_i[24];
      mem_1527_sv2v_reg <= w_data_i[23];
      mem_1526_sv2v_reg <= w_data_i[22];
      mem_1525_sv2v_reg <= w_data_i[21];
      mem_1524_sv2v_reg <= w_data_i[20];
      mem_1523_sv2v_reg <= w_data_i[19];
      mem_1522_sv2v_reg <= w_data_i[18];
      mem_1521_sv2v_reg <= w_data_i[17];
      mem_1520_sv2v_reg <= w_data_i[16];
      mem_1519_sv2v_reg <= w_data_i[15];
      mem_1518_sv2v_reg <= w_data_i[14];
      mem_1517_sv2v_reg <= w_data_i[13];
      mem_1516_sv2v_reg <= w_data_i[12];
      mem_1515_sv2v_reg <= w_data_i[11];
      mem_1514_sv2v_reg <= w_data_i[10];
      mem_1513_sv2v_reg <= w_data_i[9];
      mem_1512_sv2v_reg <= w_data_i[8];
      mem_1511_sv2v_reg <= w_data_i[7];
      mem_1510_sv2v_reg <= w_data_i[6];
      mem_1509_sv2v_reg <= w_data_i[5];
      mem_1508_sv2v_reg <= w_data_i[4];
      mem_1507_sv2v_reg <= w_data_i[3];
      mem_1506_sv2v_reg <= w_data_i[2];
      mem_1505_sv2v_reg <= w_data_i[1];
      mem_1504_sv2v_reg <= w_data_i[0];
    end 
    if(N420) begin
      mem_1503_sv2v_reg <= w_data_i[31];
      mem_1502_sv2v_reg <= w_data_i[30];
      mem_1501_sv2v_reg <= w_data_i[29];
      mem_1500_sv2v_reg <= w_data_i[28];
      mem_1499_sv2v_reg <= w_data_i[27];
      mem_1498_sv2v_reg <= w_data_i[26];
      mem_1497_sv2v_reg <= w_data_i[25];
      mem_1496_sv2v_reg <= w_data_i[24];
      mem_1495_sv2v_reg <= w_data_i[23];
      mem_1494_sv2v_reg <= w_data_i[22];
      mem_1493_sv2v_reg <= w_data_i[21];
      mem_1492_sv2v_reg <= w_data_i[20];
      mem_1491_sv2v_reg <= w_data_i[19];
      mem_1490_sv2v_reg <= w_data_i[18];
      mem_1489_sv2v_reg <= w_data_i[17];
      mem_1488_sv2v_reg <= w_data_i[16];
      mem_1487_sv2v_reg <= w_data_i[15];
      mem_1486_sv2v_reg <= w_data_i[14];
      mem_1485_sv2v_reg <= w_data_i[13];
      mem_1484_sv2v_reg <= w_data_i[12];
      mem_1483_sv2v_reg <= w_data_i[11];
      mem_1482_sv2v_reg <= w_data_i[10];
      mem_1481_sv2v_reg <= w_data_i[9];
      mem_1480_sv2v_reg <= w_data_i[8];
      mem_1479_sv2v_reg <= w_data_i[7];
      mem_1478_sv2v_reg <= w_data_i[6];
      mem_1477_sv2v_reg <= w_data_i[5];
      mem_1476_sv2v_reg <= w_data_i[4];
      mem_1475_sv2v_reg <= w_data_i[3];
      mem_1474_sv2v_reg <= w_data_i[2];
      mem_1473_sv2v_reg <= w_data_i[1];
      mem_1472_sv2v_reg <= w_data_i[0];
    end 
    if(N419) begin
      mem_1471_sv2v_reg <= w_data_i[31];
      mem_1470_sv2v_reg <= w_data_i[30];
      mem_1469_sv2v_reg <= w_data_i[29];
      mem_1468_sv2v_reg <= w_data_i[28];
      mem_1467_sv2v_reg <= w_data_i[27];
      mem_1466_sv2v_reg <= w_data_i[26];
      mem_1465_sv2v_reg <= w_data_i[25];
      mem_1464_sv2v_reg <= w_data_i[24];
      mem_1463_sv2v_reg <= w_data_i[23];
      mem_1462_sv2v_reg <= w_data_i[22];
      mem_1461_sv2v_reg <= w_data_i[21];
      mem_1460_sv2v_reg <= w_data_i[20];
      mem_1459_sv2v_reg <= w_data_i[19];
      mem_1458_sv2v_reg <= w_data_i[18];
      mem_1457_sv2v_reg <= w_data_i[17];
      mem_1456_sv2v_reg <= w_data_i[16];
      mem_1455_sv2v_reg <= w_data_i[15];
      mem_1454_sv2v_reg <= w_data_i[14];
      mem_1453_sv2v_reg <= w_data_i[13];
      mem_1452_sv2v_reg <= w_data_i[12];
      mem_1451_sv2v_reg <= w_data_i[11];
      mem_1450_sv2v_reg <= w_data_i[10];
      mem_1449_sv2v_reg <= w_data_i[9];
      mem_1448_sv2v_reg <= w_data_i[8];
      mem_1447_sv2v_reg <= w_data_i[7];
      mem_1446_sv2v_reg <= w_data_i[6];
      mem_1445_sv2v_reg <= w_data_i[5];
      mem_1444_sv2v_reg <= w_data_i[4];
      mem_1443_sv2v_reg <= w_data_i[3];
      mem_1442_sv2v_reg <= w_data_i[2];
      mem_1441_sv2v_reg <= w_data_i[1];
      mem_1440_sv2v_reg <= w_data_i[0];
    end 
    if(N418) begin
      mem_1439_sv2v_reg <= w_data_i[31];
      mem_1438_sv2v_reg <= w_data_i[30];
      mem_1437_sv2v_reg <= w_data_i[29];
      mem_1436_sv2v_reg <= w_data_i[28];
      mem_1435_sv2v_reg <= w_data_i[27];
      mem_1434_sv2v_reg <= w_data_i[26];
      mem_1433_sv2v_reg <= w_data_i[25];
      mem_1432_sv2v_reg <= w_data_i[24];
      mem_1431_sv2v_reg <= w_data_i[23];
      mem_1430_sv2v_reg <= w_data_i[22];
      mem_1429_sv2v_reg <= w_data_i[21];
      mem_1428_sv2v_reg <= w_data_i[20];
      mem_1427_sv2v_reg <= w_data_i[19];
      mem_1426_sv2v_reg <= w_data_i[18];
      mem_1425_sv2v_reg <= w_data_i[17];
      mem_1424_sv2v_reg <= w_data_i[16];
      mem_1423_sv2v_reg <= w_data_i[15];
      mem_1422_sv2v_reg <= w_data_i[14];
      mem_1421_sv2v_reg <= w_data_i[13];
      mem_1420_sv2v_reg <= w_data_i[12];
      mem_1419_sv2v_reg <= w_data_i[11];
      mem_1418_sv2v_reg <= w_data_i[10];
      mem_1417_sv2v_reg <= w_data_i[9];
      mem_1416_sv2v_reg <= w_data_i[8];
      mem_1415_sv2v_reg <= w_data_i[7];
      mem_1414_sv2v_reg <= w_data_i[6];
      mem_1413_sv2v_reg <= w_data_i[5];
      mem_1412_sv2v_reg <= w_data_i[4];
      mem_1411_sv2v_reg <= w_data_i[3];
      mem_1410_sv2v_reg <= w_data_i[2];
      mem_1409_sv2v_reg <= w_data_i[1];
      mem_1408_sv2v_reg <= w_data_i[0];
    end 
    if(N417) begin
      mem_1407_sv2v_reg <= w_data_i[31];
      mem_1406_sv2v_reg <= w_data_i[30];
      mem_1405_sv2v_reg <= w_data_i[29];
      mem_1404_sv2v_reg <= w_data_i[28];
      mem_1403_sv2v_reg <= w_data_i[27];
      mem_1402_sv2v_reg <= w_data_i[26];
      mem_1401_sv2v_reg <= w_data_i[25];
      mem_1400_sv2v_reg <= w_data_i[24];
      mem_1399_sv2v_reg <= w_data_i[23];
      mem_1398_sv2v_reg <= w_data_i[22];
      mem_1397_sv2v_reg <= w_data_i[21];
      mem_1396_sv2v_reg <= w_data_i[20];
      mem_1395_sv2v_reg <= w_data_i[19];
      mem_1394_sv2v_reg <= w_data_i[18];
      mem_1393_sv2v_reg <= w_data_i[17];
      mem_1392_sv2v_reg <= w_data_i[16];
      mem_1391_sv2v_reg <= w_data_i[15];
      mem_1390_sv2v_reg <= w_data_i[14];
      mem_1389_sv2v_reg <= w_data_i[13];
      mem_1388_sv2v_reg <= w_data_i[12];
      mem_1387_sv2v_reg <= w_data_i[11];
      mem_1386_sv2v_reg <= w_data_i[10];
      mem_1385_sv2v_reg <= w_data_i[9];
      mem_1384_sv2v_reg <= w_data_i[8];
      mem_1383_sv2v_reg <= w_data_i[7];
      mem_1382_sv2v_reg <= w_data_i[6];
      mem_1381_sv2v_reg <= w_data_i[5];
      mem_1380_sv2v_reg <= w_data_i[4];
      mem_1379_sv2v_reg <= w_data_i[3];
      mem_1378_sv2v_reg <= w_data_i[2];
      mem_1377_sv2v_reg <= w_data_i[1];
      mem_1376_sv2v_reg <= w_data_i[0];
    end 
    if(N416) begin
      mem_1375_sv2v_reg <= w_data_i[31];
      mem_1374_sv2v_reg <= w_data_i[30];
      mem_1373_sv2v_reg <= w_data_i[29];
      mem_1372_sv2v_reg <= w_data_i[28];
      mem_1371_sv2v_reg <= w_data_i[27];
      mem_1370_sv2v_reg <= w_data_i[26];
      mem_1369_sv2v_reg <= w_data_i[25];
      mem_1368_sv2v_reg <= w_data_i[24];
      mem_1367_sv2v_reg <= w_data_i[23];
      mem_1366_sv2v_reg <= w_data_i[22];
      mem_1365_sv2v_reg <= w_data_i[21];
      mem_1364_sv2v_reg <= w_data_i[20];
      mem_1363_sv2v_reg <= w_data_i[19];
      mem_1362_sv2v_reg <= w_data_i[18];
      mem_1361_sv2v_reg <= w_data_i[17];
      mem_1360_sv2v_reg <= w_data_i[16];
      mem_1359_sv2v_reg <= w_data_i[15];
      mem_1358_sv2v_reg <= w_data_i[14];
      mem_1357_sv2v_reg <= w_data_i[13];
      mem_1356_sv2v_reg <= w_data_i[12];
      mem_1355_sv2v_reg <= w_data_i[11];
      mem_1354_sv2v_reg <= w_data_i[10];
      mem_1353_sv2v_reg <= w_data_i[9];
      mem_1352_sv2v_reg <= w_data_i[8];
      mem_1351_sv2v_reg <= w_data_i[7];
      mem_1350_sv2v_reg <= w_data_i[6];
      mem_1349_sv2v_reg <= w_data_i[5];
      mem_1348_sv2v_reg <= w_data_i[4];
      mem_1347_sv2v_reg <= w_data_i[3];
      mem_1346_sv2v_reg <= w_data_i[2];
      mem_1345_sv2v_reg <= w_data_i[1];
      mem_1344_sv2v_reg <= w_data_i[0];
    end 
    if(N415) begin
      mem_1343_sv2v_reg <= w_data_i[31];
      mem_1342_sv2v_reg <= w_data_i[30];
      mem_1341_sv2v_reg <= w_data_i[29];
      mem_1340_sv2v_reg <= w_data_i[28];
      mem_1339_sv2v_reg <= w_data_i[27];
      mem_1338_sv2v_reg <= w_data_i[26];
      mem_1337_sv2v_reg <= w_data_i[25];
      mem_1336_sv2v_reg <= w_data_i[24];
      mem_1335_sv2v_reg <= w_data_i[23];
      mem_1334_sv2v_reg <= w_data_i[22];
      mem_1333_sv2v_reg <= w_data_i[21];
      mem_1332_sv2v_reg <= w_data_i[20];
      mem_1331_sv2v_reg <= w_data_i[19];
      mem_1330_sv2v_reg <= w_data_i[18];
      mem_1329_sv2v_reg <= w_data_i[17];
      mem_1328_sv2v_reg <= w_data_i[16];
      mem_1327_sv2v_reg <= w_data_i[15];
      mem_1326_sv2v_reg <= w_data_i[14];
      mem_1325_sv2v_reg <= w_data_i[13];
      mem_1324_sv2v_reg <= w_data_i[12];
      mem_1323_sv2v_reg <= w_data_i[11];
      mem_1322_sv2v_reg <= w_data_i[10];
      mem_1321_sv2v_reg <= w_data_i[9];
      mem_1320_sv2v_reg <= w_data_i[8];
      mem_1319_sv2v_reg <= w_data_i[7];
      mem_1318_sv2v_reg <= w_data_i[6];
      mem_1317_sv2v_reg <= w_data_i[5];
      mem_1316_sv2v_reg <= w_data_i[4];
      mem_1315_sv2v_reg <= w_data_i[3];
      mem_1314_sv2v_reg <= w_data_i[2];
      mem_1313_sv2v_reg <= w_data_i[1];
      mem_1312_sv2v_reg <= w_data_i[0];
    end 
    if(N414) begin
      mem_1311_sv2v_reg <= w_data_i[31];
      mem_1310_sv2v_reg <= w_data_i[30];
      mem_1309_sv2v_reg <= w_data_i[29];
      mem_1308_sv2v_reg <= w_data_i[28];
      mem_1307_sv2v_reg <= w_data_i[27];
      mem_1306_sv2v_reg <= w_data_i[26];
      mem_1305_sv2v_reg <= w_data_i[25];
      mem_1304_sv2v_reg <= w_data_i[24];
      mem_1303_sv2v_reg <= w_data_i[23];
      mem_1302_sv2v_reg <= w_data_i[22];
      mem_1301_sv2v_reg <= w_data_i[21];
      mem_1300_sv2v_reg <= w_data_i[20];
      mem_1299_sv2v_reg <= w_data_i[19];
      mem_1298_sv2v_reg <= w_data_i[18];
      mem_1297_sv2v_reg <= w_data_i[17];
      mem_1296_sv2v_reg <= w_data_i[16];
      mem_1295_sv2v_reg <= w_data_i[15];
      mem_1294_sv2v_reg <= w_data_i[14];
      mem_1293_sv2v_reg <= w_data_i[13];
      mem_1292_sv2v_reg <= w_data_i[12];
      mem_1291_sv2v_reg <= w_data_i[11];
      mem_1290_sv2v_reg <= w_data_i[10];
      mem_1289_sv2v_reg <= w_data_i[9];
      mem_1288_sv2v_reg <= w_data_i[8];
      mem_1287_sv2v_reg <= w_data_i[7];
      mem_1286_sv2v_reg <= w_data_i[6];
      mem_1285_sv2v_reg <= w_data_i[5];
      mem_1284_sv2v_reg <= w_data_i[4];
      mem_1283_sv2v_reg <= w_data_i[3];
      mem_1282_sv2v_reg <= w_data_i[2];
      mem_1281_sv2v_reg <= w_data_i[1];
      mem_1280_sv2v_reg <= w_data_i[0];
    end 
    if(N413) begin
      mem_1279_sv2v_reg <= w_data_i[31];
      mem_1278_sv2v_reg <= w_data_i[30];
      mem_1277_sv2v_reg <= w_data_i[29];
      mem_1276_sv2v_reg <= w_data_i[28];
      mem_1275_sv2v_reg <= w_data_i[27];
      mem_1274_sv2v_reg <= w_data_i[26];
      mem_1273_sv2v_reg <= w_data_i[25];
      mem_1272_sv2v_reg <= w_data_i[24];
      mem_1271_sv2v_reg <= w_data_i[23];
      mem_1270_sv2v_reg <= w_data_i[22];
      mem_1269_sv2v_reg <= w_data_i[21];
      mem_1268_sv2v_reg <= w_data_i[20];
      mem_1267_sv2v_reg <= w_data_i[19];
      mem_1266_sv2v_reg <= w_data_i[18];
      mem_1265_sv2v_reg <= w_data_i[17];
      mem_1264_sv2v_reg <= w_data_i[16];
      mem_1263_sv2v_reg <= w_data_i[15];
      mem_1262_sv2v_reg <= w_data_i[14];
      mem_1261_sv2v_reg <= w_data_i[13];
      mem_1260_sv2v_reg <= w_data_i[12];
      mem_1259_sv2v_reg <= w_data_i[11];
      mem_1258_sv2v_reg <= w_data_i[10];
      mem_1257_sv2v_reg <= w_data_i[9];
      mem_1256_sv2v_reg <= w_data_i[8];
      mem_1255_sv2v_reg <= w_data_i[7];
      mem_1254_sv2v_reg <= w_data_i[6];
      mem_1253_sv2v_reg <= w_data_i[5];
      mem_1252_sv2v_reg <= w_data_i[4];
      mem_1251_sv2v_reg <= w_data_i[3];
      mem_1250_sv2v_reg <= w_data_i[2];
      mem_1249_sv2v_reg <= w_data_i[1];
      mem_1248_sv2v_reg <= w_data_i[0];
    end 
    if(N412) begin
      mem_1247_sv2v_reg <= w_data_i[31];
      mem_1246_sv2v_reg <= w_data_i[30];
      mem_1245_sv2v_reg <= w_data_i[29];
      mem_1244_sv2v_reg <= w_data_i[28];
      mem_1243_sv2v_reg <= w_data_i[27];
      mem_1242_sv2v_reg <= w_data_i[26];
      mem_1241_sv2v_reg <= w_data_i[25];
      mem_1240_sv2v_reg <= w_data_i[24];
      mem_1239_sv2v_reg <= w_data_i[23];
      mem_1238_sv2v_reg <= w_data_i[22];
      mem_1237_sv2v_reg <= w_data_i[21];
      mem_1236_sv2v_reg <= w_data_i[20];
      mem_1235_sv2v_reg <= w_data_i[19];
      mem_1234_sv2v_reg <= w_data_i[18];
      mem_1233_sv2v_reg <= w_data_i[17];
      mem_1232_sv2v_reg <= w_data_i[16];
      mem_1231_sv2v_reg <= w_data_i[15];
      mem_1230_sv2v_reg <= w_data_i[14];
      mem_1229_sv2v_reg <= w_data_i[13];
      mem_1228_sv2v_reg <= w_data_i[12];
      mem_1227_sv2v_reg <= w_data_i[11];
      mem_1226_sv2v_reg <= w_data_i[10];
      mem_1225_sv2v_reg <= w_data_i[9];
      mem_1224_sv2v_reg <= w_data_i[8];
      mem_1223_sv2v_reg <= w_data_i[7];
      mem_1222_sv2v_reg <= w_data_i[6];
      mem_1221_sv2v_reg <= w_data_i[5];
      mem_1220_sv2v_reg <= w_data_i[4];
      mem_1219_sv2v_reg <= w_data_i[3];
      mem_1218_sv2v_reg <= w_data_i[2];
      mem_1217_sv2v_reg <= w_data_i[1];
      mem_1216_sv2v_reg <= w_data_i[0];
    end 
    if(N411) begin
      mem_1215_sv2v_reg <= w_data_i[31];
      mem_1214_sv2v_reg <= w_data_i[30];
      mem_1213_sv2v_reg <= w_data_i[29];
      mem_1212_sv2v_reg <= w_data_i[28];
      mem_1211_sv2v_reg <= w_data_i[27];
      mem_1210_sv2v_reg <= w_data_i[26];
      mem_1209_sv2v_reg <= w_data_i[25];
      mem_1208_sv2v_reg <= w_data_i[24];
      mem_1207_sv2v_reg <= w_data_i[23];
      mem_1206_sv2v_reg <= w_data_i[22];
      mem_1205_sv2v_reg <= w_data_i[21];
      mem_1204_sv2v_reg <= w_data_i[20];
      mem_1203_sv2v_reg <= w_data_i[19];
      mem_1202_sv2v_reg <= w_data_i[18];
      mem_1201_sv2v_reg <= w_data_i[17];
      mem_1200_sv2v_reg <= w_data_i[16];
      mem_1199_sv2v_reg <= w_data_i[15];
      mem_1198_sv2v_reg <= w_data_i[14];
      mem_1197_sv2v_reg <= w_data_i[13];
      mem_1196_sv2v_reg <= w_data_i[12];
      mem_1195_sv2v_reg <= w_data_i[11];
      mem_1194_sv2v_reg <= w_data_i[10];
      mem_1193_sv2v_reg <= w_data_i[9];
      mem_1192_sv2v_reg <= w_data_i[8];
      mem_1191_sv2v_reg <= w_data_i[7];
      mem_1190_sv2v_reg <= w_data_i[6];
      mem_1189_sv2v_reg <= w_data_i[5];
      mem_1188_sv2v_reg <= w_data_i[4];
      mem_1187_sv2v_reg <= w_data_i[3];
      mem_1186_sv2v_reg <= w_data_i[2];
      mem_1185_sv2v_reg <= w_data_i[1];
      mem_1184_sv2v_reg <= w_data_i[0];
    end 
    if(N410) begin
      mem_1183_sv2v_reg <= w_data_i[31];
      mem_1182_sv2v_reg <= w_data_i[30];
      mem_1181_sv2v_reg <= w_data_i[29];
      mem_1180_sv2v_reg <= w_data_i[28];
      mem_1179_sv2v_reg <= w_data_i[27];
      mem_1178_sv2v_reg <= w_data_i[26];
      mem_1177_sv2v_reg <= w_data_i[25];
      mem_1176_sv2v_reg <= w_data_i[24];
      mem_1175_sv2v_reg <= w_data_i[23];
      mem_1174_sv2v_reg <= w_data_i[22];
      mem_1173_sv2v_reg <= w_data_i[21];
      mem_1172_sv2v_reg <= w_data_i[20];
      mem_1171_sv2v_reg <= w_data_i[19];
      mem_1170_sv2v_reg <= w_data_i[18];
      mem_1169_sv2v_reg <= w_data_i[17];
      mem_1168_sv2v_reg <= w_data_i[16];
      mem_1167_sv2v_reg <= w_data_i[15];
      mem_1166_sv2v_reg <= w_data_i[14];
      mem_1165_sv2v_reg <= w_data_i[13];
      mem_1164_sv2v_reg <= w_data_i[12];
      mem_1163_sv2v_reg <= w_data_i[11];
      mem_1162_sv2v_reg <= w_data_i[10];
      mem_1161_sv2v_reg <= w_data_i[9];
      mem_1160_sv2v_reg <= w_data_i[8];
      mem_1159_sv2v_reg <= w_data_i[7];
      mem_1158_sv2v_reg <= w_data_i[6];
      mem_1157_sv2v_reg <= w_data_i[5];
      mem_1156_sv2v_reg <= w_data_i[4];
      mem_1155_sv2v_reg <= w_data_i[3];
      mem_1154_sv2v_reg <= w_data_i[2];
      mem_1153_sv2v_reg <= w_data_i[1];
      mem_1152_sv2v_reg <= w_data_i[0];
    end 
    if(N409) begin
      mem_1151_sv2v_reg <= w_data_i[31];
      mem_1150_sv2v_reg <= w_data_i[30];
      mem_1149_sv2v_reg <= w_data_i[29];
      mem_1148_sv2v_reg <= w_data_i[28];
      mem_1147_sv2v_reg <= w_data_i[27];
      mem_1146_sv2v_reg <= w_data_i[26];
      mem_1145_sv2v_reg <= w_data_i[25];
      mem_1144_sv2v_reg <= w_data_i[24];
      mem_1143_sv2v_reg <= w_data_i[23];
      mem_1142_sv2v_reg <= w_data_i[22];
      mem_1141_sv2v_reg <= w_data_i[21];
      mem_1140_sv2v_reg <= w_data_i[20];
      mem_1139_sv2v_reg <= w_data_i[19];
      mem_1138_sv2v_reg <= w_data_i[18];
      mem_1137_sv2v_reg <= w_data_i[17];
      mem_1136_sv2v_reg <= w_data_i[16];
      mem_1135_sv2v_reg <= w_data_i[15];
      mem_1134_sv2v_reg <= w_data_i[14];
      mem_1133_sv2v_reg <= w_data_i[13];
      mem_1132_sv2v_reg <= w_data_i[12];
      mem_1131_sv2v_reg <= w_data_i[11];
      mem_1130_sv2v_reg <= w_data_i[10];
      mem_1129_sv2v_reg <= w_data_i[9];
      mem_1128_sv2v_reg <= w_data_i[8];
      mem_1127_sv2v_reg <= w_data_i[7];
      mem_1126_sv2v_reg <= w_data_i[6];
      mem_1125_sv2v_reg <= w_data_i[5];
      mem_1124_sv2v_reg <= w_data_i[4];
      mem_1123_sv2v_reg <= w_data_i[3];
      mem_1122_sv2v_reg <= w_data_i[2];
      mem_1121_sv2v_reg <= w_data_i[1];
      mem_1120_sv2v_reg <= w_data_i[0];
    end 
    if(N408) begin
      mem_1119_sv2v_reg <= w_data_i[31];
      mem_1118_sv2v_reg <= w_data_i[30];
      mem_1117_sv2v_reg <= w_data_i[29];
      mem_1116_sv2v_reg <= w_data_i[28];
      mem_1115_sv2v_reg <= w_data_i[27];
      mem_1114_sv2v_reg <= w_data_i[26];
      mem_1113_sv2v_reg <= w_data_i[25];
      mem_1112_sv2v_reg <= w_data_i[24];
      mem_1111_sv2v_reg <= w_data_i[23];
      mem_1110_sv2v_reg <= w_data_i[22];
      mem_1109_sv2v_reg <= w_data_i[21];
      mem_1108_sv2v_reg <= w_data_i[20];
      mem_1107_sv2v_reg <= w_data_i[19];
      mem_1106_sv2v_reg <= w_data_i[18];
      mem_1105_sv2v_reg <= w_data_i[17];
      mem_1104_sv2v_reg <= w_data_i[16];
      mem_1103_sv2v_reg <= w_data_i[15];
      mem_1102_sv2v_reg <= w_data_i[14];
      mem_1101_sv2v_reg <= w_data_i[13];
      mem_1100_sv2v_reg <= w_data_i[12];
      mem_1099_sv2v_reg <= w_data_i[11];
      mem_1098_sv2v_reg <= w_data_i[10];
      mem_1097_sv2v_reg <= w_data_i[9];
      mem_1096_sv2v_reg <= w_data_i[8];
      mem_1095_sv2v_reg <= w_data_i[7];
      mem_1094_sv2v_reg <= w_data_i[6];
      mem_1093_sv2v_reg <= w_data_i[5];
      mem_1092_sv2v_reg <= w_data_i[4];
      mem_1091_sv2v_reg <= w_data_i[3];
      mem_1090_sv2v_reg <= w_data_i[2];
      mem_1089_sv2v_reg <= w_data_i[1];
      mem_1088_sv2v_reg <= w_data_i[0];
    end 
    if(N407) begin
      mem_1087_sv2v_reg <= w_data_i[31];
      mem_1086_sv2v_reg <= w_data_i[30];
      mem_1085_sv2v_reg <= w_data_i[29];
      mem_1084_sv2v_reg <= w_data_i[28];
      mem_1083_sv2v_reg <= w_data_i[27];
      mem_1082_sv2v_reg <= w_data_i[26];
      mem_1081_sv2v_reg <= w_data_i[25];
      mem_1080_sv2v_reg <= w_data_i[24];
      mem_1079_sv2v_reg <= w_data_i[23];
      mem_1078_sv2v_reg <= w_data_i[22];
      mem_1077_sv2v_reg <= w_data_i[21];
      mem_1076_sv2v_reg <= w_data_i[20];
      mem_1075_sv2v_reg <= w_data_i[19];
      mem_1074_sv2v_reg <= w_data_i[18];
      mem_1073_sv2v_reg <= w_data_i[17];
      mem_1072_sv2v_reg <= w_data_i[16];
      mem_1071_sv2v_reg <= w_data_i[15];
      mem_1070_sv2v_reg <= w_data_i[14];
      mem_1069_sv2v_reg <= w_data_i[13];
      mem_1068_sv2v_reg <= w_data_i[12];
      mem_1067_sv2v_reg <= w_data_i[11];
      mem_1066_sv2v_reg <= w_data_i[10];
      mem_1065_sv2v_reg <= w_data_i[9];
      mem_1064_sv2v_reg <= w_data_i[8];
      mem_1063_sv2v_reg <= w_data_i[7];
      mem_1062_sv2v_reg <= w_data_i[6];
      mem_1061_sv2v_reg <= w_data_i[5];
      mem_1060_sv2v_reg <= w_data_i[4];
      mem_1059_sv2v_reg <= w_data_i[3];
      mem_1058_sv2v_reg <= w_data_i[2];
      mem_1057_sv2v_reg <= w_data_i[1];
      mem_1056_sv2v_reg <= w_data_i[0];
    end 
    if(N406) begin
      mem_1055_sv2v_reg <= w_data_i[31];
      mem_1054_sv2v_reg <= w_data_i[30];
      mem_1053_sv2v_reg <= w_data_i[29];
      mem_1052_sv2v_reg <= w_data_i[28];
      mem_1051_sv2v_reg <= w_data_i[27];
      mem_1050_sv2v_reg <= w_data_i[26];
      mem_1049_sv2v_reg <= w_data_i[25];
      mem_1048_sv2v_reg <= w_data_i[24];
      mem_1047_sv2v_reg <= w_data_i[23];
      mem_1046_sv2v_reg <= w_data_i[22];
      mem_1045_sv2v_reg <= w_data_i[21];
      mem_1044_sv2v_reg <= w_data_i[20];
      mem_1043_sv2v_reg <= w_data_i[19];
      mem_1042_sv2v_reg <= w_data_i[18];
      mem_1041_sv2v_reg <= w_data_i[17];
      mem_1040_sv2v_reg <= w_data_i[16];
      mem_1039_sv2v_reg <= w_data_i[15];
      mem_1038_sv2v_reg <= w_data_i[14];
      mem_1037_sv2v_reg <= w_data_i[13];
      mem_1036_sv2v_reg <= w_data_i[12];
      mem_1035_sv2v_reg <= w_data_i[11];
      mem_1034_sv2v_reg <= w_data_i[10];
      mem_1033_sv2v_reg <= w_data_i[9];
      mem_1032_sv2v_reg <= w_data_i[8];
      mem_1031_sv2v_reg <= w_data_i[7];
      mem_1030_sv2v_reg <= w_data_i[6];
      mem_1029_sv2v_reg <= w_data_i[5];
      mem_1028_sv2v_reg <= w_data_i[4];
      mem_1027_sv2v_reg <= w_data_i[3];
      mem_1026_sv2v_reg <= w_data_i[2];
      mem_1025_sv2v_reg <= w_data_i[1];
      mem_1024_sv2v_reg <= w_data_i[0];
    end 
    if(N405) begin
      mem_1023_sv2v_reg <= w_data_i[31];
      mem_1022_sv2v_reg <= w_data_i[30];
      mem_1021_sv2v_reg <= w_data_i[29];
      mem_1020_sv2v_reg <= w_data_i[28];
      mem_1019_sv2v_reg <= w_data_i[27];
      mem_1018_sv2v_reg <= w_data_i[26];
      mem_1017_sv2v_reg <= w_data_i[25];
      mem_1016_sv2v_reg <= w_data_i[24];
      mem_1015_sv2v_reg <= w_data_i[23];
      mem_1014_sv2v_reg <= w_data_i[22];
      mem_1013_sv2v_reg <= w_data_i[21];
      mem_1012_sv2v_reg <= w_data_i[20];
      mem_1011_sv2v_reg <= w_data_i[19];
      mem_1010_sv2v_reg <= w_data_i[18];
      mem_1009_sv2v_reg <= w_data_i[17];
      mem_1008_sv2v_reg <= w_data_i[16];
      mem_1007_sv2v_reg <= w_data_i[15];
      mem_1006_sv2v_reg <= w_data_i[14];
      mem_1005_sv2v_reg <= w_data_i[13];
      mem_1004_sv2v_reg <= w_data_i[12];
      mem_1003_sv2v_reg <= w_data_i[11];
      mem_1002_sv2v_reg <= w_data_i[10];
      mem_1001_sv2v_reg <= w_data_i[9];
      mem_1000_sv2v_reg <= w_data_i[8];
      mem_999_sv2v_reg <= w_data_i[7];
      mem_998_sv2v_reg <= w_data_i[6];
      mem_997_sv2v_reg <= w_data_i[5];
      mem_996_sv2v_reg <= w_data_i[4];
      mem_995_sv2v_reg <= w_data_i[3];
      mem_994_sv2v_reg <= w_data_i[2];
      mem_993_sv2v_reg <= w_data_i[1];
      mem_992_sv2v_reg <= w_data_i[0];
    end 
    if(N404) begin
      mem_991_sv2v_reg <= w_data_i[31];
      mem_990_sv2v_reg <= w_data_i[30];
      mem_989_sv2v_reg <= w_data_i[29];
      mem_988_sv2v_reg <= w_data_i[28];
      mem_987_sv2v_reg <= w_data_i[27];
      mem_986_sv2v_reg <= w_data_i[26];
      mem_985_sv2v_reg <= w_data_i[25];
      mem_984_sv2v_reg <= w_data_i[24];
      mem_983_sv2v_reg <= w_data_i[23];
      mem_982_sv2v_reg <= w_data_i[22];
      mem_981_sv2v_reg <= w_data_i[21];
      mem_980_sv2v_reg <= w_data_i[20];
      mem_979_sv2v_reg <= w_data_i[19];
      mem_978_sv2v_reg <= w_data_i[18];
      mem_977_sv2v_reg <= w_data_i[17];
      mem_976_sv2v_reg <= w_data_i[16];
      mem_975_sv2v_reg <= w_data_i[15];
      mem_974_sv2v_reg <= w_data_i[14];
      mem_973_sv2v_reg <= w_data_i[13];
      mem_972_sv2v_reg <= w_data_i[12];
      mem_971_sv2v_reg <= w_data_i[11];
      mem_970_sv2v_reg <= w_data_i[10];
      mem_969_sv2v_reg <= w_data_i[9];
      mem_968_sv2v_reg <= w_data_i[8];
      mem_967_sv2v_reg <= w_data_i[7];
      mem_966_sv2v_reg <= w_data_i[6];
      mem_965_sv2v_reg <= w_data_i[5];
      mem_964_sv2v_reg <= w_data_i[4];
      mem_963_sv2v_reg <= w_data_i[3];
      mem_962_sv2v_reg <= w_data_i[2];
      mem_961_sv2v_reg <= w_data_i[1];
      mem_960_sv2v_reg <= w_data_i[0];
    end 
    if(N403) begin
      mem_959_sv2v_reg <= w_data_i[31];
      mem_958_sv2v_reg <= w_data_i[30];
      mem_957_sv2v_reg <= w_data_i[29];
      mem_956_sv2v_reg <= w_data_i[28];
      mem_955_sv2v_reg <= w_data_i[27];
      mem_954_sv2v_reg <= w_data_i[26];
      mem_953_sv2v_reg <= w_data_i[25];
      mem_952_sv2v_reg <= w_data_i[24];
      mem_951_sv2v_reg <= w_data_i[23];
      mem_950_sv2v_reg <= w_data_i[22];
      mem_949_sv2v_reg <= w_data_i[21];
      mem_948_sv2v_reg <= w_data_i[20];
      mem_947_sv2v_reg <= w_data_i[19];
      mem_946_sv2v_reg <= w_data_i[18];
      mem_945_sv2v_reg <= w_data_i[17];
      mem_944_sv2v_reg <= w_data_i[16];
      mem_943_sv2v_reg <= w_data_i[15];
      mem_942_sv2v_reg <= w_data_i[14];
      mem_941_sv2v_reg <= w_data_i[13];
      mem_940_sv2v_reg <= w_data_i[12];
      mem_939_sv2v_reg <= w_data_i[11];
      mem_938_sv2v_reg <= w_data_i[10];
      mem_937_sv2v_reg <= w_data_i[9];
      mem_936_sv2v_reg <= w_data_i[8];
      mem_935_sv2v_reg <= w_data_i[7];
      mem_934_sv2v_reg <= w_data_i[6];
      mem_933_sv2v_reg <= w_data_i[5];
      mem_932_sv2v_reg <= w_data_i[4];
      mem_931_sv2v_reg <= w_data_i[3];
      mem_930_sv2v_reg <= w_data_i[2];
      mem_929_sv2v_reg <= w_data_i[1];
      mem_928_sv2v_reg <= w_data_i[0];
    end 
    if(N402) begin
      mem_927_sv2v_reg <= w_data_i[31];
      mem_926_sv2v_reg <= w_data_i[30];
      mem_925_sv2v_reg <= w_data_i[29];
      mem_924_sv2v_reg <= w_data_i[28];
      mem_923_sv2v_reg <= w_data_i[27];
      mem_922_sv2v_reg <= w_data_i[26];
      mem_921_sv2v_reg <= w_data_i[25];
      mem_920_sv2v_reg <= w_data_i[24];
      mem_919_sv2v_reg <= w_data_i[23];
      mem_918_sv2v_reg <= w_data_i[22];
      mem_917_sv2v_reg <= w_data_i[21];
      mem_916_sv2v_reg <= w_data_i[20];
      mem_915_sv2v_reg <= w_data_i[19];
      mem_914_sv2v_reg <= w_data_i[18];
      mem_913_sv2v_reg <= w_data_i[17];
      mem_912_sv2v_reg <= w_data_i[16];
      mem_911_sv2v_reg <= w_data_i[15];
      mem_910_sv2v_reg <= w_data_i[14];
      mem_909_sv2v_reg <= w_data_i[13];
      mem_908_sv2v_reg <= w_data_i[12];
      mem_907_sv2v_reg <= w_data_i[11];
      mem_906_sv2v_reg <= w_data_i[10];
      mem_905_sv2v_reg <= w_data_i[9];
      mem_904_sv2v_reg <= w_data_i[8];
      mem_903_sv2v_reg <= w_data_i[7];
      mem_902_sv2v_reg <= w_data_i[6];
      mem_901_sv2v_reg <= w_data_i[5];
      mem_900_sv2v_reg <= w_data_i[4];
      mem_899_sv2v_reg <= w_data_i[3];
      mem_898_sv2v_reg <= w_data_i[2];
      mem_897_sv2v_reg <= w_data_i[1];
      mem_896_sv2v_reg <= w_data_i[0];
    end 
    if(N401) begin
      mem_895_sv2v_reg <= w_data_i[31];
      mem_894_sv2v_reg <= w_data_i[30];
      mem_893_sv2v_reg <= w_data_i[29];
      mem_892_sv2v_reg <= w_data_i[28];
      mem_891_sv2v_reg <= w_data_i[27];
      mem_890_sv2v_reg <= w_data_i[26];
      mem_889_sv2v_reg <= w_data_i[25];
      mem_888_sv2v_reg <= w_data_i[24];
      mem_887_sv2v_reg <= w_data_i[23];
      mem_886_sv2v_reg <= w_data_i[22];
      mem_885_sv2v_reg <= w_data_i[21];
      mem_884_sv2v_reg <= w_data_i[20];
      mem_883_sv2v_reg <= w_data_i[19];
      mem_882_sv2v_reg <= w_data_i[18];
      mem_881_sv2v_reg <= w_data_i[17];
      mem_880_sv2v_reg <= w_data_i[16];
      mem_879_sv2v_reg <= w_data_i[15];
      mem_878_sv2v_reg <= w_data_i[14];
      mem_877_sv2v_reg <= w_data_i[13];
      mem_876_sv2v_reg <= w_data_i[12];
      mem_875_sv2v_reg <= w_data_i[11];
      mem_874_sv2v_reg <= w_data_i[10];
      mem_873_sv2v_reg <= w_data_i[9];
      mem_872_sv2v_reg <= w_data_i[8];
      mem_871_sv2v_reg <= w_data_i[7];
      mem_870_sv2v_reg <= w_data_i[6];
      mem_869_sv2v_reg <= w_data_i[5];
      mem_868_sv2v_reg <= w_data_i[4];
      mem_867_sv2v_reg <= w_data_i[3];
      mem_866_sv2v_reg <= w_data_i[2];
      mem_865_sv2v_reg <= w_data_i[1];
      mem_864_sv2v_reg <= w_data_i[0];
    end 
    if(N400) begin
      mem_863_sv2v_reg <= w_data_i[31];
      mem_862_sv2v_reg <= w_data_i[30];
      mem_861_sv2v_reg <= w_data_i[29];
      mem_860_sv2v_reg <= w_data_i[28];
      mem_859_sv2v_reg <= w_data_i[27];
      mem_858_sv2v_reg <= w_data_i[26];
      mem_857_sv2v_reg <= w_data_i[25];
      mem_856_sv2v_reg <= w_data_i[24];
      mem_855_sv2v_reg <= w_data_i[23];
      mem_854_sv2v_reg <= w_data_i[22];
      mem_853_sv2v_reg <= w_data_i[21];
      mem_852_sv2v_reg <= w_data_i[20];
      mem_851_sv2v_reg <= w_data_i[19];
      mem_850_sv2v_reg <= w_data_i[18];
      mem_849_sv2v_reg <= w_data_i[17];
      mem_848_sv2v_reg <= w_data_i[16];
      mem_847_sv2v_reg <= w_data_i[15];
      mem_846_sv2v_reg <= w_data_i[14];
      mem_845_sv2v_reg <= w_data_i[13];
      mem_844_sv2v_reg <= w_data_i[12];
      mem_843_sv2v_reg <= w_data_i[11];
      mem_842_sv2v_reg <= w_data_i[10];
      mem_841_sv2v_reg <= w_data_i[9];
      mem_840_sv2v_reg <= w_data_i[8];
      mem_839_sv2v_reg <= w_data_i[7];
      mem_838_sv2v_reg <= w_data_i[6];
      mem_837_sv2v_reg <= w_data_i[5];
      mem_836_sv2v_reg <= w_data_i[4];
      mem_835_sv2v_reg <= w_data_i[3];
      mem_834_sv2v_reg <= w_data_i[2];
      mem_833_sv2v_reg <= w_data_i[1];
      mem_832_sv2v_reg <= w_data_i[0];
    end 
    if(N399) begin
      mem_831_sv2v_reg <= w_data_i[31];
      mem_830_sv2v_reg <= w_data_i[30];
      mem_829_sv2v_reg <= w_data_i[29];
      mem_828_sv2v_reg <= w_data_i[28];
      mem_827_sv2v_reg <= w_data_i[27];
      mem_826_sv2v_reg <= w_data_i[26];
      mem_825_sv2v_reg <= w_data_i[25];
      mem_824_sv2v_reg <= w_data_i[24];
      mem_823_sv2v_reg <= w_data_i[23];
      mem_822_sv2v_reg <= w_data_i[22];
      mem_821_sv2v_reg <= w_data_i[21];
      mem_820_sv2v_reg <= w_data_i[20];
      mem_819_sv2v_reg <= w_data_i[19];
      mem_818_sv2v_reg <= w_data_i[18];
      mem_817_sv2v_reg <= w_data_i[17];
      mem_816_sv2v_reg <= w_data_i[16];
      mem_815_sv2v_reg <= w_data_i[15];
      mem_814_sv2v_reg <= w_data_i[14];
      mem_813_sv2v_reg <= w_data_i[13];
      mem_812_sv2v_reg <= w_data_i[12];
      mem_811_sv2v_reg <= w_data_i[11];
      mem_810_sv2v_reg <= w_data_i[10];
      mem_809_sv2v_reg <= w_data_i[9];
      mem_808_sv2v_reg <= w_data_i[8];
      mem_807_sv2v_reg <= w_data_i[7];
      mem_806_sv2v_reg <= w_data_i[6];
      mem_805_sv2v_reg <= w_data_i[5];
      mem_804_sv2v_reg <= w_data_i[4];
      mem_803_sv2v_reg <= w_data_i[3];
      mem_802_sv2v_reg <= w_data_i[2];
      mem_801_sv2v_reg <= w_data_i[1];
      mem_800_sv2v_reg <= w_data_i[0];
    end 
    if(N398) begin
      mem_799_sv2v_reg <= w_data_i[31];
      mem_798_sv2v_reg <= w_data_i[30];
      mem_797_sv2v_reg <= w_data_i[29];
      mem_796_sv2v_reg <= w_data_i[28];
      mem_795_sv2v_reg <= w_data_i[27];
      mem_794_sv2v_reg <= w_data_i[26];
      mem_793_sv2v_reg <= w_data_i[25];
      mem_792_sv2v_reg <= w_data_i[24];
      mem_791_sv2v_reg <= w_data_i[23];
      mem_790_sv2v_reg <= w_data_i[22];
      mem_789_sv2v_reg <= w_data_i[21];
      mem_788_sv2v_reg <= w_data_i[20];
      mem_787_sv2v_reg <= w_data_i[19];
      mem_786_sv2v_reg <= w_data_i[18];
      mem_785_sv2v_reg <= w_data_i[17];
      mem_784_sv2v_reg <= w_data_i[16];
      mem_783_sv2v_reg <= w_data_i[15];
      mem_782_sv2v_reg <= w_data_i[14];
      mem_781_sv2v_reg <= w_data_i[13];
      mem_780_sv2v_reg <= w_data_i[12];
      mem_779_sv2v_reg <= w_data_i[11];
      mem_778_sv2v_reg <= w_data_i[10];
      mem_777_sv2v_reg <= w_data_i[9];
      mem_776_sv2v_reg <= w_data_i[8];
      mem_775_sv2v_reg <= w_data_i[7];
      mem_774_sv2v_reg <= w_data_i[6];
      mem_773_sv2v_reg <= w_data_i[5];
      mem_772_sv2v_reg <= w_data_i[4];
      mem_771_sv2v_reg <= w_data_i[3];
      mem_770_sv2v_reg <= w_data_i[2];
      mem_769_sv2v_reg <= w_data_i[1];
      mem_768_sv2v_reg <= w_data_i[0];
    end 
    if(N397) begin
      mem_767_sv2v_reg <= w_data_i[31];
      mem_766_sv2v_reg <= w_data_i[30];
      mem_765_sv2v_reg <= w_data_i[29];
      mem_764_sv2v_reg <= w_data_i[28];
      mem_763_sv2v_reg <= w_data_i[27];
      mem_762_sv2v_reg <= w_data_i[26];
      mem_761_sv2v_reg <= w_data_i[25];
      mem_760_sv2v_reg <= w_data_i[24];
      mem_759_sv2v_reg <= w_data_i[23];
      mem_758_sv2v_reg <= w_data_i[22];
      mem_757_sv2v_reg <= w_data_i[21];
      mem_756_sv2v_reg <= w_data_i[20];
      mem_755_sv2v_reg <= w_data_i[19];
      mem_754_sv2v_reg <= w_data_i[18];
      mem_753_sv2v_reg <= w_data_i[17];
      mem_752_sv2v_reg <= w_data_i[16];
      mem_751_sv2v_reg <= w_data_i[15];
      mem_750_sv2v_reg <= w_data_i[14];
      mem_749_sv2v_reg <= w_data_i[13];
      mem_748_sv2v_reg <= w_data_i[12];
      mem_747_sv2v_reg <= w_data_i[11];
      mem_746_sv2v_reg <= w_data_i[10];
      mem_745_sv2v_reg <= w_data_i[9];
      mem_744_sv2v_reg <= w_data_i[8];
      mem_743_sv2v_reg <= w_data_i[7];
      mem_742_sv2v_reg <= w_data_i[6];
      mem_741_sv2v_reg <= w_data_i[5];
      mem_740_sv2v_reg <= w_data_i[4];
      mem_739_sv2v_reg <= w_data_i[3];
      mem_738_sv2v_reg <= w_data_i[2];
      mem_737_sv2v_reg <= w_data_i[1];
      mem_736_sv2v_reg <= w_data_i[0];
    end 
    if(N396) begin
      mem_735_sv2v_reg <= w_data_i[31];
      mem_734_sv2v_reg <= w_data_i[30];
      mem_733_sv2v_reg <= w_data_i[29];
      mem_732_sv2v_reg <= w_data_i[28];
      mem_731_sv2v_reg <= w_data_i[27];
      mem_730_sv2v_reg <= w_data_i[26];
      mem_729_sv2v_reg <= w_data_i[25];
      mem_728_sv2v_reg <= w_data_i[24];
      mem_727_sv2v_reg <= w_data_i[23];
      mem_726_sv2v_reg <= w_data_i[22];
      mem_725_sv2v_reg <= w_data_i[21];
      mem_724_sv2v_reg <= w_data_i[20];
      mem_723_sv2v_reg <= w_data_i[19];
      mem_722_sv2v_reg <= w_data_i[18];
      mem_721_sv2v_reg <= w_data_i[17];
      mem_720_sv2v_reg <= w_data_i[16];
      mem_719_sv2v_reg <= w_data_i[15];
      mem_718_sv2v_reg <= w_data_i[14];
      mem_717_sv2v_reg <= w_data_i[13];
      mem_716_sv2v_reg <= w_data_i[12];
      mem_715_sv2v_reg <= w_data_i[11];
      mem_714_sv2v_reg <= w_data_i[10];
      mem_713_sv2v_reg <= w_data_i[9];
      mem_712_sv2v_reg <= w_data_i[8];
      mem_711_sv2v_reg <= w_data_i[7];
      mem_710_sv2v_reg <= w_data_i[6];
      mem_709_sv2v_reg <= w_data_i[5];
      mem_708_sv2v_reg <= w_data_i[4];
      mem_707_sv2v_reg <= w_data_i[3];
      mem_706_sv2v_reg <= w_data_i[2];
      mem_705_sv2v_reg <= w_data_i[1];
      mem_704_sv2v_reg <= w_data_i[0];
    end 
    if(N395) begin
      mem_703_sv2v_reg <= w_data_i[31];
      mem_702_sv2v_reg <= w_data_i[30];
      mem_701_sv2v_reg <= w_data_i[29];
      mem_700_sv2v_reg <= w_data_i[28];
      mem_699_sv2v_reg <= w_data_i[27];
      mem_698_sv2v_reg <= w_data_i[26];
      mem_697_sv2v_reg <= w_data_i[25];
      mem_696_sv2v_reg <= w_data_i[24];
      mem_695_sv2v_reg <= w_data_i[23];
      mem_694_sv2v_reg <= w_data_i[22];
      mem_693_sv2v_reg <= w_data_i[21];
      mem_692_sv2v_reg <= w_data_i[20];
      mem_691_sv2v_reg <= w_data_i[19];
      mem_690_sv2v_reg <= w_data_i[18];
      mem_689_sv2v_reg <= w_data_i[17];
      mem_688_sv2v_reg <= w_data_i[16];
      mem_687_sv2v_reg <= w_data_i[15];
      mem_686_sv2v_reg <= w_data_i[14];
      mem_685_sv2v_reg <= w_data_i[13];
      mem_684_sv2v_reg <= w_data_i[12];
      mem_683_sv2v_reg <= w_data_i[11];
      mem_682_sv2v_reg <= w_data_i[10];
      mem_681_sv2v_reg <= w_data_i[9];
      mem_680_sv2v_reg <= w_data_i[8];
      mem_679_sv2v_reg <= w_data_i[7];
      mem_678_sv2v_reg <= w_data_i[6];
      mem_677_sv2v_reg <= w_data_i[5];
      mem_676_sv2v_reg <= w_data_i[4];
      mem_675_sv2v_reg <= w_data_i[3];
      mem_674_sv2v_reg <= w_data_i[2];
      mem_673_sv2v_reg <= w_data_i[1];
      mem_672_sv2v_reg <= w_data_i[0];
    end 
    if(N394) begin
      mem_671_sv2v_reg <= w_data_i[31];
      mem_670_sv2v_reg <= w_data_i[30];
      mem_669_sv2v_reg <= w_data_i[29];
      mem_668_sv2v_reg <= w_data_i[28];
      mem_667_sv2v_reg <= w_data_i[27];
      mem_666_sv2v_reg <= w_data_i[26];
      mem_665_sv2v_reg <= w_data_i[25];
      mem_664_sv2v_reg <= w_data_i[24];
      mem_663_sv2v_reg <= w_data_i[23];
      mem_662_sv2v_reg <= w_data_i[22];
      mem_661_sv2v_reg <= w_data_i[21];
      mem_660_sv2v_reg <= w_data_i[20];
      mem_659_sv2v_reg <= w_data_i[19];
      mem_658_sv2v_reg <= w_data_i[18];
      mem_657_sv2v_reg <= w_data_i[17];
      mem_656_sv2v_reg <= w_data_i[16];
      mem_655_sv2v_reg <= w_data_i[15];
      mem_654_sv2v_reg <= w_data_i[14];
      mem_653_sv2v_reg <= w_data_i[13];
      mem_652_sv2v_reg <= w_data_i[12];
      mem_651_sv2v_reg <= w_data_i[11];
      mem_650_sv2v_reg <= w_data_i[10];
      mem_649_sv2v_reg <= w_data_i[9];
      mem_648_sv2v_reg <= w_data_i[8];
      mem_647_sv2v_reg <= w_data_i[7];
      mem_646_sv2v_reg <= w_data_i[6];
      mem_645_sv2v_reg <= w_data_i[5];
      mem_644_sv2v_reg <= w_data_i[4];
      mem_643_sv2v_reg <= w_data_i[3];
      mem_642_sv2v_reg <= w_data_i[2];
      mem_641_sv2v_reg <= w_data_i[1];
      mem_640_sv2v_reg <= w_data_i[0];
    end 
    if(N393) begin
      mem_639_sv2v_reg <= w_data_i[31];
      mem_638_sv2v_reg <= w_data_i[30];
      mem_637_sv2v_reg <= w_data_i[29];
      mem_636_sv2v_reg <= w_data_i[28];
      mem_635_sv2v_reg <= w_data_i[27];
      mem_634_sv2v_reg <= w_data_i[26];
      mem_633_sv2v_reg <= w_data_i[25];
      mem_632_sv2v_reg <= w_data_i[24];
      mem_631_sv2v_reg <= w_data_i[23];
      mem_630_sv2v_reg <= w_data_i[22];
      mem_629_sv2v_reg <= w_data_i[21];
      mem_628_sv2v_reg <= w_data_i[20];
      mem_627_sv2v_reg <= w_data_i[19];
      mem_626_sv2v_reg <= w_data_i[18];
      mem_625_sv2v_reg <= w_data_i[17];
      mem_624_sv2v_reg <= w_data_i[16];
      mem_623_sv2v_reg <= w_data_i[15];
      mem_622_sv2v_reg <= w_data_i[14];
      mem_621_sv2v_reg <= w_data_i[13];
      mem_620_sv2v_reg <= w_data_i[12];
      mem_619_sv2v_reg <= w_data_i[11];
      mem_618_sv2v_reg <= w_data_i[10];
      mem_617_sv2v_reg <= w_data_i[9];
      mem_616_sv2v_reg <= w_data_i[8];
      mem_615_sv2v_reg <= w_data_i[7];
      mem_614_sv2v_reg <= w_data_i[6];
      mem_613_sv2v_reg <= w_data_i[5];
      mem_612_sv2v_reg <= w_data_i[4];
      mem_611_sv2v_reg <= w_data_i[3];
      mem_610_sv2v_reg <= w_data_i[2];
      mem_609_sv2v_reg <= w_data_i[1];
      mem_608_sv2v_reg <= w_data_i[0];
    end 
    if(N392) begin
      mem_607_sv2v_reg <= w_data_i[31];
      mem_606_sv2v_reg <= w_data_i[30];
      mem_605_sv2v_reg <= w_data_i[29];
      mem_604_sv2v_reg <= w_data_i[28];
      mem_603_sv2v_reg <= w_data_i[27];
      mem_602_sv2v_reg <= w_data_i[26];
      mem_601_sv2v_reg <= w_data_i[25];
      mem_600_sv2v_reg <= w_data_i[24];
      mem_599_sv2v_reg <= w_data_i[23];
      mem_598_sv2v_reg <= w_data_i[22];
      mem_597_sv2v_reg <= w_data_i[21];
      mem_596_sv2v_reg <= w_data_i[20];
      mem_595_sv2v_reg <= w_data_i[19];
      mem_594_sv2v_reg <= w_data_i[18];
      mem_593_sv2v_reg <= w_data_i[17];
      mem_592_sv2v_reg <= w_data_i[16];
      mem_591_sv2v_reg <= w_data_i[15];
      mem_590_sv2v_reg <= w_data_i[14];
      mem_589_sv2v_reg <= w_data_i[13];
      mem_588_sv2v_reg <= w_data_i[12];
      mem_587_sv2v_reg <= w_data_i[11];
      mem_586_sv2v_reg <= w_data_i[10];
      mem_585_sv2v_reg <= w_data_i[9];
      mem_584_sv2v_reg <= w_data_i[8];
      mem_583_sv2v_reg <= w_data_i[7];
      mem_582_sv2v_reg <= w_data_i[6];
      mem_581_sv2v_reg <= w_data_i[5];
      mem_580_sv2v_reg <= w_data_i[4];
      mem_579_sv2v_reg <= w_data_i[3];
      mem_578_sv2v_reg <= w_data_i[2];
      mem_577_sv2v_reg <= w_data_i[1];
      mem_576_sv2v_reg <= w_data_i[0];
    end 
    if(N391) begin
      mem_575_sv2v_reg <= w_data_i[31];
      mem_574_sv2v_reg <= w_data_i[30];
      mem_573_sv2v_reg <= w_data_i[29];
      mem_572_sv2v_reg <= w_data_i[28];
      mem_571_sv2v_reg <= w_data_i[27];
      mem_570_sv2v_reg <= w_data_i[26];
      mem_569_sv2v_reg <= w_data_i[25];
      mem_568_sv2v_reg <= w_data_i[24];
      mem_567_sv2v_reg <= w_data_i[23];
      mem_566_sv2v_reg <= w_data_i[22];
      mem_565_sv2v_reg <= w_data_i[21];
      mem_564_sv2v_reg <= w_data_i[20];
      mem_563_sv2v_reg <= w_data_i[19];
      mem_562_sv2v_reg <= w_data_i[18];
      mem_561_sv2v_reg <= w_data_i[17];
      mem_560_sv2v_reg <= w_data_i[16];
      mem_559_sv2v_reg <= w_data_i[15];
      mem_558_sv2v_reg <= w_data_i[14];
      mem_557_sv2v_reg <= w_data_i[13];
      mem_556_sv2v_reg <= w_data_i[12];
      mem_555_sv2v_reg <= w_data_i[11];
      mem_554_sv2v_reg <= w_data_i[10];
      mem_553_sv2v_reg <= w_data_i[9];
      mem_552_sv2v_reg <= w_data_i[8];
      mem_551_sv2v_reg <= w_data_i[7];
      mem_550_sv2v_reg <= w_data_i[6];
      mem_549_sv2v_reg <= w_data_i[5];
      mem_548_sv2v_reg <= w_data_i[4];
      mem_547_sv2v_reg <= w_data_i[3];
      mem_546_sv2v_reg <= w_data_i[2];
      mem_545_sv2v_reg <= w_data_i[1];
      mem_544_sv2v_reg <= w_data_i[0];
    end 
    if(N390) begin
      mem_543_sv2v_reg <= w_data_i[31];
      mem_542_sv2v_reg <= w_data_i[30];
      mem_541_sv2v_reg <= w_data_i[29];
      mem_540_sv2v_reg <= w_data_i[28];
      mem_539_sv2v_reg <= w_data_i[27];
      mem_538_sv2v_reg <= w_data_i[26];
      mem_537_sv2v_reg <= w_data_i[25];
      mem_536_sv2v_reg <= w_data_i[24];
      mem_535_sv2v_reg <= w_data_i[23];
      mem_534_sv2v_reg <= w_data_i[22];
      mem_533_sv2v_reg <= w_data_i[21];
      mem_532_sv2v_reg <= w_data_i[20];
      mem_531_sv2v_reg <= w_data_i[19];
      mem_530_sv2v_reg <= w_data_i[18];
      mem_529_sv2v_reg <= w_data_i[17];
      mem_528_sv2v_reg <= w_data_i[16];
      mem_527_sv2v_reg <= w_data_i[15];
      mem_526_sv2v_reg <= w_data_i[14];
      mem_525_sv2v_reg <= w_data_i[13];
      mem_524_sv2v_reg <= w_data_i[12];
      mem_523_sv2v_reg <= w_data_i[11];
      mem_522_sv2v_reg <= w_data_i[10];
      mem_521_sv2v_reg <= w_data_i[9];
      mem_520_sv2v_reg <= w_data_i[8];
      mem_519_sv2v_reg <= w_data_i[7];
      mem_518_sv2v_reg <= w_data_i[6];
      mem_517_sv2v_reg <= w_data_i[5];
      mem_516_sv2v_reg <= w_data_i[4];
      mem_515_sv2v_reg <= w_data_i[3];
      mem_514_sv2v_reg <= w_data_i[2];
      mem_513_sv2v_reg <= w_data_i[1];
      mem_512_sv2v_reg <= w_data_i[0];
    end 
    if(N389) begin
      mem_511_sv2v_reg <= w_data_i[31];
      mem_510_sv2v_reg <= w_data_i[30];
      mem_509_sv2v_reg <= w_data_i[29];
      mem_508_sv2v_reg <= w_data_i[28];
      mem_507_sv2v_reg <= w_data_i[27];
      mem_506_sv2v_reg <= w_data_i[26];
      mem_505_sv2v_reg <= w_data_i[25];
      mem_504_sv2v_reg <= w_data_i[24];
      mem_503_sv2v_reg <= w_data_i[23];
      mem_502_sv2v_reg <= w_data_i[22];
      mem_501_sv2v_reg <= w_data_i[21];
      mem_500_sv2v_reg <= w_data_i[20];
      mem_499_sv2v_reg <= w_data_i[19];
      mem_498_sv2v_reg <= w_data_i[18];
      mem_497_sv2v_reg <= w_data_i[17];
      mem_496_sv2v_reg <= w_data_i[16];
      mem_495_sv2v_reg <= w_data_i[15];
      mem_494_sv2v_reg <= w_data_i[14];
      mem_493_sv2v_reg <= w_data_i[13];
      mem_492_sv2v_reg <= w_data_i[12];
      mem_491_sv2v_reg <= w_data_i[11];
      mem_490_sv2v_reg <= w_data_i[10];
      mem_489_sv2v_reg <= w_data_i[9];
      mem_488_sv2v_reg <= w_data_i[8];
      mem_487_sv2v_reg <= w_data_i[7];
      mem_486_sv2v_reg <= w_data_i[6];
      mem_485_sv2v_reg <= w_data_i[5];
      mem_484_sv2v_reg <= w_data_i[4];
      mem_483_sv2v_reg <= w_data_i[3];
      mem_482_sv2v_reg <= w_data_i[2];
      mem_481_sv2v_reg <= w_data_i[1];
      mem_480_sv2v_reg <= w_data_i[0];
    end 
    if(N388) begin
      mem_479_sv2v_reg <= w_data_i[31];
      mem_478_sv2v_reg <= w_data_i[30];
      mem_477_sv2v_reg <= w_data_i[29];
      mem_476_sv2v_reg <= w_data_i[28];
      mem_475_sv2v_reg <= w_data_i[27];
      mem_474_sv2v_reg <= w_data_i[26];
      mem_473_sv2v_reg <= w_data_i[25];
      mem_472_sv2v_reg <= w_data_i[24];
      mem_471_sv2v_reg <= w_data_i[23];
      mem_470_sv2v_reg <= w_data_i[22];
      mem_469_sv2v_reg <= w_data_i[21];
      mem_468_sv2v_reg <= w_data_i[20];
      mem_467_sv2v_reg <= w_data_i[19];
      mem_466_sv2v_reg <= w_data_i[18];
      mem_465_sv2v_reg <= w_data_i[17];
      mem_464_sv2v_reg <= w_data_i[16];
      mem_463_sv2v_reg <= w_data_i[15];
      mem_462_sv2v_reg <= w_data_i[14];
      mem_461_sv2v_reg <= w_data_i[13];
      mem_460_sv2v_reg <= w_data_i[12];
      mem_459_sv2v_reg <= w_data_i[11];
      mem_458_sv2v_reg <= w_data_i[10];
      mem_457_sv2v_reg <= w_data_i[9];
      mem_456_sv2v_reg <= w_data_i[8];
      mem_455_sv2v_reg <= w_data_i[7];
      mem_454_sv2v_reg <= w_data_i[6];
      mem_453_sv2v_reg <= w_data_i[5];
      mem_452_sv2v_reg <= w_data_i[4];
      mem_451_sv2v_reg <= w_data_i[3];
      mem_450_sv2v_reg <= w_data_i[2];
      mem_449_sv2v_reg <= w_data_i[1];
      mem_448_sv2v_reg <= w_data_i[0];
    end 
    if(N387) begin
      mem_447_sv2v_reg <= w_data_i[31];
      mem_446_sv2v_reg <= w_data_i[30];
      mem_445_sv2v_reg <= w_data_i[29];
      mem_444_sv2v_reg <= w_data_i[28];
      mem_443_sv2v_reg <= w_data_i[27];
      mem_442_sv2v_reg <= w_data_i[26];
      mem_441_sv2v_reg <= w_data_i[25];
      mem_440_sv2v_reg <= w_data_i[24];
      mem_439_sv2v_reg <= w_data_i[23];
      mem_438_sv2v_reg <= w_data_i[22];
      mem_437_sv2v_reg <= w_data_i[21];
      mem_436_sv2v_reg <= w_data_i[20];
      mem_435_sv2v_reg <= w_data_i[19];
      mem_434_sv2v_reg <= w_data_i[18];
      mem_433_sv2v_reg <= w_data_i[17];
      mem_432_sv2v_reg <= w_data_i[16];
      mem_431_sv2v_reg <= w_data_i[15];
      mem_430_sv2v_reg <= w_data_i[14];
      mem_429_sv2v_reg <= w_data_i[13];
      mem_428_sv2v_reg <= w_data_i[12];
      mem_427_sv2v_reg <= w_data_i[11];
      mem_426_sv2v_reg <= w_data_i[10];
      mem_425_sv2v_reg <= w_data_i[9];
      mem_424_sv2v_reg <= w_data_i[8];
      mem_423_sv2v_reg <= w_data_i[7];
      mem_422_sv2v_reg <= w_data_i[6];
      mem_421_sv2v_reg <= w_data_i[5];
      mem_420_sv2v_reg <= w_data_i[4];
      mem_419_sv2v_reg <= w_data_i[3];
      mem_418_sv2v_reg <= w_data_i[2];
      mem_417_sv2v_reg <= w_data_i[1];
      mem_416_sv2v_reg <= w_data_i[0];
    end 
    if(N386) begin
      mem_415_sv2v_reg <= w_data_i[31];
      mem_414_sv2v_reg <= w_data_i[30];
      mem_413_sv2v_reg <= w_data_i[29];
      mem_412_sv2v_reg <= w_data_i[28];
      mem_411_sv2v_reg <= w_data_i[27];
      mem_410_sv2v_reg <= w_data_i[26];
      mem_409_sv2v_reg <= w_data_i[25];
      mem_408_sv2v_reg <= w_data_i[24];
      mem_407_sv2v_reg <= w_data_i[23];
      mem_406_sv2v_reg <= w_data_i[22];
      mem_405_sv2v_reg <= w_data_i[21];
      mem_404_sv2v_reg <= w_data_i[20];
      mem_403_sv2v_reg <= w_data_i[19];
      mem_402_sv2v_reg <= w_data_i[18];
      mem_401_sv2v_reg <= w_data_i[17];
      mem_400_sv2v_reg <= w_data_i[16];
      mem_399_sv2v_reg <= w_data_i[15];
      mem_398_sv2v_reg <= w_data_i[14];
      mem_397_sv2v_reg <= w_data_i[13];
      mem_396_sv2v_reg <= w_data_i[12];
      mem_395_sv2v_reg <= w_data_i[11];
      mem_394_sv2v_reg <= w_data_i[10];
      mem_393_sv2v_reg <= w_data_i[9];
      mem_392_sv2v_reg <= w_data_i[8];
      mem_391_sv2v_reg <= w_data_i[7];
      mem_390_sv2v_reg <= w_data_i[6];
      mem_389_sv2v_reg <= w_data_i[5];
      mem_388_sv2v_reg <= w_data_i[4];
      mem_387_sv2v_reg <= w_data_i[3];
      mem_386_sv2v_reg <= w_data_i[2];
      mem_385_sv2v_reg <= w_data_i[1];
      mem_384_sv2v_reg <= w_data_i[0];
    end 
    if(N385) begin
      mem_383_sv2v_reg <= w_data_i[31];
      mem_382_sv2v_reg <= w_data_i[30];
      mem_381_sv2v_reg <= w_data_i[29];
      mem_380_sv2v_reg <= w_data_i[28];
      mem_379_sv2v_reg <= w_data_i[27];
      mem_378_sv2v_reg <= w_data_i[26];
      mem_377_sv2v_reg <= w_data_i[25];
      mem_376_sv2v_reg <= w_data_i[24];
      mem_375_sv2v_reg <= w_data_i[23];
      mem_374_sv2v_reg <= w_data_i[22];
      mem_373_sv2v_reg <= w_data_i[21];
      mem_372_sv2v_reg <= w_data_i[20];
      mem_371_sv2v_reg <= w_data_i[19];
      mem_370_sv2v_reg <= w_data_i[18];
      mem_369_sv2v_reg <= w_data_i[17];
      mem_368_sv2v_reg <= w_data_i[16];
      mem_367_sv2v_reg <= w_data_i[15];
      mem_366_sv2v_reg <= w_data_i[14];
      mem_365_sv2v_reg <= w_data_i[13];
      mem_364_sv2v_reg <= w_data_i[12];
      mem_363_sv2v_reg <= w_data_i[11];
      mem_362_sv2v_reg <= w_data_i[10];
      mem_361_sv2v_reg <= w_data_i[9];
      mem_360_sv2v_reg <= w_data_i[8];
      mem_359_sv2v_reg <= w_data_i[7];
      mem_358_sv2v_reg <= w_data_i[6];
      mem_357_sv2v_reg <= w_data_i[5];
      mem_356_sv2v_reg <= w_data_i[4];
      mem_355_sv2v_reg <= w_data_i[3];
      mem_354_sv2v_reg <= w_data_i[2];
      mem_353_sv2v_reg <= w_data_i[1];
      mem_352_sv2v_reg <= w_data_i[0];
    end 
    if(N384) begin
      mem_351_sv2v_reg <= w_data_i[31];
      mem_350_sv2v_reg <= w_data_i[30];
      mem_349_sv2v_reg <= w_data_i[29];
      mem_348_sv2v_reg <= w_data_i[28];
      mem_347_sv2v_reg <= w_data_i[27];
      mem_346_sv2v_reg <= w_data_i[26];
      mem_345_sv2v_reg <= w_data_i[25];
      mem_344_sv2v_reg <= w_data_i[24];
      mem_343_sv2v_reg <= w_data_i[23];
      mem_342_sv2v_reg <= w_data_i[22];
      mem_341_sv2v_reg <= w_data_i[21];
      mem_340_sv2v_reg <= w_data_i[20];
      mem_339_sv2v_reg <= w_data_i[19];
      mem_338_sv2v_reg <= w_data_i[18];
      mem_337_sv2v_reg <= w_data_i[17];
      mem_336_sv2v_reg <= w_data_i[16];
      mem_335_sv2v_reg <= w_data_i[15];
      mem_334_sv2v_reg <= w_data_i[14];
      mem_333_sv2v_reg <= w_data_i[13];
      mem_332_sv2v_reg <= w_data_i[12];
      mem_331_sv2v_reg <= w_data_i[11];
      mem_330_sv2v_reg <= w_data_i[10];
      mem_329_sv2v_reg <= w_data_i[9];
      mem_328_sv2v_reg <= w_data_i[8];
      mem_327_sv2v_reg <= w_data_i[7];
      mem_326_sv2v_reg <= w_data_i[6];
      mem_325_sv2v_reg <= w_data_i[5];
      mem_324_sv2v_reg <= w_data_i[4];
      mem_323_sv2v_reg <= w_data_i[3];
      mem_322_sv2v_reg <= w_data_i[2];
      mem_321_sv2v_reg <= w_data_i[1];
      mem_320_sv2v_reg <= w_data_i[0];
    end 
    if(N383) begin
      mem_319_sv2v_reg <= w_data_i[31];
      mem_318_sv2v_reg <= w_data_i[30];
      mem_317_sv2v_reg <= w_data_i[29];
      mem_316_sv2v_reg <= w_data_i[28];
      mem_315_sv2v_reg <= w_data_i[27];
      mem_314_sv2v_reg <= w_data_i[26];
      mem_313_sv2v_reg <= w_data_i[25];
      mem_312_sv2v_reg <= w_data_i[24];
      mem_311_sv2v_reg <= w_data_i[23];
      mem_310_sv2v_reg <= w_data_i[22];
      mem_309_sv2v_reg <= w_data_i[21];
      mem_308_sv2v_reg <= w_data_i[20];
      mem_307_sv2v_reg <= w_data_i[19];
      mem_306_sv2v_reg <= w_data_i[18];
      mem_305_sv2v_reg <= w_data_i[17];
      mem_304_sv2v_reg <= w_data_i[16];
      mem_303_sv2v_reg <= w_data_i[15];
      mem_302_sv2v_reg <= w_data_i[14];
      mem_301_sv2v_reg <= w_data_i[13];
      mem_300_sv2v_reg <= w_data_i[12];
      mem_299_sv2v_reg <= w_data_i[11];
      mem_298_sv2v_reg <= w_data_i[10];
      mem_297_sv2v_reg <= w_data_i[9];
      mem_296_sv2v_reg <= w_data_i[8];
      mem_295_sv2v_reg <= w_data_i[7];
      mem_294_sv2v_reg <= w_data_i[6];
      mem_293_sv2v_reg <= w_data_i[5];
      mem_292_sv2v_reg <= w_data_i[4];
      mem_291_sv2v_reg <= w_data_i[3];
      mem_290_sv2v_reg <= w_data_i[2];
      mem_289_sv2v_reg <= w_data_i[1];
      mem_288_sv2v_reg <= w_data_i[0];
    end 
    if(N382) begin
      mem_287_sv2v_reg <= w_data_i[31];
      mem_286_sv2v_reg <= w_data_i[30];
      mem_285_sv2v_reg <= w_data_i[29];
      mem_284_sv2v_reg <= w_data_i[28];
      mem_283_sv2v_reg <= w_data_i[27];
      mem_282_sv2v_reg <= w_data_i[26];
      mem_281_sv2v_reg <= w_data_i[25];
      mem_280_sv2v_reg <= w_data_i[24];
      mem_279_sv2v_reg <= w_data_i[23];
      mem_278_sv2v_reg <= w_data_i[22];
      mem_277_sv2v_reg <= w_data_i[21];
      mem_276_sv2v_reg <= w_data_i[20];
      mem_275_sv2v_reg <= w_data_i[19];
      mem_274_sv2v_reg <= w_data_i[18];
      mem_273_sv2v_reg <= w_data_i[17];
      mem_272_sv2v_reg <= w_data_i[16];
      mem_271_sv2v_reg <= w_data_i[15];
      mem_270_sv2v_reg <= w_data_i[14];
      mem_269_sv2v_reg <= w_data_i[13];
      mem_268_sv2v_reg <= w_data_i[12];
      mem_267_sv2v_reg <= w_data_i[11];
      mem_266_sv2v_reg <= w_data_i[10];
      mem_265_sv2v_reg <= w_data_i[9];
      mem_264_sv2v_reg <= w_data_i[8];
      mem_263_sv2v_reg <= w_data_i[7];
      mem_262_sv2v_reg <= w_data_i[6];
      mem_261_sv2v_reg <= w_data_i[5];
      mem_260_sv2v_reg <= w_data_i[4];
      mem_259_sv2v_reg <= w_data_i[3];
      mem_258_sv2v_reg <= w_data_i[2];
      mem_257_sv2v_reg <= w_data_i[1];
      mem_256_sv2v_reg <= w_data_i[0];
    end 
    if(N381) begin
      mem_255_sv2v_reg <= w_data_i[31];
      mem_254_sv2v_reg <= w_data_i[30];
      mem_253_sv2v_reg <= w_data_i[29];
      mem_252_sv2v_reg <= w_data_i[28];
      mem_251_sv2v_reg <= w_data_i[27];
      mem_250_sv2v_reg <= w_data_i[26];
      mem_249_sv2v_reg <= w_data_i[25];
      mem_248_sv2v_reg <= w_data_i[24];
      mem_247_sv2v_reg <= w_data_i[23];
      mem_246_sv2v_reg <= w_data_i[22];
      mem_245_sv2v_reg <= w_data_i[21];
      mem_244_sv2v_reg <= w_data_i[20];
      mem_243_sv2v_reg <= w_data_i[19];
      mem_242_sv2v_reg <= w_data_i[18];
      mem_241_sv2v_reg <= w_data_i[17];
      mem_240_sv2v_reg <= w_data_i[16];
      mem_239_sv2v_reg <= w_data_i[15];
      mem_238_sv2v_reg <= w_data_i[14];
      mem_237_sv2v_reg <= w_data_i[13];
      mem_236_sv2v_reg <= w_data_i[12];
      mem_235_sv2v_reg <= w_data_i[11];
      mem_234_sv2v_reg <= w_data_i[10];
      mem_233_sv2v_reg <= w_data_i[9];
      mem_232_sv2v_reg <= w_data_i[8];
      mem_231_sv2v_reg <= w_data_i[7];
      mem_230_sv2v_reg <= w_data_i[6];
      mem_229_sv2v_reg <= w_data_i[5];
      mem_228_sv2v_reg <= w_data_i[4];
      mem_227_sv2v_reg <= w_data_i[3];
      mem_226_sv2v_reg <= w_data_i[2];
      mem_225_sv2v_reg <= w_data_i[1];
      mem_224_sv2v_reg <= w_data_i[0];
    end 
    if(N380) begin
      mem_223_sv2v_reg <= w_data_i[31];
      mem_222_sv2v_reg <= w_data_i[30];
      mem_221_sv2v_reg <= w_data_i[29];
      mem_220_sv2v_reg <= w_data_i[28];
      mem_219_sv2v_reg <= w_data_i[27];
      mem_218_sv2v_reg <= w_data_i[26];
      mem_217_sv2v_reg <= w_data_i[25];
      mem_216_sv2v_reg <= w_data_i[24];
      mem_215_sv2v_reg <= w_data_i[23];
      mem_214_sv2v_reg <= w_data_i[22];
      mem_213_sv2v_reg <= w_data_i[21];
      mem_212_sv2v_reg <= w_data_i[20];
      mem_211_sv2v_reg <= w_data_i[19];
      mem_210_sv2v_reg <= w_data_i[18];
      mem_209_sv2v_reg <= w_data_i[17];
      mem_208_sv2v_reg <= w_data_i[16];
      mem_207_sv2v_reg <= w_data_i[15];
      mem_206_sv2v_reg <= w_data_i[14];
      mem_205_sv2v_reg <= w_data_i[13];
      mem_204_sv2v_reg <= w_data_i[12];
      mem_203_sv2v_reg <= w_data_i[11];
      mem_202_sv2v_reg <= w_data_i[10];
      mem_201_sv2v_reg <= w_data_i[9];
      mem_200_sv2v_reg <= w_data_i[8];
      mem_199_sv2v_reg <= w_data_i[7];
      mem_198_sv2v_reg <= w_data_i[6];
      mem_197_sv2v_reg <= w_data_i[5];
      mem_196_sv2v_reg <= w_data_i[4];
      mem_195_sv2v_reg <= w_data_i[3];
      mem_194_sv2v_reg <= w_data_i[2];
      mem_193_sv2v_reg <= w_data_i[1];
      mem_192_sv2v_reg <= w_data_i[0];
    end 
    if(N379) begin
      mem_191_sv2v_reg <= w_data_i[31];
      mem_190_sv2v_reg <= w_data_i[30];
      mem_189_sv2v_reg <= w_data_i[29];
      mem_188_sv2v_reg <= w_data_i[28];
      mem_187_sv2v_reg <= w_data_i[27];
      mem_186_sv2v_reg <= w_data_i[26];
      mem_185_sv2v_reg <= w_data_i[25];
      mem_184_sv2v_reg <= w_data_i[24];
      mem_183_sv2v_reg <= w_data_i[23];
      mem_182_sv2v_reg <= w_data_i[22];
      mem_181_sv2v_reg <= w_data_i[21];
      mem_180_sv2v_reg <= w_data_i[20];
      mem_179_sv2v_reg <= w_data_i[19];
      mem_178_sv2v_reg <= w_data_i[18];
      mem_177_sv2v_reg <= w_data_i[17];
      mem_176_sv2v_reg <= w_data_i[16];
      mem_175_sv2v_reg <= w_data_i[15];
      mem_174_sv2v_reg <= w_data_i[14];
      mem_173_sv2v_reg <= w_data_i[13];
      mem_172_sv2v_reg <= w_data_i[12];
      mem_171_sv2v_reg <= w_data_i[11];
      mem_170_sv2v_reg <= w_data_i[10];
      mem_169_sv2v_reg <= w_data_i[9];
      mem_168_sv2v_reg <= w_data_i[8];
      mem_167_sv2v_reg <= w_data_i[7];
      mem_166_sv2v_reg <= w_data_i[6];
      mem_165_sv2v_reg <= w_data_i[5];
      mem_164_sv2v_reg <= w_data_i[4];
      mem_163_sv2v_reg <= w_data_i[3];
      mem_162_sv2v_reg <= w_data_i[2];
      mem_161_sv2v_reg <= w_data_i[1];
      mem_160_sv2v_reg <= w_data_i[0];
    end 
    if(N378) begin
      mem_159_sv2v_reg <= w_data_i[31];
      mem_158_sv2v_reg <= w_data_i[30];
      mem_157_sv2v_reg <= w_data_i[29];
      mem_156_sv2v_reg <= w_data_i[28];
      mem_155_sv2v_reg <= w_data_i[27];
      mem_154_sv2v_reg <= w_data_i[26];
      mem_153_sv2v_reg <= w_data_i[25];
      mem_152_sv2v_reg <= w_data_i[24];
      mem_151_sv2v_reg <= w_data_i[23];
      mem_150_sv2v_reg <= w_data_i[22];
      mem_149_sv2v_reg <= w_data_i[21];
      mem_148_sv2v_reg <= w_data_i[20];
      mem_147_sv2v_reg <= w_data_i[19];
      mem_146_sv2v_reg <= w_data_i[18];
      mem_145_sv2v_reg <= w_data_i[17];
      mem_144_sv2v_reg <= w_data_i[16];
      mem_143_sv2v_reg <= w_data_i[15];
      mem_142_sv2v_reg <= w_data_i[14];
      mem_141_sv2v_reg <= w_data_i[13];
      mem_140_sv2v_reg <= w_data_i[12];
      mem_139_sv2v_reg <= w_data_i[11];
      mem_138_sv2v_reg <= w_data_i[10];
      mem_137_sv2v_reg <= w_data_i[9];
      mem_136_sv2v_reg <= w_data_i[8];
      mem_135_sv2v_reg <= w_data_i[7];
      mem_134_sv2v_reg <= w_data_i[6];
      mem_133_sv2v_reg <= w_data_i[5];
      mem_132_sv2v_reg <= w_data_i[4];
      mem_131_sv2v_reg <= w_data_i[3];
      mem_130_sv2v_reg <= w_data_i[2];
      mem_129_sv2v_reg <= w_data_i[1];
      mem_128_sv2v_reg <= w_data_i[0];
    end 
    if(N377) begin
      mem_127_sv2v_reg <= w_data_i[31];
      mem_126_sv2v_reg <= w_data_i[30];
      mem_125_sv2v_reg <= w_data_i[29];
      mem_124_sv2v_reg <= w_data_i[28];
      mem_123_sv2v_reg <= w_data_i[27];
      mem_122_sv2v_reg <= w_data_i[26];
      mem_121_sv2v_reg <= w_data_i[25];
      mem_120_sv2v_reg <= w_data_i[24];
      mem_119_sv2v_reg <= w_data_i[23];
      mem_118_sv2v_reg <= w_data_i[22];
      mem_117_sv2v_reg <= w_data_i[21];
      mem_116_sv2v_reg <= w_data_i[20];
      mem_115_sv2v_reg <= w_data_i[19];
      mem_114_sv2v_reg <= w_data_i[18];
      mem_113_sv2v_reg <= w_data_i[17];
      mem_112_sv2v_reg <= w_data_i[16];
      mem_111_sv2v_reg <= w_data_i[15];
      mem_110_sv2v_reg <= w_data_i[14];
      mem_109_sv2v_reg <= w_data_i[13];
      mem_108_sv2v_reg <= w_data_i[12];
      mem_107_sv2v_reg <= w_data_i[11];
      mem_106_sv2v_reg <= w_data_i[10];
      mem_105_sv2v_reg <= w_data_i[9];
      mem_104_sv2v_reg <= w_data_i[8];
      mem_103_sv2v_reg <= w_data_i[7];
      mem_102_sv2v_reg <= w_data_i[6];
      mem_101_sv2v_reg <= w_data_i[5];
      mem_100_sv2v_reg <= w_data_i[4];
      mem_99_sv2v_reg <= w_data_i[3];
      mem_98_sv2v_reg <= w_data_i[2];
      mem_97_sv2v_reg <= w_data_i[1];
      mem_96_sv2v_reg <= w_data_i[0];
    end 
    if(N376) begin
      mem_95_sv2v_reg <= w_data_i[31];
      mem_94_sv2v_reg <= w_data_i[30];
      mem_93_sv2v_reg <= w_data_i[29];
      mem_92_sv2v_reg <= w_data_i[28];
      mem_91_sv2v_reg <= w_data_i[27];
      mem_90_sv2v_reg <= w_data_i[26];
      mem_89_sv2v_reg <= w_data_i[25];
      mem_88_sv2v_reg <= w_data_i[24];
      mem_87_sv2v_reg <= w_data_i[23];
      mem_86_sv2v_reg <= w_data_i[22];
      mem_85_sv2v_reg <= w_data_i[21];
      mem_84_sv2v_reg <= w_data_i[20];
      mem_83_sv2v_reg <= w_data_i[19];
      mem_82_sv2v_reg <= w_data_i[18];
      mem_81_sv2v_reg <= w_data_i[17];
      mem_80_sv2v_reg <= w_data_i[16];
      mem_79_sv2v_reg <= w_data_i[15];
      mem_78_sv2v_reg <= w_data_i[14];
      mem_77_sv2v_reg <= w_data_i[13];
      mem_76_sv2v_reg <= w_data_i[12];
      mem_75_sv2v_reg <= w_data_i[11];
      mem_74_sv2v_reg <= w_data_i[10];
      mem_73_sv2v_reg <= w_data_i[9];
      mem_72_sv2v_reg <= w_data_i[8];
      mem_71_sv2v_reg <= w_data_i[7];
      mem_70_sv2v_reg <= w_data_i[6];
      mem_69_sv2v_reg <= w_data_i[5];
      mem_68_sv2v_reg <= w_data_i[4];
      mem_67_sv2v_reg <= w_data_i[3];
      mem_66_sv2v_reg <= w_data_i[2];
      mem_65_sv2v_reg <= w_data_i[1];
      mem_64_sv2v_reg <= w_data_i[0];
    end 
    if(N375) begin
      mem_63_sv2v_reg <= w_data_i[31];
      mem_62_sv2v_reg <= w_data_i[30];
      mem_61_sv2v_reg <= w_data_i[29];
      mem_60_sv2v_reg <= w_data_i[28];
      mem_59_sv2v_reg <= w_data_i[27];
      mem_58_sv2v_reg <= w_data_i[26];
      mem_57_sv2v_reg <= w_data_i[25];
      mem_56_sv2v_reg <= w_data_i[24];
      mem_55_sv2v_reg <= w_data_i[23];
      mem_54_sv2v_reg <= w_data_i[22];
      mem_53_sv2v_reg <= w_data_i[21];
      mem_52_sv2v_reg <= w_data_i[20];
      mem_51_sv2v_reg <= w_data_i[19];
      mem_50_sv2v_reg <= w_data_i[18];
      mem_49_sv2v_reg <= w_data_i[17];
      mem_48_sv2v_reg <= w_data_i[16];
      mem_47_sv2v_reg <= w_data_i[15];
      mem_46_sv2v_reg <= w_data_i[14];
      mem_45_sv2v_reg <= w_data_i[13];
      mem_44_sv2v_reg <= w_data_i[12];
      mem_43_sv2v_reg <= w_data_i[11];
      mem_42_sv2v_reg <= w_data_i[10];
      mem_41_sv2v_reg <= w_data_i[9];
      mem_40_sv2v_reg <= w_data_i[8];
      mem_39_sv2v_reg <= w_data_i[7];
      mem_38_sv2v_reg <= w_data_i[6];
      mem_37_sv2v_reg <= w_data_i[5];
      mem_36_sv2v_reg <= w_data_i[4];
      mem_35_sv2v_reg <= w_data_i[3];
      mem_34_sv2v_reg <= w_data_i[2];
      mem_33_sv2v_reg <= w_data_i[1];
      mem_32_sv2v_reg <= w_data_i[0];
    end 
    if(N374) begin
      mem_31_sv2v_reg <= w_data_i[31];
      mem_30_sv2v_reg <= w_data_i[30];
      mem_29_sv2v_reg <= w_data_i[29];
      mem_28_sv2v_reg <= w_data_i[28];
      mem_27_sv2v_reg <= w_data_i[27];
      mem_26_sv2v_reg <= w_data_i[26];
      mem_25_sv2v_reg <= w_data_i[25];
      mem_24_sv2v_reg <= w_data_i[24];
      mem_23_sv2v_reg <= w_data_i[23];
      mem_22_sv2v_reg <= w_data_i[22];
      mem_21_sv2v_reg <= w_data_i[21];
      mem_20_sv2v_reg <= w_data_i[20];
      mem_19_sv2v_reg <= w_data_i[19];
      mem_18_sv2v_reg <= w_data_i[18];
      mem_17_sv2v_reg <= w_data_i[17];
      mem_16_sv2v_reg <= w_data_i[16];
      mem_15_sv2v_reg <= w_data_i[15];
      mem_14_sv2v_reg <= w_data_i[14];
      mem_13_sv2v_reg <= w_data_i[13];
      mem_12_sv2v_reg <= w_data_i[12];
      mem_11_sv2v_reg <= w_data_i[11];
      mem_10_sv2v_reg <= w_data_i[10];
      mem_9_sv2v_reg <= w_data_i[9];
      mem_8_sv2v_reg <= w_data_i[8];
      mem_7_sv2v_reg <= w_data_i[7];
      mem_6_sv2v_reg <= w_data_i[6];
      mem_5_sv2v_reg <= w_data_i[5];
      mem_4_sv2v_reg <= w_data_i[4];
      mem_3_sv2v_reg <= w_data_i[3];
      mem_2_sv2v_reg <= w_data_i[2];
      mem_1_sv2v_reg <= w_data_i[1];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p50_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [31:0] w_data_i;
  input [5:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p50_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p32_els_p50_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2,sv2v_dc_3,sv2v_dc_4,sv2v_dc_5,
  sv2v_dc_6;
  wire [5:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p50
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2, sv2v_dc_3, sv2v_dc_4, sv2v_dc_5, sv2v_dc_6 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p32_els_p50_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p32_els_p50_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p32_els_p50_ready_THEN_valid_p0
  \unhardened.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_channel_narrow_width_in_p32_width_out_p64_lsb_to_msb_p1
(
  clk_i,
  reset_i,
  data_i,
  deque_o,
  data_o,
  deque_i
);

  input [31:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input deque_i;
  output deque_o;
  wire [63:0] data_o;
  wire deque_o,data_o_31_,data_o_30_,data_o_29_,data_o_28_,data_o_27_,data_o_26_,
  data_o_25_,data_o_24_,data_o_23_,data_o_22_,data_o_21_,data_o_20_,data_o_19_,
  data_o_18_,data_o_17_,data_o_16_,data_o_15_,data_o_14_,data_o_13_,data_o_12_,data_o_11_,
  data_o_10_,data_o_9_,data_o_8_,data_o_7_,data_o_6_,data_o_5_,data_o_4_,data_o_3_,
  data_o_2_,data_o_1_,data_o_0_;
  assign data_o[32] = 1'b0;
  assign data_o[33] = 1'b0;
  assign data_o[34] = 1'b0;
  assign data_o[35] = 1'b0;
  assign data_o[36] = 1'b0;
  assign data_o[37] = 1'b0;
  assign data_o[38] = 1'b0;
  assign data_o[39] = 1'b0;
  assign data_o[40] = 1'b0;
  assign data_o[41] = 1'b0;
  assign data_o[42] = 1'b0;
  assign data_o[43] = 1'b0;
  assign data_o[44] = 1'b0;
  assign data_o[45] = 1'b0;
  assign data_o[46] = 1'b0;
  assign data_o[47] = 1'b0;
  assign data_o[48] = 1'b0;
  assign data_o[49] = 1'b0;
  assign data_o[50] = 1'b0;
  assign data_o[51] = 1'b0;
  assign data_o[52] = 1'b0;
  assign data_o[53] = 1'b0;
  assign data_o[54] = 1'b0;
  assign data_o[55] = 1'b0;
  assign data_o[56] = 1'b0;
  assign data_o[57] = 1'b0;
  assign data_o[58] = 1'b0;
  assign data_o[59] = 1'b0;
  assign data_o[60] = 1'b0;
  assign data_o[61] = 1'b0;
  assign data_o[62] = 1'b0;
  assign data_o[63] = 1'b0;
  assign deque_o = deque_i;
  assign data_o_31_ = data_i[31];
  assign data_o[31] = data_o_31_;
  assign data_o_30_ = data_i[30];
  assign data_o[30] = data_o_30_;
  assign data_o_29_ = data_i[29];
  assign data_o[29] = data_o_29_;
  assign data_o_28_ = data_i[28];
  assign data_o[28] = data_o_28_;
  assign data_o_27_ = data_i[27];
  assign data_o[27] = data_o_27_;
  assign data_o_26_ = data_i[26];
  assign data_o[26] = data_o_26_;
  assign data_o_25_ = data_i[25];
  assign data_o[25] = data_o_25_;
  assign data_o_24_ = data_i[24];
  assign data_o[24] = data_o_24_;
  assign data_o_23_ = data_i[23];
  assign data_o[23] = data_o_23_;
  assign data_o_22_ = data_i[22];
  assign data_o[22] = data_o_22_;
  assign data_o_21_ = data_i[21];
  assign data_o[21] = data_o_21_;
  assign data_o_20_ = data_i[20];
  assign data_o[20] = data_o_20_;
  assign data_o_19_ = data_i[19];
  assign data_o[19] = data_o_19_;
  assign data_o_18_ = data_i[18];
  assign data_o[18] = data_o_18_;
  assign data_o_17_ = data_i[17];
  assign data_o[17] = data_o_17_;
  assign data_o_16_ = data_i[16];
  assign data_o[16] = data_o_16_;
  assign data_o_15_ = data_i[15];
  assign data_o[15] = data_o_15_;
  assign data_o_14_ = data_i[14];
  assign data_o[14] = data_o_14_;
  assign data_o_13_ = data_i[13];
  assign data_o[13] = data_o_13_;
  assign data_o_12_ = data_i[12];
  assign data_o[12] = data_o_12_;
  assign data_o_11_ = data_i[11];
  assign data_o[11] = data_o_11_;
  assign data_o_10_ = data_i[10];
  assign data_o[10] = data_o_10_;
  assign data_o_9_ = data_i[9];
  assign data_o[9] = data_o_9_;
  assign data_o_8_ = data_i[8];
  assign data_o[8] = data_o_8_;
  assign data_o_7_ = data_i[7];
  assign data_o[7] = data_o_7_;
  assign data_o_6_ = data_i[6];
  assign data_o[6] = data_o_6_;
  assign data_o_5_ = data_i[5];
  assign data_o[5] = data_o_5_;
  assign data_o_4_ = data_i[4];
  assign data_o[4] = data_o_4_;
  assign data_o_3_ = data_i[3];
  assign data_o[3] = data_o_3_;
  assign data_o_2_ = data_i[2];
  assign data_o[2] = data_o_2_;
  assign data_o_1_ = data_i[1];
  assign data_o[1] = data_o_1_;
  assign data_o_0_ = data_i[0];
  assign data_o[0] = data_o_0_;

endmodule



module bsg_fifo_1r1w_narrowed
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [63:0] data_o;
  wire ready_o,v_o,yumi;
  wire [31:0] data;

  bsg_fifo_1r1w_small_width_p32_els_p50_ready_THEN_valid_p0
  main_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data),
    .yumi_i(yumi)
  );


  bsg_channel_narrow_width_in_p32_width_out_p64_lsb_to_msb_p1
  output_narrower
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data),
    .deque_o(yumi),
    .data_o(data_o),
    .deque_i(yumi_i)
  );


endmodule

