

module top
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  yumi_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [69:0] cache_pkt_i;
  output [31:0] data_o;
  output [32:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output yumi_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;

  bsg_cache
  wrapper
  (
    .cache_pkt_i(cache_pkt_i),
    .data_o(data_o),
    .dma_pkt_o(dma_pkt_o),
    .dma_data_i(dma_data_i),
    .dma_data_o(dma_data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_yumi_i(dma_data_yumi_i),
    .yumi_o(yumi_o),
    .v_o(v_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_v_o(dma_data_v_o),
    .v_we_o(v_we_o)
  );


endmodule



module bsg_cache_decode
(
  opcode_i,
  decode_o
);

  input [5:0] opcode_i;
  output [20:0] decode_o;
  wire [20:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N146,N147,N148,N150,N152,
  N153,N154,N155,N156,N158,N160,N161,N163,N165,N166,N167,N168,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297;
  assign N17 = N80 | N138;
  assign N18 = opcode_i[3] | opcode_i[2];
  assign N19 = opcode_i[1] | opcode_i[0];
  assign N20 = N17 | N18;
  assign N21 = N20 | N19;
  assign N22 = opcode_i[1] | N139;
  assign N23 = N20 | N22;
  assign N24 = N146 | N139;
  assign N25 = N20 | N24;
  assign N26 = opcode_i[3] | N165;
  assign N27 = N17 | N26;
  assign N28 = N27 | N19;
  assign N29 = N146 | opcode_i[0];
  assign N30 = N20 | N29;
  assign N31 = N27 | N22;
  assign N32 = N27 | N29;
  assign N33 = N27 | N24;
  assign N34 = N152 | opcode_i[2];
  assign N35 = N17 | N34;
  assign N36 = N35 | N19;
  assign N37 = opcode_i[5] | opcode_i[4];
  assign N38 = N37 | N18;
  assign N39 = N38 | N24;
  assign N40 = N37 | N34;
  assign N41 = N40 | N24;
  assign N42 = N37 | N26;
  assign N43 = N42 | N24;
  assign N45 = N80 | opcode_i[4];
  assign N46 = N45 | N18;
  assign N47 = N46 | N19;
  assign N48 = N46 | N22;
  assign N49 = N46 | N24;
  assign N50 = N45 | N26;
  assign N51 = N50 | N19;
  assign N52 = N46 | N29;
  assign N53 = N50 | N22;
  assign N54 = N50 | N29;
  assign N55 = N50 | N24;
  assign N56 = N45 | N34;
  assign N57 = N56 | N19;
  assign N58 = N38 | N29;
  assign N59 = N40 | N29;
  assign N60 = N42 | N29;
  assign N62 = N38 | N22;
  assign N63 = N40 | N22;
  assign N64 = N42 | N22;
  assign N66 = N80 & N138;
  assign N67 = N152 & N165;
  assign N68 = N146 & N139;
  assign N69 = N66 & N67;
  assign N70 = N69 & N68;
  assign N71 = N40 | N19;
  assign N72 = N42 | N19;
  assign N74 = opcode_i[5] & opcode_i[3];
  assign N75 = N74 & opcode_i[0];
  assign N76 = N74 & opcode_i[1];
  assign N77 = opcode_i[3] & opcode_i[2];
  assign N78 = N80 & opcode_i[4];
  assign N81 = N138 & N152;
  assign N82 = N165 & N146;
  assign N83 = N81 & N82;
  assign N84 = N83 & N139;
  assign N85 = N138 | opcode_i[3];
  assign N86 = opcode_i[2] | opcode_i[1];
  assign N87 = N85 | N86;
  assign N88 = N87 | opcode_i[0];
  assign N90 = opcode_i[4] | opcode_i[3];
  assign N91 = N90 | N86;
  assign N92 = N91 | N139;
  assign N93 = N87 | N139;
  assign N95 = opcode_i[2] | N146;
  assign N96 = N90 | N95;
  assign N97 = N96 | opcode_i[0];
  assign N98 = N85 | N95;
  assign N99 = N98 | opcode_i[0];
  assign N101 = N96 | N139;
  assign N102 = N98 | N139;
  assign N104 = N165 | opcode_i[1];
  assign N105 = N90 | N104;
  assign N106 = N105 | opcode_i[0];
  assign N107 = N85 | N104;
  assign N108 = N107 | opcode_i[0];
  assign N110 = N105 | N139;
  assign N111 = N107 | N139;
  assign N113 = N165 | N146;
  assign N114 = N90 | N113;
  assign N115 = N114 | opcode_i[0];
  assign N116 = N85 | N113;
  assign N117 = N116 | opcode_i[0];
  assign N119 = N114 | N139;
  assign N120 = N116 | N139;
  assign N122 = opcode_i[4] | N152;
  assign N123 = N122 | N86;
  assign N124 = N123 | opcode_i[0];
  assign N125 = N138 | N152;
  assign N126 = N125 | N86;
  assign N127 = N126 | opcode_i[0];
  assign N129 = opcode_i[3] & opcode_i[0];
  assign N130 = opcode_i[3] & opcode_i[1];
  assign N138 = ~opcode_i[4];
  assign N139 = ~opcode_i[0];
  assign N140 = N138 | opcode_i[5];
  assign N141 = opcode_i[3] | N140;
  assign N142 = opcode_i[2] | N141;
  assign N143 = opcode_i[1] | N142;
  assign N144 = N139 | N143;
  assign decode_o[13] = ~N144;
  assign N146 = ~opcode_i[1];
  assign N147 = N146 | N142;
  assign N148 = opcode_i[0] | N147;
  assign decode_o[12] = ~N148;
  assign N150 = N139 | N147;
  assign decode_o[11] = ~N150;
  assign N152 = ~opcode_i[3];
  assign N153 = N152 | N140;
  assign N154 = opcode_i[2] | N153;
  assign N155 = opcode_i[1] | N154;
  assign N156 = opcode_i[0] | N155;
  assign decode_o[10] = ~N156;
  assign N158 = N139 | N155;
  assign decode_o[9] = ~N158;
  assign N160 = N146 | N154;
  assign N161 = opcode_i[0] | N160;
  assign decode_o[8] = ~N161;
  assign N163 = N139 | N160;
  assign decode_o[7] = ~N163;
  assign N165 = ~opcode_i[2];
  assign N166 = N165 | N153;
  assign N167 = opcode_i[1] | N166;
  assign N168 = opcode_i[0] | N167;
  assign decode_o[6] = ~N168;
  assign N170 = opcode_i[4] | opcode_i[5];
  assign N171 = opcode_i[3] | N170;
  assign N172 = opcode_i[2] | N171;
  assign N173 = opcode_i[1] | N172;
  assign N174 = opcode_i[0] | N173;
  assign N175 = ~N174;
  assign N176 = N139 | N173;
  assign N177 = ~N176;
  assign N178 = N146 | N172;
  assign N179 = opcode_i[0] | N178;
  assign N180 = ~N179;
  assign N181 = N139 | N178;
  assign N182 = ~N181;
  assign N183 = N152 | N170;
  assign N184 = N165 | N183;
  assign N185 = opcode_i[1] | N184;
  assign N186 = opcode_i[0] | N185;
  assign N187 = ~N186;
  assign N188 = N139 | N185;
  assign N189 = ~N188;
  assign N190 = N165 | N171;
  assign N191 = opcode_i[1] | N190;
  assign N192 = opcode_i[0] | N191;
  assign N193 = ~N192;
  assign N194 = N139 | N191;
  assign N195 = ~N194;
  assign N196 = N146 | N190;
  assign N197 = opcode_i[0] | N196;
  assign N198 = ~N197;
  assign N199 = N139 | N196;
  assign N200 = ~N199;
  assign N201 = opcode_i[2] | N183;
  assign N202 = opcode_i[1] | N201;
  assign N203 = opcode_i[0] | N202;
  assign N204 = ~N203;
  assign N205 = N139 | N202;
  assign N206 = ~N205;
  assign N207 = N146 | N201;
  assign N208 = opcode_i[0] | N207;
  assign N209 = ~N208;
  assign N210 = N139 | N207;
  assign N211 = ~N210;
  assign N212 = opcode_i[0] | N143;
  assign decode_o[14] = ~N212;
  assign decode_o[20:19] = (N0)? { 1'b1, 1'b1 } : 
                           (N1)? { 1'b1, 1'b0 } : 
                           (N2)? { 1'b0, 1'b1 } : 
                           (N3)? { 1'b0, 1'b0 } : 
                           (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N44;
  assign N1 = N61;
  assign N2 = N65;
  assign N3 = N73;
  assign N4 = N79;
  assign { N135, N134, N133, N132 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N6)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N7)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N8)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N9)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N10)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N11)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N12)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N13)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N14)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N89;
  assign N6 = N94;
  assign N7 = N100;
  assign N8 = N103;
  assign N9 = N109;
  assign N10 = N112;
  assign N11 = N118;
  assign N12 = N121;
  assign N13 = N128;
  assign N14 = N131;
  assign decode_o[4:0] = (N15)? { N137, N135, N134, N133, N132 } : 
                         (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = opcode_i[5];
  assign N16 = N80;
  assign N44 = N234 | N235;
  assign N234 = N232 | N233;
  assign N232 = N230 | N231;
  assign N230 = N228 | N229;
  assign N228 = N226 | N227;
  assign N226 = N224 | N225;
  assign N224 = N222 | N223;
  assign N222 = N220 | N221;
  assign N220 = N218 | N219;
  assign N218 = N216 | N217;
  assign N216 = N214 | N215;
  assign N214 = ~N21;
  assign N215 = ~N23;
  assign N217 = ~N25;
  assign N219 = ~N28;
  assign N221 = ~N30;
  assign N223 = ~N31;
  assign N225 = ~N32;
  assign N227 = ~N33;
  assign N229 = ~N36;
  assign N231 = ~N39;
  assign N233 = ~N41;
  assign N235 = ~N43;
  assign N61 = N256 | N257;
  assign N256 = N254 | N255;
  assign N254 = N252 | N253;
  assign N252 = N250 | N251;
  assign N250 = N248 | N249;
  assign N248 = N246 | N247;
  assign N246 = N244 | N245;
  assign N244 = N242 | N243;
  assign N242 = N240 | N241;
  assign N240 = N238 | N239;
  assign N238 = N236 | N237;
  assign N236 = ~N47;
  assign N237 = ~N48;
  assign N239 = ~N49;
  assign N241 = ~N51;
  assign N243 = ~N52;
  assign N245 = ~N53;
  assign N247 = ~N54;
  assign N249 = ~N55;
  assign N251 = ~N57;
  assign N253 = ~N58;
  assign N255 = ~N59;
  assign N257 = ~N60;
  assign N65 = N260 | N261;
  assign N260 = N258 | N259;
  assign N258 = ~N62;
  assign N259 = ~N63;
  assign N261 = ~N64;
  assign N73 = N263 | N264;
  assign N263 = N70 | N262;
  assign N262 = ~N71;
  assign N264 = ~N72;
  assign N79 = N75 | N266;
  assign N266 = N76 | N265;
  assign N265 = N77 | N78;
  assign decode_o[17] = N187 | N189;
  assign decode_o[18] = N269 | decode_o[4];
  assign N269 = N268 | N182;
  assign N268 = N267 | N180;
  assign N267 = N175 | N177;
  assign decode_o[16] = N276 | N187;
  assign N276 = N275 | N200;
  assign N275 = N274 | N198;
  assign N274 = N273 | N195;
  assign N273 = N272 | N193;
  assign N272 = N271 | N182;
  assign N271 = N270 | N180;
  assign N270 = N175 | N177;
  assign decode_o[15] = N279 | N189;
  assign N279 = N278 | N211;
  assign N278 = N277 | N209;
  assign N277 = N204 | N206;
  assign decode_o[5] = ~decode_o[14];
  assign N80 = ~opcode_i[5];
  assign N89 = N84 | N280;
  assign N280 = ~N88;
  assign N94 = N281 | N282;
  assign N281 = ~N92;
  assign N282 = ~N93;
  assign N100 = N283 | N284;
  assign N283 = ~N97;
  assign N284 = ~N99;
  assign N103 = N285 | N286;
  assign N285 = ~N101;
  assign N286 = ~N102;
  assign N109 = N287 | N288;
  assign N287 = ~N106;
  assign N288 = ~N108;
  assign N112 = N289 | N290;
  assign N289 = ~N110;
  assign N290 = ~N111;
  assign N118 = N291 | N292;
  assign N291 = ~N115;
  assign N292 = ~N117;
  assign N121 = N293 | N294;
  assign N293 = ~N119;
  assign N294 = ~N120;
  assign N128 = N295 | N296;
  assign N295 = ~N124;
  assign N296 = ~N127;
  assign N131 = N129 | N297;
  assign N297 = N130 | N77;
  assign N136 = ~N131;
  assign N137 = N136;

endmodule



module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p80_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [79:0] data_i;
  output [79:0] data_o;
  input clk_i;
  input en_i;
  wire [79:0] data_o;
  reg data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_79_sv2v_reg <= data_i[79];
      data_o_78_sv2v_reg <= data_i[78];
      data_o_77_sv2v_reg <= data_i[77];
      data_o_76_sv2v_reg <= data_i[76];
      data_o_75_sv2v_reg <= data_i[75];
      data_o_74_sv2v_reg <= data_i[74];
      data_o_73_sv2v_reg <= data_i[73];
      data_o_72_sv2v_reg <= data_i[72];
      data_o_71_sv2v_reg <= data_i[71];
      data_o_70_sv2v_reg <= data_i[70];
      data_o_69_sv2v_reg <= data_i[69];
      data_o_68_sv2v_reg <= data_i[68];
      data_o_67_sv2v_reg <= data_i[67];
      data_o_66_sv2v_reg <= data_i[66];
      data_o_65_sv2v_reg <= data_i[65];
      data_o_64_sv2v_reg <= data_i[64];
      data_o_63_sv2v_reg <= data_i[63];
      data_o_62_sv2v_reg <= data_i[62];
      data_o_61_sv2v_reg <= data_i[61];
      data_o_60_sv2v_reg <= data_i[60];
      data_o_59_sv2v_reg <= data_i[59];
      data_o_58_sv2v_reg <= data_i[58];
      data_o_57_sv2v_reg <= data_i[57];
      data_o_56_sv2v_reg <= data_i[56];
      data_o_55_sv2v_reg <= data_i[55];
      data_o_54_sv2v_reg <= data_i[54];
      data_o_53_sv2v_reg <= data_i[53];
      data_o_52_sv2v_reg <= data_i[52];
      data_o_51_sv2v_reg <= data_i[51];
      data_o_50_sv2v_reg <= data_i[50];
      data_o_49_sv2v_reg <= data_i[49];
      data_o_48_sv2v_reg <= data_i[48];
      data_o_47_sv2v_reg <= data_i[47];
      data_o_46_sv2v_reg <= data_i[46];
      data_o_45_sv2v_reg <= data_i[45];
      data_o_44_sv2v_reg <= data_i[44];
      data_o_43_sv2v_reg <= data_i[43];
      data_o_42_sv2v_reg <= data_i[42];
      data_o_41_sv2v_reg <= data_i[41];
      data_o_40_sv2v_reg <= data_i[40];
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p80
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [79:0] data_i;
  output [79:0] data_o;
  input clk_i;
  input en_i;
  wire [79:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p80_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p80_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [79:0] data_i;
  input [5:0] addr_i;
  input [79:0] w_mask_i;
  output [79:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [79:0] data_o,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,\nz.read_en ,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  \nz.llr.read_en_r ,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,
  N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,
  N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,
  N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,
  N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,
  N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,
  N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,
  N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
  N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,
  N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,
  N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
  N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,
  N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,
  N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
  N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,
  N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,
  N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
  N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,
  N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,
  N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
  N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,
  N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,
  N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
  N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,
  N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,
  N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
  N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,
  N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,
  N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
  N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,
  N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,
  N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
  N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,
  N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,
  N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
  N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,
  N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,
  N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
  N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,
  N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,
  N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
  N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,
  N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,
  N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
  N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,
  N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,
  N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
  N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,
  N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,
  N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
  N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,
  N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,
  N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
  N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,
  N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,
  N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
  N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,
  N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,
  N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
  N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,
  N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,
  N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
  N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,
  N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,
  N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
  N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,
  N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,
  N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
  N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,
  N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,
  N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
  N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,
  N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,
  N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
  N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,
  N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,
  N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
  N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,
  N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,
  N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
  N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,
  N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,
  N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
  N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,
  N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,
  N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
  N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,
  N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,
  N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
  N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,
  N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,
  N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
  N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
  N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,
  N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
  N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,
  N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,
  N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
  N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,
  N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,
  N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
  N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,
  N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,
  N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
  N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,
  N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,
  N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
  N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,
  N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,
  N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
  N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,
  N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,
  N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
  N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,
  N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,
  N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
  N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,
  N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,
  N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
  N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,
  N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,
  N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
  N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,
  N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,
  N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
  N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,
  N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,
  N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
  N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,
  N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,
  N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
  N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,
  N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,
  N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
  N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,
  N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,
  N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
  N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,
  N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,
  N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
  N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,
  N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,
  N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
  N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,
  N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,
  N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
  N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,
  N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,
  N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
  N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,
  N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
  N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
  N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,
  N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,
  N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
  N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,
  N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,
  N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
  N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,
  N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,
  N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
  N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,
  N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,
  N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
  N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,
  N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,
  N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
  N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,
  N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,
  N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
  N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,
  N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,
  N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
  N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,
  N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,
  N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
  N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,
  N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,
  N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
  N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,
  N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,
  N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
  N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,
  N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,
  N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
  N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,
  N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,
  N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
  N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,
  N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,
  N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
  N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,
  N4193,N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,
  N4206,N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,
  N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,
  N4233,N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,
  N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,
  N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,
  N4273,N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,
  N4286,N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,
  N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,
  N4313,N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,
  N4326,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,
  N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,
  N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,
  N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,
  N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,
  N4393,N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,
  N4406,N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,
  N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,
  N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,
  N4446,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,
  N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,
  N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,
  N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,
  N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,
  N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,
  N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,
  N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,
  N4553,N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,
  N4566,N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,
  N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,
  N4593,N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,
  N4606,N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,
  N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,
  N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,
  N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,
  N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,
  N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,
  N4686,N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,
  N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,
  N4713,N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,
  N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,
  N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,
  N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,
  N4766,N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,
  N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,
  N4793,N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,
  N4806,N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,
  N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,
  N4833,N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,
  N4846,N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,
  N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,
  N4873,N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,
  N4886,N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,
  N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,
  N4913,N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,
  N4926,N4927,N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,
  N4939,N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,
  N4953,N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,
  N4966,N4967,N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,
  N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,
  N4993,N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,
  N5006,N5007,N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,
  N5019,N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,
  N5033,N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,
  N5046,N5047,N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,
  N5059,N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,
  N5073,N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,
  N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,
  N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,
  N5113,N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,
  N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,
  N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,
  N5153,N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,
  N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,
  N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,
  N5193,N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,
  N5206,N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,
  N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,
  N5233,N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,
  N5246,N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,
  N5259,N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,
  N5273,N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,
  N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,
  N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,
  N5313,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,
  N5326,N5327,N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,
  N5339,N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,
  N5353,N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,
  N5366,N5367,N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,
  N5379,N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,
  N5393,N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,
  N5406,N5407,N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,
  N5419,N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,
  N5433,N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,
  N5446,N5447,N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,
  N5459,N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,
  N5473,N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,
  N5486,N5487,N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,
  N5499,N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,
  N5513,N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,
  N5526,N5527,N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,
  N5539,N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,
  N5553,N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,
  N5566,N5567,N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,
  N5579,N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,
  N5593,N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,
  N5606,N5607,N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,
  N5619,N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,
  N5633,N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,
  N5646,N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,
  N5659,N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,
  N5673,N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,
  N5686,N5687,N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,
  N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,
  N5713,N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,
  N5726,N5727,N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,
  N5739,N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,
  N5753,N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,
  N5766,N5767,N5768,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,
  N5779,N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,
  N5793,N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,
  N5806,N5807,N5808,N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,
  N5819,N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,
  N5833,N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,
  N5846,N5847,N5848,N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,
  N5859,N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,
  N5873,N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,
  N5886,N5887,N5888,N5889,N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,
  N5899,N5900,N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,
  N5913,N5914,N5915,N5916,N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,
  N5926,N5927,N5928,N5929,N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,
  N5939,N5940,N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,
  N5953,N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,
  N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,
  N5979,N5980,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,
  N5993,N5994,N5995,N5996,N5997,N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,
  N6006,N6007,N6008,N6009,N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,
  N6019,N6020,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,
  N6033,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,
  N6046,N6047,N6048,N6049,N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,
  N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,
  N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,
  N6086,N6087,N6088,N6089,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,
  N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,
  N6113,N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,
  N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,
  N6139,N6140,N6141,N6142,N6143,N6144,N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,
  N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,
  N6166,N6167,N6168,N6169,N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,
  N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,
  N6193,N6194,N6195,N6196,N6197,N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,
  N6206,N6207,N6208,N6209,N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,
  N6219,N6220,N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,
  N6233,N6234,N6235,N6236,N6237,N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,
  N6246,N6247,N6248,N6249,N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,
  N6259,N6260,N6261,N6262,N6263,N6264,N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,
  N6273,N6274,N6275,N6276,N6277,N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,
  N6286,N6287,N6288,N6289,N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,
  N6299,N6300,N6301,N6302,N6303,N6304,N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,
  N6313,N6314,N6315,N6316,N6317,N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,
  N6326,N6327,N6328,N6329,N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,
  N6339,N6340,N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,
  N6353,N6354,N6355,N6356,N6357,N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,
  N6366,N6367,N6368,N6369,N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,
  N6379,N6380,N6381,N6382,N6383,N6384,N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,
  N6393,N6394,N6395,N6396,N6397,N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,
  N6406,N6407,N6408,N6409,N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,
  N6419,N6420,N6421,N6422,N6423,N6424,N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,
  N6433,N6434,N6435,N6436,N6437,N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,
  N6446,N6447,N6448,N6449,N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,
  N6459,N6460,N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,
  N6473,N6474,N6475,N6476,N6477,N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,
  N6486,N6487,N6488,N6489,N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,
  N6499,N6500,N6501,N6502,N6503,N6504,N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,
  N6513,N6514,N6515,N6516,N6517,N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,
  N6526,N6527,N6528,N6529,N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,
  N6539,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,
  N6553,N6554,N6555,N6556,N6557,N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,
  N6566,N6567,N6568,N6569,N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,
  N6579,N6580,N6581,N6582,N6583,N6584,N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,
  N6593,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,
  N6606,N6607,N6608,N6609,N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,
  N6619,N6620,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,
  N6633,N6634,N6635,N6636,N6637,N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,
  N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,
  N6659,N6660,N6661,N6662,N6663,N6664,N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,
  N6673,N6674,N6675,N6676,N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,
  N6686,N6687,N6688,N6689,N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,
  N6699,N6700,N6701,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,
  N6713,N6714,N6715,N6716,N6717,N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,
  N6726,N6727,N6728,N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,
  N6739,N6740,N6741,N6742,N6743,N6744,N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,
  N6753,N6754,N6755,N6756,N6757,N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,
  N6766,N6767,N6768,N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,
  N6779,N6780,N6781,N6782,N6783,N6784,N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,
  N6793,N6794,N6795,N6796,N6797,N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,
  N6806,N6807,N6808,N6809,N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,
  N6819,N6820,N6821,N6822,N6823,N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,
  N6833,N6834,N6835,N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,
  N6846,N6847,N6848,N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,
  N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,
  N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,
  N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,
  N6899,N6900,N6901,N6902,N6903,N6904,N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,
  N6913,N6914,N6915,N6916,N6917,N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,
  N6926,N6927,N6928,N6929,N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,
  N6939,N6940,N6941,N6942,N6943,N6944,N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,
  N6953,N6954,N6955,N6956,N6957,N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,
  N6966,N6967,N6968,N6969,N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,
  N6979,N6980,N6981,N6982,N6983,N6984,N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,
  N6993,N6994,N6995,N6996,N6997,N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,
  N7006,N7007,N7008,N7009,N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,
  N7019,N7020,N7021,N7022,N7023,N7024,N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,
  N7033,N7034,N7035,N7036,N7037,N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,
  N7046,N7047,N7048,N7049,N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,
  N7059,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,
  N7073,N7074,N7075,N7076,N7077,N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,
  N7086,N7087,N7088,N7089,N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,
  N7099,N7100,N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,
  N7113,N7114,N7115,N7116,N7117,N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,
  N7126,N7127,N7128,N7129,N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,
  N7139,N7140,N7141,N7142,N7143,N7144,N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,
  N7153,N7154,N7155,N7156,N7157,N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,
  N7166,N7167,N7168,N7169,N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,
  N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,N7189,N7190,N7191,N7192,
  N7193,N7194,N7195,N7196,N7197,N7198,N7199,N7200,N7201,N7202,N7203,N7204,N7205,
  N7206,N7207,N7208,N7209,N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,
  N7219,N7220,N7221,N7222,N7223,N7224,N7225,N7226,N7227,N7228,N7229,N7230,N7231,N7232,
  N7233,N7234,N7235,N7236,N7237,N7238,N7239,N7240,N7241,N7242,N7243,N7244,N7245,
  N7246,N7247,N7248,N7249,N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,
  N7259,N7260,N7261,N7262,N7263,N7264,N7265,N7266,N7267,N7268,N7269,N7270,N7271,N7272,
  N7273,N7274,N7275,N7276,N7277,N7278,N7279,N7280,N7281,N7282,N7283,N7284,N7285,
  N7286,N7287,N7288,N7289,N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,
  N7299,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307,N7308,N7309,N7310,N7311,N7312,
  N7313,N7314,N7315,N7316,N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7324,N7325,
  N7326,N7327,N7328,N7329,N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,
  N7339,N7340,N7341,N7342,N7343,N7344,N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352,
  N7353,N7354,N7355,N7356,N7357,N7358,N7359,N7360,N7361,N7362,N7363,N7364,N7365,
  N7366,N7367,N7368,N7369,N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,
  N7379,N7380,N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388,N7389,N7390,N7391,N7392,
  N7393,N7394,N7395,N7396,N7397,N7398,N7399,N7400,N7401,N7402,N7403,N7404,N7405,
  N7406,N7407,N7408,N7409,N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,
  N7419,N7420,N7421,N7422,N7423,N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7432,
  N7433,N7434,N7435,N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,
  N7446,N7447,N7448,N7449,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,
  N7459,N7460,N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,
  N7473,N7474,N7475,N7476,N7477,N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,
  N7486,N7487,N7488,N7489,N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,
  N7499,N7500,N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,
  N7513,N7514,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,
  N7526,N7527,N7528,N7529,N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,
  N7539,N7540,N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,
  N7553,N7554,N7555,N7556,N7557,N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,
  N7566,N7567,N7568,N7569,N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,
  N7579,N7580,N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,
  N7593,N7594,N7595,N7596,N7597,N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,
  N7606,N7607,N7608,N7609,N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,
  N7619,N7620,N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,
  N7633,N7634,N7635,N7636,N7637,N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,
  N7646,N7647,N7648,N7649,N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,
  N7659,N7660,N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,
  N7673,N7674,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,
  N7686,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,
  N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,
  N7713,N7714,N7715,N7716,N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,
  N7726,N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,
  N7739,N7740,N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,
  N7753,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,
  N7766,N7767,N7768,N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,
  N7779,N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,
  N7793,N7794,N7795,N7796,N7797,N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,
  N7806,N7807,N7808,N7809,N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,
  N7819,N7820,N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,
  N7833,N7834,N7835,N7836,N7837,N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,
  N7846,N7847,N7848,N7849,N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,
  N7859,N7860,N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,
  N7873,N7874,N7875,N7876,N7877,N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,
  N7886,N7887,N7888,N7889,N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,
  N7899,N7900,N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,
  N7913,N7914,N7915,N7916,N7917,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,
  N7926,N7927,N7928,N7929,N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,
  N7939,N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,N7949,N7950,N7951,N7952,
  N7953,N7954,N7955,N7956,N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7964,N7965,
  N7966,N7967,N7968,N7969,N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,
  N7979,N7980,N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,N7989,N7990,N7991,N7992,
  N7993,N7994,N7995,N7996,N7997,N7998,N7999,N8000,N8001,N8002,N8003,N8004,N8005,
  N8006,N8007,N8008,N8009,N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,
  N8019,N8020,N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,N8029,N8030,N8031,N8032,
  N8033,N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,
  N8046,N8047,N8048,N8049,N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,
  N8059,N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,N8069,N8070,N8071,N8072,
  N8073,N8074,N8075,N8076,N8077,N8078,N8079,N8080,N8081,N8082,N8083,N8084,N8085,
  N8086,N8087,N8088,N8089,N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,
  N8099,N8100,N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111,N8112,
  N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,N8121,N8122,N8123,N8124,N8125,
  N8126,N8127,N8128,N8129,N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,
  N8139,N8140,N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,N8149,N8150,N8151,N8152,
  N8153,N8154,N8155,N8156,N8157,N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165,
  N8166,N8167,N8168,N8169,N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,
  N8179,N8180,N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,N8189,N8190,N8191,N8192,
  N8193,N8194,N8195,N8196,N8197,N8198,N8199,N8200,N8201,N8202,N8203,N8204,N8205,
  N8206,N8207,N8208,N8209,N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,
  N8219,N8220,N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,N8229,N8230,N8231,N8232,
  N8233,N8234,N8235,N8236,N8237,N8238,N8239,N8240,N8241,N8242,N8243,N8244,N8245,
  N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,
  N8259,N8260,N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,N8269,N8270,N8271,N8272,
  N8273,N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,
  N8286,N8287,N8288,N8289,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,
  N8299,N8300,N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,N8309,N8310,N8311,N8312,
  N8313,N8314,N8315,N8316,N8317,N8318,N8319,N8320,N8321,N8322,N8323,N8324,N8325,
  N8326,N8327,N8328,N8329,N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,
  N8339,N8340,N8341,N8342,N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,
  N8353,N8354,N8355,N8356,N8357,N8358,N8359,N8360,N8361,N8362,N8363,N8364,N8365,
  N8366,N8367,N8368,N8369,N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,
  N8379,N8380,N8381,N8382,N8383,N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,
  N8393,N8394,N8395,N8396,N8397,N8398,N8399,N8400,N8401,N8402,N8403,N8404,N8405,
  N8406,N8407,N8408,N8409,N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,
  N8419,N8420,N8421,N8422,N8423,N8424,N8425,N8426,N8427,N8428,N8429,N8430,N8431,N8432,
  N8433,N8434,N8435,N8436,N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445,
  N8446,N8447,N8448,N8449,N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,
  N8459,N8460,N8461,N8462,N8463,N8464,N8465,N8466,N8467,N8468,N8469,N8470,N8471,N8472,
  N8473,N8474,N8475,N8476,N8477,N8478,N8479,N8480,N8481,N8482,N8483,N8484,N8485,
  N8486,N8487,N8488,N8489,N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,
  N8499,N8500,N8501,N8502,N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,
  N8513,N8514,N8515,N8516,N8517,N8518,N8519,N8520,N8521,N8522,N8523,N8524,N8525,
  N8526,N8527,N8528,N8529,N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,
  N8539,N8540,N8541,N8542,N8543,N8544,N8545,N8546,N8547,N8548,N8549,N8550,N8551,N8552,
  N8553,N8554,N8555,N8556,N8557,N8558,N8559,N8560,N8561,N8562,N8563,N8564,N8565,
  N8566,N8567,N8568,N8569,N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,
  N8579,N8580,N8581,N8582,N8583,N8584,N8585,N8586,N8587,N8588,N8589,N8590,N8591,N8592,
  N8593,N8594,N8595,N8596,N8597,N8598,N8599,N8600,N8601,N8602,N8603,N8604,N8605,
  N8606,N8607,N8608,N8609,N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,
  N8619,N8620,N8621,N8622,N8623,N8624,N8625,N8626,N8627,N8628,N8629,N8630,N8631,N8632,
  N8633,N8634,N8635,N8636,N8637,N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645,
  N8646,N8647,N8648,N8649,N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,
  N8659,N8660,N8661,N8662,N8663,N8664,N8665,N8666,N8667,N8668,N8669,N8670,N8671,N8672,
  N8673,N8674,N8675,N8676,N8677,N8678,N8679,N8680,N8681,N8682,N8683,N8684,N8685,
  N8686,N8687,N8688,N8689,N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,
  N8699,N8700,N8701,N8702,N8703,N8704,N8705,N8706,N8707,N8708,N8709,N8710,N8711,N8712,
  N8713,N8714,N8715,N8716,N8717,N8718,N8719,N8720,N8721,N8722,N8723,N8724,N8725,
  N8726,N8727,N8728,N8729,N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,
  N8739,N8740,N8741,N8742,N8743,N8744,N8745,N8746,N8747,N8748,N8749,N8750,N8751,N8752,
  N8753,N8754,N8755,N8756,N8757,N8758,N8759,N8760,N8761,N8762,N8763,N8764,N8765,
  N8766,N8767,N8768,N8769,N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,
  N8779,N8780,N8781,N8782,N8783,N8784,N8785,N8786,N8787,N8788,N8789,N8790,N8791,N8792,
  N8793,N8794,N8795,N8796,N8797,N8798,N8799,N8800,N8801,N8802,N8803,N8804,N8805,
  N8806,N8807,N8808,N8809,N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,
  N8819,N8820,N8821,N8822,N8823,N8824,N8825,N8826,N8827,N8828,N8829,N8830,N8831,N8832,
  N8833,N8834,N8835,N8836,N8837,N8838,N8839,N8840,N8841,N8842,N8843,N8844,N8845,
  N8846,N8847,N8848,N8849,N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,
  N8859,N8860,N8861,N8862,N8863,N8864,N8865,N8866,N8867,N8868,N8869,N8870,N8871,N8872,
  N8873,N8874,N8875,N8876,N8877,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,
  N8886,N8887,N8888,N8889,N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,
  N8899,N8900,N8901,N8902,N8903,N8904,N8905,N8906,N8907,N8908,N8909,N8910,N8911,N8912,
  N8913,N8914,N8915,N8916,N8917,N8918,N8919,N8920,N8921,N8922,N8923,N8924,N8925,
  N8926,N8927,N8928,N8929,N8930,N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,
  N8939,N8940,N8941,N8942,N8943,N8944,N8945,N8946,N8947,N8948,N8949,N8950,N8951,N8952,
  N8953,N8954,N8955,N8956,N8957,N8958,N8959,N8960,N8961,N8962,N8963,N8964,N8965,
  N8966,N8967,N8968,N8969,N8970,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,
  N8979,N8980,N8981,N8982,N8983,N8984,N8985,N8986,N8987,N8988,N8989,N8990,N8991,N8992,
  N8993,N8994,N8995,N8996,N8997,N8998,N8999,N9000,N9001,N9002,N9003,N9004,N9005,
  N9006,N9007,N9008,N9009,N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,
  N9019,N9020,N9021,N9022,N9023,N9024,N9025,N9026,N9027,N9028,N9029,N9030,N9031,N9032,
  N9033,N9034,N9035,N9036,N9037,N9038,N9039,N9040,N9041,N9042,N9043,N9044,N9045,
  N9046,N9047,N9048,N9049,N9050,N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,
  N9059,N9060,N9061,N9062,N9063,N9064,N9065,N9066,N9067,N9068,N9069,N9070,N9071,N9072,
  N9073,N9074,N9075,N9076,N9077,N9078,N9079,N9080,N9081,N9082,N9083,N9084,N9085,
  N9086,N9087,N9088,N9089,N9090,N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,
  N9099,N9100,N9101,N9102,N9103,N9104,N9105,N9106,N9107,N9108,N9109,N9110,N9111,N9112,
  N9113,N9114,N9115,N9116,N9117,N9118,N9119,N9120,N9121,N9122,N9123,N9124,N9125,
  N9126,N9127,N9128,N9129,N9130,N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,
  N9139,N9140,N9141,N9142,N9143,N9144,N9145,N9146,N9147,N9148,N9149,N9150,N9151,N9152,
  N9153,N9154,N9155,N9156,N9157,N9158,N9159,N9160,N9161,N9162,N9163,N9164,N9165,
  N9166,N9167,N9168,N9169,N9170,N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,
  N9179,N9180,N9181,N9182,N9183,N9184,N9185,N9186,N9187,N9188,N9189,N9190,N9191,N9192,
  N9193,N9194,N9195,N9196,N9197,N9198,N9199,N9200,N9201,N9202,N9203,N9204,N9205,
  N9206,N9207,N9208,N9209,N9210,N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,
  N9219,N9220,N9221,N9222,N9223,N9224,N9225,N9226,N9227,N9228,N9229,N9230,N9231,N9232,
  N9233,N9234,N9235,N9236,N9237,N9238,N9239,N9240,N9241,N9242,N9243,N9244,N9245,
  N9246,N9247,N9248,N9249,N9250,N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,
  N9259,N9260,N9261,N9262,N9263,N9264,N9265,N9266,N9267,N9268,N9269,N9270,N9271,N9272,
  N9273,N9274,N9275,N9276,N9277,N9278,N9279,N9280,N9281,N9282,N9283,N9284,N9285,
  N9286,N9287,N9288,N9289,N9290,N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,
  N9299,N9300,N9301,N9302,N9303,N9304,N9305,N9306,N9307,N9308,N9309,N9310,N9311,N9312,
  N9313,N9314,N9315,N9316,N9317,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9325,
  N9326,N9327,N9328,N9329,N9330,N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,
  N9339,N9340,N9341,N9342,N9343,N9344,N9345,N9346,N9347,N9348,N9349,N9350,N9351,N9352,
  N9353,N9354,N9355,N9356,N9357,N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,
  N9366,N9367,N9368,N9369,N9370,N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,
  N9379,N9380,N9381,N9382,N9383,N9384,N9385,N9386,N9387,N9388,N9389,N9390,N9391,N9392,
  N9393,N9394,N9395,N9396,N9397,N9398,N9399,N9400,N9401,N9402,N9403,N9404,N9405,
  N9406,N9407,N9408,N9409,N9410,N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,
  N9419,N9420,N9421,N9422,N9423,N9424,N9425,N9426,N9427,N9428,N9429,N9430,N9431,N9432,
  N9433,N9434,N9435,N9436,N9437,N9438,N9439,N9440,N9441,N9442,N9443,N9444,N9445,
  N9446,N9447,N9448,N9449,N9450,N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,
  N9459,N9460,N9461,N9462,N9463,N9464,N9465,N9466,N9467,N9468,N9469,N9470,N9471,N9472,
  N9473,N9474,N9475,N9476,N9477,N9478,N9479,N9480,N9481,N9482,N9483,N9484,N9485,
  N9486,N9487,N9488,N9489,N9490,N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,
  N9499,N9500,N9501,N9502,N9503,N9504,N9505,N9506,N9507,N9508,N9509,N9510,N9511,N9512,
  N9513,N9514,N9515,N9516,N9517,N9518,N9519,N9520,N9521,N9522,N9523,N9524,N9525,
  N9526,N9527,N9528,N9529,N9530,N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,
  N9539,N9540,N9541,N9542,N9543,N9544,N9545,N9546,N9547,N9548,N9549,N9550,N9551,N9552,
  N9553,N9554,N9555,N9556,N9557,N9558,N9559,N9560,N9561,N9562,N9563,N9564,N9565,
  N9566,N9567,N9568,N9569,N9570,N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,
  N9579,N9580,N9581,N9582,N9583,N9584,N9585,N9586,N9587,N9588,N9589,N9590,N9591,N9592,
  N9593,N9594,N9595,N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,
  N9606,N9607,N9608,N9609,N9610,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,
  N9619,N9620,N9621,N9622,N9623,N9624,N9625,N9626,N9627,N9628,N9629,N9630,N9631,N9632,
  N9633,N9634,N9635,N9636,N9637,N9638,N9639,N9640,N9641,N9642,N9643,N9644,N9645,
  N9646,N9647,N9648,N9649,N9650,N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,
  N9659,N9660,N9661,N9662,N9663,N9664,N9665,N9666,N9667,N9668,N9669,N9670,N9671,N9672,
  N9673,N9674,N9675,N9676,N9677,N9678,N9679,N9680,N9681,N9682,N9683,N9684,N9685,
  N9686,N9687,N9688,N9689,N9690,N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,
  N9699,N9700,N9701,N9702,N9703,N9704,N9705,N9706,N9707,N9708,N9709,N9710,N9711,N9712,
  N9713,N9714,N9715,N9716,N9717,N9718,N9719,N9720,N9721,N9722,N9723,N9724,N9725,
  N9726,N9727,N9728,N9729,N9730,N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,
  N9739,N9740,N9741,N9742,N9743,N9744,N9745,N9746,N9747,N9748,N9749,N9750,N9751,N9752,
  N9753,N9754,N9755,N9756,N9757,N9758,N9759,N9760,N9761,N9762,N9763,N9764,N9765,
  N9766,N9767,N9768,N9769,N9770,N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,
  N9779,N9780,N9781,N9782,N9783,N9784,N9785,N9786,N9787,N9788,N9789,N9790,N9791,N9792,
  N9793,N9794,N9795,N9796,N9797,N9798,N9799,N9800,N9801,N9802,N9803,N9804,N9805,
  N9806,N9807,N9808,N9809,N9810,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,
  N9819,N9820,N9821,N9822,N9823,N9824,N9825,N9826,N9827,N9828,N9829,N9830,N9831,N9832,
  N9833,N9834,N9835,N9836,N9837,N9838,N9839,N9840,N9841,N9842,N9843,N9844,N9845,
  N9846,N9847,N9848,N9849,N9850,N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,
  N9859,N9860,N9861,N9862,N9863,N9864,N9865,N9866,N9867,N9868,N9869,N9870,N9871,N9872,
  N9873,N9874,N9875,N9876,N9877,N9878,N9879,N9880,N9881,N9882,N9883,N9884,N9885,
  N9886,N9887,N9888,N9889,N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,
  N9899,N9900,N9901,N9902,N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9912,
  N9913,N9914,N9915,N9916,N9917,N9918,N9919,N9920,N9921,N9922,N9923,N9924,N9925,
  N9926,N9927,N9928,N9929,N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,
  N9939,N9940,N9941,N9942,N9943,N9944,N9945,N9946,N9947,N9948,N9949,N9950,N9951,N9952,
  N9953,N9954,N9955,N9956,N9957,N9958,N9959,N9960,N9961,N9962,N9963,N9964,N9965,
  N9966,N9967,N9968,N9969,N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,
  N9979,N9980,N9981,N9982,N9983,N9984,N9985,N9986,N9987,N9988,N9989,N9990,N9991,N9992,
  N9993,N9994,N9995,N9996,N9997,N9998,N9999,N10000,N10001,N10002,N10003,N10004,
  N10005,N10006,N10007,N10008,N10009,N10010,N10011,N10012,N10013,N10014,N10015,
  N10016,N10017,N10018,N10019,N10020,N10021,N10022,N10023,N10024,N10025,N10026,N10027,
  N10028,N10029,N10030,N10031,N10032,N10033,N10034,N10035,N10036,N10037,N10038,
  N10039,N10040,N10041,N10042,N10043,N10044,N10045,N10046,N10047,N10048,N10049,N10050,
  N10051,N10052,N10053,N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061,
  N10062,N10063,N10064,N10065,N10066,N10067,N10068,N10069,N10070,N10071,N10072,N10073,
  N10074,N10075,N10076,N10077,N10078,N10079,N10080,N10081,N10082,N10083,N10084,
  N10085,N10086,N10087,N10088,N10089,N10090,N10091,N10092,N10093,N10094,N10095,
  N10096,N10097,N10098,N10099,N10100,N10101,N10102,N10103,N10104,N10105,N10106,N10107,
  N10108,N10109,N10110,N10111,N10112,N10113,N10114,N10115,N10116,N10117,N10118,
  N10119,N10120,N10121,N10122,N10123,N10124,N10125,N10126,N10127,N10128,N10129,N10130,
  N10131,N10132,N10133,N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,
  N10142,N10143,N10144,N10145,N10146,N10147,N10148,N10149,N10150,N10151,N10152,N10153,
  N10154,N10155,N10156,N10157,N10158,N10159,N10160,N10161,N10162,N10163,N10164,
  N10165,N10166,N10167,N10168,N10169,N10170,N10171,N10172,N10173,N10174,N10175,
  N10176,N10177,N10178,N10179,N10180,N10181,N10182,N10183,N10184,N10185,N10186,N10187,
  N10188,N10189,N10190,N10191,N10192,N10193,N10194,N10195,N10196,N10197,N10198,
  N10199,N10200,N10201,N10202,N10203,N10204,N10205,N10206,N10207,N10208,N10209,N10210,
  N10211,N10212,N10213,N10214,N10215,N10216,N10217,N10218,N10219,N10220,N10221,
  N10222,N10223,N10224,N10225,N10226,N10227,N10228,N10229,N10230,N10231,N10232,N10233,
  N10234,N10235,N10236,N10237,N10238,N10239,N10240,N10241,N10242,N10243,N10244,
  N10245,N10246,N10247,N10248,N10249,N10250,N10251,N10252,N10253,N10254,N10255,
  N10256,N10257,N10258,N10259,N10260,N10261,N10262,N10263,N10264,N10265,N10266,N10267,
  N10268,N10269,N10270,N10271,N10272,N10273,N10274,N10275,N10276,N10277,N10278,
  N10279,N10280,N10281,N10282,N10283,N10284,N10285,N10286,N10287,N10288,N10289,N10290,
  N10291,N10292,N10293,N10294,N10295,N10296,N10297,N10298,N10299,N10300,N10301,
  N10302,N10303,N10304,N10305,N10306,N10307,N10308,N10309,N10310,N10311,N10312,N10313,
  N10314,N10315,N10316,N10317,N10318,N10319,N10320,N10321,N10322,N10323,N10324,
  N10325,N10326,N10327,N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10335,
  N10336,N10337,N10338,N10339,N10340,N10341,N10342,N10343,N10344,N10345,N10346,N10347,
  N10348,N10349,N10350,N10351,N10352,N10353,N10354,N10355,N10356,N10357,N10358,
  N10359,N10360,N10361,N10362,N10363,N10364,N10365,N10366,N10367,N10368,N10369,N10370,
  N10371,N10372,N10373,N10374,N10375,N10376,N10377,N10378,N10379,N10380,N10381,
  N10382,N10383,N10384,N10385,N10386,N10387,N10388,N10389,N10390,N10391,N10392,N10393,
  N10394,N10395,N10396,N10397,N10398,N10399,N10400,N10401,N10402,N10403,N10404,
  N10405,N10406,N10407,N10408,N10409,N10410,N10411,N10412,N10413,N10414,N10415,
  N10416,N10417,N10418,N10419,N10420,N10421,N10422,N10423,N10424,N10425,N10426,N10427,
  N10428,N10429,N10430,N10431,N10432,N10433,N10434,N10435,N10436,N10437,N10438,
  N10439,N10440,N10441,N10442,N10443,N10444,N10445,N10446,N10447,N10448,N10449,N10450,
  N10451,N10452,N10453,N10454,N10455,N10456,N10457,N10458,N10459,N10460,N10461,
  N10462,N10463,N10464,N10465,N10466,N10467,N10468,N10469,N10470,N10471,N10472,N10473,
  N10474,N10475,N10476,N10477,N10478,N10479,N10480,N10481,N10482,N10483,N10484,
  N10485,N10486,N10487,N10488,N10489,N10490,N10491,N10492,N10493,N10494,N10495,
  N10496,N10497,N10498,N10499,N10500,N10501,N10502,N10503,N10504,N10505,N10506,N10507,
  N10508,N10509,N10510,N10511,N10512,N10513,N10514,N10515,N10516,N10517,N10518,
  N10519,N10520,N10521,N10522,N10523,N10524,N10525,N10526,N10527,N10528,N10529,N10530,
  N10531,N10532,N10533,N10534,N10535,N10536,N10537,N10538,N10539,N10540,N10541,
  N10542,N10543,N10544,N10545,N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,
  N10554,N10555,N10556,N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,
  N10565,N10566,N10567,N10568,N10569,N10570,N10571,N10572,N10573,N10574,N10575,
  N10576,N10577,N10578,N10579,N10580,N10581,N10582,N10583,N10584,N10585,N10586,N10587,
  N10588,N10589,N10590,N10591,N10592,N10593,N10594,N10595,N10596,N10597,N10598,
  N10599,N10600,N10601,N10602,N10603,N10604,N10605,N10606,N10607,N10608,N10609,N10610,
  N10611,N10612,N10613,N10614,N10615,N10616,N10617,N10618,N10619,N10620,N10621,
  N10622,N10623,N10624,N10625,N10626,N10627,N10628,N10629,N10630,N10631,N10632,N10633,
  N10634,N10635,N10636,N10637,N10638,N10639,N10640,N10641,N10642,N10643,N10644,
  N10645,N10646,N10647,N10648,N10649,N10650,N10651,N10652,N10653,N10654,N10655,
  N10656,N10657,N10658,N10659,N10660,N10661,N10662,N10663,N10664,N10665,N10666,N10667,
  N10668,N10669,N10670,N10671,N10672,N10673,N10674,N10675,N10676,N10677,N10678,
  N10679,N10680,N10681,N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,
  N10691,N10692,N10693,N10694,N10695,N10696,N10697,N10698,N10699,N10700,N10701,
  N10702,N10703,N10704,N10705,N10706,N10707,N10708,N10709,N10710,N10711,N10712,N10713,
  N10714,N10715,N10716,N10717,N10718,N10719,N10720,N10721,N10722,N10723,N10724,
  N10725,N10726,N10727,N10728,N10729,N10730,N10731,N10732,N10733,N10734,N10735,
  N10736,N10737,N10738,N10739,N10740,N10741,N10742,N10743,N10744,N10745,N10746,N10747,
  N10748,N10749,N10750,N10751,N10752,N10753,N10754,N10755,N10756,N10757,N10758,
  N10759,N10760,N10761,N10762,N10763,N10764,N10765,N10766,N10767,N10768,N10769,N10770,
  N10771,N10772,N10773,N10774,N10775,N10776,N10777,N10778,N10779,N10780,N10781,
  N10782,N10783,N10784,N10785,N10786,N10787,N10788,N10789,N10790,N10791,N10792,N10793,
  N10794,N10795,N10796,N10797,N10798,N10799,N10800,N10801,N10802,N10803,N10804,
  N10805,N10806,N10807,N10808,N10809,N10810,N10811,N10812,N10813,N10814,N10815,
  N10816,N10817,N10818,N10819,N10820,N10821,N10822,N10823,N10824,N10825,N10826,N10827,
  N10828,N10829,N10830,N10831,N10832,N10833,N10834,N10835,N10836,N10837,N10838,
  N10839,N10840,N10841,N10842,N10843,N10844,N10845,N10846,N10847,N10848,N10849,N10850,
  N10851,N10852,N10853,N10854,N10855,N10856,N10857,N10858,N10859,N10860,N10861,
  N10862,N10863,N10864,N10865,N10866,N10867,N10868,N10869,N10870,N10871,N10872,N10873,
  N10874,N10875,N10876,N10877,N10878,N10879,N10880,N10881,N10882,N10883,N10884,
  N10885,N10886,N10887,N10888,N10889,N10890,N10891,N10892,N10893,N10894,N10895,
  N10896,N10897,N10898,N10899,N10900,N10901,N10902,N10903,N10904,N10905,N10906,N10907,
  N10908,N10909,N10910,N10911,N10912,N10913,N10914,N10915,N10916,N10917,N10918,
  N10919,N10920,N10921,N10922,N10923,N10924,N10925,N10926,N10927,N10928,N10929,N10930,
  N10931,N10932,N10933,N10934,N10935,N10936,N10937,N10938,N10939,N10940,N10941,
  N10942,N10943,N10944,N10945,N10946,N10947,N10948,N10949,N10950,N10951,N10952,N10953,
  N10954,N10955,N10956,N10957,N10958,N10959,N10960,N10961,N10962,N10963,N10964,
  N10965,N10966,N10967,N10968,N10969,N10970,N10971,N10972,N10973,N10974,N10975,
  N10976,N10977,N10978,N10979,N10980,N10981,N10982,N10983,N10984,N10985,N10986,N10987,
  N10988,N10989,N10990,N10991,N10992,N10993,N10994,N10995,N10996,N10997,N10998,
  N10999,N11000,N11001,N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11009,N11010,
  N11011,N11012,N11013,N11014,N11015,N11016,N11017,N11018,N11019,N11020,N11021,
  N11022,N11023,N11024,N11025,N11026,N11027,N11028,N11029,N11030,N11031,N11032,N11033,
  N11034,N11035,N11036,N11037,N11038,N11039,N11040,N11041,N11042,N11043,N11044,
  N11045,N11046,N11047,N11048,N11049,N11050,N11051,N11052,N11053,N11054,N11055,
  N11056,N11057,N11058,N11059,N11060,N11061,N11062,N11063,N11064,N11065,N11066,N11067,
  N11068,N11069,N11070,N11071,N11072,N11073,N11074,N11075,N11076,N11077,N11078,
  N11079,N11080,N11081,N11082,N11083,N11084,N11085,N11086,N11087,N11088,N11089,N11090,
  N11091,N11092,N11093,N11094,N11095,N11096,N11097,N11098,N11099,N11100,N11101,
  N11102,N11103,N11104,N11105,N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,
  N11114,N11115,N11116,N11117,N11118,N11119,N11120,N11121,N11122,N11123,N11124,
  N11125,N11126,N11127,N11128,N11129,N11130,N11131,N11132,N11133,N11134,N11135,
  N11136,N11137,N11138,N11139,N11140,N11141,N11142,N11143,N11144,N11145,N11146,N11147,
  N11148,N11149,N11150,N11151,N11152,N11153,N11154,N11155,N11156,N11157,N11158,
  N11159,N11160,N11161,N11162,N11163,N11164,N11165,N11166,N11167,N11168,N11169,N11170,
  N11171,N11172,N11173,N11174,N11175,N11176,N11177,N11178,N11179,N11180,N11181,
  N11182,N11183,N11184,N11185,N11186,N11187,N11188,N11189,N11190,N11191,N11192,N11193,
  N11194,N11195,N11196,N11197,N11198,N11199,N11200,N11201,N11202,N11203,N11204,
  N11205,N11206,N11207,N11208,N11209,N11210,N11211,N11212,N11213,N11214,N11215,
  N11216,N11217,N11218,N11219,N11220,N11221,N11222,N11223,N11224,N11225,N11226,N11227,
  N11228,N11229,N11230,N11231,N11232,N11233,N11234,N11235,N11236,N11237,N11238,
  N11239,N11240,N11241,N11242,N11243,N11244,N11245,N11246,N11247,N11248,N11249,N11250,
  N11251,N11252,N11253,N11254,N11255,N11256,N11257,N11258,N11259,N11260,N11261,
  N11262,N11263,N11264,N11265,N11266,N11267,N11268,N11269,N11270,N11271,N11272,N11273,
  N11274,N11275,N11276,N11277,N11278,N11279,N11280,N11281,N11282,N11283,N11284,
  N11285,N11286,N11287,N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,
  N11296,N11297,N11298,N11299,N11300,N11301,N11302,N11303,N11304,N11305,N11306,N11307,
  N11308,N11309,N11310,N11311,N11312,N11313,N11314,N11315,N11316,N11317,N11318,
  N11319,N11320,N11321,N11322,N11323,N11324,N11325,N11326,N11327,N11328,N11329,N11330,
  N11331,N11332,N11333,N11334,N11335,N11336,N11337,N11338,N11339,N11340,N11341,
  N11342,N11343,N11344,N11345,N11346,N11347,N11348,N11349,N11350,N11351,N11352,N11353,
  N11354,N11355,N11356,N11357,N11358,N11359,N11360,N11361,N11362,N11363,N11364,
  N11365,N11366,N11367,N11368,N11369,N11370,N11371,N11372,N11373,N11374,N11375,
  N11376,N11377,N11378,N11379,N11380,N11381,N11382,N11383,N11384,N11385,N11386,N11387,
  N11388,N11389,N11390,N11391,N11392,N11393,N11394,N11395,N11396,N11397,N11398,
  N11399,N11400,N11401,N11402,N11403,N11404,N11405,N11406,N11407,N11408,N11409,N11410,
  N11411,N11412,N11413,N11414,N11415,N11416,N11417,N11418,N11419,N11420,N11421,
  N11422,N11423,N11424,N11425,N11426,N11427,N11428,N11429,N11430,N11431,N11432,N11433,
  N11434,N11435,N11436,N11437,N11438,N11439,N11440,N11441,N11442,N11443,N11444,
  N11445,N11446,N11447,N11448,N11449,N11450,N11451,N11452,N11453,N11454,N11455,
  N11456,N11457,N11458,N11459,N11460,N11461,N11462,N11463,N11464,N11465,N11466,N11467,
  N11468,N11469,N11470,N11471,N11472,N11473,N11474,N11475,N11476,N11477,N11478,
  N11479,N11480,N11481,N11482,N11483,N11484,N11485,N11486,N11487,N11488,N11489,N11490,
  N11491,N11492,N11493,N11494,N11495,N11496,N11497,N11498,N11499,N11500,N11501,
  N11502,N11503,N11504,N11505,N11506,N11507,N11508,N11509,N11510,N11511,N11512,N11513,
  N11514,N11515,N11516,N11517,N11518,N11519,N11520,N11521,N11522,N11523,N11524,
  N11525,N11526,N11527,N11528,N11529,N11530,N11531,N11532,N11533,N11534,N11535,
  N11536,N11537,N11538,N11539,N11540,N11541,N11542,N11543,N11544,N11545,N11546,N11547,
  N11548,N11549,N11550,N11551,N11552,N11553,N11554,N11555,N11556,N11557,N11558,
  N11559,N11560,N11561,N11562,N11563,N11564,N11565,N11566,N11567,N11568,N11569,N11570,
  N11571,N11572,N11573,N11574,N11575,N11576,N11577,N11578,N11579,N11580,N11581,
  N11582,N11583,N11584,N11585,N11586,N11587,N11588,N11589,N11590,N11591,N11592,N11593,
  N11594,N11595,N11596,N11597,N11598,N11599,N11600,N11601,N11602,N11603,N11604,
  N11605,N11606,N11607,N11608,N11609,N11610,N11611,N11612,N11613,N11614,N11615,
  N11616,N11617,N11618,N11619,N11620,N11621,N11622,N11623,N11624,N11625,N11626,N11627,
  N11628,N11629,N11630,N11631,N11632,N11633,N11634,N11635,N11636,N11637,N11638,
  N11639,N11640,N11641,N11642,N11643,N11644,N11645,N11646,N11647,N11648,N11649,N11650,
  N11651,N11652,N11653,N11654,N11655,N11656,N11657,N11658,N11659;
  wire [5:0] \nz.addr_r ;
  wire [5119:0] \nz.mem ;
  reg \nz.addr_r_5_sv2v_reg ,\nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,
  \nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,
  \nz.mem_5119_sv2v_reg ,\nz.mem_5118_sv2v_reg ,\nz.mem_5117_sv2v_reg ,\nz.mem_5116_sv2v_reg ,
  \nz.mem_5115_sv2v_reg ,\nz.mem_5114_sv2v_reg ,\nz.mem_5113_sv2v_reg ,
  \nz.mem_5112_sv2v_reg ,\nz.mem_5111_sv2v_reg ,\nz.mem_5110_sv2v_reg ,\nz.mem_5109_sv2v_reg ,
  \nz.mem_5108_sv2v_reg ,\nz.mem_5107_sv2v_reg ,\nz.mem_5106_sv2v_reg ,
  \nz.mem_5105_sv2v_reg ,\nz.mem_5104_sv2v_reg ,\nz.mem_5103_sv2v_reg ,\nz.mem_5102_sv2v_reg ,
  \nz.mem_5101_sv2v_reg ,\nz.mem_5100_sv2v_reg ,\nz.mem_5099_sv2v_reg ,
  \nz.mem_5098_sv2v_reg ,\nz.mem_5097_sv2v_reg ,\nz.mem_5096_sv2v_reg ,\nz.mem_5095_sv2v_reg ,
  \nz.mem_5094_sv2v_reg ,\nz.mem_5093_sv2v_reg ,\nz.mem_5092_sv2v_reg ,
  \nz.mem_5091_sv2v_reg ,\nz.mem_5090_sv2v_reg ,\nz.mem_5089_sv2v_reg ,\nz.mem_5088_sv2v_reg ,
  \nz.mem_5087_sv2v_reg ,\nz.mem_5086_sv2v_reg ,\nz.mem_5085_sv2v_reg ,
  \nz.mem_5084_sv2v_reg ,\nz.mem_5083_sv2v_reg ,\nz.mem_5082_sv2v_reg ,\nz.mem_5081_sv2v_reg ,
  \nz.mem_5080_sv2v_reg ,\nz.mem_5079_sv2v_reg ,\nz.mem_5078_sv2v_reg ,
  \nz.mem_5077_sv2v_reg ,\nz.mem_5076_sv2v_reg ,\nz.mem_5075_sv2v_reg ,\nz.mem_5074_sv2v_reg ,
  \nz.mem_5073_sv2v_reg ,\nz.mem_5072_sv2v_reg ,\nz.mem_5071_sv2v_reg ,
  \nz.mem_5070_sv2v_reg ,\nz.mem_5069_sv2v_reg ,\nz.mem_5068_sv2v_reg ,\nz.mem_5067_sv2v_reg ,
  \nz.mem_5066_sv2v_reg ,\nz.mem_5065_sv2v_reg ,\nz.mem_5064_sv2v_reg ,
  \nz.mem_5063_sv2v_reg ,\nz.mem_5062_sv2v_reg ,\nz.mem_5061_sv2v_reg ,\nz.mem_5060_sv2v_reg ,
  \nz.mem_5059_sv2v_reg ,\nz.mem_5058_sv2v_reg ,\nz.mem_5057_sv2v_reg ,
  \nz.mem_5056_sv2v_reg ,\nz.mem_5055_sv2v_reg ,\nz.mem_5054_sv2v_reg ,\nz.mem_5053_sv2v_reg ,
  \nz.mem_5052_sv2v_reg ,\nz.mem_5051_sv2v_reg ,\nz.mem_5050_sv2v_reg ,
  \nz.mem_5049_sv2v_reg ,\nz.mem_5048_sv2v_reg ,\nz.mem_5047_sv2v_reg ,\nz.mem_5046_sv2v_reg ,
  \nz.mem_5045_sv2v_reg ,\nz.mem_5044_sv2v_reg ,\nz.mem_5043_sv2v_reg ,
  \nz.mem_5042_sv2v_reg ,\nz.mem_5041_sv2v_reg ,\nz.mem_5040_sv2v_reg ,
  \nz.mem_5039_sv2v_reg ,\nz.mem_5038_sv2v_reg ,\nz.mem_5037_sv2v_reg ,\nz.mem_5036_sv2v_reg ,
  \nz.mem_5035_sv2v_reg ,\nz.mem_5034_sv2v_reg ,\nz.mem_5033_sv2v_reg ,
  \nz.mem_5032_sv2v_reg ,\nz.mem_5031_sv2v_reg ,\nz.mem_5030_sv2v_reg ,\nz.mem_5029_sv2v_reg ,
  \nz.mem_5028_sv2v_reg ,\nz.mem_5027_sv2v_reg ,\nz.mem_5026_sv2v_reg ,
  \nz.mem_5025_sv2v_reg ,\nz.mem_5024_sv2v_reg ,\nz.mem_5023_sv2v_reg ,\nz.mem_5022_sv2v_reg ,
  \nz.mem_5021_sv2v_reg ,\nz.mem_5020_sv2v_reg ,\nz.mem_5019_sv2v_reg ,
  \nz.mem_5018_sv2v_reg ,\nz.mem_5017_sv2v_reg ,\nz.mem_5016_sv2v_reg ,\nz.mem_5015_sv2v_reg ,
  \nz.mem_5014_sv2v_reg ,\nz.mem_5013_sv2v_reg ,\nz.mem_5012_sv2v_reg ,
  \nz.mem_5011_sv2v_reg ,\nz.mem_5010_sv2v_reg ,\nz.mem_5009_sv2v_reg ,\nz.mem_5008_sv2v_reg ,
  \nz.mem_5007_sv2v_reg ,\nz.mem_5006_sv2v_reg ,\nz.mem_5005_sv2v_reg ,
  \nz.mem_5004_sv2v_reg ,\nz.mem_5003_sv2v_reg ,\nz.mem_5002_sv2v_reg ,\nz.mem_5001_sv2v_reg ,
  \nz.mem_5000_sv2v_reg ,\nz.mem_4999_sv2v_reg ,\nz.mem_4998_sv2v_reg ,
  \nz.mem_4997_sv2v_reg ,\nz.mem_4996_sv2v_reg ,\nz.mem_4995_sv2v_reg ,\nz.mem_4994_sv2v_reg ,
  \nz.mem_4993_sv2v_reg ,\nz.mem_4992_sv2v_reg ,\nz.mem_4991_sv2v_reg ,
  \nz.mem_4990_sv2v_reg ,\nz.mem_4989_sv2v_reg ,\nz.mem_4988_sv2v_reg ,\nz.mem_4987_sv2v_reg ,
  \nz.mem_4986_sv2v_reg ,\nz.mem_4985_sv2v_reg ,\nz.mem_4984_sv2v_reg ,
  \nz.mem_4983_sv2v_reg ,\nz.mem_4982_sv2v_reg ,\nz.mem_4981_sv2v_reg ,\nz.mem_4980_sv2v_reg ,
  \nz.mem_4979_sv2v_reg ,\nz.mem_4978_sv2v_reg ,\nz.mem_4977_sv2v_reg ,
  \nz.mem_4976_sv2v_reg ,\nz.mem_4975_sv2v_reg ,\nz.mem_4974_sv2v_reg ,\nz.mem_4973_sv2v_reg ,
  \nz.mem_4972_sv2v_reg ,\nz.mem_4971_sv2v_reg ,\nz.mem_4970_sv2v_reg ,
  \nz.mem_4969_sv2v_reg ,\nz.mem_4968_sv2v_reg ,\nz.mem_4967_sv2v_reg ,\nz.mem_4966_sv2v_reg ,
  \nz.mem_4965_sv2v_reg ,\nz.mem_4964_sv2v_reg ,\nz.mem_4963_sv2v_reg ,
  \nz.mem_4962_sv2v_reg ,\nz.mem_4961_sv2v_reg ,\nz.mem_4960_sv2v_reg ,
  \nz.mem_4959_sv2v_reg ,\nz.mem_4958_sv2v_reg ,\nz.mem_4957_sv2v_reg ,\nz.mem_4956_sv2v_reg ,
  \nz.mem_4955_sv2v_reg ,\nz.mem_4954_sv2v_reg ,\nz.mem_4953_sv2v_reg ,
  \nz.mem_4952_sv2v_reg ,\nz.mem_4951_sv2v_reg ,\nz.mem_4950_sv2v_reg ,\nz.mem_4949_sv2v_reg ,
  \nz.mem_4948_sv2v_reg ,\nz.mem_4947_sv2v_reg ,\nz.mem_4946_sv2v_reg ,
  \nz.mem_4945_sv2v_reg ,\nz.mem_4944_sv2v_reg ,\nz.mem_4943_sv2v_reg ,\nz.mem_4942_sv2v_reg ,
  \nz.mem_4941_sv2v_reg ,\nz.mem_4940_sv2v_reg ,\nz.mem_4939_sv2v_reg ,
  \nz.mem_4938_sv2v_reg ,\nz.mem_4937_sv2v_reg ,\nz.mem_4936_sv2v_reg ,\nz.mem_4935_sv2v_reg ,
  \nz.mem_4934_sv2v_reg ,\nz.mem_4933_sv2v_reg ,\nz.mem_4932_sv2v_reg ,
  \nz.mem_4931_sv2v_reg ,\nz.mem_4930_sv2v_reg ,\nz.mem_4929_sv2v_reg ,\nz.mem_4928_sv2v_reg ,
  \nz.mem_4927_sv2v_reg ,\nz.mem_4926_sv2v_reg ,\nz.mem_4925_sv2v_reg ,
  \nz.mem_4924_sv2v_reg ,\nz.mem_4923_sv2v_reg ,\nz.mem_4922_sv2v_reg ,\nz.mem_4921_sv2v_reg ,
  \nz.mem_4920_sv2v_reg ,\nz.mem_4919_sv2v_reg ,\nz.mem_4918_sv2v_reg ,
  \nz.mem_4917_sv2v_reg ,\nz.mem_4916_sv2v_reg ,\nz.mem_4915_sv2v_reg ,\nz.mem_4914_sv2v_reg ,
  \nz.mem_4913_sv2v_reg ,\nz.mem_4912_sv2v_reg ,\nz.mem_4911_sv2v_reg ,
  \nz.mem_4910_sv2v_reg ,\nz.mem_4909_sv2v_reg ,\nz.mem_4908_sv2v_reg ,\nz.mem_4907_sv2v_reg ,
  \nz.mem_4906_sv2v_reg ,\nz.mem_4905_sv2v_reg ,\nz.mem_4904_sv2v_reg ,
  \nz.mem_4903_sv2v_reg ,\nz.mem_4902_sv2v_reg ,\nz.mem_4901_sv2v_reg ,\nz.mem_4900_sv2v_reg ,
  \nz.mem_4899_sv2v_reg ,\nz.mem_4898_sv2v_reg ,\nz.mem_4897_sv2v_reg ,
  \nz.mem_4896_sv2v_reg ,\nz.mem_4895_sv2v_reg ,\nz.mem_4894_sv2v_reg ,\nz.mem_4893_sv2v_reg ,
  \nz.mem_4892_sv2v_reg ,\nz.mem_4891_sv2v_reg ,\nz.mem_4890_sv2v_reg ,
  \nz.mem_4889_sv2v_reg ,\nz.mem_4888_sv2v_reg ,\nz.mem_4887_sv2v_reg ,\nz.mem_4886_sv2v_reg ,
  \nz.mem_4885_sv2v_reg ,\nz.mem_4884_sv2v_reg ,\nz.mem_4883_sv2v_reg ,
  \nz.mem_4882_sv2v_reg ,\nz.mem_4881_sv2v_reg ,\nz.mem_4880_sv2v_reg ,
  \nz.mem_4879_sv2v_reg ,\nz.mem_4878_sv2v_reg ,\nz.mem_4877_sv2v_reg ,\nz.mem_4876_sv2v_reg ,
  \nz.mem_4875_sv2v_reg ,\nz.mem_4874_sv2v_reg ,\nz.mem_4873_sv2v_reg ,
  \nz.mem_4872_sv2v_reg ,\nz.mem_4871_sv2v_reg ,\nz.mem_4870_sv2v_reg ,\nz.mem_4869_sv2v_reg ,
  \nz.mem_4868_sv2v_reg ,\nz.mem_4867_sv2v_reg ,\nz.mem_4866_sv2v_reg ,
  \nz.mem_4865_sv2v_reg ,\nz.mem_4864_sv2v_reg ,\nz.mem_4863_sv2v_reg ,\nz.mem_4862_sv2v_reg ,
  \nz.mem_4861_sv2v_reg ,\nz.mem_4860_sv2v_reg ,\nz.mem_4859_sv2v_reg ,
  \nz.mem_4858_sv2v_reg ,\nz.mem_4857_sv2v_reg ,\nz.mem_4856_sv2v_reg ,\nz.mem_4855_sv2v_reg ,
  \nz.mem_4854_sv2v_reg ,\nz.mem_4853_sv2v_reg ,\nz.mem_4852_sv2v_reg ,
  \nz.mem_4851_sv2v_reg ,\nz.mem_4850_sv2v_reg ,\nz.mem_4849_sv2v_reg ,\nz.mem_4848_sv2v_reg ,
  \nz.mem_4847_sv2v_reg ,\nz.mem_4846_sv2v_reg ,\nz.mem_4845_sv2v_reg ,
  \nz.mem_4844_sv2v_reg ,\nz.mem_4843_sv2v_reg ,\nz.mem_4842_sv2v_reg ,\nz.mem_4841_sv2v_reg ,
  \nz.mem_4840_sv2v_reg ,\nz.mem_4839_sv2v_reg ,\nz.mem_4838_sv2v_reg ,
  \nz.mem_4837_sv2v_reg ,\nz.mem_4836_sv2v_reg ,\nz.mem_4835_sv2v_reg ,\nz.mem_4834_sv2v_reg ,
  \nz.mem_4833_sv2v_reg ,\nz.mem_4832_sv2v_reg ,\nz.mem_4831_sv2v_reg ,
  \nz.mem_4830_sv2v_reg ,\nz.mem_4829_sv2v_reg ,\nz.mem_4828_sv2v_reg ,\nz.mem_4827_sv2v_reg ,
  \nz.mem_4826_sv2v_reg ,\nz.mem_4825_sv2v_reg ,\nz.mem_4824_sv2v_reg ,
  \nz.mem_4823_sv2v_reg ,\nz.mem_4822_sv2v_reg ,\nz.mem_4821_sv2v_reg ,\nz.mem_4820_sv2v_reg ,
  \nz.mem_4819_sv2v_reg ,\nz.mem_4818_sv2v_reg ,\nz.mem_4817_sv2v_reg ,
  \nz.mem_4816_sv2v_reg ,\nz.mem_4815_sv2v_reg ,\nz.mem_4814_sv2v_reg ,\nz.mem_4813_sv2v_reg ,
  \nz.mem_4812_sv2v_reg ,\nz.mem_4811_sv2v_reg ,\nz.mem_4810_sv2v_reg ,
  \nz.mem_4809_sv2v_reg ,\nz.mem_4808_sv2v_reg ,\nz.mem_4807_sv2v_reg ,\nz.mem_4806_sv2v_reg ,
  \nz.mem_4805_sv2v_reg ,\nz.mem_4804_sv2v_reg ,\nz.mem_4803_sv2v_reg ,
  \nz.mem_4802_sv2v_reg ,\nz.mem_4801_sv2v_reg ,\nz.mem_4800_sv2v_reg ,
  \nz.mem_4799_sv2v_reg ,\nz.mem_4798_sv2v_reg ,\nz.mem_4797_sv2v_reg ,\nz.mem_4796_sv2v_reg ,
  \nz.mem_4795_sv2v_reg ,\nz.mem_4794_sv2v_reg ,\nz.mem_4793_sv2v_reg ,
  \nz.mem_4792_sv2v_reg ,\nz.mem_4791_sv2v_reg ,\nz.mem_4790_sv2v_reg ,\nz.mem_4789_sv2v_reg ,
  \nz.mem_4788_sv2v_reg ,\nz.mem_4787_sv2v_reg ,\nz.mem_4786_sv2v_reg ,
  \nz.mem_4785_sv2v_reg ,\nz.mem_4784_sv2v_reg ,\nz.mem_4783_sv2v_reg ,\nz.mem_4782_sv2v_reg ,
  \nz.mem_4781_sv2v_reg ,\nz.mem_4780_sv2v_reg ,\nz.mem_4779_sv2v_reg ,
  \nz.mem_4778_sv2v_reg ,\nz.mem_4777_sv2v_reg ,\nz.mem_4776_sv2v_reg ,\nz.mem_4775_sv2v_reg ,
  \nz.mem_4774_sv2v_reg ,\nz.mem_4773_sv2v_reg ,\nz.mem_4772_sv2v_reg ,
  \nz.mem_4771_sv2v_reg ,\nz.mem_4770_sv2v_reg ,\nz.mem_4769_sv2v_reg ,\nz.mem_4768_sv2v_reg ,
  \nz.mem_4767_sv2v_reg ,\nz.mem_4766_sv2v_reg ,\nz.mem_4765_sv2v_reg ,
  \nz.mem_4764_sv2v_reg ,\nz.mem_4763_sv2v_reg ,\nz.mem_4762_sv2v_reg ,\nz.mem_4761_sv2v_reg ,
  \nz.mem_4760_sv2v_reg ,\nz.mem_4759_sv2v_reg ,\nz.mem_4758_sv2v_reg ,
  \nz.mem_4757_sv2v_reg ,\nz.mem_4756_sv2v_reg ,\nz.mem_4755_sv2v_reg ,\nz.mem_4754_sv2v_reg ,
  \nz.mem_4753_sv2v_reg ,\nz.mem_4752_sv2v_reg ,\nz.mem_4751_sv2v_reg ,
  \nz.mem_4750_sv2v_reg ,\nz.mem_4749_sv2v_reg ,\nz.mem_4748_sv2v_reg ,\nz.mem_4747_sv2v_reg ,
  \nz.mem_4746_sv2v_reg ,\nz.mem_4745_sv2v_reg ,\nz.mem_4744_sv2v_reg ,
  \nz.mem_4743_sv2v_reg ,\nz.mem_4742_sv2v_reg ,\nz.mem_4741_sv2v_reg ,\nz.mem_4740_sv2v_reg ,
  \nz.mem_4739_sv2v_reg ,\nz.mem_4738_sv2v_reg ,\nz.mem_4737_sv2v_reg ,
  \nz.mem_4736_sv2v_reg ,\nz.mem_4735_sv2v_reg ,\nz.mem_4734_sv2v_reg ,\nz.mem_4733_sv2v_reg ,
  \nz.mem_4732_sv2v_reg ,\nz.mem_4731_sv2v_reg ,\nz.mem_4730_sv2v_reg ,
  \nz.mem_4729_sv2v_reg ,\nz.mem_4728_sv2v_reg ,\nz.mem_4727_sv2v_reg ,\nz.mem_4726_sv2v_reg ,
  \nz.mem_4725_sv2v_reg ,\nz.mem_4724_sv2v_reg ,\nz.mem_4723_sv2v_reg ,
  \nz.mem_4722_sv2v_reg ,\nz.mem_4721_sv2v_reg ,\nz.mem_4720_sv2v_reg ,
  \nz.mem_4719_sv2v_reg ,\nz.mem_4718_sv2v_reg ,\nz.mem_4717_sv2v_reg ,\nz.mem_4716_sv2v_reg ,
  \nz.mem_4715_sv2v_reg ,\nz.mem_4714_sv2v_reg ,\nz.mem_4713_sv2v_reg ,
  \nz.mem_4712_sv2v_reg ,\nz.mem_4711_sv2v_reg ,\nz.mem_4710_sv2v_reg ,\nz.mem_4709_sv2v_reg ,
  \nz.mem_4708_sv2v_reg ,\nz.mem_4707_sv2v_reg ,\nz.mem_4706_sv2v_reg ,
  \nz.mem_4705_sv2v_reg ,\nz.mem_4704_sv2v_reg ,\nz.mem_4703_sv2v_reg ,\nz.mem_4702_sv2v_reg ,
  \nz.mem_4701_sv2v_reg ,\nz.mem_4700_sv2v_reg ,\nz.mem_4699_sv2v_reg ,
  \nz.mem_4698_sv2v_reg ,\nz.mem_4697_sv2v_reg ,\nz.mem_4696_sv2v_reg ,\nz.mem_4695_sv2v_reg ,
  \nz.mem_4694_sv2v_reg ,\nz.mem_4693_sv2v_reg ,\nz.mem_4692_sv2v_reg ,
  \nz.mem_4691_sv2v_reg ,\nz.mem_4690_sv2v_reg ,\nz.mem_4689_sv2v_reg ,\nz.mem_4688_sv2v_reg ,
  \nz.mem_4687_sv2v_reg ,\nz.mem_4686_sv2v_reg ,\nz.mem_4685_sv2v_reg ,
  \nz.mem_4684_sv2v_reg ,\nz.mem_4683_sv2v_reg ,\nz.mem_4682_sv2v_reg ,\nz.mem_4681_sv2v_reg ,
  \nz.mem_4680_sv2v_reg ,\nz.mem_4679_sv2v_reg ,\nz.mem_4678_sv2v_reg ,
  \nz.mem_4677_sv2v_reg ,\nz.mem_4676_sv2v_reg ,\nz.mem_4675_sv2v_reg ,\nz.mem_4674_sv2v_reg ,
  \nz.mem_4673_sv2v_reg ,\nz.mem_4672_sv2v_reg ,\nz.mem_4671_sv2v_reg ,
  \nz.mem_4670_sv2v_reg ,\nz.mem_4669_sv2v_reg ,\nz.mem_4668_sv2v_reg ,\nz.mem_4667_sv2v_reg ,
  \nz.mem_4666_sv2v_reg ,\nz.mem_4665_sv2v_reg ,\nz.mem_4664_sv2v_reg ,
  \nz.mem_4663_sv2v_reg ,\nz.mem_4662_sv2v_reg ,\nz.mem_4661_sv2v_reg ,\nz.mem_4660_sv2v_reg ,
  \nz.mem_4659_sv2v_reg ,\nz.mem_4658_sv2v_reg ,\nz.mem_4657_sv2v_reg ,
  \nz.mem_4656_sv2v_reg ,\nz.mem_4655_sv2v_reg ,\nz.mem_4654_sv2v_reg ,\nz.mem_4653_sv2v_reg ,
  \nz.mem_4652_sv2v_reg ,\nz.mem_4651_sv2v_reg ,\nz.mem_4650_sv2v_reg ,
  \nz.mem_4649_sv2v_reg ,\nz.mem_4648_sv2v_reg ,\nz.mem_4647_sv2v_reg ,\nz.mem_4646_sv2v_reg ,
  \nz.mem_4645_sv2v_reg ,\nz.mem_4644_sv2v_reg ,\nz.mem_4643_sv2v_reg ,
  \nz.mem_4642_sv2v_reg ,\nz.mem_4641_sv2v_reg ,\nz.mem_4640_sv2v_reg ,
  \nz.mem_4639_sv2v_reg ,\nz.mem_4638_sv2v_reg ,\nz.mem_4637_sv2v_reg ,\nz.mem_4636_sv2v_reg ,
  \nz.mem_4635_sv2v_reg ,\nz.mem_4634_sv2v_reg ,\nz.mem_4633_sv2v_reg ,
  \nz.mem_4632_sv2v_reg ,\nz.mem_4631_sv2v_reg ,\nz.mem_4630_sv2v_reg ,\nz.mem_4629_sv2v_reg ,
  \nz.mem_4628_sv2v_reg ,\nz.mem_4627_sv2v_reg ,\nz.mem_4626_sv2v_reg ,
  \nz.mem_4625_sv2v_reg ,\nz.mem_4624_sv2v_reg ,\nz.mem_4623_sv2v_reg ,\nz.mem_4622_sv2v_reg ,
  \nz.mem_4621_sv2v_reg ,\nz.mem_4620_sv2v_reg ,\nz.mem_4619_sv2v_reg ,
  \nz.mem_4618_sv2v_reg ,\nz.mem_4617_sv2v_reg ,\nz.mem_4616_sv2v_reg ,\nz.mem_4615_sv2v_reg ,
  \nz.mem_4614_sv2v_reg ,\nz.mem_4613_sv2v_reg ,\nz.mem_4612_sv2v_reg ,
  \nz.mem_4611_sv2v_reg ,\nz.mem_4610_sv2v_reg ,\nz.mem_4609_sv2v_reg ,\nz.mem_4608_sv2v_reg ,
  \nz.mem_4607_sv2v_reg ,\nz.mem_4606_sv2v_reg ,\nz.mem_4605_sv2v_reg ,
  \nz.mem_4604_sv2v_reg ,\nz.mem_4603_sv2v_reg ,\nz.mem_4602_sv2v_reg ,\nz.mem_4601_sv2v_reg ,
  \nz.mem_4600_sv2v_reg ,\nz.mem_4599_sv2v_reg ,\nz.mem_4598_sv2v_reg ,
  \nz.mem_4597_sv2v_reg ,\nz.mem_4596_sv2v_reg ,\nz.mem_4595_sv2v_reg ,\nz.mem_4594_sv2v_reg ,
  \nz.mem_4593_sv2v_reg ,\nz.mem_4592_sv2v_reg ,\nz.mem_4591_sv2v_reg ,
  \nz.mem_4590_sv2v_reg ,\nz.mem_4589_sv2v_reg ,\nz.mem_4588_sv2v_reg ,\nz.mem_4587_sv2v_reg ,
  \nz.mem_4586_sv2v_reg ,\nz.mem_4585_sv2v_reg ,\nz.mem_4584_sv2v_reg ,
  \nz.mem_4583_sv2v_reg ,\nz.mem_4582_sv2v_reg ,\nz.mem_4581_sv2v_reg ,\nz.mem_4580_sv2v_reg ,
  \nz.mem_4579_sv2v_reg ,\nz.mem_4578_sv2v_reg ,\nz.mem_4577_sv2v_reg ,
  \nz.mem_4576_sv2v_reg ,\nz.mem_4575_sv2v_reg ,\nz.mem_4574_sv2v_reg ,\nz.mem_4573_sv2v_reg ,
  \nz.mem_4572_sv2v_reg ,\nz.mem_4571_sv2v_reg ,\nz.mem_4570_sv2v_reg ,
  \nz.mem_4569_sv2v_reg ,\nz.mem_4568_sv2v_reg ,\nz.mem_4567_sv2v_reg ,\nz.mem_4566_sv2v_reg ,
  \nz.mem_4565_sv2v_reg ,\nz.mem_4564_sv2v_reg ,\nz.mem_4563_sv2v_reg ,
  \nz.mem_4562_sv2v_reg ,\nz.mem_4561_sv2v_reg ,\nz.mem_4560_sv2v_reg ,
  \nz.mem_4559_sv2v_reg ,\nz.mem_4558_sv2v_reg ,\nz.mem_4557_sv2v_reg ,\nz.mem_4556_sv2v_reg ,
  \nz.mem_4555_sv2v_reg ,\nz.mem_4554_sv2v_reg ,\nz.mem_4553_sv2v_reg ,
  \nz.mem_4552_sv2v_reg ,\nz.mem_4551_sv2v_reg ,\nz.mem_4550_sv2v_reg ,\nz.mem_4549_sv2v_reg ,
  \nz.mem_4548_sv2v_reg ,\nz.mem_4547_sv2v_reg ,\nz.mem_4546_sv2v_reg ,
  \nz.mem_4545_sv2v_reg ,\nz.mem_4544_sv2v_reg ,\nz.mem_4543_sv2v_reg ,\nz.mem_4542_sv2v_reg ,
  \nz.mem_4541_sv2v_reg ,\nz.mem_4540_sv2v_reg ,\nz.mem_4539_sv2v_reg ,
  \nz.mem_4538_sv2v_reg ,\nz.mem_4537_sv2v_reg ,\nz.mem_4536_sv2v_reg ,\nz.mem_4535_sv2v_reg ,
  \nz.mem_4534_sv2v_reg ,\nz.mem_4533_sv2v_reg ,\nz.mem_4532_sv2v_reg ,
  \nz.mem_4531_sv2v_reg ,\nz.mem_4530_sv2v_reg ,\nz.mem_4529_sv2v_reg ,\nz.mem_4528_sv2v_reg ,
  \nz.mem_4527_sv2v_reg ,\nz.mem_4526_sv2v_reg ,\nz.mem_4525_sv2v_reg ,
  \nz.mem_4524_sv2v_reg ,\nz.mem_4523_sv2v_reg ,\nz.mem_4522_sv2v_reg ,\nz.mem_4521_sv2v_reg ,
  \nz.mem_4520_sv2v_reg ,\nz.mem_4519_sv2v_reg ,\nz.mem_4518_sv2v_reg ,
  \nz.mem_4517_sv2v_reg ,\nz.mem_4516_sv2v_reg ,\nz.mem_4515_sv2v_reg ,\nz.mem_4514_sv2v_reg ,
  \nz.mem_4513_sv2v_reg ,\nz.mem_4512_sv2v_reg ,\nz.mem_4511_sv2v_reg ,
  \nz.mem_4510_sv2v_reg ,\nz.mem_4509_sv2v_reg ,\nz.mem_4508_sv2v_reg ,\nz.mem_4507_sv2v_reg ,
  \nz.mem_4506_sv2v_reg ,\nz.mem_4505_sv2v_reg ,\nz.mem_4504_sv2v_reg ,
  \nz.mem_4503_sv2v_reg ,\nz.mem_4502_sv2v_reg ,\nz.mem_4501_sv2v_reg ,\nz.mem_4500_sv2v_reg ,
  \nz.mem_4499_sv2v_reg ,\nz.mem_4498_sv2v_reg ,\nz.mem_4497_sv2v_reg ,
  \nz.mem_4496_sv2v_reg ,\nz.mem_4495_sv2v_reg ,\nz.mem_4494_sv2v_reg ,\nz.mem_4493_sv2v_reg ,
  \nz.mem_4492_sv2v_reg ,\nz.mem_4491_sv2v_reg ,\nz.mem_4490_sv2v_reg ,
  \nz.mem_4489_sv2v_reg ,\nz.mem_4488_sv2v_reg ,\nz.mem_4487_sv2v_reg ,\nz.mem_4486_sv2v_reg ,
  \nz.mem_4485_sv2v_reg ,\nz.mem_4484_sv2v_reg ,\nz.mem_4483_sv2v_reg ,
  \nz.mem_4482_sv2v_reg ,\nz.mem_4481_sv2v_reg ,\nz.mem_4480_sv2v_reg ,
  \nz.mem_4479_sv2v_reg ,\nz.mem_4478_sv2v_reg ,\nz.mem_4477_sv2v_reg ,\nz.mem_4476_sv2v_reg ,
  \nz.mem_4475_sv2v_reg ,\nz.mem_4474_sv2v_reg ,\nz.mem_4473_sv2v_reg ,
  \nz.mem_4472_sv2v_reg ,\nz.mem_4471_sv2v_reg ,\nz.mem_4470_sv2v_reg ,\nz.mem_4469_sv2v_reg ,
  \nz.mem_4468_sv2v_reg ,\nz.mem_4467_sv2v_reg ,\nz.mem_4466_sv2v_reg ,
  \nz.mem_4465_sv2v_reg ,\nz.mem_4464_sv2v_reg ,\nz.mem_4463_sv2v_reg ,\nz.mem_4462_sv2v_reg ,
  \nz.mem_4461_sv2v_reg ,\nz.mem_4460_sv2v_reg ,\nz.mem_4459_sv2v_reg ,
  \nz.mem_4458_sv2v_reg ,\nz.mem_4457_sv2v_reg ,\nz.mem_4456_sv2v_reg ,\nz.mem_4455_sv2v_reg ,
  \nz.mem_4454_sv2v_reg ,\nz.mem_4453_sv2v_reg ,\nz.mem_4452_sv2v_reg ,
  \nz.mem_4451_sv2v_reg ,\nz.mem_4450_sv2v_reg ,\nz.mem_4449_sv2v_reg ,\nz.mem_4448_sv2v_reg ,
  \nz.mem_4447_sv2v_reg ,\nz.mem_4446_sv2v_reg ,\nz.mem_4445_sv2v_reg ,
  \nz.mem_4444_sv2v_reg ,\nz.mem_4443_sv2v_reg ,\nz.mem_4442_sv2v_reg ,\nz.mem_4441_sv2v_reg ,
  \nz.mem_4440_sv2v_reg ,\nz.mem_4439_sv2v_reg ,\nz.mem_4438_sv2v_reg ,
  \nz.mem_4437_sv2v_reg ,\nz.mem_4436_sv2v_reg ,\nz.mem_4435_sv2v_reg ,\nz.mem_4434_sv2v_reg ,
  \nz.mem_4433_sv2v_reg ,\nz.mem_4432_sv2v_reg ,\nz.mem_4431_sv2v_reg ,
  \nz.mem_4430_sv2v_reg ,\nz.mem_4429_sv2v_reg ,\nz.mem_4428_sv2v_reg ,\nz.mem_4427_sv2v_reg ,
  \nz.mem_4426_sv2v_reg ,\nz.mem_4425_sv2v_reg ,\nz.mem_4424_sv2v_reg ,
  \nz.mem_4423_sv2v_reg ,\nz.mem_4422_sv2v_reg ,\nz.mem_4421_sv2v_reg ,\nz.mem_4420_sv2v_reg ,
  \nz.mem_4419_sv2v_reg ,\nz.mem_4418_sv2v_reg ,\nz.mem_4417_sv2v_reg ,
  \nz.mem_4416_sv2v_reg ,\nz.mem_4415_sv2v_reg ,\nz.mem_4414_sv2v_reg ,\nz.mem_4413_sv2v_reg ,
  \nz.mem_4412_sv2v_reg ,\nz.mem_4411_sv2v_reg ,\nz.mem_4410_sv2v_reg ,
  \nz.mem_4409_sv2v_reg ,\nz.mem_4408_sv2v_reg ,\nz.mem_4407_sv2v_reg ,\nz.mem_4406_sv2v_reg ,
  \nz.mem_4405_sv2v_reg ,\nz.mem_4404_sv2v_reg ,\nz.mem_4403_sv2v_reg ,
  \nz.mem_4402_sv2v_reg ,\nz.mem_4401_sv2v_reg ,\nz.mem_4400_sv2v_reg ,
  \nz.mem_4399_sv2v_reg ,\nz.mem_4398_sv2v_reg ,\nz.mem_4397_sv2v_reg ,\nz.mem_4396_sv2v_reg ,
  \nz.mem_4395_sv2v_reg ,\nz.mem_4394_sv2v_reg ,\nz.mem_4393_sv2v_reg ,
  \nz.mem_4392_sv2v_reg ,\nz.mem_4391_sv2v_reg ,\nz.mem_4390_sv2v_reg ,\nz.mem_4389_sv2v_reg ,
  \nz.mem_4388_sv2v_reg ,\nz.mem_4387_sv2v_reg ,\nz.mem_4386_sv2v_reg ,
  \nz.mem_4385_sv2v_reg ,\nz.mem_4384_sv2v_reg ,\nz.mem_4383_sv2v_reg ,\nz.mem_4382_sv2v_reg ,
  \nz.mem_4381_sv2v_reg ,\nz.mem_4380_sv2v_reg ,\nz.mem_4379_sv2v_reg ,
  \nz.mem_4378_sv2v_reg ,\nz.mem_4377_sv2v_reg ,\nz.mem_4376_sv2v_reg ,\nz.mem_4375_sv2v_reg ,
  \nz.mem_4374_sv2v_reg ,\nz.mem_4373_sv2v_reg ,\nz.mem_4372_sv2v_reg ,
  \nz.mem_4371_sv2v_reg ,\nz.mem_4370_sv2v_reg ,\nz.mem_4369_sv2v_reg ,\nz.mem_4368_sv2v_reg ,
  \nz.mem_4367_sv2v_reg ,\nz.mem_4366_sv2v_reg ,\nz.mem_4365_sv2v_reg ,
  \nz.mem_4364_sv2v_reg ,\nz.mem_4363_sv2v_reg ,\nz.mem_4362_sv2v_reg ,\nz.mem_4361_sv2v_reg ,
  \nz.mem_4360_sv2v_reg ,\nz.mem_4359_sv2v_reg ,\nz.mem_4358_sv2v_reg ,
  \nz.mem_4357_sv2v_reg ,\nz.mem_4356_sv2v_reg ,\nz.mem_4355_sv2v_reg ,\nz.mem_4354_sv2v_reg ,
  \nz.mem_4353_sv2v_reg ,\nz.mem_4352_sv2v_reg ,\nz.mem_4351_sv2v_reg ,
  \nz.mem_4350_sv2v_reg ,\nz.mem_4349_sv2v_reg ,\nz.mem_4348_sv2v_reg ,\nz.mem_4347_sv2v_reg ,
  \nz.mem_4346_sv2v_reg ,\nz.mem_4345_sv2v_reg ,\nz.mem_4344_sv2v_reg ,
  \nz.mem_4343_sv2v_reg ,\nz.mem_4342_sv2v_reg ,\nz.mem_4341_sv2v_reg ,\nz.mem_4340_sv2v_reg ,
  \nz.mem_4339_sv2v_reg ,\nz.mem_4338_sv2v_reg ,\nz.mem_4337_sv2v_reg ,
  \nz.mem_4336_sv2v_reg ,\nz.mem_4335_sv2v_reg ,\nz.mem_4334_sv2v_reg ,\nz.mem_4333_sv2v_reg ,
  \nz.mem_4332_sv2v_reg ,\nz.mem_4331_sv2v_reg ,\nz.mem_4330_sv2v_reg ,
  \nz.mem_4329_sv2v_reg ,\nz.mem_4328_sv2v_reg ,\nz.mem_4327_sv2v_reg ,\nz.mem_4326_sv2v_reg ,
  \nz.mem_4325_sv2v_reg ,\nz.mem_4324_sv2v_reg ,\nz.mem_4323_sv2v_reg ,
  \nz.mem_4322_sv2v_reg ,\nz.mem_4321_sv2v_reg ,\nz.mem_4320_sv2v_reg ,
  \nz.mem_4319_sv2v_reg ,\nz.mem_4318_sv2v_reg ,\nz.mem_4317_sv2v_reg ,\nz.mem_4316_sv2v_reg ,
  \nz.mem_4315_sv2v_reg ,\nz.mem_4314_sv2v_reg ,\nz.mem_4313_sv2v_reg ,
  \nz.mem_4312_sv2v_reg ,\nz.mem_4311_sv2v_reg ,\nz.mem_4310_sv2v_reg ,\nz.mem_4309_sv2v_reg ,
  \nz.mem_4308_sv2v_reg ,\nz.mem_4307_sv2v_reg ,\nz.mem_4306_sv2v_reg ,
  \nz.mem_4305_sv2v_reg ,\nz.mem_4304_sv2v_reg ,\nz.mem_4303_sv2v_reg ,\nz.mem_4302_sv2v_reg ,
  \nz.mem_4301_sv2v_reg ,\nz.mem_4300_sv2v_reg ,\nz.mem_4299_sv2v_reg ,
  \nz.mem_4298_sv2v_reg ,\nz.mem_4297_sv2v_reg ,\nz.mem_4296_sv2v_reg ,\nz.mem_4295_sv2v_reg ,
  \nz.mem_4294_sv2v_reg ,\nz.mem_4293_sv2v_reg ,\nz.mem_4292_sv2v_reg ,
  \nz.mem_4291_sv2v_reg ,\nz.mem_4290_sv2v_reg ,\nz.mem_4289_sv2v_reg ,\nz.mem_4288_sv2v_reg ,
  \nz.mem_4287_sv2v_reg ,\nz.mem_4286_sv2v_reg ,\nz.mem_4285_sv2v_reg ,
  \nz.mem_4284_sv2v_reg ,\nz.mem_4283_sv2v_reg ,\nz.mem_4282_sv2v_reg ,\nz.mem_4281_sv2v_reg ,
  \nz.mem_4280_sv2v_reg ,\nz.mem_4279_sv2v_reg ,\nz.mem_4278_sv2v_reg ,
  \nz.mem_4277_sv2v_reg ,\nz.mem_4276_sv2v_reg ,\nz.mem_4275_sv2v_reg ,\nz.mem_4274_sv2v_reg ,
  \nz.mem_4273_sv2v_reg ,\nz.mem_4272_sv2v_reg ,\nz.mem_4271_sv2v_reg ,
  \nz.mem_4270_sv2v_reg ,\nz.mem_4269_sv2v_reg ,\nz.mem_4268_sv2v_reg ,\nz.mem_4267_sv2v_reg ,
  \nz.mem_4266_sv2v_reg ,\nz.mem_4265_sv2v_reg ,\nz.mem_4264_sv2v_reg ,
  \nz.mem_4263_sv2v_reg ,\nz.mem_4262_sv2v_reg ,\nz.mem_4261_sv2v_reg ,\nz.mem_4260_sv2v_reg ,
  \nz.mem_4259_sv2v_reg ,\nz.mem_4258_sv2v_reg ,\nz.mem_4257_sv2v_reg ,
  \nz.mem_4256_sv2v_reg ,\nz.mem_4255_sv2v_reg ,\nz.mem_4254_sv2v_reg ,\nz.mem_4253_sv2v_reg ,
  \nz.mem_4252_sv2v_reg ,\nz.mem_4251_sv2v_reg ,\nz.mem_4250_sv2v_reg ,
  \nz.mem_4249_sv2v_reg ,\nz.mem_4248_sv2v_reg ,\nz.mem_4247_sv2v_reg ,\nz.mem_4246_sv2v_reg ,
  \nz.mem_4245_sv2v_reg ,\nz.mem_4244_sv2v_reg ,\nz.mem_4243_sv2v_reg ,
  \nz.mem_4242_sv2v_reg ,\nz.mem_4241_sv2v_reg ,\nz.mem_4240_sv2v_reg ,
  \nz.mem_4239_sv2v_reg ,\nz.mem_4238_sv2v_reg ,\nz.mem_4237_sv2v_reg ,\nz.mem_4236_sv2v_reg ,
  \nz.mem_4235_sv2v_reg ,\nz.mem_4234_sv2v_reg ,\nz.mem_4233_sv2v_reg ,
  \nz.mem_4232_sv2v_reg ,\nz.mem_4231_sv2v_reg ,\nz.mem_4230_sv2v_reg ,\nz.mem_4229_sv2v_reg ,
  \nz.mem_4228_sv2v_reg ,\nz.mem_4227_sv2v_reg ,\nz.mem_4226_sv2v_reg ,
  \nz.mem_4225_sv2v_reg ,\nz.mem_4224_sv2v_reg ,\nz.mem_4223_sv2v_reg ,\nz.mem_4222_sv2v_reg ,
  \nz.mem_4221_sv2v_reg ,\nz.mem_4220_sv2v_reg ,\nz.mem_4219_sv2v_reg ,
  \nz.mem_4218_sv2v_reg ,\nz.mem_4217_sv2v_reg ,\nz.mem_4216_sv2v_reg ,\nz.mem_4215_sv2v_reg ,
  \nz.mem_4214_sv2v_reg ,\nz.mem_4213_sv2v_reg ,\nz.mem_4212_sv2v_reg ,
  \nz.mem_4211_sv2v_reg ,\nz.mem_4210_sv2v_reg ,\nz.mem_4209_sv2v_reg ,\nz.mem_4208_sv2v_reg ,
  \nz.mem_4207_sv2v_reg ,\nz.mem_4206_sv2v_reg ,\nz.mem_4205_sv2v_reg ,
  \nz.mem_4204_sv2v_reg ,\nz.mem_4203_sv2v_reg ,\nz.mem_4202_sv2v_reg ,\nz.mem_4201_sv2v_reg ,
  \nz.mem_4200_sv2v_reg ,\nz.mem_4199_sv2v_reg ,\nz.mem_4198_sv2v_reg ,
  \nz.mem_4197_sv2v_reg ,\nz.mem_4196_sv2v_reg ,\nz.mem_4195_sv2v_reg ,\nz.mem_4194_sv2v_reg ,
  \nz.mem_4193_sv2v_reg ,\nz.mem_4192_sv2v_reg ,\nz.mem_4191_sv2v_reg ,
  \nz.mem_4190_sv2v_reg ,\nz.mem_4189_sv2v_reg ,\nz.mem_4188_sv2v_reg ,\nz.mem_4187_sv2v_reg ,
  \nz.mem_4186_sv2v_reg ,\nz.mem_4185_sv2v_reg ,\nz.mem_4184_sv2v_reg ,
  \nz.mem_4183_sv2v_reg ,\nz.mem_4182_sv2v_reg ,\nz.mem_4181_sv2v_reg ,\nz.mem_4180_sv2v_reg ,
  \nz.mem_4179_sv2v_reg ,\nz.mem_4178_sv2v_reg ,\nz.mem_4177_sv2v_reg ,
  \nz.mem_4176_sv2v_reg ,\nz.mem_4175_sv2v_reg ,\nz.mem_4174_sv2v_reg ,\nz.mem_4173_sv2v_reg ,
  \nz.mem_4172_sv2v_reg ,\nz.mem_4171_sv2v_reg ,\nz.mem_4170_sv2v_reg ,
  \nz.mem_4169_sv2v_reg ,\nz.mem_4168_sv2v_reg ,\nz.mem_4167_sv2v_reg ,\nz.mem_4166_sv2v_reg ,
  \nz.mem_4165_sv2v_reg ,\nz.mem_4164_sv2v_reg ,\nz.mem_4163_sv2v_reg ,
  \nz.mem_4162_sv2v_reg ,\nz.mem_4161_sv2v_reg ,\nz.mem_4160_sv2v_reg ,
  \nz.mem_4159_sv2v_reg ,\nz.mem_4158_sv2v_reg ,\nz.mem_4157_sv2v_reg ,\nz.mem_4156_sv2v_reg ,
  \nz.mem_4155_sv2v_reg ,\nz.mem_4154_sv2v_reg ,\nz.mem_4153_sv2v_reg ,
  \nz.mem_4152_sv2v_reg ,\nz.mem_4151_sv2v_reg ,\nz.mem_4150_sv2v_reg ,\nz.mem_4149_sv2v_reg ,
  \nz.mem_4148_sv2v_reg ,\nz.mem_4147_sv2v_reg ,\nz.mem_4146_sv2v_reg ,
  \nz.mem_4145_sv2v_reg ,\nz.mem_4144_sv2v_reg ,\nz.mem_4143_sv2v_reg ,\nz.mem_4142_sv2v_reg ,
  \nz.mem_4141_sv2v_reg ,\nz.mem_4140_sv2v_reg ,\nz.mem_4139_sv2v_reg ,
  \nz.mem_4138_sv2v_reg ,\nz.mem_4137_sv2v_reg ,\nz.mem_4136_sv2v_reg ,\nz.mem_4135_sv2v_reg ,
  \nz.mem_4134_sv2v_reg ,\nz.mem_4133_sv2v_reg ,\nz.mem_4132_sv2v_reg ,
  \nz.mem_4131_sv2v_reg ,\nz.mem_4130_sv2v_reg ,\nz.mem_4129_sv2v_reg ,\nz.mem_4128_sv2v_reg ,
  \nz.mem_4127_sv2v_reg ,\nz.mem_4126_sv2v_reg ,\nz.mem_4125_sv2v_reg ,
  \nz.mem_4124_sv2v_reg ,\nz.mem_4123_sv2v_reg ,\nz.mem_4122_sv2v_reg ,\nz.mem_4121_sv2v_reg ,
  \nz.mem_4120_sv2v_reg ,\nz.mem_4119_sv2v_reg ,\nz.mem_4118_sv2v_reg ,
  \nz.mem_4117_sv2v_reg ,\nz.mem_4116_sv2v_reg ,\nz.mem_4115_sv2v_reg ,\nz.mem_4114_sv2v_reg ,
  \nz.mem_4113_sv2v_reg ,\nz.mem_4112_sv2v_reg ,\nz.mem_4111_sv2v_reg ,
  \nz.mem_4110_sv2v_reg ,\nz.mem_4109_sv2v_reg ,\nz.mem_4108_sv2v_reg ,\nz.mem_4107_sv2v_reg ,
  \nz.mem_4106_sv2v_reg ,\nz.mem_4105_sv2v_reg ,\nz.mem_4104_sv2v_reg ,
  \nz.mem_4103_sv2v_reg ,\nz.mem_4102_sv2v_reg ,\nz.mem_4101_sv2v_reg ,\nz.mem_4100_sv2v_reg ,
  \nz.mem_4099_sv2v_reg ,\nz.mem_4098_sv2v_reg ,\nz.mem_4097_sv2v_reg ,
  \nz.mem_4096_sv2v_reg ,\nz.mem_4095_sv2v_reg ,\nz.mem_4094_sv2v_reg ,\nz.mem_4093_sv2v_reg ,
  \nz.mem_4092_sv2v_reg ,\nz.mem_4091_sv2v_reg ,\nz.mem_4090_sv2v_reg ,
  \nz.mem_4089_sv2v_reg ,\nz.mem_4088_sv2v_reg ,\nz.mem_4087_sv2v_reg ,\nz.mem_4086_sv2v_reg ,
  \nz.mem_4085_sv2v_reg ,\nz.mem_4084_sv2v_reg ,\nz.mem_4083_sv2v_reg ,
  \nz.mem_4082_sv2v_reg ,\nz.mem_4081_sv2v_reg ,\nz.mem_4080_sv2v_reg ,
  \nz.mem_4079_sv2v_reg ,\nz.mem_4078_sv2v_reg ,\nz.mem_4077_sv2v_reg ,\nz.mem_4076_sv2v_reg ,
  \nz.mem_4075_sv2v_reg ,\nz.mem_4074_sv2v_reg ,\nz.mem_4073_sv2v_reg ,
  \nz.mem_4072_sv2v_reg ,\nz.mem_4071_sv2v_reg ,\nz.mem_4070_sv2v_reg ,\nz.mem_4069_sv2v_reg ,
  \nz.mem_4068_sv2v_reg ,\nz.mem_4067_sv2v_reg ,\nz.mem_4066_sv2v_reg ,
  \nz.mem_4065_sv2v_reg ,\nz.mem_4064_sv2v_reg ,\nz.mem_4063_sv2v_reg ,\nz.mem_4062_sv2v_reg ,
  \nz.mem_4061_sv2v_reg ,\nz.mem_4060_sv2v_reg ,\nz.mem_4059_sv2v_reg ,
  \nz.mem_4058_sv2v_reg ,\nz.mem_4057_sv2v_reg ,\nz.mem_4056_sv2v_reg ,\nz.mem_4055_sv2v_reg ,
  \nz.mem_4054_sv2v_reg ,\nz.mem_4053_sv2v_reg ,\nz.mem_4052_sv2v_reg ,
  \nz.mem_4051_sv2v_reg ,\nz.mem_4050_sv2v_reg ,\nz.mem_4049_sv2v_reg ,\nz.mem_4048_sv2v_reg ,
  \nz.mem_4047_sv2v_reg ,\nz.mem_4046_sv2v_reg ,\nz.mem_4045_sv2v_reg ,
  \nz.mem_4044_sv2v_reg ,\nz.mem_4043_sv2v_reg ,\nz.mem_4042_sv2v_reg ,\nz.mem_4041_sv2v_reg ,
  \nz.mem_4040_sv2v_reg ,\nz.mem_4039_sv2v_reg ,\nz.mem_4038_sv2v_reg ,
  \nz.mem_4037_sv2v_reg ,\nz.mem_4036_sv2v_reg ,\nz.mem_4035_sv2v_reg ,\nz.mem_4034_sv2v_reg ,
  \nz.mem_4033_sv2v_reg ,\nz.mem_4032_sv2v_reg ,\nz.mem_4031_sv2v_reg ,
  \nz.mem_4030_sv2v_reg ,\nz.mem_4029_sv2v_reg ,\nz.mem_4028_sv2v_reg ,\nz.mem_4027_sv2v_reg ,
  \nz.mem_4026_sv2v_reg ,\nz.mem_4025_sv2v_reg ,\nz.mem_4024_sv2v_reg ,
  \nz.mem_4023_sv2v_reg ,\nz.mem_4022_sv2v_reg ,\nz.mem_4021_sv2v_reg ,\nz.mem_4020_sv2v_reg ,
  \nz.mem_4019_sv2v_reg ,\nz.mem_4018_sv2v_reg ,\nz.mem_4017_sv2v_reg ,
  \nz.mem_4016_sv2v_reg ,\nz.mem_4015_sv2v_reg ,\nz.mem_4014_sv2v_reg ,\nz.mem_4013_sv2v_reg ,
  \nz.mem_4012_sv2v_reg ,\nz.mem_4011_sv2v_reg ,\nz.mem_4010_sv2v_reg ,
  \nz.mem_4009_sv2v_reg ,\nz.mem_4008_sv2v_reg ,\nz.mem_4007_sv2v_reg ,\nz.mem_4006_sv2v_reg ,
  \nz.mem_4005_sv2v_reg ,\nz.mem_4004_sv2v_reg ,\nz.mem_4003_sv2v_reg ,
  \nz.mem_4002_sv2v_reg ,\nz.mem_4001_sv2v_reg ,\nz.mem_4000_sv2v_reg ,
  \nz.mem_3999_sv2v_reg ,\nz.mem_3998_sv2v_reg ,\nz.mem_3997_sv2v_reg ,\nz.mem_3996_sv2v_reg ,
  \nz.mem_3995_sv2v_reg ,\nz.mem_3994_sv2v_reg ,\nz.mem_3993_sv2v_reg ,
  \nz.mem_3992_sv2v_reg ,\nz.mem_3991_sv2v_reg ,\nz.mem_3990_sv2v_reg ,\nz.mem_3989_sv2v_reg ,
  \nz.mem_3988_sv2v_reg ,\nz.mem_3987_sv2v_reg ,\nz.mem_3986_sv2v_reg ,
  \nz.mem_3985_sv2v_reg ,\nz.mem_3984_sv2v_reg ,\nz.mem_3983_sv2v_reg ,\nz.mem_3982_sv2v_reg ,
  \nz.mem_3981_sv2v_reg ,\nz.mem_3980_sv2v_reg ,\nz.mem_3979_sv2v_reg ,
  \nz.mem_3978_sv2v_reg ,\nz.mem_3977_sv2v_reg ,\nz.mem_3976_sv2v_reg ,\nz.mem_3975_sv2v_reg ,
  \nz.mem_3974_sv2v_reg ,\nz.mem_3973_sv2v_reg ,\nz.mem_3972_sv2v_reg ,
  \nz.mem_3971_sv2v_reg ,\nz.mem_3970_sv2v_reg ,\nz.mem_3969_sv2v_reg ,\nz.mem_3968_sv2v_reg ,
  \nz.mem_3967_sv2v_reg ,\nz.mem_3966_sv2v_reg ,\nz.mem_3965_sv2v_reg ,
  \nz.mem_3964_sv2v_reg ,\nz.mem_3963_sv2v_reg ,\nz.mem_3962_sv2v_reg ,\nz.mem_3961_sv2v_reg ,
  \nz.mem_3960_sv2v_reg ,\nz.mem_3959_sv2v_reg ,\nz.mem_3958_sv2v_reg ,
  \nz.mem_3957_sv2v_reg ,\nz.mem_3956_sv2v_reg ,\nz.mem_3955_sv2v_reg ,\nz.mem_3954_sv2v_reg ,
  \nz.mem_3953_sv2v_reg ,\nz.mem_3952_sv2v_reg ,\nz.mem_3951_sv2v_reg ,
  \nz.mem_3950_sv2v_reg ,\nz.mem_3949_sv2v_reg ,\nz.mem_3948_sv2v_reg ,\nz.mem_3947_sv2v_reg ,
  \nz.mem_3946_sv2v_reg ,\nz.mem_3945_sv2v_reg ,\nz.mem_3944_sv2v_reg ,
  \nz.mem_3943_sv2v_reg ,\nz.mem_3942_sv2v_reg ,\nz.mem_3941_sv2v_reg ,\nz.mem_3940_sv2v_reg ,
  \nz.mem_3939_sv2v_reg ,\nz.mem_3938_sv2v_reg ,\nz.mem_3937_sv2v_reg ,
  \nz.mem_3936_sv2v_reg ,\nz.mem_3935_sv2v_reg ,\nz.mem_3934_sv2v_reg ,\nz.mem_3933_sv2v_reg ,
  \nz.mem_3932_sv2v_reg ,\nz.mem_3931_sv2v_reg ,\nz.mem_3930_sv2v_reg ,
  \nz.mem_3929_sv2v_reg ,\nz.mem_3928_sv2v_reg ,\nz.mem_3927_sv2v_reg ,\nz.mem_3926_sv2v_reg ,
  \nz.mem_3925_sv2v_reg ,\nz.mem_3924_sv2v_reg ,\nz.mem_3923_sv2v_reg ,
  \nz.mem_3922_sv2v_reg ,\nz.mem_3921_sv2v_reg ,\nz.mem_3920_sv2v_reg ,
  \nz.mem_3919_sv2v_reg ,\nz.mem_3918_sv2v_reg ,\nz.mem_3917_sv2v_reg ,\nz.mem_3916_sv2v_reg ,
  \nz.mem_3915_sv2v_reg ,\nz.mem_3914_sv2v_reg ,\nz.mem_3913_sv2v_reg ,
  \nz.mem_3912_sv2v_reg ,\nz.mem_3911_sv2v_reg ,\nz.mem_3910_sv2v_reg ,\nz.mem_3909_sv2v_reg ,
  \nz.mem_3908_sv2v_reg ,\nz.mem_3907_sv2v_reg ,\nz.mem_3906_sv2v_reg ,
  \nz.mem_3905_sv2v_reg ,\nz.mem_3904_sv2v_reg ,\nz.mem_3903_sv2v_reg ,\nz.mem_3902_sv2v_reg ,
  \nz.mem_3901_sv2v_reg ,\nz.mem_3900_sv2v_reg ,\nz.mem_3899_sv2v_reg ,
  \nz.mem_3898_sv2v_reg ,\nz.mem_3897_sv2v_reg ,\nz.mem_3896_sv2v_reg ,\nz.mem_3895_sv2v_reg ,
  \nz.mem_3894_sv2v_reg ,\nz.mem_3893_sv2v_reg ,\nz.mem_3892_sv2v_reg ,
  \nz.mem_3891_sv2v_reg ,\nz.mem_3890_sv2v_reg ,\nz.mem_3889_sv2v_reg ,\nz.mem_3888_sv2v_reg ,
  \nz.mem_3887_sv2v_reg ,\nz.mem_3886_sv2v_reg ,\nz.mem_3885_sv2v_reg ,
  \nz.mem_3884_sv2v_reg ,\nz.mem_3883_sv2v_reg ,\nz.mem_3882_sv2v_reg ,\nz.mem_3881_sv2v_reg ,
  \nz.mem_3880_sv2v_reg ,\nz.mem_3879_sv2v_reg ,\nz.mem_3878_sv2v_reg ,
  \nz.mem_3877_sv2v_reg ,\nz.mem_3876_sv2v_reg ,\nz.mem_3875_sv2v_reg ,\nz.mem_3874_sv2v_reg ,
  \nz.mem_3873_sv2v_reg ,\nz.mem_3872_sv2v_reg ,\nz.mem_3871_sv2v_reg ,
  \nz.mem_3870_sv2v_reg ,\nz.mem_3869_sv2v_reg ,\nz.mem_3868_sv2v_reg ,\nz.mem_3867_sv2v_reg ,
  \nz.mem_3866_sv2v_reg ,\nz.mem_3865_sv2v_reg ,\nz.mem_3864_sv2v_reg ,
  \nz.mem_3863_sv2v_reg ,\nz.mem_3862_sv2v_reg ,\nz.mem_3861_sv2v_reg ,\nz.mem_3860_sv2v_reg ,
  \nz.mem_3859_sv2v_reg ,\nz.mem_3858_sv2v_reg ,\nz.mem_3857_sv2v_reg ,
  \nz.mem_3856_sv2v_reg ,\nz.mem_3855_sv2v_reg ,\nz.mem_3854_sv2v_reg ,\nz.mem_3853_sv2v_reg ,
  \nz.mem_3852_sv2v_reg ,\nz.mem_3851_sv2v_reg ,\nz.mem_3850_sv2v_reg ,
  \nz.mem_3849_sv2v_reg ,\nz.mem_3848_sv2v_reg ,\nz.mem_3847_sv2v_reg ,\nz.mem_3846_sv2v_reg ,
  \nz.mem_3845_sv2v_reg ,\nz.mem_3844_sv2v_reg ,\nz.mem_3843_sv2v_reg ,
  \nz.mem_3842_sv2v_reg ,\nz.mem_3841_sv2v_reg ,\nz.mem_3840_sv2v_reg ,
  \nz.mem_3839_sv2v_reg ,\nz.mem_3838_sv2v_reg ,\nz.mem_3837_sv2v_reg ,\nz.mem_3836_sv2v_reg ,
  \nz.mem_3835_sv2v_reg ,\nz.mem_3834_sv2v_reg ,\nz.mem_3833_sv2v_reg ,
  \nz.mem_3832_sv2v_reg ,\nz.mem_3831_sv2v_reg ,\nz.mem_3830_sv2v_reg ,\nz.mem_3829_sv2v_reg ,
  \nz.mem_3828_sv2v_reg ,\nz.mem_3827_sv2v_reg ,\nz.mem_3826_sv2v_reg ,
  \nz.mem_3825_sv2v_reg ,\nz.mem_3824_sv2v_reg ,\nz.mem_3823_sv2v_reg ,\nz.mem_3822_sv2v_reg ,
  \nz.mem_3821_sv2v_reg ,\nz.mem_3820_sv2v_reg ,\nz.mem_3819_sv2v_reg ,
  \nz.mem_3818_sv2v_reg ,\nz.mem_3817_sv2v_reg ,\nz.mem_3816_sv2v_reg ,\nz.mem_3815_sv2v_reg ,
  \nz.mem_3814_sv2v_reg ,\nz.mem_3813_sv2v_reg ,\nz.mem_3812_sv2v_reg ,
  \nz.mem_3811_sv2v_reg ,\nz.mem_3810_sv2v_reg ,\nz.mem_3809_sv2v_reg ,\nz.mem_3808_sv2v_reg ,
  \nz.mem_3807_sv2v_reg ,\nz.mem_3806_sv2v_reg ,\nz.mem_3805_sv2v_reg ,
  \nz.mem_3804_sv2v_reg ,\nz.mem_3803_sv2v_reg ,\nz.mem_3802_sv2v_reg ,\nz.mem_3801_sv2v_reg ,
  \nz.mem_3800_sv2v_reg ,\nz.mem_3799_sv2v_reg ,\nz.mem_3798_sv2v_reg ,
  \nz.mem_3797_sv2v_reg ,\nz.mem_3796_sv2v_reg ,\nz.mem_3795_sv2v_reg ,\nz.mem_3794_sv2v_reg ,
  \nz.mem_3793_sv2v_reg ,\nz.mem_3792_sv2v_reg ,\nz.mem_3791_sv2v_reg ,
  \nz.mem_3790_sv2v_reg ,\nz.mem_3789_sv2v_reg ,\nz.mem_3788_sv2v_reg ,\nz.mem_3787_sv2v_reg ,
  \nz.mem_3786_sv2v_reg ,\nz.mem_3785_sv2v_reg ,\nz.mem_3784_sv2v_reg ,
  \nz.mem_3783_sv2v_reg ,\nz.mem_3782_sv2v_reg ,\nz.mem_3781_sv2v_reg ,\nz.mem_3780_sv2v_reg ,
  \nz.mem_3779_sv2v_reg ,\nz.mem_3778_sv2v_reg ,\nz.mem_3777_sv2v_reg ,
  \nz.mem_3776_sv2v_reg ,\nz.mem_3775_sv2v_reg ,\nz.mem_3774_sv2v_reg ,\nz.mem_3773_sv2v_reg ,
  \nz.mem_3772_sv2v_reg ,\nz.mem_3771_sv2v_reg ,\nz.mem_3770_sv2v_reg ,
  \nz.mem_3769_sv2v_reg ,\nz.mem_3768_sv2v_reg ,\nz.mem_3767_sv2v_reg ,\nz.mem_3766_sv2v_reg ,
  \nz.mem_3765_sv2v_reg ,\nz.mem_3764_sv2v_reg ,\nz.mem_3763_sv2v_reg ,
  \nz.mem_3762_sv2v_reg ,\nz.mem_3761_sv2v_reg ,\nz.mem_3760_sv2v_reg ,
  \nz.mem_3759_sv2v_reg ,\nz.mem_3758_sv2v_reg ,\nz.mem_3757_sv2v_reg ,\nz.mem_3756_sv2v_reg ,
  \nz.mem_3755_sv2v_reg ,\nz.mem_3754_sv2v_reg ,\nz.mem_3753_sv2v_reg ,
  \nz.mem_3752_sv2v_reg ,\nz.mem_3751_sv2v_reg ,\nz.mem_3750_sv2v_reg ,\nz.mem_3749_sv2v_reg ,
  \nz.mem_3748_sv2v_reg ,\nz.mem_3747_sv2v_reg ,\nz.mem_3746_sv2v_reg ,
  \nz.mem_3745_sv2v_reg ,\nz.mem_3744_sv2v_reg ,\nz.mem_3743_sv2v_reg ,\nz.mem_3742_sv2v_reg ,
  \nz.mem_3741_sv2v_reg ,\nz.mem_3740_sv2v_reg ,\nz.mem_3739_sv2v_reg ,
  \nz.mem_3738_sv2v_reg ,\nz.mem_3737_sv2v_reg ,\nz.mem_3736_sv2v_reg ,\nz.mem_3735_sv2v_reg ,
  \nz.mem_3734_sv2v_reg ,\nz.mem_3733_sv2v_reg ,\nz.mem_3732_sv2v_reg ,
  \nz.mem_3731_sv2v_reg ,\nz.mem_3730_sv2v_reg ,\nz.mem_3729_sv2v_reg ,\nz.mem_3728_sv2v_reg ,
  \nz.mem_3727_sv2v_reg ,\nz.mem_3726_sv2v_reg ,\nz.mem_3725_sv2v_reg ,
  \nz.mem_3724_sv2v_reg ,\nz.mem_3723_sv2v_reg ,\nz.mem_3722_sv2v_reg ,\nz.mem_3721_sv2v_reg ,
  \nz.mem_3720_sv2v_reg ,\nz.mem_3719_sv2v_reg ,\nz.mem_3718_sv2v_reg ,
  \nz.mem_3717_sv2v_reg ,\nz.mem_3716_sv2v_reg ,\nz.mem_3715_sv2v_reg ,\nz.mem_3714_sv2v_reg ,
  \nz.mem_3713_sv2v_reg ,\nz.mem_3712_sv2v_reg ,\nz.mem_3711_sv2v_reg ,
  \nz.mem_3710_sv2v_reg ,\nz.mem_3709_sv2v_reg ,\nz.mem_3708_sv2v_reg ,\nz.mem_3707_sv2v_reg ,
  \nz.mem_3706_sv2v_reg ,\nz.mem_3705_sv2v_reg ,\nz.mem_3704_sv2v_reg ,
  \nz.mem_3703_sv2v_reg ,\nz.mem_3702_sv2v_reg ,\nz.mem_3701_sv2v_reg ,\nz.mem_3700_sv2v_reg ,
  \nz.mem_3699_sv2v_reg ,\nz.mem_3698_sv2v_reg ,\nz.mem_3697_sv2v_reg ,
  \nz.mem_3696_sv2v_reg ,\nz.mem_3695_sv2v_reg ,\nz.mem_3694_sv2v_reg ,\nz.mem_3693_sv2v_reg ,
  \nz.mem_3692_sv2v_reg ,\nz.mem_3691_sv2v_reg ,\nz.mem_3690_sv2v_reg ,
  \nz.mem_3689_sv2v_reg ,\nz.mem_3688_sv2v_reg ,\nz.mem_3687_sv2v_reg ,\nz.mem_3686_sv2v_reg ,
  \nz.mem_3685_sv2v_reg ,\nz.mem_3684_sv2v_reg ,\nz.mem_3683_sv2v_reg ,
  \nz.mem_3682_sv2v_reg ,\nz.mem_3681_sv2v_reg ,\nz.mem_3680_sv2v_reg ,
  \nz.mem_3679_sv2v_reg ,\nz.mem_3678_sv2v_reg ,\nz.mem_3677_sv2v_reg ,\nz.mem_3676_sv2v_reg ,
  \nz.mem_3675_sv2v_reg ,\nz.mem_3674_sv2v_reg ,\nz.mem_3673_sv2v_reg ,
  \nz.mem_3672_sv2v_reg ,\nz.mem_3671_sv2v_reg ,\nz.mem_3670_sv2v_reg ,\nz.mem_3669_sv2v_reg ,
  \nz.mem_3668_sv2v_reg ,\nz.mem_3667_sv2v_reg ,\nz.mem_3666_sv2v_reg ,
  \nz.mem_3665_sv2v_reg ,\nz.mem_3664_sv2v_reg ,\nz.mem_3663_sv2v_reg ,\nz.mem_3662_sv2v_reg ,
  \nz.mem_3661_sv2v_reg ,\nz.mem_3660_sv2v_reg ,\nz.mem_3659_sv2v_reg ,
  \nz.mem_3658_sv2v_reg ,\nz.mem_3657_sv2v_reg ,\nz.mem_3656_sv2v_reg ,\nz.mem_3655_sv2v_reg ,
  \nz.mem_3654_sv2v_reg ,\nz.mem_3653_sv2v_reg ,\nz.mem_3652_sv2v_reg ,
  \nz.mem_3651_sv2v_reg ,\nz.mem_3650_sv2v_reg ,\nz.mem_3649_sv2v_reg ,\nz.mem_3648_sv2v_reg ,
  \nz.mem_3647_sv2v_reg ,\nz.mem_3646_sv2v_reg ,\nz.mem_3645_sv2v_reg ,
  \nz.mem_3644_sv2v_reg ,\nz.mem_3643_sv2v_reg ,\nz.mem_3642_sv2v_reg ,\nz.mem_3641_sv2v_reg ,
  \nz.mem_3640_sv2v_reg ,\nz.mem_3639_sv2v_reg ,\nz.mem_3638_sv2v_reg ,
  \nz.mem_3637_sv2v_reg ,\nz.mem_3636_sv2v_reg ,\nz.mem_3635_sv2v_reg ,\nz.mem_3634_sv2v_reg ,
  \nz.mem_3633_sv2v_reg ,\nz.mem_3632_sv2v_reg ,\nz.mem_3631_sv2v_reg ,
  \nz.mem_3630_sv2v_reg ,\nz.mem_3629_sv2v_reg ,\nz.mem_3628_sv2v_reg ,\nz.mem_3627_sv2v_reg ,
  \nz.mem_3626_sv2v_reg ,\nz.mem_3625_sv2v_reg ,\nz.mem_3624_sv2v_reg ,
  \nz.mem_3623_sv2v_reg ,\nz.mem_3622_sv2v_reg ,\nz.mem_3621_sv2v_reg ,\nz.mem_3620_sv2v_reg ,
  \nz.mem_3619_sv2v_reg ,\nz.mem_3618_sv2v_reg ,\nz.mem_3617_sv2v_reg ,
  \nz.mem_3616_sv2v_reg ,\nz.mem_3615_sv2v_reg ,\nz.mem_3614_sv2v_reg ,\nz.mem_3613_sv2v_reg ,
  \nz.mem_3612_sv2v_reg ,\nz.mem_3611_sv2v_reg ,\nz.mem_3610_sv2v_reg ,
  \nz.mem_3609_sv2v_reg ,\nz.mem_3608_sv2v_reg ,\nz.mem_3607_sv2v_reg ,\nz.mem_3606_sv2v_reg ,
  \nz.mem_3605_sv2v_reg ,\nz.mem_3604_sv2v_reg ,\nz.mem_3603_sv2v_reg ,
  \nz.mem_3602_sv2v_reg ,\nz.mem_3601_sv2v_reg ,\nz.mem_3600_sv2v_reg ,
  \nz.mem_3599_sv2v_reg ,\nz.mem_3598_sv2v_reg ,\nz.mem_3597_sv2v_reg ,\nz.mem_3596_sv2v_reg ,
  \nz.mem_3595_sv2v_reg ,\nz.mem_3594_sv2v_reg ,\nz.mem_3593_sv2v_reg ,
  \nz.mem_3592_sv2v_reg ,\nz.mem_3591_sv2v_reg ,\nz.mem_3590_sv2v_reg ,\nz.mem_3589_sv2v_reg ,
  \nz.mem_3588_sv2v_reg ,\nz.mem_3587_sv2v_reg ,\nz.mem_3586_sv2v_reg ,
  \nz.mem_3585_sv2v_reg ,\nz.mem_3584_sv2v_reg ,\nz.mem_3583_sv2v_reg ,\nz.mem_3582_sv2v_reg ,
  \nz.mem_3581_sv2v_reg ,\nz.mem_3580_sv2v_reg ,\nz.mem_3579_sv2v_reg ,
  \nz.mem_3578_sv2v_reg ,\nz.mem_3577_sv2v_reg ,\nz.mem_3576_sv2v_reg ,\nz.mem_3575_sv2v_reg ,
  \nz.mem_3574_sv2v_reg ,\nz.mem_3573_sv2v_reg ,\nz.mem_3572_sv2v_reg ,
  \nz.mem_3571_sv2v_reg ,\nz.mem_3570_sv2v_reg ,\nz.mem_3569_sv2v_reg ,\nz.mem_3568_sv2v_reg ,
  \nz.mem_3567_sv2v_reg ,\nz.mem_3566_sv2v_reg ,\nz.mem_3565_sv2v_reg ,
  \nz.mem_3564_sv2v_reg ,\nz.mem_3563_sv2v_reg ,\nz.mem_3562_sv2v_reg ,\nz.mem_3561_sv2v_reg ,
  \nz.mem_3560_sv2v_reg ,\nz.mem_3559_sv2v_reg ,\nz.mem_3558_sv2v_reg ,
  \nz.mem_3557_sv2v_reg ,\nz.mem_3556_sv2v_reg ,\nz.mem_3555_sv2v_reg ,\nz.mem_3554_sv2v_reg ,
  \nz.mem_3553_sv2v_reg ,\nz.mem_3552_sv2v_reg ,\nz.mem_3551_sv2v_reg ,
  \nz.mem_3550_sv2v_reg ,\nz.mem_3549_sv2v_reg ,\nz.mem_3548_sv2v_reg ,\nz.mem_3547_sv2v_reg ,
  \nz.mem_3546_sv2v_reg ,\nz.mem_3545_sv2v_reg ,\nz.mem_3544_sv2v_reg ,
  \nz.mem_3543_sv2v_reg ,\nz.mem_3542_sv2v_reg ,\nz.mem_3541_sv2v_reg ,\nz.mem_3540_sv2v_reg ,
  \nz.mem_3539_sv2v_reg ,\nz.mem_3538_sv2v_reg ,\nz.mem_3537_sv2v_reg ,
  \nz.mem_3536_sv2v_reg ,\nz.mem_3535_sv2v_reg ,\nz.mem_3534_sv2v_reg ,\nz.mem_3533_sv2v_reg ,
  \nz.mem_3532_sv2v_reg ,\nz.mem_3531_sv2v_reg ,\nz.mem_3530_sv2v_reg ,
  \nz.mem_3529_sv2v_reg ,\nz.mem_3528_sv2v_reg ,\nz.mem_3527_sv2v_reg ,\nz.mem_3526_sv2v_reg ,
  \nz.mem_3525_sv2v_reg ,\nz.mem_3524_sv2v_reg ,\nz.mem_3523_sv2v_reg ,
  \nz.mem_3522_sv2v_reg ,\nz.mem_3521_sv2v_reg ,\nz.mem_3520_sv2v_reg ,
  \nz.mem_3519_sv2v_reg ,\nz.mem_3518_sv2v_reg ,\nz.mem_3517_sv2v_reg ,\nz.mem_3516_sv2v_reg ,
  \nz.mem_3515_sv2v_reg ,\nz.mem_3514_sv2v_reg ,\nz.mem_3513_sv2v_reg ,
  \nz.mem_3512_sv2v_reg ,\nz.mem_3511_sv2v_reg ,\nz.mem_3510_sv2v_reg ,\nz.mem_3509_sv2v_reg ,
  \nz.mem_3508_sv2v_reg ,\nz.mem_3507_sv2v_reg ,\nz.mem_3506_sv2v_reg ,
  \nz.mem_3505_sv2v_reg ,\nz.mem_3504_sv2v_reg ,\nz.mem_3503_sv2v_reg ,\nz.mem_3502_sv2v_reg ,
  \nz.mem_3501_sv2v_reg ,\nz.mem_3500_sv2v_reg ,\nz.mem_3499_sv2v_reg ,
  \nz.mem_3498_sv2v_reg ,\nz.mem_3497_sv2v_reg ,\nz.mem_3496_sv2v_reg ,\nz.mem_3495_sv2v_reg ,
  \nz.mem_3494_sv2v_reg ,\nz.mem_3493_sv2v_reg ,\nz.mem_3492_sv2v_reg ,
  \nz.mem_3491_sv2v_reg ,\nz.mem_3490_sv2v_reg ,\nz.mem_3489_sv2v_reg ,\nz.mem_3488_sv2v_reg ,
  \nz.mem_3487_sv2v_reg ,\nz.mem_3486_sv2v_reg ,\nz.mem_3485_sv2v_reg ,
  \nz.mem_3484_sv2v_reg ,\nz.mem_3483_sv2v_reg ,\nz.mem_3482_sv2v_reg ,\nz.mem_3481_sv2v_reg ,
  \nz.mem_3480_sv2v_reg ,\nz.mem_3479_sv2v_reg ,\nz.mem_3478_sv2v_reg ,
  \nz.mem_3477_sv2v_reg ,\nz.mem_3476_sv2v_reg ,\nz.mem_3475_sv2v_reg ,\nz.mem_3474_sv2v_reg ,
  \nz.mem_3473_sv2v_reg ,\nz.mem_3472_sv2v_reg ,\nz.mem_3471_sv2v_reg ,
  \nz.mem_3470_sv2v_reg ,\nz.mem_3469_sv2v_reg ,\nz.mem_3468_sv2v_reg ,\nz.mem_3467_sv2v_reg ,
  \nz.mem_3466_sv2v_reg ,\nz.mem_3465_sv2v_reg ,\nz.mem_3464_sv2v_reg ,
  \nz.mem_3463_sv2v_reg ,\nz.mem_3462_sv2v_reg ,\nz.mem_3461_sv2v_reg ,\nz.mem_3460_sv2v_reg ,
  \nz.mem_3459_sv2v_reg ,\nz.mem_3458_sv2v_reg ,\nz.mem_3457_sv2v_reg ,
  \nz.mem_3456_sv2v_reg ,\nz.mem_3455_sv2v_reg ,\nz.mem_3454_sv2v_reg ,\nz.mem_3453_sv2v_reg ,
  \nz.mem_3452_sv2v_reg ,\nz.mem_3451_sv2v_reg ,\nz.mem_3450_sv2v_reg ,
  \nz.mem_3449_sv2v_reg ,\nz.mem_3448_sv2v_reg ,\nz.mem_3447_sv2v_reg ,\nz.mem_3446_sv2v_reg ,
  \nz.mem_3445_sv2v_reg ,\nz.mem_3444_sv2v_reg ,\nz.mem_3443_sv2v_reg ,
  \nz.mem_3442_sv2v_reg ,\nz.mem_3441_sv2v_reg ,\nz.mem_3440_sv2v_reg ,
  \nz.mem_3439_sv2v_reg ,\nz.mem_3438_sv2v_reg ,\nz.mem_3437_sv2v_reg ,\nz.mem_3436_sv2v_reg ,
  \nz.mem_3435_sv2v_reg ,\nz.mem_3434_sv2v_reg ,\nz.mem_3433_sv2v_reg ,
  \nz.mem_3432_sv2v_reg ,\nz.mem_3431_sv2v_reg ,\nz.mem_3430_sv2v_reg ,\nz.mem_3429_sv2v_reg ,
  \nz.mem_3428_sv2v_reg ,\nz.mem_3427_sv2v_reg ,\nz.mem_3426_sv2v_reg ,
  \nz.mem_3425_sv2v_reg ,\nz.mem_3424_sv2v_reg ,\nz.mem_3423_sv2v_reg ,\nz.mem_3422_sv2v_reg ,
  \nz.mem_3421_sv2v_reg ,\nz.mem_3420_sv2v_reg ,\nz.mem_3419_sv2v_reg ,
  \nz.mem_3418_sv2v_reg ,\nz.mem_3417_sv2v_reg ,\nz.mem_3416_sv2v_reg ,\nz.mem_3415_sv2v_reg ,
  \nz.mem_3414_sv2v_reg ,\nz.mem_3413_sv2v_reg ,\nz.mem_3412_sv2v_reg ,
  \nz.mem_3411_sv2v_reg ,\nz.mem_3410_sv2v_reg ,\nz.mem_3409_sv2v_reg ,\nz.mem_3408_sv2v_reg ,
  \nz.mem_3407_sv2v_reg ,\nz.mem_3406_sv2v_reg ,\nz.mem_3405_sv2v_reg ,
  \nz.mem_3404_sv2v_reg ,\nz.mem_3403_sv2v_reg ,\nz.mem_3402_sv2v_reg ,\nz.mem_3401_sv2v_reg ,
  \nz.mem_3400_sv2v_reg ,\nz.mem_3399_sv2v_reg ,\nz.mem_3398_sv2v_reg ,
  \nz.mem_3397_sv2v_reg ,\nz.mem_3396_sv2v_reg ,\nz.mem_3395_sv2v_reg ,\nz.mem_3394_sv2v_reg ,
  \nz.mem_3393_sv2v_reg ,\nz.mem_3392_sv2v_reg ,\nz.mem_3391_sv2v_reg ,
  \nz.mem_3390_sv2v_reg ,\nz.mem_3389_sv2v_reg ,\nz.mem_3388_sv2v_reg ,\nz.mem_3387_sv2v_reg ,
  \nz.mem_3386_sv2v_reg ,\nz.mem_3385_sv2v_reg ,\nz.mem_3384_sv2v_reg ,
  \nz.mem_3383_sv2v_reg ,\nz.mem_3382_sv2v_reg ,\nz.mem_3381_sv2v_reg ,\nz.mem_3380_sv2v_reg ,
  \nz.mem_3379_sv2v_reg ,\nz.mem_3378_sv2v_reg ,\nz.mem_3377_sv2v_reg ,
  \nz.mem_3376_sv2v_reg ,\nz.mem_3375_sv2v_reg ,\nz.mem_3374_sv2v_reg ,\nz.mem_3373_sv2v_reg ,
  \nz.mem_3372_sv2v_reg ,\nz.mem_3371_sv2v_reg ,\nz.mem_3370_sv2v_reg ,
  \nz.mem_3369_sv2v_reg ,\nz.mem_3368_sv2v_reg ,\nz.mem_3367_sv2v_reg ,\nz.mem_3366_sv2v_reg ,
  \nz.mem_3365_sv2v_reg ,\nz.mem_3364_sv2v_reg ,\nz.mem_3363_sv2v_reg ,
  \nz.mem_3362_sv2v_reg ,\nz.mem_3361_sv2v_reg ,\nz.mem_3360_sv2v_reg ,
  \nz.mem_3359_sv2v_reg ,\nz.mem_3358_sv2v_reg ,\nz.mem_3357_sv2v_reg ,\nz.mem_3356_sv2v_reg ,
  \nz.mem_3355_sv2v_reg ,\nz.mem_3354_sv2v_reg ,\nz.mem_3353_sv2v_reg ,
  \nz.mem_3352_sv2v_reg ,\nz.mem_3351_sv2v_reg ,\nz.mem_3350_sv2v_reg ,\nz.mem_3349_sv2v_reg ,
  \nz.mem_3348_sv2v_reg ,\nz.mem_3347_sv2v_reg ,\nz.mem_3346_sv2v_reg ,
  \nz.mem_3345_sv2v_reg ,\nz.mem_3344_sv2v_reg ,\nz.mem_3343_sv2v_reg ,\nz.mem_3342_sv2v_reg ,
  \nz.mem_3341_sv2v_reg ,\nz.mem_3340_sv2v_reg ,\nz.mem_3339_sv2v_reg ,
  \nz.mem_3338_sv2v_reg ,\nz.mem_3337_sv2v_reg ,\nz.mem_3336_sv2v_reg ,\nz.mem_3335_sv2v_reg ,
  \nz.mem_3334_sv2v_reg ,\nz.mem_3333_sv2v_reg ,\nz.mem_3332_sv2v_reg ,
  \nz.mem_3331_sv2v_reg ,\nz.mem_3330_sv2v_reg ,\nz.mem_3329_sv2v_reg ,\nz.mem_3328_sv2v_reg ,
  \nz.mem_3327_sv2v_reg ,\nz.mem_3326_sv2v_reg ,\nz.mem_3325_sv2v_reg ,
  \nz.mem_3324_sv2v_reg ,\nz.mem_3323_sv2v_reg ,\nz.mem_3322_sv2v_reg ,\nz.mem_3321_sv2v_reg ,
  \nz.mem_3320_sv2v_reg ,\nz.mem_3319_sv2v_reg ,\nz.mem_3318_sv2v_reg ,
  \nz.mem_3317_sv2v_reg ,\nz.mem_3316_sv2v_reg ,\nz.mem_3315_sv2v_reg ,\nz.mem_3314_sv2v_reg ,
  \nz.mem_3313_sv2v_reg ,\nz.mem_3312_sv2v_reg ,\nz.mem_3311_sv2v_reg ,
  \nz.mem_3310_sv2v_reg ,\nz.mem_3309_sv2v_reg ,\nz.mem_3308_sv2v_reg ,\nz.mem_3307_sv2v_reg ,
  \nz.mem_3306_sv2v_reg ,\nz.mem_3305_sv2v_reg ,\nz.mem_3304_sv2v_reg ,
  \nz.mem_3303_sv2v_reg ,\nz.mem_3302_sv2v_reg ,\nz.mem_3301_sv2v_reg ,\nz.mem_3300_sv2v_reg ,
  \nz.mem_3299_sv2v_reg ,\nz.mem_3298_sv2v_reg ,\nz.mem_3297_sv2v_reg ,
  \nz.mem_3296_sv2v_reg ,\nz.mem_3295_sv2v_reg ,\nz.mem_3294_sv2v_reg ,\nz.mem_3293_sv2v_reg ,
  \nz.mem_3292_sv2v_reg ,\nz.mem_3291_sv2v_reg ,\nz.mem_3290_sv2v_reg ,
  \nz.mem_3289_sv2v_reg ,\nz.mem_3288_sv2v_reg ,\nz.mem_3287_sv2v_reg ,\nz.mem_3286_sv2v_reg ,
  \nz.mem_3285_sv2v_reg ,\nz.mem_3284_sv2v_reg ,\nz.mem_3283_sv2v_reg ,
  \nz.mem_3282_sv2v_reg ,\nz.mem_3281_sv2v_reg ,\nz.mem_3280_sv2v_reg ,
  \nz.mem_3279_sv2v_reg ,\nz.mem_3278_sv2v_reg ,\nz.mem_3277_sv2v_reg ,\nz.mem_3276_sv2v_reg ,
  \nz.mem_3275_sv2v_reg ,\nz.mem_3274_sv2v_reg ,\nz.mem_3273_sv2v_reg ,
  \nz.mem_3272_sv2v_reg ,\nz.mem_3271_sv2v_reg ,\nz.mem_3270_sv2v_reg ,\nz.mem_3269_sv2v_reg ,
  \nz.mem_3268_sv2v_reg ,\nz.mem_3267_sv2v_reg ,\nz.mem_3266_sv2v_reg ,
  \nz.mem_3265_sv2v_reg ,\nz.mem_3264_sv2v_reg ,\nz.mem_3263_sv2v_reg ,\nz.mem_3262_sv2v_reg ,
  \nz.mem_3261_sv2v_reg ,\nz.mem_3260_sv2v_reg ,\nz.mem_3259_sv2v_reg ,
  \nz.mem_3258_sv2v_reg ,\nz.mem_3257_sv2v_reg ,\nz.mem_3256_sv2v_reg ,\nz.mem_3255_sv2v_reg ,
  \nz.mem_3254_sv2v_reg ,\nz.mem_3253_sv2v_reg ,\nz.mem_3252_sv2v_reg ,
  \nz.mem_3251_sv2v_reg ,\nz.mem_3250_sv2v_reg ,\nz.mem_3249_sv2v_reg ,\nz.mem_3248_sv2v_reg ,
  \nz.mem_3247_sv2v_reg ,\nz.mem_3246_sv2v_reg ,\nz.mem_3245_sv2v_reg ,
  \nz.mem_3244_sv2v_reg ,\nz.mem_3243_sv2v_reg ,\nz.mem_3242_sv2v_reg ,\nz.mem_3241_sv2v_reg ,
  \nz.mem_3240_sv2v_reg ,\nz.mem_3239_sv2v_reg ,\nz.mem_3238_sv2v_reg ,
  \nz.mem_3237_sv2v_reg ,\nz.mem_3236_sv2v_reg ,\nz.mem_3235_sv2v_reg ,\nz.mem_3234_sv2v_reg ,
  \nz.mem_3233_sv2v_reg ,\nz.mem_3232_sv2v_reg ,\nz.mem_3231_sv2v_reg ,
  \nz.mem_3230_sv2v_reg ,\nz.mem_3229_sv2v_reg ,\nz.mem_3228_sv2v_reg ,\nz.mem_3227_sv2v_reg ,
  \nz.mem_3226_sv2v_reg ,\nz.mem_3225_sv2v_reg ,\nz.mem_3224_sv2v_reg ,
  \nz.mem_3223_sv2v_reg ,\nz.mem_3222_sv2v_reg ,\nz.mem_3221_sv2v_reg ,\nz.mem_3220_sv2v_reg ,
  \nz.mem_3219_sv2v_reg ,\nz.mem_3218_sv2v_reg ,\nz.mem_3217_sv2v_reg ,
  \nz.mem_3216_sv2v_reg ,\nz.mem_3215_sv2v_reg ,\nz.mem_3214_sv2v_reg ,\nz.mem_3213_sv2v_reg ,
  \nz.mem_3212_sv2v_reg ,\nz.mem_3211_sv2v_reg ,\nz.mem_3210_sv2v_reg ,
  \nz.mem_3209_sv2v_reg ,\nz.mem_3208_sv2v_reg ,\nz.mem_3207_sv2v_reg ,\nz.mem_3206_sv2v_reg ,
  \nz.mem_3205_sv2v_reg ,\nz.mem_3204_sv2v_reg ,\nz.mem_3203_sv2v_reg ,
  \nz.mem_3202_sv2v_reg ,\nz.mem_3201_sv2v_reg ,\nz.mem_3200_sv2v_reg ,
  \nz.mem_3199_sv2v_reg ,\nz.mem_3198_sv2v_reg ,\nz.mem_3197_sv2v_reg ,\nz.mem_3196_sv2v_reg ,
  \nz.mem_3195_sv2v_reg ,\nz.mem_3194_sv2v_reg ,\nz.mem_3193_sv2v_reg ,
  \nz.mem_3192_sv2v_reg ,\nz.mem_3191_sv2v_reg ,\nz.mem_3190_sv2v_reg ,\nz.mem_3189_sv2v_reg ,
  \nz.mem_3188_sv2v_reg ,\nz.mem_3187_sv2v_reg ,\nz.mem_3186_sv2v_reg ,
  \nz.mem_3185_sv2v_reg ,\nz.mem_3184_sv2v_reg ,\nz.mem_3183_sv2v_reg ,\nz.mem_3182_sv2v_reg ,
  \nz.mem_3181_sv2v_reg ,\nz.mem_3180_sv2v_reg ,\nz.mem_3179_sv2v_reg ,
  \nz.mem_3178_sv2v_reg ,\nz.mem_3177_sv2v_reg ,\nz.mem_3176_sv2v_reg ,\nz.mem_3175_sv2v_reg ,
  \nz.mem_3174_sv2v_reg ,\nz.mem_3173_sv2v_reg ,\nz.mem_3172_sv2v_reg ,
  \nz.mem_3171_sv2v_reg ,\nz.mem_3170_sv2v_reg ,\nz.mem_3169_sv2v_reg ,\nz.mem_3168_sv2v_reg ,
  \nz.mem_3167_sv2v_reg ,\nz.mem_3166_sv2v_reg ,\nz.mem_3165_sv2v_reg ,
  \nz.mem_3164_sv2v_reg ,\nz.mem_3163_sv2v_reg ,\nz.mem_3162_sv2v_reg ,\nz.mem_3161_sv2v_reg ,
  \nz.mem_3160_sv2v_reg ,\nz.mem_3159_sv2v_reg ,\nz.mem_3158_sv2v_reg ,
  \nz.mem_3157_sv2v_reg ,\nz.mem_3156_sv2v_reg ,\nz.mem_3155_sv2v_reg ,\nz.mem_3154_sv2v_reg ,
  \nz.mem_3153_sv2v_reg ,\nz.mem_3152_sv2v_reg ,\nz.mem_3151_sv2v_reg ,
  \nz.mem_3150_sv2v_reg ,\nz.mem_3149_sv2v_reg ,\nz.mem_3148_sv2v_reg ,\nz.mem_3147_sv2v_reg ,
  \nz.mem_3146_sv2v_reg ,\nz.mem_3145_sv2v_reg ,\nz.mem_3144_sv2v_reg ,
  \nz.mem_3143_sv2v_reg ,\nz.mem_3142_sv2v_reg ,\nz.mem_3141_sv2v_reg ,\nz.mem_3140_sv2v_reg ,
  \nz.mem_3139_sv2v_reg ,\nz.mem_3138_sv2v_reg ,\nz.mem_3137_sv2v_reg ,
  \nz.mem_3136_sv2v_reg ,\nz.mem_3135_sv2v_reg ,\nz.mem_3134_sv2v_reg ,\nz.mem_3133_sv2v_reg ,
  \nz.mem_3132_sv2v_reg ,\nz.mem_3131_sv2v_reg ,\nz.mem_3130_sv2v_reg ,
  \nz.mem_3129_sv2v_reg ,\nz.mem_3128_sv2v_reg ,\nz.mem_3127_sv2v_reg ,\nz.mem_3126_sv2v_reg ,
  \nz.mem_3125_sv2v_reg ,\nz.mem_3124_sv2v_reg ,\nz.mem_3123_sv2v_reg ,
  \nz.mem_3122_sv2v_reg ,\nz.mem_3121_sv2v_reg ,\nz.mem_3120_sv2v_reg ,
  \nz.mem_3119_sv2v_reg ,\nz.mem_3118_sv2v_reg ,\nz.mem_3117_sv2v_reg ,\nz.mem_3116_sv2v_reg ,
  \nz.mem_3115_sv2v_reg ,\nz.mem_3114_sv2v_reg ,\nz.mem_3113_sv2v_reg ,
  \nz.mem_3112_sv2v_reg ,\nz.mem_3111_sv2v_reg ,\nz.mem_3110_sv2v_reg ,\nz.mem_3109_sv2v_reg ,
  \nz.mem_3108_sv2v_reg ,\nz.mem_3107_sv2v_reg ,\nz.mem_3106_sv2v_reg ,
  \nz.mem_3105_sv2v_reg ,\nz.mem_3104_sv2v_reg ,\nz.mem_3103_sv2v_reg ,\nz.mem_3102_sv2v_reg ,
  \nz.mem_3101_sv2v_reg ,\nz.mem_3100_sv2v_reg ,\nz.mem_3099_sv2v_reg ,
  \nz.mem_3098_sv2v_reg ,\nz.mem_3097_sv2v_reg ,\nz.mem_3096_sv2v_reg ,\nz.mem_3095_sv2v_reg ,
  \nz.mem_3094_sv2v_reg ,\nz.mem_3093_sv2v_reg ,\nz.mem_3092_sv2v_reg ,
  \nz.mem_3091_sv2v_reg ,\nz.mem_3090_sv2v_reg ,\nz.mem_3089_sv2v_reg ,\nz.mem_3088_sv2v_reg ,
  \nz.mem_3087_sv2v_reg ,\nz.mem_3086_sv2v_reg ,\nz.mem_3085_sv2v_reg ,
  \nz.mem_3084_sv2v_reg ,\nz.mem_3083_sv2v_reg ,\nz.mem_3082_sv2v_reg ,\nz.mem_3081_sv2v_reg ,
  \nz.mem_3080_sv2v_reg ,\nz.mem_3079_sv2v_reg ,\nz.mem_3078_sv2v_reg ,
  \nz.mem_3077_sv2v_reg ,\nz.mem_3076_sv2v_reg ,\nz.mem_3075_sv2v_reg ,\nz.mem_3074_sv2v_reg ,
  \nz.mem_3073_sv2v_reg ,\nz.mem_3072_sv2v_reg ,\nz.mem_3071_sv2v_reg ,
  \nz.mem_3070_sv2v_reg ,\nz.mem_3069_sv2v_reg ,\nz.mem_3068_sv2v_reg ,\nz.mem_3067_sv2v_reg ,
  \nz.mem_3066_sv2v_reg ,\nz.mem_3065_sv2v_reg ,\nz.mem_3064_sv2v_reg ,
  \nz.mem_3063_sv2v_reg ,\nz.mem_3062_sv2v_reg ,\nz.mem_3061_sv2v_reg ,\nz.mem_3060_sv2v_reg ,
  \nz.mem_3059_sv2v_reg ,\nz.mem_3058_sv2v_reg ,\nz.mem_3057_sv2v_reg ,
  \nz.mem_3056_sv2v_reg ,\nz.mem_3055_sv2v_reg ,\nz.mem_3054_sv2v_reg ,\nz.mem_3053_sv2v_reg ,
  \nz.mem_3052_sv2v_reg ,\nz.mem_3051_sv2v_reg ,\nz.mem_3050_sv2v_reg ,
  \nz.mem_3049_sv2v_reg ,\nz.mem_3048_sv2v_reg ,\nz.mem_3047_sv2v_reg ,\nz.mem_3046_sv2v_reg ,
  \nz.mem_3045_sv2v_reg ,\nz.mem_3044_sv2v_reg ,\nz.mem_3043_sv2v_reg ,
  \nz.mem_3042_sv2v_reg ,\nz.mem_3041_sv2v_reg ,\nz.mem_3040_sv2v_reg ,
  \nz.mem_3039_sv2v_reg ,\nz.mem_3038_sv2v_reg ,\nz.mem_3037_sv2v_reg ,\nz.mem_3036_sv2v_reg ,
  \nz.mem_3035_sv2v_reg ,\nz.mem_3034_sv2v_reg ,\nz.mem_3033_sv2v_reg ,
  \nz.mem_3032_sv2v_reg ,\nz.mem_3031_sv2v_reg ,\nz.mem_3030_sv2v_reg ,\nz.mem_3029_sv2v_reg ,
  \nz.mem_3028_sv2v_reg ,\nz.mem_3027_sv2v_reg ,\nz.mem_3026_sv2v_reg ,
  \nz.mem_3025_sv2v_reg ,\nz.mem_3024_sv2v_reg ,\nz.mem_3023_sv2v_reg ,\nz.mem_3022_sv2v_reg ,
  \nz.mem_3021_sv2v_reg ,\nz.mem_3020_sv2v_reg ,\nz.mem_3019_sv2v_reg ,
  \nz.mem_3018_sv2v_reg ,\nz.mem_3017_sv2v_reg ,\nz.mem_3016_sv2v_reg ,\nz.mem_3015_sv2v_reg ,
  \nz.mem_3014_sv2v_reg ,\nz.mem_3013_sv2v_reg ,\nz.mem_3012_sv2v_reg ,
  \nz.mem_3011_sv2v_reg ,\nz.mem_3010_sv2v_reg ,\nz.mem_3009_sv2v_reg ,\nz.mem_3008_sv2v_reg ,
  \nz.mem_3007_sv2v_reg ,\nz.mem_3006_sv2v_reg ,\nz.mem_3005_sv2v_reg ,
  \nz.mem_3004_sv2v_reg ,\nz.mem_3003_sv2v_reg ,\nz.mem_3002_sv2v_reg ,\nz.mem_3001_sv2v_reg ,
  \nz.mem_3000_sv2v_reg ,\nz.mem_2999_sv2v_reg ,\nz.mem_2998_sv2v_reg ,
  \nz.mem_2997_sv2v_reg ,\nz.mem_2996_sv2v_reg ,\nz.mem_2995_sv2v_reg ,\nz.mem_2994_sv2v_reg ,
  \nz.mem_2993_sv2v_reg ,\nz.mem_2992_sv2v_reg ,\nz.mem_2991_sv2v_reg ,
  \nz.mem_2990_sv2v_reg ,\nz.mem_2989_sv2v_reg ,\nz.mem_2988_sv2v_reg ,\nz.mem_2987_sv2v_reg ,
  \nz.mem_2986_sv2v_reg ,\nz.mem_2985_sv2v_reg ,\nz.mem_2984_sv2v_reg ,
  \nz.mem_2983_sv2v_reg ,\nz.mem_2982_sv2v_reg ,\nz.mem_2981_sv2v_reg ,\nz.mem_2980_sv2v_reg ,
  \nz.mem_2979_sv2v_reg ,\nz.mem_2978_sv2v_reg ,\nz.mem_2977_sv2v_reg ,
  \nz.mem_2976_sv2v_reg ,\nz.mem_2975_sv2v_reg ,\nz.mem_2974_sv2v_reg ,\nz.mem_2973_sv2v_reg ,
  \nz.mem_2972_sv2v_reg ,\nz.mem_2971_sv2v_reg ,\nz.mem_2970_sv2v_reg ,
  \nz.mem_2969_sv2v_reg ,\nz.mem_2968_sv2v_reg ,\nz.mem_2967_sv2v_reg ,\nz.mem_2966_sv2v_reg ,
  \nz.mem_2965_sv2v_reg ,\nz.mem_2964_sv2v_reg ,\nz.mem_2963_sv2v_reg ,
  \nz.mem_2962_sv2v_reg ,\nz.mem_2961_sv2v_reg ,\nz.mem_2960_sv2v_reg ,
  \nz.mem_2959_sv2v_reg ,\nz.mem_2958_sv2v_reg ,\nz.mem_2957_sv2v_reg ,\nz.mem_2956_sv2v_reg ,
  \nz.mem_2955_sv2v_reg ,\nz.mem_2954_sv2v_reg ,\nz.mem_2953_sv2v_reg ,
  \nz.mem_2952_sv2v_reg ,\nz.mem_2951_sv2v_reg ,\nz.mem_2950_sv2v_reg ,\nz.mem_2949_sv2v_reg ,
  \nz.mem_2948_sv2v_reg ,\nz.mem_2947_sv2v_reg ,\nz.mem_2946_sv2v_reg ,
  \nz.mem_2945_sv2v_reg ,\nz.mem_2944_sv2v_reg ,\nz.mem_2943_sv2v_reg ,\nz.mem_2942_sv2v_reg ,
  \nz.mem_2941_sv2v_reg ,\nz.mem_2940_sv2v_reg ,\nz.mem_2939_sv2v_reg ,
  \nz.mem_2938_sv2v_reg ,\nz.mem_2937_sv2v_reg ,\nz.mem_2936_sv2v_reg ,\nz.mem_2935_sv2v_reg ,
  \nz.mem_2934_sv2v_reg ,\nz.mem_2933_sv2v_reg ,\nz.mem_2932_sv2v_reg ,
  \nz.mem_2931_sv2v_reg ,\nz.mem_2930_sv2v_reg ,\nz.mem_2929_sv2v_reg ,\nz.mem_2928_sv2v_reg ,
  \nz.mem_2927_sv2v_reg ,\nz.mem_2926_sv2v_reg ,\nz.mem_2925_sv2v_reg ,
  \nz.mem_2924_sv2v_reg ,\nz.mem_2923_sv2v_reg ,\nz.mem_2922_sv2v_reg ,\nz.mem_2921_sv2v_reg ,
  \nz.mem_2920_sv2v_reg ,\nz.mem_2919_sv2v_reg ,\nz.mem_2918_sv2v_reg ,
  \nz.mem_2917_sv2v_reg ,\nz.mem_2916_sv2v_reg ,\nz.mem_2915_sv2v_reg ,\nz.mem_2914_sv2v_reg ,
  \nz.mem_2913_sv2v_reg ,\nz.mem_2912_sv2v_reg ,\nz.mem_2911_sv2v_reg ,
  \nz.mem_2910_sv2v_reg ,\nz.mem_2909_sv2v_reg ,\nz.mem_2908_sv2v_reg ,\nz.mem_2907_sv2v_reg ,
  \nz.mem_2906_sv2v_reg ,\nz.mem_2905_sv2v_reg ,\nz.mem_2904_sv2v_reg ,
  \nz.mem_2903_sv2v_reg ,\nz.mem_2902_sv2v_reg ,\nz.mem_2901_sv2v_reg ,\nz.mem_2900_sv2v_reg ,
  \nz.mem_2899_sv2v_reg ,\nz.mem_2898_sv2v_reg ,\nz.mem_2897_sv2v_reg ,
  \nz.mem_2896_sv2v_reg ,\nz.mem_2895_sv2v_reg ,\nz.mem_2894_sv2v_reg ,\nz.mem_2893_sv2v_reg ,
  \nz.mem_2892_sv2v_reg ,\nz.mem_2891_sv2v_reg ,\nz.mem_2890_sv2v_reg ,
  \nz.mem_2889_sv2v_reg ,\nz.mem_2888_sv2v_reg ,\nz.mem_2887_sv2v_reg ,\nz.mem_2886_sv2v_reg ,
  \nz.mem_2885_sv2v_reg ,\nz.mem_2884_sv2v_reg ,\nz.mem_2883_sv2v_reg ,
  \nz.mem_2882_sv2v_reg ,\nz.mem_2881_sv2v_reg ,\nz.mem_2880_sv2v_reg ,
  \nz.mem_2879_sv2v_reg ,\nz.mem_2878_sv2v_reg ,\nz.mem_2877_sv2v_reg ,\nz.mem_2876_sv2v_reg ,
  \nz.mem_2875_sv2v_reg ,\nz.mem_2874_sv2v_reg ,\nz.mem_2873_sv2v_reg ,
  \nz.mem_2872_sv2v_reg ,\nz.mem_2871_sv2v_reg ,\nz.mem_2870_sv2v_reg ,\nz.mem_2869_sv2v_reg ,
  \nz.mem_2868_sv2v_reg ,\nz.mem_2867_sv2v_reg ,\nz.mem_2866_sv2v_reg ,
  \nz.mem_2865_sv2v_reg ,\nz.mem_2864_sv2v_reg ,\nz.mem_2863_sv2v_reg ,\nz.mem_2862_sv2v_reg ,
  \nz.mem_2861_sv2v_reg ,\nz.mem_2860_sv2v_reg ,\nz.mem_2859_sv2v_reg ,
  \nz.mem_2858_sv2v_reg ,\nz.mem_2857_sv2v_reg ,\nz.mem_2856_sv2v_reg ,\nz.mem_2855_sv2v_reg ,
  \nz.mem_2854_sv2v_reg ,\nz.mem_2853_sv2v_reg ,\nz.mem_2852_sv2v_reg ,
  \nz.mem_2851_sv2v_reg ,\nz.mem_2850_sv2v_reg ,\nz.mem_2849_sv2v_reg ,\nz.mem_2848_sv2v_reg ,
  \nz.mem_2847_sv2v_reg ,\nz.mem_2846_sv2v_reg ,\nz.mem_2845_sv2v_reg ,
  \nz.mem_2844_sv2v_reg ,\nz.mem_2843_sv2v_reg ,\nz.mem_2842_sv2v_reg ,\nz.mem_2841_sv2v_reg ,
  \nz.mem_2840_sv2v_reg ,\nz.mem_2839_sv2v_reg ,\nz.mem_2838_sv2v_reg ,
  \nz.mem_2837_sv2v_reg ,\nz.mem_2836_sv2v_reg ,\nz.mem_2835_sv2v_reg ,\nz.mem_2834_sv2v_reg ,
  \nz.mem_2833_sv2v_reg ,\nz.mem_2832_sv2v_reg ,\nz.mem_2831_sv2v_reg ,
  \nz.mem_2830_sv2v_reg ,\nz.mem_2829_sv2v_reg ,\nz.mem_2828_sv2v_reg ,\nz.mem_2827_sv2v_reg ,
  \nz.mem_2826_sv2v_reg ,\nz.mem_2825_sv2v_reg ,\nz.mem_2824_sv2v_reg ,
  \nz.mem_2823_sv2v_reg ,\nz.mem_2822_sv2v_reg ,\nz.mem_2821_sv2v_reg ,\nz.mem_2820_sv2v_reg ,
  \nz.mem_2819_sv2v_reg ,\nz.mem_2818_sv2v_reg ,\nz.mem_2817_sv2v_reg ,
  \nz.mem_2816_sv2v_reg ,\nz.mem_2815_sv2v_reg ,\nz.mem_2814_sv2v_reg ,\nz.mem_2813_sv2v_reg ,
  \nz.mem_2812_sv2v_reg ,\nz.mem_2811_sv2v_reg ,\nz.mem_2810_sv2v_reg ,
  \nz.mem_2809_sv2v_reg ,\nz.mem_2808_sv2v_reg ,\nz.mem_2807_sv2v_reg ,\nz.mem_2806_sv2v_reg ,
  \nz.mem_2805_sv2v_reg ,\nz.mem_2804_sv2v_reg ,\nz.mem_2803_sv2v_reg ,
  \nz.mem_2802_sv2v_reg ,\nz.mem_2801_sv2v_reg ,\nz.mem_2800_sv2v_reg ,
  \nz.mem_2799_sv2v_reg ,\nz.mem_2798_sv2v_reg ,\nz.mem_2797_sv2v_reg ,\nz.mem_2796_sv2v_reg ,
  \nz.mem_2795_sv2v_reg ,\nz.mem_2794_sv2v_reg ,\nz.mem_2793_sv2v_reg ,
  \nz.mem_2792_sv2v_reg ,\nz.mem_2791_sv2v_reg ,\nz.mem_2790_sv2v_reg ,\nz.mem_2789_sv2v_reg ,
  \nz.mem_2788_sv2v_reg ,\nz.mem_2787_sv2v_reg ,\nz.mem_2786_sv2v_reg ,
  \nz.mem_2785_sv2v_reg ,\nz.mem_2784_sv2v_reg ,\nz.mem_2783_sv2v_reg ,\nz.mem_2782_sv2v_reg ,
  \nz.mem_2781_sv2v_reg ,\nz.mem_2780_sv2v_reg ,\nz.mem_2779_sv2v_reg ,
  \nz.mem_2778_sv2v_reg ,\nz.mem_2777_sv2v_reg ,\nz.mem_2776_sv2v_reg ,\nz.mem_2775_sv2v_reg ,
  \nz.mem_2774_sv2v_reg ,\nz.mem_2773_sv2v_reg ,\nz.mem_2772_sv2v_reg ,
  \nz.mem_2771_sv2v_reg ,\nz.mem_2770_sv2v_reg ,\nz.mem_2769_sv2v_reg ,\nz.mem_2768_sv2v_reg ,
  \nz.mem_2767_sv2v_reg ,\nz.mem_2766_sv2v_reg ,\nz.mem_2765_sv2v_reg ,
  \nz.mem_2764_sv2v_reg ,\nz.mem_2763_sv2v_reg ,\nz.mem_2762_sv2v_reg ,\nz.mem_2761_sv2v_reg ,
  \nz.mem_2760_sv2v_reg ,\nz.mem_2759_sv2v_reg ,\nz.mem_2758_sv2v_reg ,
  \nz.mem_2757_sv2v_reg ,\nz.mem_2756_sv2v_reg ,\nz.mem_2755_sv2v_reg ,\nz.mem_2754_sv2v_reg ,
  \nz.mem_2753_sv2v_reg ,\nz.mem_2752_sv2v_reg ,\nz.mem_2751_sv2v_reg ,
  \nz.mem_2750_sv2v_reg ,\nz.mem_2749_sv2v_reg ,\nz.mem_2748_sv2v_reg ,\nz.mem_2747_sv2v_reg ,
  \nz.mem_2746_sv2v_reg ,\nz.mem_2745_sv2v_reg ,\nz.mem_2744_sv2v_reg ,
  \nz.mem_2743_sv2v_reg ,\nz.mem_2742_sv2v_reg ,\nz.mem_2741_sv2v_reg ,\nz.mem_2740_sv2v_reg ,
  \nz.mem_2739_sv2v_reg ,\nz.mem_2738_sv2v_reg ,\nz.mem_2737_sv2v_reg ,
  \nz.mem_2736_sv2v_reg ,\nz.mem_2735_sv2v_reg ,\nz.mem_2734_sv2v_reg ,\nz.mem_2733_sv2v_reg ,
  \nz.mem_2732_sv2v_reg ,\nz.mem_2731_sv2v_reg ,\nz.mem_2730_sv2v_reg ,
  \nz.mem_2729_sv2v_reg ,\nz.mem_2728_sv2v_reg ,\nz.mem_2727_sv2v_reg ,\nz.mem_2726_sv2v_reg ,
  \nz.mem_2725_sv2v_reg ,\nz.mem_2724_sv2v_reg ,\nz.mem_2723_sv2v_reg ,
  \nz.mem_2722_sv2v_reg ,\nz.mem_2721_sv2v_reg ,\nz.mem_2720_sv2v_reg ,
  \nz.mem_2719_sv2v_reg ,\nz.mem_2718_sv2v_reg ,\nz.mem_2717_sv2v_reg ,\nz.mem_2716_sv2v_reg ,
  \nz.mem_2715_sv2v_reg ,\nz.mem_2714_sv2v_reg ,\nz.mem_2713_sv2v_reg ,
  \nz.mem_2712_sv2v_reg ,\nz.mem_2711_sv2v_reg ,\nz.mem_2710_sv2v_reg ,\nz.mem_2709_sv2v_reg ,
  \nz.mem_2708_sv2v_reg ,\nz.mem_2707_sv2v_reg ,\nz.mem_2706_sv2v_reg ,
  \nz.mem_2705_sv2v_reg ,\nz.mem_2704_sv2v_reg ,\nz.mem_2703_sv2v_reg ,\nz.mem_2702_sv2v_reg ,
  \nz.mem_2701_sv2v_reg ,\nz.mem_2700_sv2v_reg ,\nz.mem_2699_sv2v_reg ,
  \nz.mem_2698_sv2v_reg ,\nz.mem_2697_sv2v_reg ,\nz.mem_2696_sv2v_reg ,\nz.mem_2695_sv2v_reg ,
  \nz.mem_2694_sv2v_reg ,\nz.mem_2693_sv2v_reg ,\nz.mem_2692_sv2v_reg ,
  \nz.mem_2691_sv2v_reg ,\nz.mem_2690_sv2v_reg ,\nz.mem_2689_sv2v_reg ,\nz.mem_2688_sv2v_reg ,
  \nz.mem_2687_sv2v_reg ,\nz.mem_2686_sv2v_reg ,\nz.mem_2685_sv2v_reg ,
  \nz.mem_2684_sv2v_reg ,\nz.mem_2683_sv2v_reg ,\nz.mem_2682_sv2v_reg ,\nz.mem_2681_sv2v_reg ,
  \nz.mem_2680_sv2v_reg ,\nz.mem_2679_sv2v_reg ,\nz.mem_2678_sv2v_reg ,
  \nz.mem_2677_sv2v_reg ,\nz.mem_2676_sv2v_reg ,\nz.mem_2675_sv2v_reg ,\nz.mem_2674_sv2v_reg ,
  \nz.mem_2673_sv2v_reg ,\nz.mem_2672_sv2v_reg ,\nz.mem_2671_sv2v_reg ,
  \nz.mem_2670_sv2v_reg ,\nz.mem_2669_sv2v_reg ,\nz.mem_2668_sv2v_reg ,\nz.mem_2667_sv2v_reg ,
  \nz.mem_2666_sv2v_reg ,\nz.mem_2665_sv2v_reg ,\nz.mem_2664_sv2v_reg ,
  \nz.mem_2663_sv2v_reg ,\nz.mem_2662_sv2v_reg ,\nz.mem_2661_sv2v_reg ,\nz.mem_2660_sv2v_reg ,
  \nz.mem_2659_sv2v_reg ,\nz.mem_2658_sv2v_reg ,\nz.mem_2657_sv2v_reg ,
  \nz.mem_2656_sv2v_reg ,\nz.mem_2655_sv2v_reg ,\nz.mem_2654_sv2v_reg ,\nz.mem_2653_sv2v_reg ,
  \nz.mem_2652_sv2v_reg ,\nz.mem_2651_sv2v_reg ,\nz.mem_2650_sv2v_reg ,
  \nz.mem_2649_sv2v_reg ,\nz.mem_2648_sv2v_reg ,\nz.mem_2647_sv2v_reg ,\nz.mem_2646_sv2v_reg ,
  \nz.mem_2645_sv2v_reg ,\nz.mem_2644_sv2v_reg ,\nz.mem_2643_sv2v_reg ,
  \nz.mem_2642_sv2v_reg ,\nz.mem_2641_sv2v_reg ,\nz.mem_2640_sv2v_reg ,
  \nz.mem_2639_sv2v_reg ,\nz.mem_2638_sv2v_reg ,\nz.mem_2637_sv2v_reg ,\nz.mem_2636_sv2v_reg ,
  \nz.mem_2635_sv2v_reg ,\nz.mem_2634_sv2v_reg ,\nz.mem_2633_sv2v_reg ,
  \nz.mem_2632_sv2v_reg ,\nz.mem_2631_sv2v_reg ,\nz.mem_2630_sv2v_reg ,\nz.mem_2629_sv2v_reg ,
  \nz.mem_2628_sv2v_reg ,\nz.mem_2627_sv2v_reg ,\nz.mem_2626_sv2v_reg ,
  \nz.mem_2625_sv2v_reg ,\nz.mem_2624_sv2v_reg ,\nz.mem_2623_sv2v_reg ,\nz.mem_2622_sv2v_reg ,
  \nz.mem_2621_sv2v_reg ,\nz.mem_2620_sv2v_reg ,\nz.mem_2619_sv2v_reg ,
  \nz.mem_2618_sv2v_reg ,\nz.mem_2617_sv2v_reg ,\nz.mem_2616_sv2v_reg ,\nz.mem_2615_sv2v_reg ,
  \nz.mem_2614_sv2v_reg ,\nz.mem_2613_sv2v_reg ,\nz.mem_2612_sv2v_reg ,
  \nz.mem_2611_sv2v_reg ,\nz.mem_2610_sv2v_reg ,\nz.mem_2609_sv2v_reg ,\nz.mem_2608_sv2v_reg ,
  \nz.mem_2607_sv2v_reg ,\nz.mem_2606_sv2v_reg ,\nz.mem_2605_sv2v_reg ,
  \nz.mem_2604_sv2v_reg ,\nz.mem_2603_sv2v_reg ,\nz.mem_2602_sv2v_reg ,\nz.mem_2601_sv2v_reg ,
  \nz.mem_2600_sv2v_reg ,\nz.mem_2599_sv2v_reg ,\nz.mem_2598_sv2v_reg ,
  \nz.mem_2597_sv2v_reg ,\nz.mem_2596_sv2v_reg ,\nz.mem_2595_sv2v_reg ,\nz.mem_2594_sv2v_reg ,
  \nz.mem_2593_sv2v_reg ,\nz.mem_2592_sv2v_reg ,\nz.mem_2591_sv2v_reg ,
  \nz.mem_2590_sv2v_reg ,\nz.mem_2589_sv2v_reg ,\nz.mem_2588_sv2v_reg ,\nz.mem_2587_sv2v_reg ,
  \nz.mem_2586_sv2v_reg ,\nz.mem_2585_sv2v_reg ,\nz.mem_2584_sv2v_reg ,
  \nz.mem_2583_sv2v_reg ,\nz.mem_2582_sv2v_reg ,\nz.mem_2581_sv2v_reg ,\nz.mem_2580_sv2v_reg ,
  \nz.mem_2579_sv2v_reg ,\nz.mem_2578_sv2v_reg ,\nz.mem_2577_sv2v_reg ,
  \nz.mem_2576_sv2v_reg ,\nz.mem_2575_sv2v_reg ,\nz.mem_2574_sv2v_reg ,\nz.mem_2573_sv2v_reg ,
  \nz.mem_2572_sv2v_reg ,\nz.mem_2571_sv2v_reg ,\nz.mem_2570_sv2v_reg ,
  \nz.mem_2569_sv2v_reg ,\nz.mem_2568_sv2v_reg ,\nz.mem_2567_sv2v_reg ,\nz.mem_2566_sv2v_reg ,
  \nz.mem_2565_sv2v_reg ,\nz.mem_2564_sv2v_reg ,\nz.mem_2563_sv2v_reg ,
  \nz.mem_2562_sv2v_reg ,\nz.mem_2561_sv2v_reg ,\nz.mem_2560_sv2v_reg ,
  \nz.mem_2559_sv2v_reg ,\nz.mem_2558_sv2v_reg ,\nz.mem_2557_sv2v_reg ,\nz.mem_2556_sv2v_reg ,
  \nz.mem_2555_sv2v_reg ,\nz.mem_2554_sv2v_reg ,\nz.mem_2553_sv2v_reg ,
  \nz.mem_2552_sv2v_reg ,\nz.mem_2551_sv2v_reg ,\nz.mem_2550_sv2v_reg ,\nz.mem_2549_sv2v_reg ,
  \nz.mem_2548_sv2v_reg ,\nz.mem_2547_sv2v_reg ,\nz.mem_2546_sv2v_reg ,
  \nz.mem_2545_sv2v_reg ,\nz.mem_2544_sv2v_reg ,\nz.mem_2543_sv2v_reg ,\nz.mem_2542_sv2v_reg ,
  \nz.mem_2541_sv2v_reg ,\nz.mem_2540_sv2v_reg ,\nz.mem_2539_sv2v_reg ,
  \nz.mem_2538_sv2v_reg ,\nz.mem_2537_sv2v_reg ,\nz.mem_2536_sv2v_reg ,\nz.mem_2535_sv2v_reg ,
  \nz.mem_2534_sv2v_reg ,\nz.mem_2533_sv2v_reg ,\nz.mem_2532_sv2v_reg ,
  \nz.mem_2531_sv2v_reg ,\nz.mem_2530_sv2v_reg ,\nz.mem_2529_sv2v_reg ,\nz.mem_2528_sv2v_reg ,
  \nz.mem_2527_sv2v_reg ,\nz.mem_2526_sv2v_reg ,\nz.mem_2525_sv2v_reg ,
  \nz.mem_2524_sv2v_reg ,\nz.mem_2523_sv2v_reg ,\nz.mem_2522_sv2v_reg ,\nz.mem_2521_sv2v_reg ,
  \nz.mem_2520_sv2v_reg ,\nz.mem_2519_sv2v_reg ,\nz.mem_2518_sv2v_reg ,
  \nz.mem_2517_sv2v_reg ,\nz.mem_2516_sv2v_reg ,\nz.mem_2515_sv2v_reg ,\nz.mem_2514_sv2v_reg ,
  \nz.mem_2513_sv2v_reg ,\nz.mem_2512_sv2v_reg ,\nz.mem_2511_sv2v_reg ,
  \nz.mem_2510_sv2v_reg ,\nz.mem_2509_sv2v_reg ,\nz.mem_2508_sv2v_reg ,\nz.mem_2507_sv2v_reg ,
  \nz.mem_2506_sv2v_reg ,\nz.mem_2505_sv2v_reg ,\nz.mem_2504_sv2v_reg ,
  \nz.mem_2503_sv2v_reg ,\nz.mem_2502_sv2v_reg ,\nz.mem_2501_sv2v_reg ,\nz.mem_2500_sv2v_reg ,
  \nz.mem_2499_sv2v_reg ,\nz.mem_2498_sv2v_reg ,\nz.mem_2497_sv2v_reg ,
  \nz.mem_2496_sv2v_reg ,\nz.mem_2495_sv2v_reg ,\nz.mem_2494_sv2v_reg ,\nz.mem_2493_sv2v_reg ,
  \nz.mem_2492_sv2v_reg ,\nz.mem_2491_sv2v_reg ,\nz.mem_2490_sv2v_reg ,
  \nz.mem_2489_sv2v_reg ,\nz.mem_2488_sv2v_reg ,\nz.mem_2487_sv2v_reg ,\nz.mem_2486_sv2v_reg ,
  \nz.mem_2485_sv2v_reg ,\nz.mem_2484_sv2v_reg ,\nz.mem_2483_sv2v_reg ,
  \nz.mem_2482_sv2v_reg ,\nz.mem_2481_sv2v_reg ,\nz.mem_2480_sv2v_reg ,
  \nz.mem_2479_sv2v_reg ,\nz.mem_2478_sv2v_reg ,\nz.mem_2477_sv2v_reg ,\nz.mem_2476_sv2v_reg ,
  \nz.mem_2475_sv2v_reg ,\nz.mem_2474_sv2v_reg ,\nz.mem_2473_sv2v_reg ,
  \nz.mem_2472_sv2v_reg ,\nz.mem_2471_sv2v_reg ,\nz.mem_2470_sv2v_reg ,\nz.mem_2469_sv2v_reg ,
  \nz.mem_2468_sv2v_reg ,\nz.mem_2467_sv2v_reg ,\nz.mem_2466_sv2v_reg ,
  \nz.mem_2465_sv2v_reg ,\nz.mem_2464_sv2v_reg ,\nz.mem_2463_sv2v_reg ,\nz.mem_2462_sv2v_reg ,
  \nz.mem_2461_sv2v_reg ,\nz.mem_2460_sv2v_reg ,\nz.mem_2459_sv2v_reg ,
  \nz.mem_2458_sv2v_reg ,\nz.mem_2457_sv2v_reg ,\nz.mem_2456_sv2v_reg ,\nz.mem_2455_sv2v_reg ,
  \nz.mem_2454_sv2v_reg ,\nz.mem_2453_sv2v_reg ,\nz.mem_2452_sv2v_reg ,
  \nz.mem_2451_sv2v_reg ,\nz.mem_2450_sv2v_reg ,\nz.mem_2449_sv2v_reg ,\nz.mem_2448_sv2v_reg ,
  \nz.mem_2447_sv2v_reg ,\nz.mem_2446_sv2v_reg ,\nz.mem_2445_sv2v_reg ,
  \nz.mem_2444_sv2v_reg ,\nz.mem_2443_sv2v_reg ,\nz.mem_2442_sv2v_reg ,\nz.mem_2441_sv2v_reg ,
  \nz.mem_2440_sv2v_reg ,\nz.mem_2439_sv2v_reg ,\nz.mem_2438_sv2v_reg ,
  \nz.mem_2437_sv2v_reg ,\nz.mem_2436_sv2v_reg ,\nz.mem_2435_sv2v_reg ,\nz.mem_2434_sv2v_reg ,
  \nz.mem_2433_sv2v_reg ,\nz.mem_2432_sv2v_reg ,\nz.mem_2431_sv2v_reg ,
  \nz.mem_2430_sv2v_reg ,\nz.mem_2429_sv2v_reg ,\nz.mem_2428_sv2v_reg ,\nz.mem_2427_sv2v_reg ,
  \nz.mem_2426_sv2v_reg ,\nz.mem_2425_sv2v_reg ,\nz.mem_2424_sv2v_reg ,
  \nz.mem_2423_sv2v_reg ,\nz.mem_2422_sv2v_reg ,\nz.mem_2421_sv2v_reg ,\nz.mem_2420_sv2v_reg ,
  \nz.mem_2419_sv2v_reg ,\nz.mem_2418_sv2v_reg ,\nz.mem_2417_sv2v_reg ,
  \nz.mem_2416_sv2v_reg ,\nz.mem_2415_sv2v_reg ,\nz.mem_2414_sv2v_reg ,\nz.mem_2413_sv2v_reg ,
  \nz.mem_2412_sv2v_reg ,\nz.mem_2411_sv2v_reg ,\nz.mem_2410_sv2v_reg ,
  \nz.mem_2409_sv2v_reg ,\nz.mem_2408_sv2v_reg ,\nz.mem_2407_sv2v_reg ,\nz.mem_2406_sv2v_reg ,
  \nz.mem_2405_sv2v_reg ,\nz.mem_2404_sv2v_reg ,\nz.mem_2403_sv2v_reg ,
  \nz.mem_2402_sv2v_reg ,\nz.mem_2401_sv2v_reg ,\nz.mem_2400_sv2v_reg ,
  \nz.mem_2399_sv2v_reg ,\nz.mem_2398_sv2v_reg ,\nz.mem_2397_sv2v_reg ,\nz.mem_2396_sv2v_reg ,
  \nz.mem_2395_sv2v_reg ,\nz.mem_2394_sv2v_reg ,\nz.mem_2393_sv2v_reg ,
  \nz.mem_2392_sv2v_reg ,\nz.mem_2391_sv2v_reg ,\nz.mem_2390_sv2v_reg ,\nz.mem_2389_sv2v_reg ,
  \nz.mem_2388_sv2v_reg ,\nz.mem_2387_sv2v_reg ,\nz.mem_2386_sv2v_reg ,
  \nz.mem_2385_sv2v_reg ,\nz.mem_2384_sv2v_reg ,\nz.mem_2383_sv2v_reg ,\nz.mem_2382_sv2v_reg ,
  \nz.mem_2381_sv2v_reg ,\nz.mem_2380_sv2v_reg ,\nz.mem_2379_sv2v_reg ,
  \nz.mem_2378_sv2v_reg ,\nz.mem_2377_sv2v_reg ,\nz.mem_2376_sv2v_reg ,\nz.mem_2375_sv2v_reg ,
  \nz.mem_2374_sv2v_reg ,\nz.mem_2373_sv2v_reg ,\nz.mem_2372_sv2v_reg ,
  \nz.mem_2371_sv2v_reg ,\nz.mem_2370_sv2v_reg ,\nz.mem_2369_sv2v_reg ,\nz.mem_2368_sv2v_reg ,
  \nz.mem_2367_sv2v_reg ,\nz.mem_2366_sv2v_reg ,\nz.mem_2365_sv2v_reg ,
  \nz.mem_2364_sv2v_reg ,\nz.mem_2363_sv2v_reg ,\nz.mem_2362_sv2v_reg ,\nz.mem_2361_sv2v_reg ,
  \nz.mem_2360_sv2v_reg ,\nz.mem_2359_sv2v_reg ,\nz.mem_2358_sv2v_reg ,
  \nz.mem_2357_sv2v_reg ,\nz.mem_2356_sv2v_reg ,\nz.mem_2355_sv2v_reg ,\nz.mem_2354_sv2v_reg ,
  \nz.mem_2353_sv2v_reg ,\nz.mem_2352_sv2v_reg ,\nz.mem_2351_sv2v_reg ,
  \nz.mem_2350_sv2v_reg ,\nz.mem_2349_sv2v_reg ,\nz.mem_2348_sv2v_reg ,\nz.mem_2347_sv2v_reg ,
  \nz.mem_2346_sv2v_reg ,\nz.mem_2345_sv2v_reg ,\nz.mem_2344_sv2v_reg ,
  \nz.mem_2343_sv2v_reg ,\nz.mem_2342_sv2v_reg ,\nz.mem_2341_sv2v_reg ,\nz.mem_2340_sv2v_reg ,
  \nz.mem_2339_sv2v_reg ,\nz.mem_2338_sv2v_reg ,\nz.mem_2337_sv2v_reg ,
  \nz.mem_2336_sv2v_reg ,\nz.mem_2335_sv2v_reg ,\nz.mem_2334_sv2v_reg ,\nz.mem_2333_sv2v_reg ,
  \nz.mem_2332_sv2v_reg ,\nz.mem_2331_sv2v_reg ,\nz.mem_2330_sv2v_reg ,
  \nz.mem_2329_sv2v_reg ,\nz.mem_2328_sv2v_reg ,\nz.mem_2327_sv2v_reg ,\nz.mem_2326_sv2v_reg ,
  \nz.mem_2325_sv2v_reg ,\nz.mem_2324_sv2v_reg ,\nz.mem_2323_sv2v_reg ,
  \nz.mem_2322_sv2v_reg ,\nz.mem_2321_sv2v_reg ,\nz.mem_2320_sv2v_reg ,
  \nz.mem_2319_sv2v_reg ,\nz.mem_2318_sv2v_reg ,\nz.mem_2317_sv2v_reg ,\nz.mem_2316_sv2v_reg ,
  \nz.mem_2315_sv2v_reg ,\nz.mem_2314_sv2v_reg ,\nz.mem_2313_sv2v_reg ,
  \nz.mem_2312_sv2v_reg ,\nz.mem_2311_sv2v_reg ,\nz.mem_2310_sv2v_reg ,\nz.mem_2309_sv2v_reg ,
  \nz.mem_2308_sv2v_reg ,\nz.mem_2307_sv2v_reg ,\nz.mem_2306_sv2v_reg ,
  \nz.mem_2305_sv2v_reg ,\nz.mem_2304_sv2v_reg ,\nz.mem_2303_sv2v_reg ,\nz.mem_2302_sv2v_reg ,
  \nz.mem_2301_sv2v_reg ,\nz.mem_2300_sv2v_reg ,\nz.mem_2299_sv2v_reg ,
  \nz.mem_2298_sv2v_reg ,\nz.mem_2297_sv2v_reg ,\nz.mem_2296_sv2v_reg ,\nz.mem_2295_sv2v_reg ,
  \nz.mem_2294_sv2v_reg ,\nz.mem_2293_sv2v_reg ,\nz.mem_2292_sv2v_reg ,
  \nz.mem_2291_sv2v_reg ,\nz.mem_2290_sv2v_reg ,\nz.mem_2289_sv2v_reg ,\nz.mem_2288_sv2v_reg ,
  \nz.mem_2287_sv2v_reg ,\nz.mem_2286_sv2v_reg ,\nz.mem_2285_sv2v_reg ,
  \nz.mem_2284_sv2v_reg ,\nz.mem_2283_sv2v_reg ,\nz.mem_2282_sv2v_reg ,\nz.mem_2281_sv2v_reg ,
  \nz.mem_2280_sv2v_reg ,\nz.mem_2279_sv2v_reg ,\nz.mem_2278_sv2v_reg ,
  \nz.mem_2277_sv2v_reg ,\nz.mem_2276_sv2v_reg ,\nz.mem_2275_sv2v_reg ,\nz.mem_2274_sv2v_reg ,
  \nz.mem_2273_sv2v_reg ,\nz.mem_2272_sv2v_reg ,\nz.mem_2271_sv2v_reg ,
  \nz.mem_2270_sv2v_reg ,\nz.mem_2269_sv2v_reg ,\nz.mem_2268_sv2v_reg ,\nz.mem_2267_sv2v_reg ,
  \nz.mem_2266_sv2v_reg ,\nz.mem_2265_sv2v_reg ,\nz.mem_2264_sv2v_reg ,
  \nz.mem_2263_sv2v_reg ,\nz.mem_2262_sv2v_reg ,\nz.mem_2261_sv2v_reg ,\nz.mem_2260_sv2v_reg ,
  \nz.mem_2259_sv2v_reg ,\nz.mem_2258_sv2v_reg ,\nz.mem_2257_sv2v_reg ,
  \nz.mem_2256_sv2v_reg ,\nz.mem_2255_sv2v_reg ,\nz.mem_2254_sv2v_reg ,\nz.mem_2253_sv2v_reg ,
  \nz.mem_2252_sv2v_reg ,\nz.mem_2251_sv2v_reg ,\nz.mem_2250_sv2v_reg ,
  \nz.mem_2249_sv2v_reg ,\nz.mem_2248_sv2v_reg ,\nz.mem_2247_sv2v_reg ,\nz.mem_2246_sv2v_reg ,
  \nz.mem_2245_sv2v_reg ,\nz.mem_2244_sv2v_reg ,\nz.mem_2243_sv2v_reg ,
  \nz.mem_2242_sv2v_reg ,\nz.mem_2241_sv2v_reg ,\nz.mem_2240_sv2v_reg ,
  \nz.mem_2239_sv2v_reg ,\nz.mem_2238_sv2v_reg ,\nz.mem_2237_sv2v_reg ,\nz.mem_2236_sv2v_reg ,
  \nz.mem_2235_sv2v_reg ,\nz.mem_2234_sv2v_reg ,\nz.mem_2233_sv2v_reg ,
  \nz.mem_2232_sv2v_reg ,\nz.mem_2231_sv2v_reg ,\nz.mem_2230_sv2v_reg ,\nz.mem_2229_sv2v_reg ,
  \nz.mem_2228_sv2v_reg ,\nz.mem_2227_sv2v_reg ,\nz.mem_2226_sv2v_reg ,
  \nz.mem_2225_sv2v_reg ,\nz.mem_2224_sv2v_reg ,\nz.mem_2223_sv2v_reg ,\nz.mem_2222_sv2v_reg ,
  \nz.mem_2221_sv2v_reg ,\nz.mem_2220_sv2v_reg ,\nz.mem_2219_sv2v_reg ,
  \nz.mem_2218_sv2v_reg ,\nz.mem_2217_sv2v_reg ,\nz.mem_2216_sv2v_reg ,\nz.mem_2215_sv2v_reg ,
  \nz.mem_2214_sv2v_reg ,\nz.mem_2213_sv2v_reg ,\nz.mem_2212_sv2v_reg ,
  \nz.mem_2211_sv2v_reg ,\nz.mem_2210_sv2v_reg ,\nz.mem_2209_sv2v_reg ,\nz.mem_2208_sv2v_reg ,
  \nz.mem_2207_sv2v_reg ,\nz.mem_2206_sv2v_reg ,\nz.mem_2205_sv2v_reg ,
  \nz.mem_2204_sv2v_reg ,\nz.mem_2203_sv2v_reg ,\nz.mem_2202_sv2v_reg ,\nz.mem_2201_sv2v_reg ,
  \nz.mem_2200_sv2v_reg ,\nz.mem_2199_sv2v_reg ,\nz.mem_2198_sv2v_reg ,
  \nz.mem_2197_sv2v_reg ,\nz.mem_2196_sv2v_reg ,\nz.mem_2195_sv2v_reg ,\nz.mem_2194_sv2v_reg ,
  \nz.mem_2193_sv2v_reg ,\nz.mem_2192_sv2v_reg ,\nz.mem_2191_sv2v_reg ,
  \nz.mem_2190_sv2v_reg ,\nz.mem_2189_sv2v_reg ,\nz.mem_2188_sv2v_reg ,\nz.mem_2187_sv2v_reg ,
  \nz.mem_2186_sv2v_reg ,\nz.mem_2185_sv2v_reg ,\nz.mem_2184_sv2v_reg ,
  \nz.mem_2183_sv2v_reg ,\nz.mem_2182_sv2v_reg ,\nz.mem_2181_sv2v_reg ,\nz.mem_2180_sv2v_reg ,
  \nz.mem_2179_sv2v_reg ,\nz.mem_2178_sv2v_reg ,\nz.mem_2177_sv2v_reg ,
  \nz.mem_2176_sv2v_reg ,\nz.mem_2175_sv2v_reg ,\nz.mem_2174_sv2v_reg ,\nz.mem_2173_sv2v_reg ,
  \nz.mem_2172_sv2v_reg ,\nz.mem_2171_sv2v_reg ,\nz.mem_2170_sv2v_reg ,
  \nz.mem_2169_sv2v_reg ,\nz.mem_2168_sv2v_reg ,\nz.mem_2167_sv2v_reg ,\nz.mem_2166_sv2v_reg ,
  \nz.mem_2165_sv2v_reg ,\nz.mem_2164_sv2v_reg ,\nz.mem_2163_sv2v_reg ,
  \nz.mem_2162_sv2v_reg ,\nz.mem_2161_sv2v_reg ,\nz.mem_2160_sv2v_reg ,
  \nz.mem_2159_sv2v_reg ,\nz.mem_2158_sv2v_reg ,\nz.mem_2157_sv2v_reg ,\nz.mem_2156_sv2v_reg ,
  \nz.mem_2155_sv2v_reg ,\nz.mem_2154_sv2v_reg ,\nz.mem_2153_sv2v_reg ,
  \nz.mem_2152_sv2v_reg ,\nz.mem_2151_sv2v_reg ,\nz.mem_2150_sv2v_reg ,\nz.mem_2149_sv2v_reg ,
  \nz.mem_2148_sv2v_reg ,\nz.mem_2147_sv2v_reg ,\nz.mem_2146_sv2v_reg ,
  \nz.mem_2145_sv2v_reg ,\nz.mem_2144_sv2v_reg ,\nz.mem_2143_sv2v_reg ,\nz.mem_2142_sv2v_reg ,
  \nz.mem_2141_sv2v_reg ,\nz.mem_2140_sv2v_reg ,\nz.mem_2139_sv2v_reg ,
  \nz.mem_2138_sv2v_reg ,\nz.mem_2137_sv2v_reg ,\nz.mem_2136_sv2v_reg ,\nz.mem_2135_sv2v_reg ,
  \nz.mem_2134_sv2v_reg ,\nz.mem_2133_sv2v_reg ,\nz.mem_2132_sv2v_reg ,
  \nz.mem_2131_sv2v_reg ,\nz.mem_2130_sv2v_reg ,\nz.mem_2129_sv2v_reg ,\nz.mem_2128_sv2v_reg ,
  \nz.mem_2127_sv2v_reg ,\nz.mem_2126_sv2v_reg ,\nz.mem_2125_sv2v_reg ,
  \nz.mem_2124_sv2v_reg ,\nz.mem_2123_sv2v_reg ,\nz.mem_2122_sv2v_reg ,\nz.mem_2121_sv2v_reg ,
  \nz.mem_2120_sv2v_reg ,\nz.mem_2119_sv2v_reg ,\nz.mem_2118_sv2v_reg ,
  \nz.mem_2117_sv2v_reg ,\nz.mem_2116_sv2v_reg ,\nz.mem_2115_sv2v_reg ,\nz.mem_2114_sv2v_reg ,
  \nz.mem_2113_sv2v_reg ,\nz.mem_2112_sv2v_reg ,\nz.mem_2111_sv2v_reg ,
  \nz.mem_2110_sv2v_reg ,\nz.mem_2109_sv2v_reg ,\nz.mem_2108_sv2v_reg ,\nz.mem_2107_sv2v_reg ,
  \nz.mem_2106_sv2v_reg ,\nz.mem_2105_sv2v_reg ,\nz.mem_2104_sv2v_reg ,
  \nz.mem_2103_sv2v_reg ,\nz.mem_2102_sv2v_reg ,\nz.mem_2101_sv2v_reg ,\nz.mem_2100_sv2v_reg ,
  \nz.mem_2099_sv2v_reg ,\nz.mem_2098_sv2v_reg ,\nz.mem_2097_sv2v_reg ,
  \nz.mem_2096_sv2v_reg ,\nz.mem_2095_sv2v_reg ,\nz.mem_2094_sv2v_reg ,\nz.mem_2093_sv2v_reg ,
  \nz.mem_2092_sv2v_reg ,\nz.mem_2091_sv2v_reg ,\nz.mem_2090_sv2v_reg ,
  \nz.mem_2089_sv2v_reg ,\nz.mem_2088_sv2v_reg ,\nz.mem_2087_sv2v_reg ,\nz.mem_2086_sv2v_reg ,
  \nz.mem_2085_sv2v_reg ,\nz.mem_2084_sv2v_reg ,\nz.mem_2083_sv2v_reg ,
  \nz.mem_2082_sv2v_reg ,\nz.mem_2081_sv2v_reg ,\nz.mem_2080_sv2v_reg ,
  \nz.mem_2079_sv2v_reg ,\nz.mem_2078_sv2v_reg ,\nz.mem_2077_sv2v_reg ,\nz.mem_2076_sv2v_reg ,
  \nz.mem_2075_sv2v_reg ,\nz.mem_2074_sv2v_reg ,\nz.mem_2073_sv2v_reg ,
  \nz.mem_2072_sv2v_reg ,\nz.mem_2071_sv2v_reg ,\nz.mem_2070_sv2v_reg ,\nz.mem_2069_sv2v_reg ,
  \nz.mem_2068_sv2v_reg ,\nz.mem_2067_sv2v_reg ,\nz.mem_2066_sv2v_reg ,
  \nz.mem_2065_sv2v_reg ,\nz.mem_2064_sv2v_reg ,\nz.mem_2063_sv2v_reg ,\nz.mem_2062_sv2v_reg ,
  \nz.mem_2061_sv2v_reg ,\nz.mem_2060_sv2v_reg ,\nz.mem_2059_sv2v_reg ,
  \nz.mem_2058_sv2v_reg ,\nz.mem_2057_sv2v_reg ,\nz.mem_2056_sv2v_reg ,\nz.mem_2055_sv2v_reg ,
  \nz.mem_2054_sv2v_reg ,\nz.mem_2053_sv2v_reg ,\nz.mem_2052_sv2v_reg ,
  \nz.mem_2051_sv2v_reg ,\nz.mem_2050_sv2v_reg ,\nz.mem_2049_sv2v_reg ,\nz.mem_2048_sv2v_reg ,
  \nz.mem_2047_sv2v_reg ,\nz.mem_2046_sv2v_reg ,\nz.mem_2045_sv2v_reg ,
  \nz.mem_2044_sv2v_reg ,\nz.mem_2043_sv2v_reg ,\nz.mem_2042_sv2v_reg ,\nz.mem_2041_sv2v_reg ,
  \nz.mem_2040_sv2v_reg ,\nz.mem_2039_sv2v_reg ,\nz.mem_2038_sv2v_reg ,
  \nz.mem_2037_sv2v_reg ,\nz.mem_2036_sv2v_reg ,\nz.mem_2035_sv2v_reg ,\nz.mem_2034_sv2v_reg ,
  \nz.mem_2033_sv2v_reg ,\nz.mem_2032_sv2v_reg ,\nz.mem_2031_sv2v_reg ,
  \nz.mem_2030_sv2v_reg ,\nz.mem_2029_sv2v_reg ,\nz.mem_2028_sv2v_reg ,\nz.mem_2027_sv2v_reg ,
  \nz.mem_2026_sv2v_reg ,\nz.mem_2025_sv2v_reg ,\nz.mem_2024_sv2v_reg ,
  \nz.mem_2023_sv2v_reg ,\nz.mem_2022_sv2v_reg ,\nz.mem_2021_sv2v_reg ,\nz.mem_2020_sv2v_reg ,
  \nz.mem_2019_sv2v_reg ,\nz.mem_2018_sv2v_reg ,\nz.mem_2017_sv2v_reg ,
  \nz.mem_2016_sv2v_reg ,\nz.mem_2015_sv2v_reg ,\nz.mem_2014_sv2v_reg ,\nz.mem_2013_sv2v_reg ,
  \nz.mem_2012_sv2v_reg ,\nz.mem_2011_sv2v_reg ,\nz.mem_2010_sv2v_reg ,
  \nz.mem_2009_sv2v_reg ,\nz.mem_2008_sv2v_reg ,\nz.mem_2007_sv2v_reg ,\nz.mem_2006_sv2v_reg ,
  \nz.mem_2005_sv2v_reg ,\nz.mem_2004_sv2v_reg ,\nz.mem_2003_sv2v_reg ,
  \nz.mem_2002_sv2v_reg ,\nz.mem_2001_sv2v_reg ,\nz.mem_2000_sv2v_reg ,
  \nz.mem_1999_sv2v_reg ,\nz.mem_1998_sv2v_reg ,\nz.mem_1997_sv2v_reg ,\nz.mem_1996_sv2v_reg ,
  \nz.mem_1995_sv2v_reg ,\nz.mem_1994_sv2v_reg ,\nz.mem_1993_sv2v_reg ,
  \nz.mem_1992_sv2v_reg ,\nz.mem_1991_sv2v_reg ,\nz.mem_1990_sv2v_reg ,\nz.mem_1989_sv2v_reg ,
  \nz.mem_1988_sv2v_reg ,\nz.mem_1987_sv2v_reg ,\nz.mem_1986_sv2v_reg ,
  \nz.mem_1985_sv2v_reg ,\nz.mem_1984_sv2v_reg ,\nz.mem_1983_sv2v_reg ,\nz.mem_1982_sv2v_reg ,
  \nz.mem_1981_sv2v_reg ,\nz.mem_1980_sv2v_reg ,\nz.mem_1979_sv2v_reg ,
  \nz.mem_1978_sv2v_reg ,\nz.mem_1977_sv2v_reg ,\nz.mem_1976_sv2v_reg ,\nz.mem_1975_sv2v_reg ,
  \nz.mem_1974_sv2v_reg ,\nz.mem_1973_sv2v_reg ,\nz.mem_1972_sv2v_reg ,
  \nz.mem_1971_sv2v_reg ,\nz.mem_1970_sv2v_reg ,\nz.mem_1969_sv2v_reg ,\nz.mem_1968_sv2v_reg ,
  \nz.mem_1967_sv2v_reg ,\nz.mem_1966_sv2v_reg ,\nz.mem_1965_sv2v_reg ,
  \nz.mem_1964_sv2v_reg ,\nz.mem_1963_sv2v_reg ,\nz.mem_1962_sv2v_reg ,\nz.mem_1961_sv2v_reg ,
  \nz.mem_1960_sv2v_reg ,\nz.mem_1959_sv2v_reg ,\nz.mem_1958_sv2v_reg ,
  \nz.mem_1957_sv2v_reg ,\nz.mem_1956_sv2v_reg ,\nz.mem_1955_sv2v_reg ,\nz.mem_1954_sv2v_reg ,
  \nz.mem_1953_sv2v_reg ,\nz.mem_1952_sv2v_reg ,\nz.mem_1951_sv2v_reg ,
  \nz.mem_1950_sv2v_reg ,\nz.mem_1949_sv2v_reg ,\nz.mem_1948_sv2v_reg ,\nz.mem_1947_sv2v_reg ,
  \nz.mem_1946_sv2v_reg ,\nz.mem_1945_sv2v_reg ,\nz.mem_1944_sv2v_reg ,
  \nz.mem_1943_sv2v_reg ,\nz.mem_1942_sv2v_reg ,\nz.mem_1941_sv2v_reg ,\nz.mem_1940_sv2v_reg ,
  \nz.mem_1939_sv2v_reg ,\nz.mem_1938_sv2v_reg ,\nz.mem_1937_sv2v_reg ,
  \nz.mem_1936_sv2v_reg ,\nz.mem_1935_sv2v_reg ,\nz.mem_1934_sv2v_reg ,\nz.mem_1933_sv2v_reg ,
  \nz.mem_1932_sv2v_reg ,\nz.mem_1931_sv2v_reg ,\nz.mem_1930_sv2v_reg ,
  \nz.mem_1929_sv2v_reg ,\nz.mem_1928_sv2v_reg ,\nz.mem_1927_sv2v_reg ,\nz.mem_1926_sv2v_reg ,
  \nz.mem_1925_sv2v_reg ,\nz.mem_1924_sv2v_reg ,\nz.mem_1923_sv2v_reg ,
  \nz.mem_1922_sv2v_reg ,\nz.mem_1921_sv2v_reg ,\nz.mem_1920_sv2v_reg ,
  \nz.mem_1919_sv2v_reg ,\nz.mem_1918_sv2v_reg ,\nz.mem_1917_sv2v_reg ,\nz.mem_1916_sv2v_reg ,
  \nz.mem_1915_sv2v_reg ,\nz.mem_1914_sv2v_reg ,\nz.mem_1913_sv2v_reg ,
  \nz.mem_1912_sv2v_reg ,\nz.mem_1911_sv2v_reg ,\nz.mem_1910_sv2v_reg ,\nz.mem_1909_sv2v_reg ,
  \nz.mem_1908_sv2v_reg ,\nz.mem_1907_sv2v_reg ,\nz.mem_1906_sv2v_reg ,
  \nz.mem_1905_sv2v_reg ,\nz.mem_1904_sv2v_reg ,\nz.mem_1903_sv2v_reg ,\nz.mem_1902_sv2v_reg ,
  \nz.mem_1901_sv2v_reg ,\nz.mem_1900_sv2v_reg ,\nz.mem_1899_sv2v_reg ,
  \nz.mem_1898_sv2v_reg ,\nz.mem_1897_sv2v_reg ,\nz.mem_1896_sv2v_reg ,\nz.mem_1895_sv2v_reg ,
  \nz.mem_1894_sv2v_reg ,\nz.mem_1893_sv2v_reg ,\nz.mem_1892_sv2v_reg ,
  \nz.mem_1891_sv2v_reg ,\nz.mem_1890_sv2v_reg ,\nz.mem_1889_sv2v_reg ,\nz.mem_1888_sv2v_reg ,
  \nz.mem_1887_sv2v_reg ,\nz.mem_1886_sv2v_reg ,\nz.mem_1885_sv2v_reg ,
  \nz.mem_1884_sv2v_reg ,\nz.mem_1883_sv2v_reg ,\nz.mem_1882_sv2v_reg ,\nz.mem_1881_sv2v_reg ,
  \nz.mem_1880_sv2v_reg ,\nz.mem_1879_sv2v_reg ,\nz.mem_1878_sv2v_reg ,
  \nz.mem_1877_sv2v_reg ,\nz.mem_1876_sv2v_reg ,\nz.mem_1875_sv2v_reg ,\nz.mem_1874_sv2v_reg ,
  \nz.mem_1873_sv2v_reg ,\nz.mem_1872_sv2v_reg ,\nz.mem_1871_sv2v_reg ,
  \nz.mem_1870_sv2v_reg ,\nz.mem_1869_sv2v_reg ,\nz.mem_1868_sv2v_reg ,\nz.mem_1867_sv2v_reg ,
  \nz.mem_1866_sv2v_reg ,\nz.mem_1865_sv2v_reg ,\nz.mem_1864_sv2v_reg ,
  \nz.mem_1863_sv2v_reg ,\nz.mem_1862_sv2v_reg ,\nz.mem_1861_sv2v_reg ,\nz.mem_1860_sv2v_reg ,
  \nz.mem_1859_sv2v_reg ,\nz.mem_1858_sv2v_reg ,\nz.mem_1857_sv2v_reg ,
  \nz.mem_1856_sv2v_reg ,\nz.mem_1855_sv2v_reg ,\nz.mem_1854_sv2v_reg ,\nz.mem_1853_sv2v_reg ,
  \nz.mem_1852_sv2v_reg ,\nz.mem_1851_sv2v_reg ,\nz.mem_1850_sv2v_reg ,
  \nz.mem_1849_sv2v_reg ,\nz.mem_1848_sv2v_reg ,\nz.mem_1847_sv2v_reg ,\nz.mem_1846_sv2v_reg ,
  \nz.mem_1845_sv2v_reg ,\nz.mem_1844_sv2v_reg ,\nz.mem_1843_sv2v_reg ,
  \nz.mem_1842_sv2v_reg ,\nz.mem_1841_sv2v_reg ,\nz.mem_1840_sv2v_reg ,
  \nz.mem_1839_sv2v_reg ,\nz.mem_1838_sv2v_reg ,\nz.mem_1837_sv2v_reg ,\nz.mem_1836_sv2v_reg ,
  \nz.mem_1835_sv2v_reg ,\nz.mem_1834_sv2v_reg ,\nz.mem_1833_sv2v_reg ,
  \nz.mem_1832_sv2v_reg ,\nz.mem_1831_sv2v_reg ,\nz.mem_1830_sv2v_reg ,\nz.mem_1829_sv2v_reg ,
  \nz.mem_1828_sv2v_reg ,\nz.mem_1827_sv2v_reg ,\nz.mem_1826_sv2v_reg ,
  \nz.mem_1825_sv2v_reg ,\nz.mem_1824_sv2v_reg ,\nz.mem_1823_sv2v_reg ,\nz.mem_1822_sv2v_reg ,
  \nz.mem_1821_sv2v_reg ,\nz.mem_1820_sv2v_reg ,\nz.mem_1819_sv2v_reg ,
  \nz.mem_1818_sv2v_reg ,\nz.mem_1817_sv2v_reg ,\nz.mem_1816_sv2v_reg ,\nz.mem_1815_sv2v_reg ,
  \nz.mem_1814_sv2v_reg ,\nz.mem_1813_sv2v_reg ,\nz.mem_1812_sv2v_reg ,
  \nz.mem_1811_sv2v_reg ,\nz.mem_1810_sv2v_reg ,\nz.mem_1809_sv2v_reg ,\nz.mem_1808_sv2v_reg ,
  \nz.mem_1807_sv2v_reg ,\nz.mem_1806_sv2v_reg ,\nz.mem_1805_sv2v_reg ,
  \nz.mem_1804_sv2v_reg ,\nz.mem_1803_sv2v_reg ,\nz.mem_1802_sv2v_reg ,\nz.mem_1801_sv2v_reg ,
  \nz.mem_1800_sv2v_reg ,\nz.mem_1799_sv2v_reg ,\nz.mem_1798_sv2v_reg ,
  \nz.mem_1797_sv2v_reg ,\nz.mem_1796_sv2v_reg ,\nz.mem_1795_sv2v_reg ,\nz.mem_1794_sv2v_reg ,
  \nz.mem_1793_sv2v_reg ,\nz.mem_1792_sv2v_reg ,\nz.mem_1791_sv2v_reg ,
  \nz.mem_1790_sv2v_reg ,\nz.mem_1789_sv2v_reg ,\nz.mem_1788_sv2v_reg ,\nz.mem_1787_sv2v_reg ,
  \nz.mem_1786_sv2v_reg ,\nz.mem_1785_sv2v_reg ,\nz.mem_1784_sv2v_reg ,
  \nz.mem_1783_sv2v_reg ,\nz.mem_1782_sv2v_reg ,\nz.mem_1781_sv2v_reg ,\nz.mem_1780_sv2v_reg ,
  \nz.mem_1779_sv2v_reg ,\nz.mem_1778_sv2v_reg ,\nz.mem_1777_sv2v_reg ,
  \nz.mem_1776_sv2v_reg ,\nz.mem_1775_sv2v_reg ,\nz.mem_1774_sv2v_reg ,\nz.mem_1773_sv2v_reg ,
  \nz.mem_1772_sv2v_reg ,\nz.mem_1771_sv2v_reg ,\nz.mem_1770_sv2v_reg ,
  \nz.mem_1769_sv2v_reg ,\nz.mem_1768_sv2v_reg ,\nz.mem_1767_sv2v_reg ,\nz.mem_1766_sv2v_reg ,
  \nz.mem_1765_sv2v_reg ,\nz.mem_1764_sv2v_reg ,\nz.mem_1763_sv2v_reg ,
  \nz.mem_1762_sv2v_reg ,\nz.mem_1761_sv2v_reg ,\nz.mem_1760_sv2v_reg ,
  \nz.mem_1759_sv2v_reg ,\nz.mem_1758_sv2v_reg ,\nz.mem_1757_sv2v_reg ,\nz.mem_1756_sv2v_reg ,
  \nz.mem_1755_sv2v_reg ,\nz.mem_1754_sv2v_reg ,\nz.mem_1753_sv2v_reg ,
  \nz.mem_1752_sv2v_reg ,\nz.mem_1751_sv2v_reg ,\nz.mem_1750_sv2v_reg ,\nz.mem_1749_sv2v_reg ,
  \nz.mem_1748_sv2v_reg ,\nz.mem_1747_sv2v_reg ,\nz.mem_1746_sv2v_reg ,
  \nz.mem_1745_sv2v_reg ,\nz.mem_1744_sv2v_reg ,\nz.mem_1743_sv2v_reg ,\nz.mem_1742_sv2v_reg ,
  \nz.mem_1741_sv2v_reg ,\nz.mem_1740_sv2v_reg ,\nz.mem_1739_sv2v_reg ,
  \nz.mem_1738_sv2v_reg ,\nz.mem_1737_sv2v_reg ,\nz.mem_1736_sv2v_reg ,\nz.mem_1735_sv2v_reg ,
  \nz.mem_1734_sv2v_reg ,\nz.mem_1733_sv2v_reg ,\nz.mem_1732_sv2v_reg ,
  \nz.mem_1731_sv2v_reg ,\nz.mem_1730_sv2v_reg ,\nz.mem_1729_sv2v_reg ,\nz.mem_1728_sv2v_reg ,
  \nz.mem_1727_sv2v_reg ,\nz.mem_1726_sv2v_reg ,\nz.mem_1725_sv2v_reg ,
  \nz.mem_1724_sv2v_reg ,\nz.mem_1723_sv2v_reg ,\nz.mem_1722_sv2v_reg ,\nz.mem_1721_sv2v_reg ,
  \nz.mem_1720_sv2v_reg ,\nz.mem_1719_sv2v_reg ,\nz.mem_1718_sv2v_reg ,
  \nz.mem_1717_sv2v_reg ,\nz.mem_1716_sv2v_reg ,\nz.mem_1715_sv2v_reg ,\nz.mem_1714_sv2v_reg ,
  \nz.mem_1713_sv2v_reg ,\nz.mem_1712_sv2v_reg ,\nz.mem_1711_sv2v_reg ,
  \nz.mem_1710_sv2v_reg ,\nz.mem_1709_sv2v_reg ,\nz.mem_1708_sv2v_reg ,\nz.mem_1707_sv2v_reg ,
  \nz.mem_1706_sv2v_reg ,\nz.mem_1705_sv2v_reg ,\nz.mem_1704_sv2v_reg ,
  \nz.mem_1703_sv2v_reg ,\nz.mem_1702_sv2v_reg ,\nz.mem_1701_sv2v_reg ,\nz.mem_1700_sv2v_reg ,
  \nz.mem_1699_sv2v_reg ,\nz.mem_1698_sv2v_reg ,\nz.mem_1697_sv2v_reg ,
  \nz.mem_1696_sv2v_reg ,\nz.mem_1695_sv2v_reg ,\nz.mem_1694_sv2v_reg ,\nz.mem_1693_sv2v_reg ,
  \nz.mem_1692_sv2v_reg ,\nz.mem_1691_sv2v_reg ,\nz.mem_1690_sv2v_reg ,
  \nz.mem_1689_sv2v_reg ,\nz.mem_1688_sv2v_reg ,\nz.mem_1687_sv2v_reg ,\nz.mem_1686_sv2v_reg ,
  \nz.mem_1685_sv2v_reg ,\nz.mem_1684_sv2v_reg ,\nz.mem_1683_sv2v_reg ,
  \nz.mem_1682_sv2v_reg ,\nz.mem_1681_sv2v_reg ,\nz.mem_1680_sv2v_reg ,
  \nz.mem_1679_sv2v_reg ,\nz.mem_1678_sv2v_reg ,\nz.mem_1677_sv2v_reg ,\nz.mem_1676_sv2v_reg ,
  \nz.mem_1675_sv2v_reg ,\nz.mem_1674_sv2v_reg ,\nz.mem_1673_sv2v_reg ,
  \nz.mem_1672_sv2v_reg ,\nz.mem_1671_sv2v_reg ,\nz.mem_1670_sv2v_reg ,\nz.mem_1669_sv2v_reg ,
  \nz.mem_1668_sv2v_reg ,\nz.mem_1667_sv2v_reg ,\nz.mem_1666_sv2v_reg ,
  \nz.mem_1665_sv2v_reg ,\nz.mem_1664_sv2v_reg ,\nz.mem_1663_sv2v_reg ,\nz.mem_1662_sv2v_reg ,
  \nz.mem_1661_sv2v_reg ,\nz.mem_1660_sv2v_reg ,\nz.mem_1659_sv2v_reg ,
  \nz.mem_1658_sv2v_reg ,\nz.mem_1657_sv2v_reg ,\nz.mem_1656_sv2v_reg ,\nz.mem_1655_sv2v_reg ,
  \nz.mem_1654_sv2v_reg ,\nz.mem_1653_sv2v_reg ,\nz.mem_1652_sv2v_reg ,
  \nz.mem_1651_sv2v_reg ,\nz.mem_1650_sv2v_reg ,\nz.mem_1649_sv2v_reg ,\nz.mem_1648_sv2v_reg ,
  \nz.mem_1647_sv2v_reg ,\nz.mem_1646_sv2v_reg ,\nz.mem_1645_sv2v_reg ,
  \nz.mem_1644_sv2v_reg ,\nz.mem_1643_sv2v_reg ,\nz.mem_1642_sv2v_reg ,\nz.mem_1641_sv2v_reg ,
  \nz.mem_1640_sv2v_reg ,\nz.mem_1639_sv2v_reg ,\nz.mem_1638_sv2v_reg ,
  \nz.mem_1637_sv2v_reg ,\nz.mem_1636_sv2v_reg ,\nz.mem_1635_sv2v_reg ,\nz.mem_1634_sv2v_reg ,
  \nz.mem_1633_sv2v_reg ,\nz.mem_1632_sv2v_reg ,\nz.mem_1631_sv2v_reg ,
  \nz.mem_1630_sv2v_reg ,\nz.mem_1629_sv2v_reg ,\nz.mem_1628_sv2v_reg ,\nz.mem_1627_sv2v_reg ,
  \nz.mem_1626_sv2v_reg ,\nz.mem_1625_sv2v_reg ,\nz.mem_1624_sv2v_reg ,
  \nz.mem_1623_sv2v_reg ,\nz.mem_1622_sv2v_reg ,\nz.mem_1621_sv2v_reg ,\nz.mem_1620_sv2v_reg ,
  \nz.mem_1619_sv2v_reg ,\nz.mem_1618_sv2v_reg ,\nz.mem_1617_sv2v_reg ,
  \nz.mem_1616_sv2v_reg ,\nz.mem_1615_sv2v_reg ,\nz.mem_1614_sv2v_reg ,\nz.mem_1613_sv2v_reg ,
  \nz.mem_1612_sv2v_reg ,\nz.mem_1611_sv2v_reg ,\nz.mem_1610_sv2v_reg ,
  \nz.mem_1609_sv2v_reg ,\nz.mem_1608_sv2v_reg ,\nz.mem_1607_sv2v_reg ,\nz.mem_1606_sv2v_reg ,
  \nz.mem_1605_sv2v_reg ,\nz.mem_1604_sv2v_reg ,\nz.mem_1603_sv2v_reg ,
  \nz.mem_1602_sv2v_reg ,\nz.mem_1601_sv2v_reg ,\nz.mem_1600_sv2v_reg ,
  \nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,\nz.mem_1596_sv2v_reg ,
  \nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,\nz.mem_1593_sv2v_reg ,
  \nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,\nz.mem_1589_sv2v_reg ,
  \nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,\nz.mem_1586_sv2v_reg ,
  \nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,\nz.mem_1582_sv2v_reg ,
  \nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,\nz.mem_1579_sv2v_reg ,
  \nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,\nz.mem_1575_sv2v_reg ,
  \nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,\nz.mem_1572_sv2v_reg ,
  \nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,\nz.mem_1569_sv2v_reg ,\nz.mem_1568_sv2v_reg ,
  \nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,\nz.mem_1565_sv2v_reg ,
  \nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,\nz.mem_1562_sv2v_reg ,\nz.mem_1561_sv2v_reg ,
  \nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,\nz.mem_1558_sv2v_reg ,
  \nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,\nz.mem_1555_sv2v_reg ,\nz.mem_1554_sv2v_reg ,
  \nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,\nz.mem_1551_sv2v_reg ,
  \nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,\nz.mem_1548_sv2v_reg ,\nz.mem_1547_sv2v_reg ,
  \nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,\nz.mem_1544_sv2v_reg ,
  \nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,\nz.mem_1541_sv2v_reg ,\nz.mem_1540_sv2v_reg ,
  \nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,\nz.mem_1537_sv2v_reg ,
  \nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,\nz.mem_1534_sv2v_reg ,\nz.mem_1533_sv2v_reg ,
  \nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,\nz.mem_1530_sv2v_reg ,
  \nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,\nz.mem_1527_sv2v_reg ,\nz.mem_1526_sv2v_reg ,
  \nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,\nz.mem_1523_sv2v_reg ,
  \nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,\nz.mem_1520_sv2v_reg ,
  \nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,\nz.mem_1516_sv2v_reg ,
  \nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,\nz.mem_1513_sv2v_reg ,
  \nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,\nz.mem_1509_sv2v_reg ,
  \nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,\nz.mem_1506_sv2v_reg ,
  \nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,\nz.mem_1502_sv2v_reg ,
  \nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,\nz.mem_1499_sv2v_reg ,
  \nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,\nz.mem_1495_sv2v_reg ,
  \nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,\nz.mem_1492_sv2v_reg ,
  \nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,\nz.mem_1489_sv2v_reg ,\nz.mem_1488_sv2v_reg ,
  \nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,\nz.mem_1485_sv2v_reg ,
  \nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,\nz.mem_1482_sv2v_reg ,\nz.mem_1481_sv2v_reg ,
  \nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,\nz.mem_1478_sv2v_reg ,
  \nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,\nz.mem_1475_sv2v_reg ,\nz.mem_1474_sv2v_reg ,
  \nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,\nz.mem_1471_sv2v_reg ,
  \nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,\nz.mem_1468_sv2v_reg ,\nz.mem_1467_sv2v_reg ,
  \nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,\nz.mem_1464_sv2v_reg ,
  \nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,\nz.mem_1461_sv2v_reg ,\nz.mem_1460_sv2v_reg ,
  \nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,\nz.mem_1457_sv2v_reg ,
  \nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,\nz.mem_1454_sv2v_reg ,\nz.mem_1453_sv2v_reg ,
  \nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,\nz.mem_1450_sv2v_reg ,
  \nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,\nz.mem_1447_sv2v_reg ,\nz.mem_1446_sv2v_reg ,
  \nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,\nz.mem_1443_sv2v_reg ,
  \nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,\nz.mem_1440_sv2v_reg ,
  \nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,\nz.mem_1436_sv2v_reg ,
  \nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,\nz.mem_1433_sv2v_reg ,
  \nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,\nz.mem_1429_sv2v_reg ,
  \nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,\nz.mem_1426_sv2v_reg ,
  \nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,\nz.mem_1422_sv2v_reg ,
  \nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,\nz.mem_1419_sv2v_reg ,
  \nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,\nz.mem_1415_sv2v_reg ,
  \nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,\nz.mem_1412_sv2v_reg ,
  \nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,\nz.mem_1409_sv2v_reg ,\nz.mem_1408_sv2v_reg ,
  \nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,\nz.mem_1405_sv2v_reg ,
  \nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,\nz.mem_1402_sv2v_reg ,\nz.mem_1401_sv2v_reg ,
  \nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,\nz.mem_1398_sv2v_reg ,
  \nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,\nz.mem_1395_sv2v_reg ,\nz.mem_1394_sv2v_reg ,
  \nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,\nz.mem_1391_sv2v_reg ,
  \nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,\nz.mem_1388_sv2v_reg ,\nz.mem_1387_sv2v_reg ,
  \nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,\nz.mem_1384_sv2v_reg ,
  \nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,\nz.mem_1381_sv2v_reg ,\nz.mem_1380_sv2v_reg ,
  \nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,\nz.mem_1377_sv2v_reg ,
  \nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,\nz.mem_1374_sv2v_reg ,\nz.mem_1373_sv2v_reg ,
  \nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,\nz.mem_1370_sv2v_reg ,
  \nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,\nz.mem_1367_sv2v_reg ,\nz.mem_1366_sv2v_reg ,
  \nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,\nz.mem_1363_sv2v_reg ,
  \nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,\nz.mem_1360_sv2v_reg ,
  \nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,\nz.mem_1356_sv2v_reg ,
  \nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,\nz.mem_1353_sv2v_reg ,
  \nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,\nz.mem_1349_sv2v_reg ,
  \nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,\nz.mem_1346_sv2v_reg ,
  \nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,\nz.mem_1342_sv2v_reg ,
  \nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,\nz.mem_1339_sv2v_reg ,
  \nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,\nz.mem_1335_sv2v_reg ,
  \nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,\nz.mem_1332_sv2v_reg ,
  \nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,\nz.mem_1329_sv2v_reg ,\nz.mem_1328_sv2v_reg ,
  \nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,\nz.mem_1325_sv2v_reg ,
  \nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,\nz.mem_1322_sv2v_reg ,\nz.mem_1321_sv2v_reg ,
  \nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,\nz.mem_1318_sv2v_reg ,
  \nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,\nz.mem_1315_sv2v_reg ,\nz.mem_1314_sv2v_reg ,
  \nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,\nz.mem_1311_sv2v_reg ,
  \nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,\nz.mem_1308_sv2v_reg ,\nz.mem_1307_sv2v_reg ,
  \nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,\nz.mem_1304_sv2v_reg ,
  \nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,\nz.mem_1301_sv2v_reg ,\nz.mem_1300_sv2v_reg ,
  \nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,\nz.mem_1297_sv2v_reg ,
  \nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,\nz.mem_1294_sv2v_reg ,\nz.mem_1293_sv2v_reg ,
  \nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,\nz.mem_1290_sv2v_reg ,
  \nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,\nz.mem_1287_sv2v_reg ,\nz.mem_1286_sv2v_reg ,
  \nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,\nz.mem_1283_sv2v_reg ,
  \nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,\nz.mem_1280_sv2v_reg ,
  \nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,\nz.mem_1276_sv2v_reg ,
  \nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,\nz.mem_1273_sv2v_reg ,
  \nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,\nz.mem_1269_sv2v_reg ,
  \nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,\nz.mem_1266_sv2v_reg ,
  \nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,\nz.mem_1262_sv2v_reg ,
  \nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,\nz.mem_1259_sv2v_reg ,
  \nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,\nz.mem_1255_sv2v_reg ,
  \nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,\nz.mem_1252_sv2v_reg ,
  \nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,\nz.mem_1249_sv2v_reg ,\nz.mem_1248_sv2v_reg ,
  \nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,\nz.mem_1245_sv2v_reg ,
  \nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,\nz.mem_1242_sv2v_reg ,\nz.mem_1241_sv2v_reg ,
  \nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,\nz.mem_1238_sv2v_reg ,
  \nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,\nz.mem_1235_sv2v_reg ,\nz.mem_1234_sv2v_reg ,
  \nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,\nz.mem_1231_sv2v_reg ,
  \nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,\nz.mem_1228_sv2v_reg ,\nz.mem_1227_sv2v_reg ,
  \nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,\nz.mem_1224_sv2v_reg ,
  \nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,\nz.mem_1221_sv2v_reg ,\nz.mem_1220_sv2v_reg ,
  \nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,\nz.mem_1217_sv2v_reg ,
  \nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,\nz.mem_1214_sv2v_reg ,\nz.mem_1213_sv2v_reg ,
  \nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,\nz.mem_1210_sv2v_reg ,
  \nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,\nz.mem_1207_sv2v_reg ,\nz.mem_1206_sv2v_reg ,
  \nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,\nz.mem_1203_sv2v_reg ,
  \nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,\nz.mem_1200_sv2v_reg ,
  \nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,\nz.mem_1196_sv2v_reg ,
  \nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,\nz.mem_1193_sv2v_reg ,
  \nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,\nz.mem_1189_sv2v_reg ,
  \nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,\nz.mem_1186_sv2v_reg ,
  \nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,\nz.mem_1182_sv2v_reg ,
  \nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,\nz.mem_1179_sv2v_reg ,
  \nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,\nz.mem_1175_sv2v_reg ,
  \nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,\nz.mem_1172_sv2v_reg ,
  \nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,\nz.mem_1169_sv2v_reg ,\nz.mem_1168_sv2v_reg ,
  \nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,\nz.mem_1165_sv2v_reg ,
  \nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,\nz.mem_1162_sv2v_reg ,\nz.mem_1161_sv2v_reg ,
  \nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,\nz.mem_1158_sv2v_reg ,
  \nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,\nz.mem_1155_sv2v_reg ,\nz.mem_1154_sv2v_reg ,
  \nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,\nz.mem_1151_sv2v_reg ,
  \nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,\nz.mem_1148_sv2v_reg ,\nz.mem_1147_sv2v_reg ,
  \nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,\nz.mem_1144_sv2v_reg ,
  \nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,\nz.mem_1141_sv2v_reg ,\nz.mem_1140_sv2v_reg ,
  \nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,\nz.mem_1137_sv2v_reg ,
  \nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,\nz.mem_1134_sv2v_reg ,\nz.mem_1133_sv2v_reg ,
  \nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,\nz.mem_1130_sv2v_reg ,
  \nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,\nz.mem_1127_sv2v_reg ,\nz.mem_1126_sv2v_reg ,
  \nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,\nz.mem_1123_sv2v_reg ,
  \nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,\nz.mem_1120_sv2v_reg ,
  \nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,\nz.mem_1116_sv2v_reg ,
  \nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,\nz.mem_1113_sv2v_reg ,
  \nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,\nz.mem_1109_sv2v_reg ,
  \nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,\nz.mem_1106_sv2v_reg ,
  \nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,\nz.mem_1102_sv2v_reg ,
  \nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,\nz.mem_1099_sv2v_reg ,
  \nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,\nz.mem_1095_sv2v_reg ,
  \nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,\nz.mem_1092_sv2v_reg ,
  \nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,\nz.mem_1089_sv2v_reg ,\nz.mem_1088_sv2v_reg ,
  \nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,\nz.mem_1085_sv2v_reg ,
  \nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,\nz.mem_1082_sv2v_reg ,\nz.mem_1081_sv2v_reg ,
  \nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,\nz.mem_1078_sv2v_reg ,
  \nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,\nz.mem_1075_sv2v_reg ,\nz.mem_1074_sv2v_reg ,
  \nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,\nz.mem_1071_sv2v_reg ,
  \nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,\nz.mem_1068_sv2v_reg ,\nz.mem_1067_sv2v_reg ,
  \nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,\nz.mem_1064_sv2v_reg ,
  \nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,\nz.mem_1061_sv2v_reg ,\nz.mem_1060_sv2v_reg ,
  \nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,\nz.mem_1057_sv2v_reg ,
  \nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,\nz.mem_1054_sv2v_reg ,\nz.mem_1053_sv2v_reg ,
  \nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,\nz.mem_1050_sv2v_reg ,
  \nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,\nz.mem_1047_sv2v_reg ,\nz.mem_1046_sv2v_reg ,
  \nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,\nz.mem_1043_sv2v_reg ,
  \nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,\nz.mem_1040_sv2v_reg ,
  \nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,\nz.mem_1036_sv2v_reg ,
  \nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,\nz.mem_1033_sv2v_reg ,
  \nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,\nz.mem_1029_sv2v_reg ,
  \nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,\nz.mem_1026_sv2v_reg ,
  \nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,\nz.mem_1022_sv2v_reg ,
  \nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,\nz.mem_1019_sv2v_reg ,
  \nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,\nz.mem_1015_sv2v_reg ,
  \nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,\nz.mem_1012_sv2v_reg ,
  \nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,\nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,
  \nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,\nz.mem_1005_sv2v_reg ,
  \nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,\nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,
  \nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,\nz.mem_998_sv2v_reg ,
  \nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,\nz.mem_994_sv2v_reg ,
  \nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,\nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,
  \nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,\nz.mem_987_sv2v_reg ,
  \nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,\nz.mem_983_sv2v_reg ,
  \nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,\nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,
  \nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,\nz.mem_976_sv2v_reg ,
  \nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,\nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,
  \nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,\nz.mem_969_sv2v_reg ,
  \nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,\nz.mem_965_sv2v_reg ,
  \nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,\nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,
  \nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,\nz.mem_958_sv2v_reg ,
  \nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,\nz.mem_954_sv2v_reg ,
  \nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,\nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,
  \nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,\nz.mem_947_sv2v_reg ,
  \nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,\nz.mem_943_sv2v_reg ,
  \nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,\nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,
  \nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,\nz.mem_936_sv2v_reg ,
  \nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,\nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,
  \nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,\nz.mem_929_sv2v_reg ,
  \nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,\nz.mem_925_sv2v_reg ,
  \nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,\nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,
  \nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,\nz.mem_918_sv2v_reg ,
  \nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,\nz.mem_914_sv2v_reg ,
  \nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,\nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,
  \nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,\nz.mem_907_sv2v_reg ,
  \nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,\nz.mem_903_sv2v_reg ,
  \nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,\nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,
  \nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,\nz.mem_896_sv2v_reg ,
  \nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,\nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,
  \nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,\nz.mem_889_sv2v_reg ,
  \nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,\nz.mem_885_sv2v_reg ,
  \nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,\nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,
  \nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,\nz.mem_878_sv2v_reg ,
  \nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,\nz.mem_874_sv2v_reg ,
  \nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,\nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,
  \nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,\nz.mem_867_sv2v_reg ,
  \nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,\nz.mem_863_sv2v_reg ,
  \nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,\nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,
  \nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,\nz.mem_856_sv2v_reg ,
  \nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,\nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,
  \nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,\nz.mem_849_sv2v_reg ,
  \nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,\nz.mem_845_sv2v_reg ,
  \nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,\nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,
  \nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,\nz.mem_838_sv2v_reg ,
  \nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,\nz.mem_834_sv2v_reg ,
  \nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,\nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,
  \nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,\nz.mem_827_sv2v_reg ,
  \nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,\nz.mem_823_sv2v_reg ,
  \nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,\nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,
  \nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,\nz.mem_816_sv2v_reg ,
  \nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,\nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,
  \nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,\nz.mem_809_sv2v_reg ,
  \nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,\nz.mem_805_sv2v_reg ,
  \nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,\nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,
  \nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,\nz.mem_798_sv2v_reg ,
  \nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,\nz.mem_794_sv2v_reg ,
  \nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,\nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,
  \nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,\nz.mem_787_sv2v_reg ,
  \nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,\nz.mem_783_sv2v_reg ,
  \nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,\nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,
  \nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,\nz.mem_776_sv2v_reg ,
  \nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,\nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,
  \nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,\nz.mem_769_sv2v_reg ,
  \nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,\nz.mem_765_sv2v_reg ,
  \nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,\nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,
  \nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,\nz.mem_758_sv2v_reg ,
  \nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,\nz.mem_754_sv2v_reg ,
  \nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,\nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,
  \nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,\nz.mem_747_sv2v_reg ,
  \nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,\nz.mem_743_sv2v_reg ,
  \nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,\nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,
  \nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,\nz.mem_736_sv2v_reg ,
  \nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,\nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,
  \nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,\nz.mem_729_sv2v_reg ,
  \nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,\nz.mem_725_sv2v_reg ,
  \nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,\nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,
  \nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,\nz.mem_718_sv2v_reg ,
  \nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,\nz.mem_714_sv2v_reg ,
  \nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,\nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,
  \nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,\nz.mem_707_sv2v_reg ,
  \nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,\nz.mem_703_sv2v_reg ,
  \nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,\nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,
  \nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,\nz.mem_696_sv2v_reg ,
  \nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,\nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,
  \nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,\nz.mem_689_sv2v_reg ,
  \nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,\nz.mem_685_sv2v_reg ,
  \nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,
  \nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,\nz.mem_678_sv2v_reg ,
  \nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,\nz.mem_674_sv2v_reg ,
  \nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,
  \nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,\nz.mem_667_sv2v_reg ,
  \nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,
  \nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,
  \nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,\nz.mem_656_sv2v_reg ,
  \nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,
  \nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,\nz.mem_649_sv2v_reg ,
  \nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,\nz.mem_645_sv2v_reg ,
  \nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,
  \nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,\nz.mem_638_sv2v_reg ,
  \nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,
  \nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,
  \nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,\nz.mem_627_sv2v_reg ,
  \nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,
  \nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,
  \nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,
  \nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,
  \nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,\nz.mem_609_sv2v_reg ,
  \nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,
  \nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,
  \nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,\nz.mem_598_sv2v_reg ,
  \nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,
  \nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,
  \nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,\nz.mem_587_sv2v_reg ,
  \nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,
  \nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,
  \nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,
  \nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,
  \nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,\nz.mem_569_sv2v_reg ,
  \nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,
  \nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,
  \nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,\nz.mem_558_sv2v_reg ,
  \nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,
  \nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,
  \nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,\nz.mem_547_sv2v_reg ,
  \nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,
  \nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,
  \nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,
  \nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,
  \nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,\nz.mem_529_sv2v_reg ,
  \nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,
  \nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,
  \nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,\nz.mem_518_sv2v_reg ,
  \nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,
  \nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,
  \nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,\nz.mem_507_sv2v_reg ,
  \nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,
  \nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,
  \nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,
  \nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,
  \nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,\nz.mem_489_sv2v_reg ,
  \nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,
  \nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,
  \nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,\nz.mem_478_sv2v_reg ,
  \nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,
  \nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,
  \nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,\nz.mem_467_sv2v_reg ,
  \nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,
  \nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,
  \nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,
  \nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,
  \nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,
  \nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,
  \nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,
  \nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,
  \nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,
  \nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,
  \nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,
  \nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,
  \nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,
  \nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,
  \nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,
  \nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,
  \nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,
  \nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,
  \nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,
  \nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,
  \nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,
  \nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,
  \nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,
  \nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,
  \nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,
  \nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,
  \nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,
  \nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,
  \nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,
  \nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,
  \nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,
  \nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,
  \nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,
  \nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,
  \nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,
  \nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,
  \nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,
  \nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,
  \nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,
  \nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,
  \nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,
  \nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,
  \nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,
  \nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,
  \nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,
  \nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,
  \nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,
  \nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,
  \nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,
  \nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,
  \nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,
  \nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,
  \nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,
  \nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,
  \nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,
  \nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,
  \nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,
  \nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,
  \nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,
  \nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,
  \nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,
  \nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,
  \nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,
  \nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,
  \nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,
  \nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,
  \nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,
  \nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,
  \nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,
  \nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,
  \nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,
  \nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,
  \nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,
  \nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,
  \nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,
  \nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,
  \nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,
  \nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,
  \nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,
  \nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,
  \nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,
  \nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,
  \nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,
  \nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,
  \nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,
  \nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,
  \nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,
  \nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,
  \nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,
  \nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [5119] = \nz.mem_5119_sv2v_reg ;
  assign \nz.mem [5118] = \nz.mem_5118_sv2v_reg ;
  assign \nz.mem [5117] = \nz.mem_5117_sv2v_reg ;
  assign \nz.mem [5116] = \nz.mem_5116_sv2v_reg ;
  assign \nz.mem [5115] = \nz.mem_5115_sv2v_reg ;
  assign \nz.mem [5114] = \nz.mem_5114_sv2v_reg ;
  assign \nz.mem [5113] = \nz.mem_5113_sv2v_reg ;
  assign \nz.mem [5112] = \nz.mem_5112_sv2v_reg ;
  assign \nz.mem [5111] = \nz.mem_5111_sv2v_reg ;
  assign \nz.mem [5110] = \nz.mem_5110_sv2v_reg ;
  assign \nz.mem [5109] = \nz.mem_5109_sv2v_reg ;
  assign \nz.mem [5108] = \nz.mem_5108_sv2v_reg ;
  assign \nz.mem [5107] = \nz.mem_5107_sv2v_reg ;
  assign \nz.mem [5106] = \nz.mem_5106_sv2v_reg ;
  assign \nz.mem [5105] = \nz.mem_5105_sv2v_reg ;
  assign \nz.mem [5104] = \nz.mem_5104_sv2v_reg ;
  assign \nz.mem [5103] = \nz.mem_5103_sv2v_reg ;
  assign \nz.mem [5102] = \nz.mem_5102_sv2v_reg ;
  assign \nz.mem [5101] = \nz.mem_5101_sv2v_reg ;
  assign \nz.mem [5100] = \nz.mem_5100_sv2v_reg ;
  assign \nz.mem [5099] = \nz.mem_5099_sv2v_reg ;
  assign \nz.mem [5098] = \nz.mem_5098_sv2v_reg ;
  assign \nz.mem [5097] = \nz.mem_5097_sv2v_reg ;
  assign \nz.mem [5096] = \nz.mem_5096_sv2v_reg ;
  assign \nz.mem [5095] = \nz.mem_5095_sv2v_reg ;
  assign \nz.mem [5094] = \nz.mem_5094_sv2v_reg ;
  assign \nz.mem [5093] = \nz.mem_5093_sv2v_reg ;
  assign \nz.mem [5092] = \nz.mem_5092_sv2v_reg ;
  assign \nz.mem [5091] = \nz.mem_5091_sv2v_reg ;
  assign \nz.mem [5090] = \nz.mem_5090_sv2v_reg ;
  assign \nz.mem [5089] = \nz.mem_5089_sv2v_reg ;
  assign \nz.mem [5088] = \nz.mem_5088_sv2v_reg ;
  assign \nz.mem [5087] = \nz.mem_5087_sv2v_reg ;
  assign \nz.mem [5086] = \nz.mem_5086_sv2v_reg ;
  assign \nz.mem [5085] = \nz.mem_5085_sv2v_reg ;
  assign \nz.mem [5084] = \nz.mem_5084_sv2v_reg ;
  assign \nz.mem [5083] = \nz.mem_5083_sv2v_reg ;
  assign \nz.mem [5082] = \nz.mem_5082_sv2v_reg ;
  assign \nz.mem [5081] = \nz.mem_5081_sv2v_reg ;
  assign \nz.mem [5080] = \nz.mem_5080_sv2v_reg ;
  assign \nz.mem [5079] = \nz.mem_5079_sv2v_reg ;
  assign \nz.mem [5078] = \nz.mem_5078_sv2v_reg ;
  assign \nz.mem [5077] = \nz.mem_5077_sv2v_reg ;
  assign \nz.mem [5076] = \nz.mem_5076_sv2v_reg ;
  assign \nz.mem [5075] = \nz.mem_5075_sv2v_reg ;
  assign \nz.mem [5074] = \nz.mem_5074_sv2v_reg ;
  assign \nz.mem [5073] = \nz.mem_5073_sv2v_reg ;
  assign \nz.mem [5072] = \nz.mem_5072_sv2v_reg ;
  assign \nz.mem [5071] = \nz.mem_5071_sv2v_reg ;
  assign \nz.mem [5070] = \nz.mem_5070_sv2v_reg ;
  assign \nz.mem [5069] = \nz.mem_5069_sv2v_reg ;
  assign \nz.mem [5068] = \nz.mem_5068_sv2v_reg ;
  assign \nz.mem [5067] = \nz.mem_5067_sv2v_reg ;
  assign \nz.mem [5066] = \nz.mem_5066_sv2v_reg ;
  assign \nz.mem [5065] = \nz.mem_5065_sv2v_reg ;
  assign \nz.mem [5064] = \nz.mem_5064_sv2v_reg ;
  assign \nz.mem [5063] = \nz.mem_5063_sv2v_reg ;
  assign \nz.mem [5062] = \nz.mem_5062_sv2v_reg ;
  assign \nz.mem [5061] = \nz.mem_5061_sv2v_reg ;
  assign \nz.mem [5060] = \nz.mem_5060_sv2v_reg ;
  assign \nz.mem [5059] = \nz.mem_5059_sv2v_reg ;
  assign \nz.mem [5058] = \nz.mem_5058_sv2v_reg ;
  assign \nz.mem [5057] = \nz.mem_5057_sv2v_reg ;
  assign \nz.mem [5056] = \nz.mem_5056_sv2v_reg ;
  assign \nz.mem [5055] = \nz.mem_5055_sv2v_reg ;
  assign \nz.mem [5054] = \nz.mem_5054_sv2v_reg ;
  assign \nz.mem [5053] = \nz.mem_5053_sv2v_reg ;
  assign \nz.mem [5052] = \nz.mem_5052_sv2v_reg ;
  assign \nz.mem [5051] = \nz.mem_5051_sv2v_reg ;
  assign \nz.mem [5050] = \nz.mem_5050_sv2v_reg ;
  assign \nz.mem [5049] = \nz.mem_5049_sv2v_reg ;
  assign \nz.mem [5048] = \nz.mem_5048_sv2v_reg ;
  assign \nz.mem [5047] = \nz.mem_5047_sv2v_reg ;
  assign \nz.mem [5046] = \nz.mem_5046_sv2v_reg ;
  assign \nz.mem [5045] = \nz.mem_5045_sv2v_reg ;
  assign \nz.mem [5044] = \nz.mem_5044_sv2v_reg ;
  assign \nz.mem [5043] = \nz.mem_5043_sv2v_reg ;
  assign \nz.mem [5042] = \nz.mem_5042_sv2v_reg ;
  assign \nz.mem [5041] = \nz.mem_5041_sv2v_reg ;
  assign \nz.mem [5040] = \nz.mem_5040_sv2v_reg ;
  assign \nz.mem [5039] = \nz.mem_5039_sv2v_reg ;
  assign \nz.mem [5038] = \nz.mem_5038_sv2v_reg ;
  assign \nz.mem [5037] = \nz.mem_5037_sv2v_reg ;
  assign \nz.mem [5036] = \nz.mem_5036_sv2v_reg ;
  assign \nz.mem [5035] = \nz.mem_5035_sv2v_reg ;
  assign \nz.mem [5034] = \nz.mem_5034_sv2v_reg ;
  assign \nz.mem [5033] = \nz.mem_5033_sv2v_reg ;
  assign \nz.mem [5032] = \nz.mem_5032_sv2v_reg ;
  assign \nz.mem [5031] = \nz.mem_5031_sv2v_reg ;
  assign \nz.mem [5030] = \nz.mem_5030_sv2v_reg ;
  assign \nz.mem [5029] = \nz.mem_5029_sv2v_reg ;
  assign \nz.mem [5028] = \nz.mem_5028_sv2v_reg ;
  assign \nz.mem [5027] = \nz.mem_5027_sv2v_reg ;
  assign \nz.mem [5026] = \nz.mem_5026_sv2v_reg ;
  assign \nz.mem [5025] = \nz.mem_5025_sv2v_reg ;
  assign \nz.mem [5024] = \nz.mem_5024_sv2v_reg ;
  assign \nz.mem [5023] = \nz.mem_5023_sv2v_reg ;
  assign \nz.mem [5022] = \nz.mem_5022_sv2v_reg ;
  assign \nz.mem [5021] = \nz.mem_5021_sv2v_reg ;
  assign \nz.mem [5020] = \nz.mem_5020_sv2v_reg ;
  assign \nz.mem [5019] = \nz.mem_5019_sv2v_reg ;
  assign \nz.mem [5018] = \nz.mem_5018_sv2v_reg ;
  assign \nz.mem [5017] = \nz.mem_5017_sv2v_reg ;
  assign \nz.mem [5016] = \nz.mem_5016_sv2v_reg ;
  assign \nz.mem [5015] = \nz.mem_5015_sv2v_reg ;
  assign \nz.mem [5014] = \nz.mem_5014_sv2v_reg ;
  assign \nz.mem [5013] = \nz.mem_5013_sv2v_reg ;
  assign \nz.mem [5012] = \nz.mem_5012_sv2v_reg ;
  assign \nz.mem [5011] = \nz.mem_5011_sv2v_reg ;
  assign \nz.mem [5010] = \nz.mem_5010_sv2v_reg ;
  assign \nz.mem [5009] = \nz.mem_5009_sv2v_reg ;
  assign \nz.mem [5008] = \nz.mem_5008_sv2v_reg ;
  assign \nz.mem [5007] = \nz.mem_5007_sv2v_reg ;
  assign \nz.mem [5006] = \nz.mem_5006_sv2v_reg ;
  assign \nz.mem [5005] = \nz.mem_5005_sv2v_reg ;
  assign \nz.mem [5004] = \nz.mem_5004_sv2v_reg ;
  assign \nz.mem [5003] = \nz.mem_5003_sv2v_reg ;
  assign \nz.mem [5002] = \nz.mem_5002_sv2v_reg ;
  assign \nz.mem [5001] = \nz.mem_5001_sv2v_reg ;
  assign \nz.mem [5000] = \nz.mem_5000_sv2v_reg ;
  assign \nz.mem [4999] = \nz.mem_4999_sv2v_reg ;
  assign \nz.mem [4998] = \nz.mem_4998_sv2v_reg ;
  assign \nz.mem [4997] = \nz.mem_4997_sv2v_reg ;
  assign \nz.mem [4996] = \nz.mem_4996_sv2v_reg ;
  assign \nz.mem [4995] = \nz.mem_4995_sv2v_reg ;
  assign \nz.mem [4994] = \nz.mem_4994_sv2v_reg ;
  assign \nz.mem [4993] = \nz.mem_4993_sv2v_reg ;
  assign \nz.mem [4992] = \nz.mem_4992_sv2v_reg ;
  assign \nz.mem [4991] = \nz.mem_4991_sv2v_reg ;
  assign \nz.mem [4990] = \nz.mem_4990_sv2v_reg ;
  assign \nz.mem [4989] = \nz.mem_4989_sv2v_reg ;
  assign \nz.mem [4988] = \nz.mem_4988_sv2v_reg ;
  assign \nz.mem [4987] = \nz.mem_4987_sv2v_reg ;
  assign \nz.mem [4986] = \nz.mem_4986_sv2v_reg ;
  assign \nz.mem [4985] = \nz.mem_4985_sv2v_reg ;
  assign \nz.mem [4984] = \nz.mem_4984_sv2v_reg ;
  assign \nz.mem [4983] = \nz.mem_4983_sv2v_reg ;
  assign \nz.mem [4982] = \nz.mem_4982_sv2v_reg ;
  assign \nz.mem [4981] = \nz.mem_4981_sv2v_reg ;
  assign \nz.mem [4980] = \nz.mem_4980_sv2v_reg ;
  assign \nz.mem [4979] = \nz.mem_4979_sv2v_reg ;
  assign \nz.mem [4978] = \nz.mem_4978_sv2v_reg ;
  assign \nz.mem [4977] = \nz.mem_4977_sv2v_reg ;
  assign \nz.mem [4976] = \nz.mem_4976_sv2v_reg ;
  assign \nz.mem [4975] = \nz.mem_4975_sv2v_reg ;
  assign \nz.mem [4974] = \nz.mem_4974_sv2v_reg ;
  assign \nz.mem [4973] = \nz.mem_4973_sv2v_reg ;
  assign \nz.mem [4972] = \nz.mem_4972_sv2v_reg ;
  assign \nz.mem [4971] = \nz.mem_4971_sv2v_reg ;
  assign \nz.mem [4970] = \nz.mem_4970_sv2v_reg ;
  assign \nz.mem [4969] = \nz.mem_4969_sv2v_reg ;
  assign \nz.mem [4968] = \nz.mem_4968_sv2v_reg ;
  assign \nz.mem [4967] = \nz.mem_4967_sv2v_reg ;
  assign \nz.mem [4966] = \nz.mem_4966_sv2v_reg ;
  assign \nz.mem [4965] = \nz.mem_4965_sv2v_reg ;
  assign \nz.mem [4964] = \nz.mem_4964_sv2v_reg ;
  assign \nz.mem [4963] = \nz.mem_4963_sv2v_reg ;
  assign \nz.mem [4962] = \nz.mem_4962_sv2v_reg ;
  assign \nz.mem [4961] = \nz.mem_4961_sv2v_reg ;
  assign \nz.mem [4960] = \nz.mem_4960_sv2v_reg ;
  assign \nz.mem [4959] = \nz.mem_4959_sv2v_reg ;
  assign \nz.mem [4958] = \nz.mem_4958_sv2v_reg ;
  assign \nz.mem [4957] = \nz.mem_4957_sv2v_reg ;
  assign \nz.mem [4956] = \nz.mem_4956_sv2v_reg ;
  assign \nz.mem [4955] = \nz.mem_4955_sv2v_reg ;
  assign \nz.mem [4954] = \nz.mem_4954_sv2v_reg ;
  assign \nz.mem [4953] = \nz.mem_4953_sv2v_reg ;
  assign \nz.mem [4952] = \nz.mem_4952_sv2v_reg ;
  assign \nz.mem [4951] = \nz.mem_4951_sv2v_reg ;
  assign \nz.mem [4950] = \nz.mem_4950_sv2v_reg ;
  assign \nz.mem [4949] = \nz.mem_4949_sv2v_reg ;
  assign \nz.mem [4948] = \nz.mem_4948_sv2v_reg ;
  assign \nz.mem [4947] = \nz.mem_4947_sv2v_reg ;
  assign \nz.mem [4946] = \nz.mem_4946_sv2v_reg ;
  assign \nz.mem [4945] = \nz.mem_4945_sv2v_reg ;
  assign \nz.mem [4944] = \nz.mem_4944_sv2v_reg ;
  assign \nz.mem [4943] = \nz.mem_4943_sv2v_reg ;
  assign \nz.mem [4942] = \nz.mem_4942_sv2v_reg ;
  assign \nz.mem [4941] = \nz.mem_4941_sv2v_reg ;
  assign \nz.mem [4940] = \nz.mem_4940_sv2v_reg ;
  assign \nz.mem [4939] = \nz.mem_4939_sv2v_reg ;
  assign \nz.mem [4938] = \nz.mem_4938_sv2v_reg ;
  assign \nz.mem [4937] = \nz.mem_4937_sv2v_reg ;
  assign \nz.mem [4936] = \nz.mem_4936_sv2v_reg ;
  assign \nz.mem [4935] = \nz.mem_4935_sv2v_reg ;
  assign \nz.mem [4934] = \nz.mem_4934_sv2v_reg ;
  assign \nz.mem [4933] = \nz.mem_4933_sv2v_reg ;
  assign \nz.mem [4932] = \nz.mem_4932_sv2v_reg ;
  assign \nz.mem [4931] = \nz.mem_4931_sv2v_reg ;
  assign \nz.mem [4930] = \nz.mem_4930_sv2v_reg ;
  assign \nz.mem [4929] = \nz.mem_4929_sv2v_reg ;
  assign \nz.mem [4928] = \nz.mem_4928_sv2v_reg ;
  assign \nz.mem [4927] = \nz.mem_4927_sv2v_reg ;
  assign \nz.mem [4926] = \nz.mem_4926_sv2v_reg ;
  assign \nz.mem [4925] = \nz.mem_4925_sv2v_reg ;
  assign \nz.mem [4924] = \nz.mem_4924_sv2v_reg ;
  assign \nz.mem [4923] = \nz.mem_4923_sv2v_reg ;
  assign \nz.mem [4922] = \nz.mem_4922_sv2v_reg ;
  assign \nz.mem [4921] = \nz.mem_4921_sv2v_reg ;
  assign \nz.mem [4920] = \nz.mem_4920_sv2v_reg ;
  assign \nz.mem [4919] = \nz.mem_4919_sv2v_reg ;
  assign \nz.mem [4918] = \nz.mem_4918_sv2v_reg ;
  assign \nz.mem [4917] = \nz.mem_4917_sv2v_reg ;
  assign \nz.mem [4916] = \nz.mem_4916_sv2v_reg ;
  assign \nz.mem [4915] = \nz.mem_4915_sv2v_reg ;
  assign \nz.mem [4914] = \nz.mem_4914_sv2v_reg ;
  assign \nz.mem [4913] = \nz.mem_4913_sv2v_reg ;
  assign \nz.mem [4912] = \nz.mem_4912_sv2v_reg ;
  assign \nz.mem [4911] = \nz.mem_4911_sv2v_reg ;
  assign \nz.mem [4910] = \nz.mem_4910_sv2v_reg ;
  assign \nz.mem [4909] = \nz.mem_4909_sv2v_reg ;
  assign \nz.mem [4908] = \nz.mem_4908_sv2v_reg ;
  assign \nz.mem [4907] = \nz.mem_4907_sv2v_reg ;
  assign \nz.mem [4906] = \nz.mem_4906_sv2v_reg ;
  assign \nz.mem [4905] = \nz.mem_4905_sv2v_reg ;
  assign \nz.mem [4904] = \nz.mem_4904_sv2v_reg ;
  assign \nz.mem [4903] = \nz.mem_4903_sv2v_reg ;
  assign \nz.mem [4902] = \nz.mem_4902_sv2v_reg ;
  assign \nz.mem [4901] = \nz.mem_4901_sv2v_reg ;
  assign \nz.mem [4900] = \nz.mem_4900_sv2v_reg ;
  assign \nz.mem [4899] = \nz.mem_4899_sv2v_reg ;
  assign \nz.mem [4898] = \nz.mem_4898_sv2v_reg ;
  assign \nz.mem [4897] = \nz.mem_4897_sv2v_reg ;
  assign \nz.mem [4896] = \nz.mem_4896_sv2v_reg ;
  assign \nz.mem [4895] = \nz.mem_4895_sv2v_reg ;
  assign \nz.mem [4894] = \nz.mem_4894_sv2v_reg ;
  assign \nz.mem [4893] = \nz.mem_4893_sv2v_reg ;
  assign \nz.mem [4892] = \nz.mem_4892_sv2v_reg ;
  assign \nz.mem [4891] = \nz.mem_4891_sv2v_reg ;
  assign \nz.mem [4890] = \nz.mem_4890_sv2v_reg ;
  assign \nz.mem [4889] = \nz.mem_4889_sv2v_reg ;
  assign \nz.mem [4888] = \nz.mem_4888_sv2v_reg ;
  assign \nz.mem [4887] = \nz.mem_4887_sv2v_reg ;
  assign \nz.mem [4886] = \nz.mem_4886_sv2v_reg ;
  assign \nz.mem [4885] = \nz.mem_4885_sv2v_reg ;
  assign \nz.mem [4884] = \nz.mem_4884_sv2v_reg ;
  assign \nz.mem [4883] = \nz.mem_4883_sv2v_reg ;
  assign \nz.mem [4882] = \nz.mem_4882_sv2v_reg ;
  assign \nz.mem [4881] = \nz.mem_4881_sv2v_reg ;
  assign \nz.mem [4880] = \nz.mem_4880_sv2v_reg ;
  assign \nz.mem [4879] = \nz.mem_4879_sv2v_reg ;
  assign \nz.mem [4878] = \nz.mem_4878_sv2v_reg ;
  assign \nz.mem [4877] = \nz.mem_4877_sv2v_reg ;
  assign \nz.mem [4876] = \nz.mem_4876_sv2v_reg ;
  assign \nz.mem [4875] = \nz.mem_4875_sv2v_reg ;
  assign \nz.mem [4874] = \nz.mem_4874_sv2v_reg ;
  assign \nz.mem [4873] = \nz.mem_4873_sv2v_reg ;
  assign \nz.mem [4872] = \nz.mem_4872_sv2v_reg ;
  assign \nz.mem [4871] = \nz.mem_4871_sv2v_reg ;
  assign \nz.mem [4870] = \nz.mem_4870_sv2v_reg ;
  assign \nz.mem [4869] = \nz.mem_4869_sv2v_reg ;
  assign \nz.mem [4868] = \nz.mem_4868_sv2v_reg ;
  assign \nz.mem [4867] = \nz.mem_4867_sv2v_reg ;
  assign \nz.mem [4866] = \nz.mem_4866_sv2v_reg ;
  assign \nz.mem [4865] = \nz.mem_4865_sv2v_reg ;
  assign \nz.mem [4864] = \nz.mem_4864_sv2v_reg ;
  assign \nz.mem [4863] = \nz.mem_4863_sv2v_reg ;
  assign \nz.mem [4862] = \nz.mem_4862_sv2v_reg ;
  assign \nz.mem [4861] = \nz.mem_4861_sv2v_reg ;
  assign \nz.mem [4860] = \nz.mem_4860_sv2v_reg ;
  assign \nz.mem [4859] = \nz.mem_4859_sv2v_reg ;
  assign \nz.mem [4858] = \nz.mem_4858_sv2v_reg ;
  assign \nz.mem [4857] = \nz.mem_4857_sv2v_reg ;
  assign \nz.mem [4856] = \nz.mem_4856_sv2v_reg ;
  assign \nz.mem [4855] = \nz.mem_4855_sv2v_reg ;
  assign \nz.mem [4854] = \nz.mem_4854_sv2v_reg ;
  assign \nz.mem [4853] = \nz.mem_4853_sv2v_reg ;
  assign \nz.mem [4852] = \nz.mem_4852_sv2v_reg ;
  assign \nz.mem [4851] = \nz.mem_4851_sv2v_reg ;
  assign \nz.mem [4850] = \nz.mem_4850_sv2v_reg ;
  assign \nz.mem [4849] = \nz.mem_4849_sv2v_reg ;
  assign \nz.mem [4848] = \nz.mem_4848_sv2v_reg ;
  assign \nz.mem [4847] = \nz.mem_4847_sv2v_reg ;
  assign \nz.mem [4846] = \nz.mem_4846_sv2v_reg ;
  assign \nz.mem [4845] = \nz.mem_4845_sv2v_reg ;
  assign \nz.mem [4844] = \nz.mem_4844_sv2v_reg ;
  assign \nz.mem [4843] = \nz.mem_4843_sv2v_reg ;
  assign \nz.mem [4842] = \nz.mem_4842_sv2v_reg ;
  assign \nz.mem [4841] = \nz.mem_4841_sv2v_reg ;
  assign \nz.mem [4840] = \nz.mem_4840_sv2v_reg ;
  assign \nz.mem [4839] = \nz.mem_4839_sv2v_reg ;
  assign \nz.mem [4838] = \nz.mem_4838_sv2v_reg ;
  assign \nz.mem [4837] = \nz.mem_4837_sv2v_reg ;
  assign \nz.mem [4836] = \nz.mem_4836_sv2v_reg ;
  assign \nz.mem [4835] = \nz.mem_4835_sv2v_reg ;
  assign \nz.mem [4834] = \nz.mem_4834_sv2v_reg ;
  assign \nz.mem [4833] = \nz.mem_4833_sv2v_reg ;
  assign \nz.mem [4832] = \nz.mem_4832_sv2v_reg ;
  assign \nz.mem [4831] = \nz.mem_4831_sv2v_reg ;
  assign \nz.mem [4830] = \nz.mem_4830_sv2v_reg ;
  assign \nz.mem [4829] = \nz.mem_4829_sv2v_reg ;
  assign \nz.mem [4828] = \nz.mem_4828_sv2v_reg ;
  assign \nz.mem [4827] = \nz.mem_4827_sv2v_reg ;
  assign \nz.mem [4826] = \nz.mem_4826_sv2v_reg ;
  assign \nz.mem [4825] = \nz.mem_4825_sv2v_reg ;
  assign \nz.mem [4824] = \nz.mem_4824_sv2v_reg ;
  assign \nz.mem [4823] = \nz.mem_4823_sv2v_reg ;
  assign \nz.mem [4822] = \nz.mem_4822_sv2v_reg ;
  assign \nz.mem [4821] = \nz.mem_4821_sv2v_reg ;
  assign \nz.mem [4820] = \nz.mem_4820_sv2v_reg ;
  assign \nz.mem [4819] = \nz.mem_4819_sv2v_reg ;
  assign \nz.mem [4818] = \nz.mem_4818_sv2v_reg ;
  assign \nz.mem [4817] = \nz.mem_4817_sv2v_reg ;
  assign \nz.mem [4816] = \nz.mem_4816_sv2v_reg ;
  assign \nz.mem [4815] = \nz.mem_4815_sv2v_reg ;
  assign \nz.mem [4814] = \nz.mem_4814_sv2v_reg ;
  assign \nz.mem [4813] = \nz.mem_4813_sv2v_reg ;
  assign \nz.mem [4812] = \nz.mem_4812_sv2v_reg ;
  assign \nz.mem [4811] = \nz.mem_4811_sv2v_reg ;
  assign \nz.mem [4810] = \nz.mem_4810_sv2v_reg ;
  assign \nz.mem [4809] = \nz.mem_4809_sv2v_reg ;
  assign \nz.mem [4808] = \nz.mem_4808_sv2v_reg ;
  assign \nz.mem [4807] = \nz.mem_4807_sv2v_reg ;
  assign \nz.mem [4806] = \nz.mem_4806_sv2v_reg ;
  assign \nz.mem [4805] = \nz.mem_4805_sv2v_reg ;
  assign \nz.mem [4804] = \nz.mem_4804_sv2v_reg ;
  assign \nz.mem [4803] = \nz.mem_4803_sv2v_reg ;
  assign \nz.mem [4802] = \nz.mem_4802_sv2v_reg ;
  assign \nz.mem [4801] = \nz.mem_4801_sv2v_reg ;
  assign \nz.mem [4800] = \nz.mem_4800_sv2v_reg ;
  assign \nz.mem [4799] = \nz.mem_4799_sv2v_reg ;
  assign \nz.mem [4798] = \nz.mem_4798_sv2v_reg ;
  assign \nz.mem [4797] = \nz.mem_4797_sv2v_reg ;
  assign \nz.mem [4796] = \nz.mem_4796_sv2v_reg ;
  assign \nz.mem [4795] = \nz.mem_4795_sv2v_reg ;
  assign \nz.mem [4794] = \nz.mem_4794_sv2v_reg ;
  assign \nz.mem [4793] = \nz.mem_4793_sv2v_reg ;
  assign \nz.mem [4792] = \nz.mem_4792_sv2v_reg ;
  assign \nz.mem [4791] = \nz.mem_4791_sv2v_reg ;
  assign \nz.mem [4790] = \nz.mem_4790_sv2v_reg ;
  assign \nz.mem [4789] = \nz.mem_4789_sv2v_reg ;
  assign \nz.mem [4788] = \nz.mem_4788_sv2v_reg ;
  assign \nz.mem [4787] = \nz.mem_4787_sv2v_reg ;
  assign \nz.mem [4786] = \nz.mem_4786_sv2v_reg ;
  assign \nz.mem [4785] = \nz.mem_4785_sv2v_reg ;
  assign \nz.mem [4784] = \nz.mem_4784_sv2v_reg ;
  assign \nz.mem [4783] = \nz.mem_4783_sv2v_reg ;
  assign \nz.mem [4782] = \nz.mem_4782_sv2v_reg ;
  assign \nz.mem [4781] = \nz.mem_4781_sv2v_reg ;
  assign \nz.mem [4780] = \nz.mem_4780_sv2v_reg ;
  assign \nz.mem [4779] = \nz.mem_4779_sv2v_reg ;
  assign \nz.mem [4778] = \nz.mem_4778_sv2v_reg ;
  assign \nz.mem [4777] = \nz.mem_4777_sv2v_reg ;
  assign \nz.mem [4776] = \nz.mem_4776_sv2v_reg ;
  assign \nz.mem [4775] = \nz.mem_4775_sv2v_reg ;
  assign \nz.mem [4774] = \nz.mem_4774_sv2v_reg ;
  assign \nz.mem [4773] = \nz.mem_4773_sv2v_reg ;
  assign \nz.mem [4772] = \nz.mem_4772_sv2v_reg ;
  assign \nz.mem [4771] = \nz.mem_4771_sv2v_reg ;
  assign \nz.mem [4770] = \nz.mem_4770_sv2v_reg ;
  assign \nz.mem [4769] = \nz.mem_4769_sv2v_reg ;
  assign \nz.mem [4768] = \nz.mem_4768_sv2v_reg ;
  assign \nz.mem [4767] = \nz.mem_4767_sv2v_reg ;
  assign \nz.mem [4766] = \nz.mem_4766_sv2v_reg ;
  assign \nz.mem [4765] = \nz.mem_4765_sv2v_reg ;
  assign \nz.mem [4764] = \nz.mem_4764_sv2v_reg ;
  assign \nz.mem [4763] = \nz.mem_4763_sv2v_reg ;
  assign \nz.mem [4762] = \nz.mem_4762_sv2v_reg ;
  assign \nz.mem [4761] = \nz.mem_4761_sv2v_reg ;
  assign \nz.mem [4760] = \nz.mem_4760_sv2v_reg ;
  assign \nz.mem [4759] = \nz.mem_4759_sv2v_reg ;
  assign \nz.mem [4758] = \nz.mem_4758_sv2v_reg ;
  assign \nz.mem [4757] = \nz.mem_4757_sv2v_reg ;
  assign \nz.mem [4756] = \nz.mem_4756_sv2v_reg ;
  assign \nz.mem [4755] = \nz.mem_4755_sv2v_reg ;
  assign \nz.mem [4754] = \nz.mem_4754_sv2v_reg ;
  assign \nz.mem [4753] = \nz.mem_4753_sv2v_reg ;
  assign \nz.mem [4752] = \nz.mem_4752_sv2v_reg ;
  assign \nz.mem [4751] = \nz.mem_4751_sv2v_reg ;
  assign \nz.mem [4750] = \nz.mem_4750_sv2v_reg ;
  assign \nz.mem [4749] = \nz.mem_4749_sv2v_reg ;
  assign \nz.mem [4748] = \nz.mem_4748_sv2v_reg ;
  assign \nz.mem [4747] = \nz.mem_4747_sv2v_reg ;
  assign \nz.mem [4746] = \nz.mem_4746_sv2v_reg ;
  assign \nz.mem [4745] = \nz.mem_4745_sv2v_reg ;
  assign \nz.mem [4744] = \nz.mem_4744_sv2v_reg ;
  assign \nz.mem [4743] = \nz.mem_4743_sv2v_reg ;
  assign \nz.mem [4742] = \nz.mem_4742_sv2v_reg ;
  assign \nz.mem [4741] = \nz.mem_4741_sv2v_reg ;
  assign \nz.mem [4740] = \nz.mem_4740_sv2v_reg ;
  assign \nz.mem [4739] = \nz.mem_4739_sv2v_reg ;
  assign \nz.mem [4738] = \nz.mem_4738_sv2v_reg ;
  assign \nz.mem [4737] = \nz.mem_4737_sv2v_reg ;
  assign \nz.mem [4736] = \nz.mem_4736_sv2v_reg ;
  assign \nz.mem [4735] = \nz.mem_4735_sv2v_reg ;
  assign \nz.mem [4734] = \nz.mem_4734_sv2v_reg ;
  assign \nz.mem [4733] = \nz.mem_4733_sv2v_reg ;
  assign \nz.mem [4732] = \nz.mem_4732_sv2v_reg ;
  assign \nz.mem [4731] = \nz.mem_4731_sv2v_reg ;
  assign \nz.mem [4730] = \nz.mem_4730_sv2v_reg ;
  assign \nz.mem [4729] = \nz.mem_4729_sv2v_reg ;
  assign \nz.mem [4728] = \nz.mem_4728_sv2v_reg ;
  assign \nz.mem [4727] = \nz.mem_4727_sv2v_reg ;
  assign \nz.mem [4726] = \nz.mem_4726_sv2v_reg ;
  assign \nz.mem [4725] = \nz.mem_4725_sv2v_reg ;
  assign \nz.mem [4724] = \nz.mem_4724_sv2v_reg ;
  assign \nz.mem [4723] = \nz.mem_4723_sv2v_reg ;
  assign \nz.mem [4722] = \nz.mem_4722_sv2v_reg ;
  assign \nz.mem [4721] = \nz.mem_4721_sv2v_reg ;
  assign \nz.mem [4720] = \nz.mem_4720_sv2v_reg ;
  assign \nz.mem [4719] = \nz.mem_4719_sv2v_reg ;
  assign \nz.mem [4718] = \nz.mem_4718_sv2v_reg ;
  assign \nz.mem [4717] = \nz.mem_4717_sv2v_reg ;
  assign \nz.mem [4716] = \nz.mem_4716_sv2v_reg ;
  assign \nz.mem [4715] = \nz.mem_4715_sv2v_reg ;
  assign \nz.mem [4714] = \nz.mem_4714_sv2v_reg ;
  assign \nz.mem [4713] = \nz.mem_4713_sv2v_reg ;
  assign \nz.mem [4712] = \nz.mem_4712_sv2v_reg ;
  assign \nz.mem [4711] = \nz.mem_4711_sv2v_reg ;
  assign \nz.mem [4710] = \nz.mem_4710_sv2v_reg ;
  assign \nz.mem [4709] = \nz.mem_4709_sv2v_reg ;
  assign \nz.mem [4708] = \nz.mem_4708_sv2v_reg ;
  assign \nz.mem [4707] = \nz.mem_4707_sv2v_reg ;
  assign \nz.mem [4706] = \nz.mem_4706_sv2v_reg ;
  assign \nz.mem [4705] = \nz.mem_4705_sv2v_reg ;
  assign \nz.mem [4704] = \nz.mem_4704_sv2v_reg ;
  assign \nz.mem [4703] = \nz.mem_4703_sv2v_reg ;
  assign \nz.mem [4702] = \nz.mem_4702_sv2v_reg ;
  assign \nz.mem [4701] = \nz.mem_4701_sv2v_reg ;
  assign \nz.mem [4700] = \nz.mem_4700_sv2v_reg ;
  assign \nz.mem [4699] = \nz.mem_4699_sv2v_reg ;
  assign \nz.mem [4698] = \nz.mem_4698_sv2v_reg ;
  assign \nz.mem [4697] = \nz.mem_4697_sv2v_reg ;
  assign \nz.mem [4696] = \nz.mem_4696_sv2v_reg ;
  assign \nz.mem [4695] = \nz.mem_4695_sv2v_reg ;
  assign \nz.mem [4694] = \nz.mem_4694_sv2v_reg ;
  assign \nz.mem [4693] = \nz.mem_4693_sv2v_reg ;
  assign \nz.mem [4692] = \nz.mem_4692_sv2v_reg ;
  assign \nz.mem [4691] = \nz.mem_4691_sv2v_reg ;
  assign \nz.mem [4690] = \nz.mem_4690_sv2v_reg ;
  assign \nz.mem [4689] = \nz.mem_4689_sv2v_reg ;
  assign \nz.mem [4688] = \nz.mem_4688_sv2v_reg ;
  assign \nz.mem [4687] = \nz.mem_4687_sv2v_reg ;
  assign \nz.mem [4686] = \nz.mem_4686_sv2v_reg ;
  assign \nz.mem [4685] = \nz.mem_4685_sv2v_reg ;
  assign \nz.mem [4684] = \nz.mem_4684_sv2v_reg ;
  assign \nz.mem [4683] = \nz.mem_4683_sv2v_reg ;
  assign \nz.mem [4682] = \nz.mem_4682_sv2v_reg ;
  assign \nz.mem [4681] = \nz.mem_4681_sv2v_reg ;
  assign \nz.mem [4680] = \nz.mem_4680_sv2v_reg ;
  assign \nz.mem [4679] = \nz.mem_4679_sv2v_reg ;
  assign \nz.mem [4678] = \nz.mem_4678_sv2v_reg ;
  assign \nz.mem [4677] = \nz.mem_4677_sv2v_reg ;
  assign \nz.mem [4676] = \nz.mem_4676_sv2v_reg ;
  assign \nz.mem [4675] = \nz.mem_4675_sv2v_reg ;
  assign \nz.mem [4674] = \nz.mem_4674_sv2v_reg ;
  assign \nz.mem [4673] = \nz.mem_4673_sv2v_reg ;
  assign \nz.mem [4672] = \nz.mem_4672_sv2v_reg ;
  assign \nz.mem [4671] = \nz.mem_4671_sv2v_reg ;
  assign \nz.mem [4670] = \nz.mem_4670_sv2v_reg ;
  assign \nz.mem [4669] = \nz.mem_4669_sv2v_reg ;
  assign \nz.mem [4668] = \nz.mem_4668_sv2v_reg ;
  assign \nz.mem [4667] = \nz.mem_4667_sv2v_reg ;
  assign \nz.mem [4666] = \nz.mem_4666_sv2v_reg ;
  assign \nz.mem [4665] = \nz.mem_4665_sv2v_reg ;
  assign \nz.mem [4664] = \nz.mem_4664_sv2v_reg ;
  assign \nz.mem [4663] = \nz.mem_4663_sv2v_reg ;
  assign \nz.mem [4662] = \nz.mem_4662_sv2v_reg ;
  assign \nz.mem [4661] = \nz.mem_4661_sv2v_reg ;
  assign \nz.mem [4660] = \nz.mem_4660_sv2v_reg ;
  assign \nz.mem [4659] = \nz.mem_4659_sv2v_reg ;
  assign \nz.mem [4658] = \nz.mem_4658_sv2v_reg ;
  assign \nz.mem [4657] = \nz.mem_4657_sv2v_reg ;
  assign \nz.mem [4656] = \nz.mem_4656_sv2v_reg ;
  assign \nz.mem [4655] = \nz.mem_4655_sv2v_reg ;
  assign \nz.mem [4654] = \nz.mem_4654_sv2v_reg ;
  assign \nz.mem [4653] = \nz.mem_4653_sv2v_reg ;
  assign \nz.mem [4652] = \nz.mem_4652_sv2v_reg ;
  assign \nz.mem [4651] = \nz.mem_4651_sv2v_reg ;
  assign \nz.mem [4650] = \nz.mem_4650_sv2v_reg ;
  assign \nz.mem [4649] = \nz.mem_4649_sv2v_reg ;
  assign \nz.mem [4648] = \nz.mem_4648_sv2v_reg ;
  assign \nz.mem [4647] = \nz.mem_4647_sv2v_reg ;
  assign \nz.mem [4646] = \nz.mem_4646_sv2v_reg ;
  assign \nz.mem [4645] = \nz.mem_4645_sv2v_reg ;
  assign \nz.mem [4644] = \nz.mem_4644_sv2v_reg ;
  assign \nz.mem [4643] = \nz.mem_4643_sv2v_reg ;
  assign \nz.mem [4642] = \nz.mem_4642_sv2v_reg ;
  assign \nz.mem [4641] = \nz.mem_4641_sv2v_reg ;
  assign \nz.mem [4640] = \nz.mem_4640_sv2v_reg ;
  assign \nz.mem [4639] = \nz.mem_4639_sv2v_reg ;
  assign \nz.mem [4638] = \nz.mem_4638_sv2v_reg ;
  assign \nz.mem [4637] = \nz.mem_4637_sv2v_reg ;
  assign \nz.mem [4636] = \nz.mem_4636_sv2v_reg ;
  assign \nz.mem [4635] = \nz.mem_4635_sv2v_reg ;
  assign \nz.mem [4634] = \nz.mem_4634_sv2v_reg ;
  assign \nz.mem [4633] = \nz.mem_4633_sv2v_reg ;
  assign \nz.mem [4632] = \nz.mem_4632_sv2v_reg ;
  assign \nz.mem [4631] = \nz.mem_4631_sv2v_reg ;
  assign \nz.mem [4630] = \nz.mem_4630_sv2v_reg ;
  assign \nz.mem [4629] = \nz.mem_4629_sv2v_reg ;
  assign \nz.mem [4628] = \nz.mem_4628_sv2v_reg ;
  assign \nz.mem [4627] = \nz.mem_4627_sv2v_reg ;
  assign \nz.mem [4626] = \nz.mem_4626_sv2v_reg ;
  assign \nz.mem [4625] = \nz.mem_4625_sv2v_reg ;
  assign \nz.mem [4624] = \nz.mem_4624_sv2v_reg ;
  assign \nz.mem [4623] = \nz.mem_4623_sv2v_reg ;
  assign \nz.mem [4622] = \nz.mem_4622_sv2v_reg ;
  assign \nz.mem [4621] = \nz.mem_4621_sv2v_reg ;
  assign \nz.mem [4620] = \nz.mem_4620_sv2v_reg ;
  assign \nz.mem [4619] = \nz.mem_4619_sv2v_reg ;
  assign \nz.mem [4618] = \nz.mem_4618_sv2v_reg ;
  assign \nz.mem [4617] = \nz.mem_4617_sv2v_reg ;
  assign \nz.mem [4616] = \nz.mem_4616_sv2v_reg ;
  assign \nz.mem [4615] = \nz.mem_4615_sv2v_reg ;
  assign \nz.mem [4614] = \nz.mem_4614_sv2v_reg ;
  assign \nz.mem [4613] = \nz.mem_4613_sv2v_reg ;
  assign \nz.mem [4612] = \nz.mem_4612_sv2v_reg ;
  assign \nz.mem [4611] = \nz.mem_4611_sv2v_reg ;
  assign \nz.mem [4610] = \nz.mem_4610_sv2v_reg ;
  assign \nz.mem [4609] = \nz.mem_4609_sv2v_reg ;
  assign \nz.mem [4608] = \nz.mem_4608_sv2v_reg ;
  assign \nz.mem [4607] = \nz.mem_4607_sv2v_reg ;
  assign \nz.mem [4606] = \nz.mem_4606_sv2v_reg ;
  assign \nz.mem [4605] = \nz.mem_4605_sv2v_reg ;
  assign \nz.mem [4604] = \nz.mem_4604_sv2v_reg ;
  assign \nz.mem [4603] = \nz.mem_4603_sv2v_reg ;
  assign \nz.mem [4602] = \nz.mem_4602_sv2v_reg ;
  assign \nz.mem [4601] = \nz.mem_4601_sv2v_reg ;
  assign \nz.mem [4600] = \nz.mem_4600_sv2v_reg ;
  assign \nz.mem [4599] = \nz.mem_4599_sv2v_reg ;
  assign \nz.mem [4598] = \nz.mem_4598_sv2v_reg ;
  assign \nz.mem [4597] = \nz.mem_4597_sv2v_reg ;
  assign \nz.mem [4596] = \nz.mem_4596_sv2v_reg ;
  assign \nz.mem [4595] = \nz.mem_4595_sv2v_reg ;
  assign \nz.mem [4594] = \nz.mem_4594_sv2v_reg ;
  assign \nz.mem [4593] = \nz.mem_4593_sv2v_reg ;
  assign \nz.mem [4592] = \nz.mem_4592_sv2v_reg ;
  assign \nz.mem [4591] = \nz.mem_4591_sv2v_reg ;
  assign \nz.mem [4590] = \nz.mem_4590_sv2v_reg ;
  assign \nz.mem [4589] = \nz.mem_4589_sv2v_reg ;
  assign \nz.mem [4588] = \nz.mem_4588_sv2v_reg ;
  assign \nz.mem [4587] = \nz.mem_4587_sv2v_reg ;
  assign \nz.mem [4586] = \nz.mem_4586_sv2v_reg ;
  assign \nz.mem [4585] = \nz.mem_4585_sv2v_reg ;
  assign \nz.mem [4584] = \nz.mem_4584_sv2v_reg ;
  assign \nz.mem [4583] = \nz.mem_4583_sv2v_reg ;
  assign \nz.mem [4582] = \nz.mem_4582_sv2v_reg ;
  assign \nz.mem [4581] = \nz.mem_4581_sv2v_reg ;
  assign \nz.mem [4580] = \nz.mem_4580_sv2v_reg ;
  assign \nz.mem [4579] = \nz.mem_4579_sv2v_reg ;
  assign \nz.mem [4578] = \nz.mem_4578_sv2v_reg ;
  assign \nz.mem [4577] = \nz.mem_4577_sv2v_reg ;
  assign \nz.mem [4576] = \nz.mem_4576_sv2v_reg ;
  assign \nz.mem [4575] = \nz.mem_4575_sv2v_reg ;
  assign \nz.mem [4574] = \nz.mem_4574_sv2v_reg ;
  assign \nz.mem [4573] = \nz.mem_4573_sv2v_reg ;
  assign \nz.mem [4572] = \nz.mem_4572_sv2v_reg ;
  assign \nz.mem [4571] = \nz.mem_4571_sv2v_reg ;
  assign \nz.mem [4570] = \nz.mem_4570_sv2v_reg ;
  assign \nz.mem [4569] = \nz.mem_4569_sv2v_reg ;
  assign \nz.mem [4568] = \nz.mem_4568_sv2v_reg ;
  assign \nz.mem [4567] = \nz.mem_4567_sv2v_reg ;
  assign \nz.mem [4566] = \nz.mem_4566_sv2v_reg ;
  assign \nz.mem [4565] = \nz.mem_4565_sv2v_reg ;
  assign \nz.mem [4564] = \nz.mem_4564_sv2v_reg ;
  assign \nz.mem [4563] = \nz.mem_4563_sv2v_reg ;
  assign \nz.mem [4562] = \nz.mem_4562_sv2v_reg ;
  assign \nz.mem [4561] = \nz.mem_4561_sv2v_reg ;
  assign \nz.mem [4560] = \nz.mem_4560_sv2v_reg ;
  assign \nz.mem [4559] = \nz.mem_4559_sv2v_reg ;
  assign \nz.mem [4558] = \nz.mem_4558_sv2v_reg ;
  assign \nz.mem [4557] = \nz.mem_4557_sv2v_reg ;
  assign \nz.mem [4556] = \nz.mem_4556_sv2v_reg ;
  assign \nz.mem [4555] = \nz.mem_4555_sv2v_reg ;
  assign \nz.mem [4554] = \nz.mem_4554_sv2v_reg ;
  assign \nz.mem [4553] = \nz.mem_4553_sv2v_reg ;
  assign \nz.mem [4552] = \nz.mem_4552_sv2v_reg ;
  assign \nz.mem [4551] = \nz.mem_4551_sv2v_reg ;
  assign \nz.mem [4550] = \nz.mem_4550_sv2v_reg ;
  assign \nz.mem [4549] = \nz.mem_4549_sv2v_reg ;
  assign \nz.mem [4548] = \nz.mem_4548_sv2v_reg ;
  assign \nz.mem [4547] = \nz.mem_4547_sv2v_reg ;
  assign \nz.mem [4546] = \nz.mem_4546_sv2v_reg ;
  assign \nz.mem [4545] = \nz.mem_4545_sv2v_reg ;
  assign \nz.mem [4544] = \nz.mem_4544_sv2v_reg ;
  assign \nz.mem [4543] = \nz.mem_4543_sv2v_reg ;
  assign \nz.mem [4542] = \nz.mem_4542_sv2v_reg ;
  assign \nz.mem [4541] = \nz.mem_4541_sv2v_reg ;
  assign \nz.mem [4540] = \nz.mem_4540_sv2v_reg ;
  assign \nz.mem [4539] = \nz.mem_4539_sv2v_reg ;
  assign \nz.mem [4538] = \nz.mem_4538_sv2v_reg ;
  assign \nz.mem [4537] = \nz.mem_4537_sv2v_reg ;
  assign \nz.mem [4536] = \nz.mem_4536_sv2v_reg ;
  assign \nz.mem [4535] = \nz.mem_4535_sv2v_reg ;
  assign \nz.mem [4534] = \nz.mem_4534_sv2v_reg ;
  assign \nz.mem [4533] = \nz.mem_4533_sv2v_reg ;
  assign \nz.mem [4532] = \nz.mem_4532_sv2v_reg ;
  assign \nz.mem [4531] = \nz.mem_4531_sv2v_reg ;
  assign \nz.mem [4530] = \nz.mem_4530_sv2v_reg ;
  assign \nz.mem [4529] = \nz.mem_4529_sv2v_reg ;
  assign \nz.mem [4528] = \nz.mem_4528_sv2v_reg ;
  assign \nz.mem [4527] = \nz.mem_4527_sv2v_reg ;
  assign \nz.mem [4526] = \nz.mem_4526_sv2v_reg ;
  assign \nz.mem [4525] = \nz.mem_4525_sv2v_reg ;
  assign \nz.mem [4524] = \nz.mem_4524_sv2v_reg ;
  assign \nz.mem [4523] = \nz.mem_4523_sv2v_reg ;
  assign \nz.mem [4522] = \nz.mem_4522_sv2v_reg ;
  assign \nz.mem [4521] = \nz.mem_4521_sv2v_reg ;
  assign \nz.mem [4520] = \nz.mem_4520_sv2v_reg ;
  assign \nz.mem [4519] = \nz.mem_4519_sv2v_reg ;
  assign \nz.mem [4518] = \nz.mem_4518_sv2v_reg ;
  assign \nz.mem [4517] = \nz.mem_4517_sv2v_reg ;
  assign \nz.mem [4516] = \nz.mem_4516_sv2v_reg ;
  assign \nz.mem [4515] = \nz.mem_4515_sv2v_reg ;
  assign \nz.mem [4514] = \nz.mem_4514_sv2v_reg ;
  assign \nz.mem [4513] = \nz.mem_4513_sv2v_reg ;
  assign \nz.mem [4512] = \nz.mem_4512_sv2v_reg ;
  assign \nz.mem [4511] = \nz.mem_4511_sv2v_reg ;
  assign \nz.mem [4510] = \nz.mem_4510_sv2v_reg ;
  assign \nz.mem [4509] = \nz.mem_4509_sv2v_reg ;
  assign \nz.mem [4508] = \nz.mem_4508_sv2v_reg ;
  assign \nz.mem [4507] = \nz.mem_4507_sv2v_reg ;
  assign \nz.mem [4506] = \nz.mem_4506_sv2v_reg ;
  assign \nz.mem [4505] = \nz.mem_4505_sv2v_reg ;
  assign \nz.mem [4504] = \nz.mem_4504_sv2v_reg ;
  assign \nz.mem [4503] = \nz.mem_4503_sv2v_reg ;
  assign \nz.mem [4502] = \nz.mem_4502_sv2v_reg ;
  assign \nz.mem [4501] = \nz.mem_4501_sv2v_reg ;
  assign \nz.mem [4500] = \nz.mem_4500_sv2v_reg ;
  assign \nz.mem [4499] = \nz.mem_4499_sv2v_reg ;
  assign \nz.mem [4498] = \nz.mem_4498_sv2v_reg ;
  assign \nz.mem [4497] = \nz.mem_4497_sv2v_reg ;
  assign \nz.mem [4496] = \nz.mem_4496_sv2v_reg ;
  assign \nz.mem [4495] = \nz.mem_4495_sv2v_reg ;
  assign \nz.mem [4494] = \nz.mem_4494_sv2v_reg ;
  assign \nz.mem [4493] = \nz.mem_4493_sv2v_reg ;
  assign \nz.mem [4492] = \nz.mem_4492_sv2v_reg ;
  assign \nz.mem [4491] = \nz.mem_4491_sv2v_reg ;
  assign \nz.mem [4490] = \nz.mem_4490_sv2v_reg ;
  assign \nz.mem [4489] = \nz.mem_4489_sv2v_reg ;
  assign \nz.mem [4488] = \nz.mem_4488_sv2v_reg ;
  assign \nz.mem [4487] = \nz.mem_4487_sv2v_reg ;
  assign \nz.mem [4486] = \nz.mem_4486_sv2v_reg ;
  assign \nz.mem [4485] = \nz.mem_4485_sv2v_reg ;
  assign \nz.mem [4484] = \nz.mem_4484_sv2v_reg ;
  assign \nz.mem [4483] = \nz.mem_4483_sv2v_reg ;
  assign \nz.mem [4482] = \nz.mem_4482_sv2v_reg ;
  assign \nz.mem [4481] = \nz.mem_4481_sv2v_reg ;
  assign \nz.mem [4480] = \nz.mem_4480_sv2v_reg ;
  assign \nz.mem [4479] = \nz.mem_4479_sv2v_reg ;
  assign \nz.mem [4478] = \nz.mem_4478_sv2v_reg ;
  assign \nz.mem [4477] = \nz.mem_4477_sv2v_reg ;
  assign \nz.mem [4476] = \nz.mem_4476_sv2v_reg ;
  assign \nz.mem [4475] = \nz.mem_4475_sv2v_reg ;
  assign \nz.mem [4474] = \nz.mem_4474_sv2v_reg ;
  assign \nz.mem [4473] = \nz.mem_4473_sv2v_reg ;
  assign \nz.mem [4472] = \nz.mem_4472_sv2v_reg ;
  assign \nz.mem [4471] = \nz.mem_4471_sv2v_reg ;
  assign \nz.mem [4470] = \nz.mem_4470_sv2v_reg ;
  assign \nz.mem [4469] = \nz.mem_4469_sv2v_reg ;
  assign \nz.mem [4468] = \nz.mem_4468_sv2v_reg ;
  assign \nz.mem [4467] = \nz.mem_4467_sv2v_reg ;
  assign \nz.mem [4466] = \nz.mem_4466_sv2v_reg ;
  assign \nz.mem [4465] = \nz.mem_4465_sv2v_reg ;
  assign \nz.mem [4464] = \nz.mem_4464_sv2v_reg ;
  assign \nz.mem [4463] = \nz.mem_4463_sv2v_reg ;
  assign \nz.mem [4462] = \nz.mem_4462_sv2v_reg ;
  assign \nz.mem [4461] = \nz.mem_4461_sv2v_reg ;
  assign \nz.mem [4460] = \nz.mem_4460_sv2v_reg ;
  assign \nz.mem [4459] = \nz.mem_4459_sv2v_reg ;
  assign \nz.mem [4458] = \nz.mem_4458_sv2v_reg ;
  assign \nz.mem [4457] = \nz.mem_4457_sv2v_reg ;
  assign \nz.mem [4456] = \nz.mem_4456_sv2v_reg ;
  assign \nz.mem [4455] = \nz.mem_4455_sv2v_reg ;
  assign \nz.mem [4454] = \nz.mem_4454_sv2v_reg ;
  assign \nz.mem [4453] = \nz.mem_4453_sv2v_reg ;
  assign \nz.mem [4452] = \nz.mem_4452_sv2v_reg ;
  assign \nz.mem [4451] = \nz.mem_4451_sv2v_reg ;
  assign \nz.mem [4450] = \nz.mem_4450_sv2v_reg ;
  assign \nz.mem [4449] = \nz.mem_4449_sv2v_reg ;
  assign \nz.mem [4448] = \nz.mem_4448_sv2v_reg ;
  assign \nz.mem [4447] = \nz.mem_4447_sv2v_reg ;
  assign \nz.mem [4446] = \nz.mem_4446_sv2v_reg ;
  assign \nz.mem [4445] = \nz.mem_4445_sv2v_reg ;
  assign \nz.mem [4444] = \nz.mem_4444_sv2v_reg ;
  assign \nz.mem [4443] = \nz.mem_4443_sv2v_reg ;
  assign \nz.mem [4442] = \nz.mem_4442_sv2v_reg ;
  assign \nz.mem [4441] = \nz.mem_4441_sv2v_reg ;
  assign \nz.mem [4440] = \nz.mem_4440_sv2v_reg ;
  assign \nz.mem [4439] = \nz.mem_4439_sv2v_reg ;
  assign \nz.mem [4438] = \nz.mem_4438_sv2v_reg ;
  assign \nz.mem [4437] = \nz.mem_4437_sv2v_reg ;
  assign \nz.mem [4436] = \nz.mem_4436_sv2v_reg ;
  assign \nz.mem [4435] = \nz.mem_4435_sv2v_reg ;
  assign \nz.mem [4434] = \nz.mem_4434_sv2v_reg ;
  assign \nz.mem [4433] = \nz.mem_4433_sv2v_reg ;
  assign \nz.mem [4432] = \nz.mem_4432_sv2v_reg ;
  assign \nz.mem [4431] = \nz.mem_4431_sv2v_reg ;
  assign \nz.mem [4430] = \nz.mem_4430_sv2v_reg ;
  assign \nz.mem [4429] = \nz.mem_4429_sv2v_reg ;
  assign \nz.mem [4428] = \nz.mem_4428_sv2v_reg ;
  assign \nz.mem [4427] = \nz.mem_4427_sv2v_reg ;
  assign \nz.mem [4426] = \nz.mem_4426_sv2v_reg ;
  assign \nz.mem [4425] = \nz.mem_4425_sv2v_reg ;
  assign \nz.mem [4424] = \nz.mem_4424_sv2v_reg ;
  assign \nz.mem [4423] = \nz.mem_4423_sv2v_reg ;
  assign \nz.mem [4422] = \nz.mem_4422_sv2v_reg ;
  assign \nz.mem [4421] = \nz.mem_4421_sv2v_reg ;
  assign \nz.mem [4420] = \nz.mem_4420_sv2v_reg ;
  assign \nz.mem [4419] = \nz.mem_4419_sv2v_reg ;
  assign \nz.mem [4418] = \nz.mem_4418_sv2v_reg ;
  assign \nz.mem [4417] = \nz.mem_4417_sv2v_reg ;
  assign \nz.mem [4416] = \nz.mem_4416_sv2v_reg ;
  assign \nz.mem [4415] = \nz.mem_4415_sv2v_reg ;
  assign \nz.mem [4414] = \nz.mem_4414_sv2v_reg ;
  assign \nz.mem [4413] = \nz.mem_4413_sv2v_reg ;
  assign \nz.mem [4412] = \nz.mem_4412_sv2v_reg ;
  assign \nz.mem [4411] = \nz.mem_4411_sv2v_reg ;
  assign \nz.mem [4410] = \nz.mem_4410_sv2v_reg ;
  assign \nz.mem [4409] = \nz.mem_4409_sv2v_reg ;
  assign \nz.mem [4408] = \nz.mem_4408_sv2v_reg ;
  assign \nz.mem [4407] = \nz.mem_4407_sv2v_reg ;
  assign \nz.mem [4406] = \nz.mem_4406_sv2v_reg ;
  assign \nz.mem [4405] = \nz.mem_4405_sv2v_reg ;
  assign \nz.mem [4404] = \nz.mem_4404_sv2v_reg ;
  assign \nz.mem [4403] = \nz.mem_4403_sv2v_reg ;
  assign \nz.mem [4402] = \nz.mem_4402_sv2v_reg ;
  assign \nz.mem [4401] = \nz.mem_4401_sv2v_reg ;
  assign \nz.mem [4400] = \nz.mem_4400_sv2v_reg ;
  assign \nz.mem [4399] = \nz.mem_4399_sv2v_reg ;
  assign \nz.mem [4398] = \nz.mem_4398_sv2v_reg ;
  assign \nz.mem [4397] = \nz.mem_4397_sv2v_reg ;
  assign \nz.mem [4396] = \nz.mem_4396_sv2v_reg ;
  assign \nz.mem [4395] = \nz.mem_4395_sv2v_reg ;
  assign \nz.mem [4394] = \nz.mem_4394_sv2v_reg ;
  assign \nz.mem [4393] = \nz.mem_4393_sv2v_reg ;
  assign \nz.mem [4392] = \nz.mem_4392_sv2v_reg ;
  assign \nz.mem [4391] = \nz.mem_4391_sv2v_reg ;
  assign \nz.mem [4390] = \nz.mem_4390_sv2v_reg ;
  assign \nz.mem [4389] = \nz.mem_4389_sv2v_reg ;
  assign \nz.mem [4388] = \nz.mem_4388_sv2v_reg ;
  assign \nz.mem [4387] = \nz.mem_4387_sv2v_reg ;
  assign \nz.mem [4386] = \nz.mem_4386_sv2v_reg ;
  assign \nz.mem [4385] = \nz.mem_4385_sv2v_reg ;
  assign \nz.mem [4384] = \nz.mem_4384_sv2v_reg ;
  assign \nz.mem [4383] = \nz.mem_4383_sv2v_reg ;
  assign \nz.mem [4382] = \nz.mem_4382_sv2v_reg ;
  assign \nz.mem [4381] = \nz.mem_4381_sv2v_reg ;
  assign \nz.mem [4380] = \nz.mem_4380_sv2v_reg ;
  assign \nz.mem [4379] = \nz.mem_4379_sv2v_reg ;
  assign \nz.mem [4378] = \nz.mem_4378_sv2v_reg ;
  assign \nz.mem [4377] = \nz.mem_4377_sv2v_reg ;
  assign \nz.mem [4376] = \nz.mem_4376_sv2v_reg ;
  assign \nz.mem [4375] = \nz.mem_4375_sv2v_reg ;
  assign \nz.mem [4374] = \nz.mem_4374_sv2v_reg ;
  assign \nz.mem [4373] = \nz.mem_4373_sv2v_reg ;
  assign \nz.mem [4372] = \nz.mem_4372_sv2v_reg ;
  assign \nz.mem [4371] = \nz.mem_4371_sv2v_reg ;
  assign \nz.mem [4370] = \nz.mem_4370_sv2v_reg ;
  assign \nz.mem [4369] = \nz.mem_4369_sv2v_reg ;
  assign \nz.mem [4368] = \nz.mem_4368_sv2v_reg ;
  assign \nz.mem [4367] = \nz.mem_4367_sv2v_reg ;
  assign \nz.mem [4366] = \nz.mem_4366_sv2v_reg ;
  assign \nz.mem [4365] = \nz.mem_4365_sv2v_reg ;
  assign \nz.mem [4364] = \nz.mem_4364_sv2v_reg ;
  assign \nz.mem [4363] = \nz.mem_4363_sv2v_reg ;
  assign \nz.mem [4362] = \nz.mem_4362_sv2v_reg ;
  assign \nz.mem [4361] = \nz.mem_4361_sv2v_reg ;
  assign \nz.mem [4360] = \nz.mem_4360_sv2v_reg ;
  assign \nz.mem [4359] = \nz.mem_4359_sv2v_reg ;
  assign \nz.mem [4358] = \nz.mem_4358_sv2v_reg ;
  assign \nz.mem [4357] = \nz.mem_4357_sv2v_reg ;
  assign \nz.mem [4356] = \nz.mem_4356_sv2v_reg ;
  assign \nz.mem [4355] = \nz.mem_4355_sv2v_reg ;
  assign \nz.mem [4354] = \nz.mem_4354_sv2v_reg ;
  assign \nz.mem [4353] = \nz.mem_4353_sv2v_reg ;
  assign \nz.mem [4352] = \nz.mem_4352_sv2v_reg ;
  assign \nz.mem [4351] = \nz.mem_4351_sv2v_reg ;
  assign \nz.mem [4350] = \nz.mem_4350_sv2v_reg ;
  assign \nz.mem [4349] = \nz.mem_4349_sv2v_reg ;
  assign \nz.mem [4348] = \nz.mem_4348_sv2v_reg ;
  assign \nz.mem [4347] = \nz.mem_4347_sv2v_reg ;
  assign \nz.mem [4346] = \nz.mem_4346_sv2v_reg ;
  assign \nz.mem [4345] = \nz.mem_4345_sv2v_reg ;
  assign \nz.mem [4344] = \nz.mem_4344_sv2v_reg ;
  assign \nz.mem [4343] = \nz.mem_4343_sv2v_reg ;
  assign \nz.mem [4342] = \nz.mem_4342_sv2v_reg ;
  assign \nz.mem [4341] = \nz.mem_4341_sv2v_reg ;
  assign \nz.mem [4340] = \nz.mem_4340_sv2v_reg ;
  assign \nz.mem [4339] = \nz.mem_4339_sv2v_reg ;
  assign \nz.mem [4338] = \nz.mem_4338_sv2v_reg ;
  assign \nz.mem [4337] = \nz.mem_4337_sv2v_reg ;
  assign \nz.mem [4336] = \nz.mem_4336_sv2v_reg ;
  assign \nz.mem [4335] = \nz.mem_4335_sv2v_reg ;
  assign \nz.mem [4334] = \nz.mem_4334_sv2v_reg ;
  assign \nz.mem [4333] = \nz.mem_4333_sv2v_reg ;
  assign \nz.mem [4332] = \nz.mem_4332_sv2v_reg ;
  assign \nz.mem [4331] = \nz.mem_4331_sv2v_reg ;
  assign \nz.mem [4330] = \nz.mem_4330_sv2v_reg ;
  assign \nz.mem [4329] = \nz.mem_4329_sv2v_reg ;
  assign \nz.mem [4328] = \nz.mem_4328_sv2v_reg ;
  assign \nz.mem [4327] = \nz.mem_4327_sv2v_reg ;
  assign \nz.mem [4326] = \nz.mem_4326_sv2v_reg ;
  assign \nz.mem [4325] = \nz.mem_4325_sv2v_reg ;
  assign \nz.mem [4324] = \nz.mem_4324_sv2v_reg ;
  assign \nz.mem [4323] = \nz.mem_4323_sv2v_reg ;
  assign \nz.mem [4322] = \nz.mem_4322_sv2v_reg ;
  assign \nz.mem [4321] = \nz.mem_4321_sv2v_reg ;
  assign \nz.mem [4320] = \nz.mem_4320_sv2v_reg ;
  assign \nz.mem [4319] = \nz.mem_4319_sv2v_reg ;
  assign \nz.mem [4318] = \nz.mem_4318_sv2v_reg ;
  assign \nz.mem [4317] = \nz.mem_4317_sv2v_reg ;
  assign \nz.mem [4316] = \nz.mem_4316_sv2v_reg ;
  assign \nz.mem [4315] = \nz.mem_4315_sv2v_reg ;
  assign \nz.mem [4314] = \nz.mem_4314_sv2v_reg ;
  assign \nz.mem [4313] = \nz.mem_4313_sv2v_reg ;
  assign \nz.mem [4312] = \nz.mem_4312_sv2v_reg ;
  assign \nz.mem [4311] = \nz.mem_4311_sv2v_reg ;
  assign \nz.mem [4310] = \nz.mem_4310_sv2v_reg ;
  assign \nz.mem [4309] = \nz.mem_4309_sv2v_reg ;
  assign \nz.mem [4308] = \nz.mem_4308_sv2v_reg ;
  assign \nz.mem [4307] = \nz.mem_4307_sv2v_reg ;
  assign \nz.mem [4306] = \nz.mem_4306_sv2v_reg ;
  assign \nz.mem [4305] = \nz.mem_4305_sv2v_reg ;
  assign \nz.mem [4304] = \nz.mem_4304_sv2v_reg ;
  assign \nz.mem [4303] = \nz.mem_4303_sv2v_reg ;
  assign \nz.mem [4302] = \nz.mem_4302_sv2v_reg ;
  assign \nz.mem [4301] = \nz.mem_4301_sv2v_reg ;
  assign \nz.mem [4300] = \nz.mem_4300_sv2v_reg ;
  assign \nz.mem [4299] = \nz.mem_4299_sv2v_reg ;
  assign \nz.mem [4298] = \nz.mem_4298_sv2v_reg ;
  assign \nz.mem [4297] = \nz.mem_4297_sv2v_reg ;
  assign \nz.mem [4296] = \nz.mem_4296_sv2v_reg ;
  assign \nz.mem [4295] = \nz.mem_4295_sv2v_reg ;
  assign \nz.mem [4294] = \nz.mem_4294_sv2v_reg ;
  assign \nz.mem [4293] = \nz.mem_4293_sv2v_reg ;
  assign \nz.mem [4292] = \nz.mem_4292_sv2v_reg ;
  assign \nz.mem [4291] = \nz.mem_4291_sv2v_reg ;
  assign \nz.mem [4290] = \nz.mem_4290_sv2v_reg ;
  assign \nz.mem [4289] = \nz.mem_4289_sv2v_reg ;
  assign \nz.mem [4288] = \nz.mem_4288_sv2v_reg ;
  assign \nz.mem [4287] = \nz.mem_4287_sv2v_reg ;
  assign \nz.mem [4286] = \nz.mem_4286_sv2v_reg ;
  assign \nz.mem [4285] = \nz.mem_4285_sv2v_reg ;
  assign \nz.mem [4284] = \nz.mem_4284_sv2v_reg ;
  assign \nz.mem [4283] = \nz.mem_4283_sv2v_reg ;
  assign \nz.mem [4282] = \nz.mem_4282_sv2v_reg ;
  assign \nz.mem [4281] = \nz.mem_4281_sv2v_reg ;
  assign \nz.mem [4280] = \nz.mem_4280_sv2v_reg ;
  assign \nz.mem [4279] = \nz.mem_4279_sv2v_reg ;
  assign \nz.mem [4278] = \nz.mem_4278_sv2v_reg ;
  assign \nz.mem [4277] = \nz.mem_4277_sv2v_reg ;
  assign \nz.mem [4276] = \nz.mem_4276_sv2v_reg ;
  assign \nz.mem [4275] = \nz.mem_4275_sv2v_reg ;
  assign \nz.mem [4274] = \nz.mem_4274_sv2v_reg ;
  assign \nz.mem [4273] = \nz.mem_4273_sv2v_reg ;
  assign \nz.mem [4272] = \nz.mem_4272_sv2v_reg ;
  assign \nz.mem [4271] = \nz.mem_4271_sv2v_reg ;
  assign \nz.mem [4270] = \nz.mem_4270_sv2v_reg ;
  assign \nz.mem [4269] = \nz.mem_4269_sv2v_reg ;
  assign \nz.mem [4268] = \nz.mem_4268_sv2v_reg ;
  assign \nz.mem [4267] = \nz.mem_4267_sv2v_reg ;
  assign \nz.mem [4266] = \nz.mem_4266_sv2v_reg ;
  assign \nz.mem [4265] = \nz.mem_4265_sv2v_reg ;
  assign \nz.mem [4264] = \nz.mem_4264_sv2v_reg ;
  assign \nz.mem [4263] = \nz.mem_4263_sv2v_reg ;
  assign \nz.mem [4262] = \nz.mem_4262_sv2v_reg ;
  assign \nz.mem [4261] = \nz.mem_4261_sv2v_reg ;
  assign \nz.mem [4260] = \nz.mem_4260_sv2v_reg ;
  assign \nz.mem [4259] = \nz.mem_4259_sv2v_reg ;
  assign \nz.mem [4258] = \nz.mem_4258_sv2v_reg ;
  assign \nz.mem [4257] = \nz.mem_4257_sv2v_reg ;
  assign \nz.mem [4256] = \nz.mem_4256_sv2v_reg ;
  assign \nz.mem [4255] = \nz.mem_4255_sv2v_reg ;
  assign \nz.mem [4254] = \nz.mem_4254_sv2v_reg ;
  assign \nz.mem [4253] = \nz.mem_4253_sv2v_reg ;
  assign \nz.mem [4252] = \nz.mem_4252_sv2v_reg ;
  assign \nz.mem [4251] = \nz.mem_4251_sv2v_reg ;
  assign \nz.mem [4250] = \nz.mem_4250_sv2v_reg ;
  assign \nz.mem [4249] = \nz.mem_4249_sv2v_reg ;
  assign \nz.mem [4248] = \nz.mem_4248_sv2v_reg ;
  assign \nz.mem [4247] = \nz.mem_4247_sv2v_reg ;
  assign \nz.mem [4246] = \nz.mem_4246_sv2v_reg ;
  assign \nz.mem [4245] = \nz.mem_4245_sv2v_reg ;
  assign \nz.mem [4244] = \nz.mem_4244_sv2v_reg ;
  assign \nz.mem [4243] = \nz.mem_4243_sv2v_reg ;
  assign \nz.mem [4242] = \nz.mem_4242_sv2v_reg ;
  assign \nz.mem [4241] = \nz.mem_4241_sv2v_reg ;
  assign \nz.mem [4240] = \nz.mem_4240_sv2v_reg ;
  assign \nz.mem [4239] = \nz.mem_4239_sv2v_reg ;
  assign \nz.mem [4238] = \nz.mem_4238_sv2v_reg ;
  assign \nz.mem [4237] = \nz.mem_4237_sv2v_reg ;
  assign \nz.mem [4236] = \nz.mem_4236_sv2v_reg ;
  assign \nz.mem [4235] = \nz.mem_4235_sv2v_reg ;
  assign \nz.mem [4234] = \nz.mem_4234_sv2v_reg ;
  assign \nz.mem [4233] = \nz.mem_4233_sv2v_reg ;
  assign \nz.mem [4232] = \nz.mem_4232_sv2v_reg ;
  assign \nz.mem [4231] = \nz.mem_4231_sv2v_reg ;
  assign \nz.mem [4230] = \nz.mem_4230_sv2v_reg ;
  assign \nz.mem [4229] = \nz.mem_4229_sv2v_reg ;
  assign \nz.mem [4228] = \nz.mem_4228_sv2v_reg ;
  assign \nz.mem [4227] = \nz.mem_4227_sv2v_reg ;
  assign \nz.mem [4226] = \nz.mem_4226_sv2v_reg ;
  assign \nz.mem [4225] = \nz.mem_4225_sv2v_reg ;
  assign \nz.mem [4224] = \nz.mem_4224_sv2v_reg ;
  assign \nz.mem [4223] = \nz.mem_4223_sv2v_reg ;
  assign \nz.mem [4222] = \nz.mem_4222_sv2v_reg ;
  assign \nz.mem [4221] = \nz.mem_4221_sv2v_reg ;
  assign \nz.mem [4220] = \nz.mem_4220_sv2v_reg ;
  assign \nz.mem [4219] = \nz.mem_4219_sv2v_reg ;
  assign \nz.mem [4218] = \nz.mem_4218_sv2v_reg ;
  assign \nz.mem [4217] = \nz.mem_4217_sv2v_reg ;
  assign \nz.mem [4216] = \nz.mem_4216_sv2v_reg ;
  assign \nz.mem [4215] = \nz.mem_4215_sv2v_reg ;
  assign \nz.mem [4214] = \nz.mem_4214_sv2v_reg ;
  assign \nz.mem [4213] = \nz.mem_4213_sv2v_reg ;
  assign \nz.mem [4212] = \nz.mem_4212_sv2v_reg ;
  assign \nz.mem [4211] = \nz.mem_4211_sv2v_reg ;
  assign \nz.mem [4210] = \nz.mem_4210_sv2v_reg ;
  assign \nz.mem [4209] = \nz.mem_4209_sv2v_reg ;
  assign \nz.mem [4208] = \nz.mem_4208_sv2v_reg ;
  assign \nz.mem [4207] = \nz.mem_4207_sv2v_reg ;
  assign \nz.mem [4206] = \nz.mem_4206_sv2v_reg ;
  assign \nz.mem [4205] = \nz.mem_4205_sv2v_reg ;
  assign \nz.mem [4204] = \nz.mem_4204_sv2v_reg ;
  assign \nz.mem [4203] = \nz.mem_4203_sv2v_reg ;
  assign \nz.mem [4202] = \nz.mem_4202_sv2v_reg ;
  assign \nz.mem [4201] = \nz.mem_4201_sv2v_reg ;
  assign \nz.mem [4200] = \nz.mem_4200_sv2v_reg ;
  assign \nz.mem [4199] = \nz.mem_4199_sv2v_reg ;
  assign \nz.mem [4198] = \nz.mem_4198_sv2v_reg ;
  assign \nz.mem [4197] = \nz.mem_4197_sv2v_reg ;
  assign \nz.mem [4196] = \nz.mem_4196_sv2v_reg ;
  assign \nz.mem [4195] = \nz.mem_4195_sv2v_reg ;
  assign \nz.mem [4194] = \nz.mem_4194_sv2v_reg ;
  assign \nz.mem [4193] = \nz.mem_4193_sv2v_reg ;
  assign \nz.mem [4192] = \nz.mem_4192_sv2v_reg ;
  assign \nz.mem [4191] = \nz.mem_4191_sv2v_reg ;
  assign \nz.mem [4190] = \nz.mem_4190_sv2v_reg ;
  assign \nz.mem [4189] = \nz.mem_4189_sv2v_reg ;
  assign \nz.mem [4188] = \nz.mem_4188_sv2v_reg ;
  assign \nz.mem [4187] = \nz.mem_4187_sv2v_reg ;
  assign \nz.mem [4186] = \nz.mem_4186_sv2v_reg ;
  assign \nz.mem [4185] = \nz.mem_4185_sv2v_reg ;
  assign \nz.mem [4184] = \nz.mem_4184_sv2v_reg ;
  assign \nz.mem [4183] = \nz.mem_4183_sv2v_reg ;
  assign \nz.mem [4182] = \nz.mem_4182_sv2v_reg ;
  assign \nz.mem [4181] = \nz.mem_4181_sv2v_reg ;
  assign \nz.mem [4180] = \nz.mem_4180_sv2v_reg ;
  assign \nz.mem [4179] = \nz.mem_4179_sv2v_reg ;
  assign \nz.mem [4178] = \nz.mem_4178_sv2v_reg ;
  assign \nz.mem [4177] = \nz.mem_4177_sv2v_reg ;
  assign \nz.mem [4176] = \nz.mem_4176_sv2v_reg ;
  assign \nz.mem [4175] = \nz.mem_4175_sv2v_reg ;
  assign \nz.mem [4174] = \nz.mem_4174_sv2v_reg ;
  assign \nz.mem [4173] = \nz.mem_4173_sv2v_reg ;
  assign \nz.mem [4172] = \nz.mem_4172_sv2v_reg ;
  assign \nz.mem [4171] = \nz.mem_4171_sv2v_reg ;
  assign \nz.mem [4170] = \nz.mem_4170_sv2v_reg ;
  assign \nz.mem [4169] = \nz.mem_4169_sv2v_reg ;
  assign \nz.mem [4168] = \nz.mem_4168_sv2v_reg ;
  assign \nz.mem [4167] = \nz.mem_4167_sv2v_reg ;
  assign \nz.mem [4166] = \nz.mem_4166_sv2v_reg ;
  assign \nz.mem [4165] = \nz.mem_4165_sv2v_reg ;
  assign \nz.mem [4164] = \nz.mem_4164_sv2v_reg ;
  assign \nz.mem [4163] = \nz.mem_4163_sv2v_reg ;
  assign \nz.mem [4162] = \nz.mem_4162_sv2v_reg ;
  assign \nz.mem [4161] = \nz.mem_4161_sv2v_reg ;
  assign \nz.mem [4160] = \nz.mem_4160_sv2v_reg ;
  assign \nz.mem [4159] = \nz.mem_4159_sv2v_reg ;
  assign \nz.mem [4158] = \nz.mem_4158_sv2v_reg ;
  assign \nz.mem [4157] = \nz.mem_4157_sv2v_reg ;
  assign \nz.mem [4156] = \nz.mem_4156_sv2v_reg ;
  assign \nz.mem [4155] = \nz.mem_4155_sv2v_reg ;
  assign \nz.mem [4154] = \nz.mem_4154_sv2v_reg ;
  assign \nz.mem [4153] = \nz.mem_4153_sv2v_reg ;
  assign \nz.mem [4152] = \nz.mem_4152_sv2v_reg ;
  assign \nz.mem [4151] = \nz.mem_4151_sv2v_reg ;
  assign \nz.mem [4150] = \nz.mem_4150_sv2v_reg ;
  assign \nz.mem [4149] = \nz.mem_4149_sv2v_reg ;
  assign \nz.mem [4148] = \nz.mem_4148_sv2v_reg ;
  assign \nz.mem [4147] = \nz.mem_4147_sv2v_reg ;
  assign \nz.mem [4146] = \nz.mem_4146_sv2v_reg ;
  assign \nz.mem [4145] = \nz.mem_4145_sv2v_reg ;
  assign \nz.mem [4144] = \nz.mem_4144_sv2v_reg ;
  assign \nz.mem [4143] = \nz.mem_4143_sv2v_reg ;
  assign \nz.mem [4142] = \nz.mem_4142_sv2v_reg ;
  assign \nz.mem [4141] = \nz.mem_4141_sv2v_reg ;
  assign \nz.mem [4140] = \nz.mem_4140_sv2v_reg ;
  assign \nz.mem [4139] = \nz.mem_4139_sv2v_reg ;
  assign \nz.mem [4138] = \nz.mem_4138_sv2v_reg ;
  assign \nz.mem [4137] = \nz.mem_4137_sv2v_reg ;
  assign \nz.mem [4136] = \nz.mem_4136_sv2v_reg ;
  assign \nz.mem [4135] = \nz.mem_4135_sv2v_reg ;
  assign \nz.mem [4134] = \nz.mem_4134_sv2v_reg ;
  assign \nz.mem [4133] = \nz.mem_4133_sv2v_reg ;
  assign \nz.mem [4132] = \nz.mem_4132_sv2v_reg ;
  assign \nz.mem [4131] = \nz.mem_4131_sv2v_reg ;
  assign \nz.mem [4130] = \nz.mem_4130_sv2v_reg ;
  assign \nz.mem [4129] = \nz.mem_4129_sv2v_reg ;
  assign \nz.mem [4128] = \nz.mem_4128_sv2v_reg ;
  assign \nz.mem [4127] = \nz.mem_4127_sv2v_reg ;
  assign \nz.mem [4126] = \nz.mem_4126_sv2v_reg ;
  assign \nz.mem [4125] = \nz.mem_4125_sv2v_reg ;
  assign \nz.mem [4124] = \nz.mem_4124_sv2v_reg ;
  assign \nz.mem [4123] = \nz.mem_4123_sv2v_reg ;
  assign \nz.mem [4122] = \nz.mem_4122_sv2v_reg ;
  assign \nz.mem [4121] = \nz.mem_4121_sv2v_reg ;
  assign \nz.mem [4120] = \nz.mem_4120_sv2v_reg ;
  assign \nz.mem [4119] = \nz.mem_4119_sv2v_reg ;
  assign \nz.mem [4118] = \nz.mem_4118_sv2v_reg ;
  assign \nz.mem [4117] = \nz.mem_4117_sv2v_reg ;
  assign \nz.mem [4116] = \nz.mem_4116_sv2v_reg ;
  assign \nz.mem [4115] = \nz.mem_4115_sv2v_reg ;
  assign \nz.mem [4114] = \nz.mem_4114_sv2v_reg ;
  assign \nz.mem [4113] = \nz.mem_4113_sv2v_reg ;
  assign \nz.mem [4112] = \nz.mem_4112_sv2v_reg ;
  assign \nz.mem [4111] = \nz.mem_4111_sv2v_reg ;
  assign \nz.mem [4110] = \nz.mem_4110_sv2v_reg ;
  assign \nz.mem [4109] = \nz.mem_4109_sv2v_reg ;
  assign \nz.mem [4108] = \nz.mem_4108_sv2v_reg ;
  assign \nz.mem [4107] = \nz.mem_4107_sv2v_reg ;
  assign \nz.mem [4106] = \nz.mem_4106_sv2v_reg ;
  assign \nz.mem [4105] = \nz.mem_4105_sv2v_reg ;
  assign \nz.mem [4104] = \nz.mem_4104_sv2v_reg ;
  assign \nz.mem [4103] = \nz.mem_4103_sv2v_reg ;
  assign \nz.mem [4102] = \nz.mem_4102_sv2v_reg ;
  assign \nz.mem [4101] = \nz.mem_4101_sv2v_reg ;
  assign \nz.mem [4100] = \nz.mem_4100_sv2v_reg ;
  assign \nz.mem [4099] = \nz.mem_4099_sv2v_reg ;
  assign \nz.mem [4098] = \nz.mem_4098_sv2v_reg ;
  assign \nz.mem [4097] = \nz.mem_4097_sv2v_reg ;
  assign \nz.mem [4096] = \nz.mem_4096_sv2v_reg ;
  assign \nz.mem [4095] = \nz.mem_4095_sv2v_reg ;
  assign \nz.mem [4094] = \nz.mem_4094_sv2v_reg ;
  assign \nz.mem [4093] = \nz.mem_4093_sv2v_reg ;
  assign \nz.mem [4092] = \nz.mem_4092_sv2v_reg ;
  assign \nz.mem [4091] = \nz.mem_4091_sv2v_reg ;
  assign \nz.mem [4090] = \nz.mem_4090_sv2v_reg ;
  assign \nz.mem [4089] = \nz.mem_4089_sv2v_reg ;
  assign \nz.mem [4088] = \nz.mem_4088_sv2v_reg ;
  assign \nz.mem [4087] = \nz.mem_4087_sv2v_reg ;
  assign \nz.mem [4086] = \nz.mem_4086_sv2v_reg ;
  assign \nz.mem [4085] = \nz.mem_4085_sv2v_reg ;
  assign \nz.mem [4084] = \nz.mem_4084_sv2v_reg ;
  assign \nz.mem [4083] = \nz.mem_4083_sv2v_reg ;
  assign \nz.mem [4082] = \nz.mem_4082_sv2v_reg ;
  assign \nz.mem [4081] = \nz.mem_4081_sv2v_reg ;
  assign \nz.mem [4080] = \nz.mem_4080_sv2v_reg ;
  assign \nz.mem [4079] = \nz.mem_4079_sv2v_reg ;
  assign \nz.mem [4078] = \nz.mem_4078_sv2v_reg ;
  assign \nz.mem [4077] = \nz.mem_4077_sv2v_reg ;
  assign \nz.mem [4076] = \nz.mem_4076_sv2v_reg ;
  assign \nz.mem [4075] = \nz.mem_4075_sv2v_reg ;
  assign \nz.mem [4074] = \nz.mem_4074_sv2v_reg ;
  assign \nz.mem [4073] = \nz.mem_4073_sv2v_reg ;
  assign \nz.mem [4072] = \nz.mem_4072_sv2v_reg ;
  assign \nz.mem [4071] = \nz.mem_4071_sv2v_reg ;
  assign \nz.mem [4070] = \nz.mem_4070_sv2v_reg ;
  assign \nz.mem [4069] = \nz.mem_4069_sv2v_reg ;
  assign \nz.mem [4068] = \nz.mem_4068_sv2v_reg ;
  assign \nz.mem [4067] = \nz.mem_4067_sv2v_reg ;
  assign \nz.mem [4066] = \nz.mem_4066_sv2v_reg ;
  assign \nz.mem [4065] = \nz.mem_4065_sv2v_reg ;
  assign \nz.mem [4064] = \nz.mem_4064_sv2v_reg ;
  assign \nz.mem [4063] = \nz.mem_4063_sv2v_reg ;
  assign \nz.mem [4062] = \nz.mem_4062_sv2v_reg ;
  assign \nz.mem [4061] = \nz.mem_4061_sv2v_reg ;
  assign \nz.mem [4060] = \nz.mem_4060_sv2v_reg ;
  assign \nz.mem [4059] = \nz.mem_4059_sv2v_reg ;
  assign \nz.mem [4058] = \nz.mem_4058_sv2v_reg ;
  assign \nz.mem [4057] = \nz.mem_4057_sv2v_reg ;
  assign \nz.mem [4056] = \nz.mem_4056_sv2v_reg ;
  assign \nz.mem [4055] = \nz.mem_4055_sv2v_reg ;
  assign \nz.mem [4054] = \nz.mem_4054_sv2v_reg ;
  assign \nz.mem [4053] = \nz.mem_4053_sv2v_reg ;
  assign \nz.mem [4052] = \nz.mem_4052_sv2v_reg ;
  assign \nz.mem [4051] = \nz.mem_4051_sv2v_reg ;
  assign \nz.mem [4050] = \nz.mem_4050_sv2v_reg ;
  assign \nz.mem [4049] = \nz.mem_4049_sv2v_reg ;
  assign \nz.mem [4048] = \nz.mem_4048_sv2v_reg ;
  assign \nz.mem [4047] = \nz.mem_4047_sv2v_reg ;
  assign \nz.mem [4046] = \nz.mem_4046_sv2v_reg ;
  assign \nz.mem [4045] = \nz.mem_4045_sv2v_reg ;
  assign \nz.mem [4044] = \nz.mem_4044_sv2v_reg ;
  assign \nz.mem [4043] = \nz.mem_4043_sv2v_reg ;
  assign \nz.mem [4042] = \nz.mem_4042_sv2v_reg ;
  assign \nz.mem [4041] = \nz.mem_4041_sv2v_reg ;
  assign \nz.mem [4040] = \nz.mem_4040_sv2v_reg ;
  assign \nz.mem [4039] = \nz.mem_4039_sv2v_reg ;
  assign \nz.mem [4038] = \nz.mem_4038_sv2v_reg ;
  assign \nz.mem [4037] = \nz.mem_4037_sv2v_reg ;
  assign \nz.mem [4036] = \nz.mem_4036_sv2v_reg ;
  assign \nz.mem [4035] = \nz.mem_4035_sv2v_reg ;
  assign \nz.mem [4034] = \nz.mem_4034_sv2v_reg ;
  assign \nz.mem [4033] = \nz.mem_4033_sv2v_reg ;
  assign \nz.mem [4032] = \nz.mem_4032_sv2v_reg ;
  assign \nz.mem [4031] = \nz.mem_4031_sv2v_reg ;
  assign \nz.mem [4030] = \nz.mem_4030_sv2v_reg ;
  assign \nz.mem [4029] = \nz.mem_4029_sv2v_reg ;
  assign \nz.mem [4028] = \nz.mem_4028_sv2v_reg ;
  assign \nz.mem [4027] = \nz.mem_4027_sv2v_reg ;
  assign \nz.mem [4026] = \nz.mem_4026_sv2v_reg ;
  assign \nz.mem [4025] = \nz.mem_4025_sv2v_reg ;
  assign \nz.mem [4024] = \nz.mem_4024_sv2v_reg ;
  assign \nz.mem [4023] = \nz.mem_4023_sv2v_reg ;
  assign \nz.mem [4022] = \nz.mem_4022_sv2v_reg ;
  assign \nz.mem [4021] = \nz.mem_4021_sv2v_reg ;
  assign \nz.mem [4020] = \nz.mem_4020_sv2v_reg ;
  assign \nz.mem [4019] = \nz.mem_4019_sv2v_reg ;
  assign \nz.mem [4018] = \nz.mem_4018_sv2v_reg ;
  assign \nz.mem [4017] = \nz.mem_4017_sv2v_reg ;
  assign \nz.mem [4016] = \nz.mem_4016_sv2v_reg ;
  assign \nz.mem [4015] = \nz.mem_4015_sv2v_reg ;
  assign \nz.mem [4014] = \nz.mem_4014_sv2v_reg ;
  assign \nz.mem [4013] = \nz.mem_4013_sv2v_reg ;
  assign \nz.mem [4012] = \nz.mem_4012_sv2v_reg ;
  assign \nz.mem [4011] = \nz.mem_4011_sv2v_reg ;
  assign \nz.mem [4010] = \nz.mem_4010_sv2v_reg ;
  assign \nz.mem [4009] = \nz.mem_4009_sv2v_reg ;
  assign \nz.mem [4008] = \nz.mem_4008_sv2v_reg ;
  assign \nz.mem [4007] = \nz.mem_4007_sv2v_reg ;
  assign \nz.mem [4006] = \nz.mem_4006_sv2v_reg ;
  assign \nz.mem [4005] = \nz.mem_4005_sv2v_reg ;
  assign \nz.mem [4004] = \nz.mem_4004_sv2v_reg ;
  assign \nz.mem [4003] = \nz.mem_4003_sv2v_reg ;
  assign \nz.mem [4002] = \nz.mem_4002_sv2v_reg ;
  assign \nz.mem [4001] = \nz.mem_4001_sv2v_reg ;
  assign \nz.mem [4000] = \nz.mem_4000_sv2v_reg ;
  assign \nz.mem [3999] = \nz.mem_3999_sv2v_reg ;
  assign \nz.mem [3998] = \nz.mem_3998_sv2v_reg ;
  assign \nz.mem [3997] = \nz.mem_3997_sv2v_reg ;
  assign \nz.mem [3996] = \nz.mem_3996_sv2v_reg ;
  assign \nz.mem [3995] = \nz.mem_3995_sv2v_reg ;
  assign \nz.mem [3994] = \nz.mem_3994_sv2v_reg ;
  assign \nz.mem [3993] = \nz.mem_3993_sv2v_reg ;
  assign \nz.mem [3992] = \nz.mem_3992_sv2v_reg ;
  assign \nz.mem [3991] = \nz.mem_3991_sv2v_reg ;
  assign \nz.mem [3990] = \nz.mem_3990_sv2v_reg ;
  assign \nz.mem [3989] = \nz.mem_3989_sv2v_reg ;
  assign \nz.mem [3988] = \nz.mem_3988_sv2v_reg ;
  assign \nz.mem [3987] = \nz.mem_3987_sv2v_reg ;
  assign \nz.mem [3986] = \nz.mem_3986_sv2v_reg ;
  assign \nz.mem [3985] = \nz.mem_3985_sv2v_reg ;
  assign \nz.mem [3984] = \nz.mem_3984_sv2v_reg ;
  assign \nz.mem [3983] = \nz.mem_3983_sv2v_reg ;
  assign \nz.mem [3982] = \nz.mem_3982_sv2v_reg ;
  assign \nz.mem [3981] = \nz.mem_3981_sv2v_reg ;
  assign \nz.mem [3980] = \nz.mem_3980_sv2v_reg ;
  assign \nz.mem [3979] = \nz.mem_3979_sv2v_reg ;
  assign \nz.mem [3978] = \nz.mem_3978_sv2v_reg ;
  assign \nz.mem [3977] = \nz.mem_3977_sv2v_reg ;
  assign \nz.mem [3976] = \nz.mem_3976_sv2v_reg ;
  assign \nz.mem [3975] = \nz.mem_3975_sv2v_reg ;
  assign \nz.mem [3974] = \nz.mem_3974_sv2v_reg ;
  assign \nz.mem [3973] = \nz.mem_3973_sv2v_reg ;
  assign \nz.mem [3972] = \nz.mem_3972_sv2v_reg ;
  assign \nz.mem [3971] = \nz.mem_3971_sv2v_reg ;
  assign \nz.mem [3970] = \nz.mem_3970_sv2v_reg ;
  assign \nz.mem [3969] = \nz.mem_3969_sv2v_reg ;
  assign \nz.mem [3968] = \nz.mem_3968_sv2v_reg ;
  assign \nz.mem [3967] = \nz.mem_3967_sv2v_reg ;
  assign \nz.mem [3966] = \nz.mem_3966_sv2v_reg ;
  assign \nz.mem [3965] = \nz.mem_3965_sv2v_reg ;
  assign \nz.mem [3964] = \nz.mem_3964_sv2v_reg ;
  assign \nz.mem [3963] = \nz.mem_3963_sv2v_reg ;
  assign \nz.mem [3962] = \nz.mem_3962_sv2v_reg ;
  assign \nz.mem [3961] = \nz.mem_3961_sv2v_reg ;
  assign \nz.mem [3960] = \nz.mem_3960_sv2v_reg ;
  assign \nz.mem [3959] = \nz.mem_3959_sv2v_reg ;
  assign \nz.mem [3958] = \nz.mem_3958_sv2v_reg ;
  assign \nz.mem [3957] = \nz.mem_3957_sv2v_reg ;
  assign \nz.mem [3956] = \nz.mem_3956_sv2v_reg ;
  assign \nz.mem [3955] = \nz.mem_3955_sv2v_reg ;
  assign \nz.mem [3954] = \nz.mem_3954_sv2v_reg ;
  assign \nz.mem [3953] = \nz.mem_3953_sv2v_reg ;
  assign \nz.mem [3952] = \nz.mem_3952_sv2v_reg ;
  assign \nz.mem [3951] = \nz.mem_3951_sv2v_reg ;
  assign \nz.mem [3950] = \nz.mem_3950_sv2v_reg ;
  assign \nz.mem [3949] = \nz.mem_3949_sv2v_reg ;
  assign \nz.mem [3948] = \nz.mem_3948_sv2v_reg ;
  assign \nz.mem [3947] = \nz.mem_3947_sv2v_reg ;
  assign \nz.mem [3946] = \nz.mem_3946_sv2v_reg ;
  assign \nz.mem [3945] = \nz.mem_3945_sv2v_reg ;
  assign \nz.mem [3944] = \nz.mem_3944_sv2v_reg ;
  assign \nz.mem [3943] = \nz.mem_3943_sv2v_reg ;
  assign \nz.mem [3942] = \nz.mem_3942_sv2v_reg ;
  assign \nz.mem [3941] = \nz.mem_3941_sv2v_reg ;
  assign \nz.mem [3940] = \nz.mem_3940_sv2v_reg ;
  assign \nz.mem [3939] = \nz.mem_3939_sv2v_reg ;
  assign \nz.mem [3938] = \nz.mem_3938_sv2v_reg ;
  assign \nz.mem [3937] = \nz.mem_3937_sv2v_reg ;
  assign \nz.mem [3936] = \nz.mem_3936_sv2v_reg ;
  assign \nz.mem [3935] = \nz.mem_3935_sv2v_reg ;
  assign \nz.mem [3934] = \nz.mem_3934_sv2v_reg ;
  assign \nz.mem [3933] = \nz.mem_3933_sv2v_reg ;
  assign \nz.mem [3932] = \nz.mem_3932_sv2v_reg ;
  assign \nz.mem [3931] = \nz.mem_3931_sv2v_reg ;
  assign \nz.mem [3930] = \nz.mem_3930_sv2v_reg ;
  assign \nz.mem [3929] = \nz.mem_3929_sv2v_reg ;
  assign \nz.mem [3928] = \nz.mem_3928_sv2v_reg ;
  assign \nz.mem [3927] = \nz.mem_3927_sv2v_reg ;
  assign \nz.mem [3926] = \nz.mem_3926_sv2v_reg ;
  assign \nz.mem [3925] = \nz.mem_3925_sv2v_reg ;
  assign \nz.mem [3924] = \nz.mem_3924_sv2v_reg ;
  assign \nz.mem [3923] = \nz.mem_3923_sv2v_reg ;
  assign \nz.mem [3922] = \nz.mem_3922_sv2v_reg ;
  assign \nz.mem [3921] = \nz.mem_3921_sv2v_reg ;
  assign \nz.mem [3920] = \nz.mem_3920_sv2v_reg ;
  assign \nz.mem [3919] = \nz.mem_3919_sv2v_reg ;
  assign \nz.mem [3918] = \nz.mem_3918_sv2v_reg ;
  assign \nz.mem [3917] = \nz.mem_3917_sv2v_reg ;
  assign \nz.mem [3916] = \nz.mem_3916_sv2v_reg ;
  assign \nz.mem [3915] = \nz.mem_3915_sv2v_reg ;
  assign \nz.mem [3914] = \nz.mem_3914_sv2v_reg ;
  assign \nz.mem [3913] = \nz.mem_3913_sv2v_reg ;
  assign \nz.mem [3912] = \nz.mem_3912_sv2v_reg ;
  assign \nz.mem [3911] = \nz.mem_3911_sv2v_reg ;
  assign \nz.mem [3910] = \nz.mem_3910_sv2v_reg ;
  assign \nz.mem [3909] = \nz.mem_3909_sv2v_reg ;
  assign \nz.mem [3908] = \nz.mem_3908_sv2v_reg ;
  assign \nz.mem [3907] = \nz.mem_3907_sv2v_reg ;
  assign \nz.mem [3906] = \nz.mem_3906_sv2v_reg ;
  assign \nz.mem [3905] = \nz.mem_3905_sv2v_reg ;
  assign \nz.mem [3904] = \nz.mem_3904_sv2v_reg ;
  assign \nz.mem [3903] = \nz.mem_3903_sv2v_reg ;
  assign \nz.mem [3902] = \nz.mem_3902_sv2v_reg ;
  assign \nz.mem [3901] = \nz.mem_3901_sv2v_reg ;
  assign \nz.mem [3900] = \nz.mem_3900_sv2v_reg ;
  assign \nz.mem [3899] = \nz.mem_3899_sv2v_reg ;
  assign \nz.mem [3898] = \nz.mem_3898_sv2v_reg ;
  assign \nz.mem [3897] = \nz.mem_3897_sv2v_reg ;
  assign \nz.mem [3896] = \nz.mem_3896_sv2v_reg ;
  assign \nz.mem [3895] = \nz.mem_3895_sv2v_reg ;
  assign \nz.mem [3894] = \nz.mem_3894_sv2v_reg ;
  assign \nz.mem [3893] = \nz.mem_3893_sv2v_reg ;
  assign \nz.mem [3892] = \nz.mem_3892_sv2v_reg ;
  assign \nz.mem [3891] = \nz.mem_3891_sv2v_reg ;
  assign \nz.mem [3890] = \nz.mem_3890_sv2v_reg ;
  assign \nz.mem [3889] = \nz.mem_3889_sv2v_reg ;
  assign \nz.mem [3888] = \nz.mem_3888_sv2v_reg ;
  assign \nz.mem [3887] = \nz.mem_3887_sv2v_reg ;
  assign \nz.mem [3886] = \nz.mem_3886_sv2v_reg ;
  assign \nz.mem [3885] = \nz.mem_3885_sv2v_reg ;
  assign \nz.mem [3884] = \nz.mem_3884_sv2v_reg ;
  assign \nz.mem [3883] = \nz.mem_3883_sv2v_reg ;
  assign \nz.mem [3882] = \nz.mem_3882_sv2v_reg ;
  assign \nz.mem [3881] = \nz.mem_3881_sv2v_reg ;
  assign \nz.mem [3880] = \nz.mem_3880_sv2v_reg ;
  assign \nz.mem [3879] = \nz.mem_3879_sv2v_reg ;
  assign \nz.mem [3878] = \nz.mem_3878_sv2v_reg ;
  assign \nz.mem [3877] = \nz.mem_3877_sv2v_reg ;
  assign \nz.mem [3876] = \nz.mem_3876_sv2v_reg ;
  assign \nz.mem [3875] = \nz.mem_3875_sv2v_reg ;
  assign \nz.mem [3874] = \nz.mem_3874_sv2v_reg ;
  assign \nz.mem [3873] = \nz.mem_3873_sv2v_reg ;
  assign \nz.mem [3872] = \nz.mem_3872_sv2v_reg ;
  assign \nz.mem [3871] = \nz.mem_3871_sv2v_reg ;
  assign \nz.mem [3870] = \nz.mem_3870_sv2v_reg ;
  assign \nz.mem [3869] = \nz.mem_3869_sv2v_reg ;
  assign \nz.mem [3868] = \nz.mem_3868_sv2v_reg ;
  assign \nz.mem [3867] = \nz.mem_3867_sv2v_reg ;
  assign \nz.mem [3866] = \nz.mem_3866_sv2v_reg ;
  assign \nz.mem [3865] = \nz.mem_3865_sv2v_reg ;
  assign \nz.mem [3864] = \nz.mem_3864_sv2v_reg ;
  assign \nz.mem [3863] = \nz.mem_3863_sv2v_reg ;
  assign \nz.mem [3862] = \nz.mem_3862_sv2v_reg ;
  assign \nz.mem [3861] = \nz.mem_3861_sv2v_reg ;
  assign \nz.mem [3860] = \nz.mem_3860_sv2v_reg ;
  assign \nz.mem [3859] = \nz.mem_3859_sv2v_reg ;
  assign \nz.mem [3858] = \nz.mem_3858_sv2v_reg ;
  assign \nz.mem [3857] = \nz.mem_3857_sv2v_reg ;
  assign \nz.mem [3856] = \nz.mem_3856_sv2v_reg ;
  assign \nz.mem [3855] = \nz.mem_3855_sv2v_reg ;
  assign \nz.mem [3854] = \nz.mem_3854_sv2v_reg ;
  assign \nz.mem [3853] = \nz.mem_3853_sv2v_reg ;
  assign \nz.mem [3852] = \nz.mem_3852_sv2v_reg ;
  assign \nz.mem [3851] = \nz.mem_3851_sv2v_reg ;
  assign \nz.mem [3850] = \nz.mem_3850_sv2v_reg ;
  assign \nz.mem [3849] = \nz.mem_3849_sv2v_reg ;
  assign \nz.mem [3848] = \nz.mem_3848_sv2v_reg ;
  assign \nz.mem [3847] = \nz.mem_3847_sv2v_reg ;
  assign \nz.mem [3846] = \nz.mem_3846_sv2v_reg ;
  assign \nz.mem [3845] = \nz.mem_3845_sv2v_reg ;
  assign \nz.mem [3844] = \nz.mem_3844_sv2v_reg ;
  assign \nz.mem [3843] = \nz.mem_3843_sv2v_reg ;
  assign \nz.mem [3842] = \nz.mem_3842_sv2v_reg ;
  assign \nz.mem [3841] = \nz.mem_3841_sv2v_reg ;
  assign \nz.mem [3840] = \nz.mem_3840_sv2v_reg ;
  assign \nz.mem [3839] = \nz.mem_3839_sv2v_reg ;
  assign \nz.mem [3838] = \nz.mem_3838_sv2v_reg ;
  assign \nz.mem [3837] = \nz.mem_3837_sv2v_reg ;
  assign \nz.mem [3836] = \nz.mem_3836_sv2v_reg ;
  assign \nz.mem [3835] = \nz.mem_3835_sv2v_reg ;
  assign \nz.mem [3834] = \nz.mem_3834_sv2v_reg ;
  assign \nz.mem [3833] = \nz.mem_3833_sv2v_reg ;
  assign \nz.mem [3832] = \nz.mem_3832_sv2v_reg ;
  assign \nz.mem [3831] = \nz.mem_3831_sv2v_reg ;
  assign \nz.mem [3830] = \nz.mem_3830_sv2v_reg ;
  assign \nz.mem [3829] = \nz.mem_3829_sv2v_reg ;
  assign \nz.mem [3828] = \nz.mem_3828_sv2v_reg ;
  assign \nz.mem [3827] = \nz.mem_3827_sv2v_reg ;
  assign \nz.mem [3826] = \nz.mem_3826_sv2v_reg ;
  assign \nz.mem [3825] = \nz.mem_3825_sv2v_reg ;
  assign \nz.mem [3824] = \nz.mem_3824_sv2v_reg ;
  assign \nz.mem [3823] = \nz.mem_3823_sv2v_reg ;
  assign \nz.mem [3822] = \nz.mem_3822_sv2v_reg ;
  assign \nz.mem [3821] = \nz.mem_3821_sv2v_reg ;
  assign \nz.mem [3820] = \nz.mem_3820_sv2v_reg ;
  assign \nz.mem [3819] = \nz.mem_3819_sv2v_reg ;
  assign \nz.mem [3818] = \nz.mem_3818_sv2v_reg ;
  assign \nz.mem [3817] = \nz.mem_3817_sv2v_reg ;
  assign \nz.mem [3816] = \nz.mem_3816_sv2v_reg ;
  assign \nz.mem [3815] = \nz.mem_3815_sv2v_reg ;
  assign \nz.mem [3814] = \nz.mem_3814_sv2v_reg ;
  assign \nz.mem [3813] = \nz.mem_3813_sv2v_reg ;
  assign \nz.mem [3812] = \nz.mem_3812_sv2v_reg ;
  assign \nz.mem [3811] = \nz.mem_3811_sv2v_reg ;
  assign \nz.mem [3810] = \nz.mem_3810_sv2v_reg ;
  assign \nz.mem [3809] = \nz.mem_3809_sv2v_reg ;
  assign \nz.mem [3808] = \nz.mem_3808_sv2v_reg ;
  assign \nz.mem [3807] = \nz.mem_3807_sv2v_reg ;
  assign \nz.mem [3806] = \nz.mem_3806_sv2v_reg ;
  assign \nz.mem [3805] = \nz.mem_3805_sv2v_reg ;
  assign \nz.mem [3804] = \nz.mem_3804_sv2v_reg ;
  assign \nz.mem [3803] = \nz.mem_3803_sv2v_reg ;
  assign \nz.mem [3802] = \nz.mem_3802_sv2v_reg ;
  assign \nz.mem [3801] = \nz.mem_3801_sv2v_reg ;
  assign \nz.mem [3800] = \nz.mem_3800_sv2v_reg ;
  assign \nz.mem [3799] = \nz.mem_3799_sv2v_reg ;
  assign \nz.mem [3798] = \nz.mem_3798_sv2v_reg ;
  assign \nz.mem [3797] = \nz.mem_3797_sv2v_reg ;
  assign \nz.mem [3796] = \nz.mem_3796_sv2v_reg ;
  assign \nz.mem [3795] = \nz.mem_3795_sv2v_reg ;
  assign \nz.mem [3794] = \nz.mem_3794_sv2v_reg ;
  assign \nz.mem [3793] = \nz.mem_3793_sv2v_reg ;
  assign \nz.mem [3792] = \nz.mem_3792_sv2v_reg ;
  assign \nz.mem [3791] = \nz.mem_3791_sv2v_reg ;
  assign \nz.mem [3790] = \nz.mem_3790_sv2v_reg ;
  assign \nz.mem [3789] = \nz.mem_3789_sv2v_reg ;
  assign \nz.mem [3788] = \nz.mem_3788_sv2v_reg ;
  assign \nz.mem [3787] = \nz.mem_3787_sv2v_reg ;
  assign \nz.mem [3786] = \nz.mem_3786_sv2v_reg ;
  assign \nz.mem [3785] = \nz.mem_3785_sv2v_reg ;
  assign \nz.mem [3784] = \nz.mem_3784_sv2v_reg ;
  assign \nz.mem [3783] = \nz.mem_3783_sv2v_reg ;
  assign \nz.mem [3782] = \nz.mem_3782_sv2v_reg ;
  assign \nz.mem [3781] = \nz.mem_3781_sv2v_reg ;
  assign \nz.mem [3780] = \nz.mem_3780_sv2v_reg ;
  assign \nz.mem [3779] = \nz.mem_3779_sv2v_reg ;
  assign \nz.mem [3778] = \nz.mem_3778_sv2v_reg ;
  assign \nz.mem [3777] = \nz.mem_3777_sv2v_reg ;
  assign \nz.mem [3776] = \nz.mem_3776_sv2v_reg ;
  assign \nz.mem [3775] = \nz.mem_3775_sv2v_reg ;
  assign \nz.mem [3774] = \nz.mem_3774_sv2v_reg ;
  assign \nz.mem [3773] = \nz.mem_3773_sv2v_reg ;
  assign \nz.mem [3772] = \nz.mem_3772_sv2v_reg ;
  assign \nz.mem [3771] = \nz.mem_3771_sv2v_reg ;
  assign \nz.mem [3770] = \nz.mem_3770_sv2v_reg ;
  assign \nz.mem [3769] = \nz.mem_3769_sv2v_reg ;
  assign \nz.mem [3768] = \nz.mem_3768_sv2v_reg ;
  assign \nz.mem [3767] = \nz.mem_3767_sv2v_reg ;
  assign \nz.mem [3766] = \nz.mem_3766_sv2v_reg ;
  assign \nz.mem [3765] = \nz.mem_3765_sv2v_reg ;
  assign \nz.mem [3764] = \nz.mem_3764_sv2v_reg ;
  assign \nz.mem [3763] = \nz.mem_3763_sv2v_reg ;
  assign \nz.mem [3762] = \nz.mem_3762_sv2v_reg ;
  assign \nz.mem [3761] = \nz.mem_3761_sv2v_reg ;
  assign \nz.mem [3760] = \nz.mem_3760_sv2v_reg ;
  assign \nz.mem [3759] = \nz.mem_3759_sv2v_reg ;
  assign \nz.mem [3758] = \nz.mem_3758_sv2v_reg ;
  assign \nz.mem [3757] = \nz.mem_3757_sv2v_reg ;
  assign \nz.mem [3756] = \nz.mem_3756_sv2v_reg ;
  assign \nz.mem [3755] = \nz.mem_3755_sv2v_reg ;
  assign \nz.mem [3754] = \nz.mem_3754_sv2v_reg ;
  assign \nz.mem [3753] = \nz.mem_3753_sv2v_reg ;
  assign \nz.mem [3752] = \nz.mem_3752_sv2v_reg ;
  assign \nz.mem [3751] = \nz.mem_3751_sv2v_reg ;
  assign \nz.mem [3750] = \nz.mem_3750_sv2v_reg ;
  assign \nz.mem [3749] = \nz.mem_3749_sv2v_reg ;
  assign \nz.mem [3748] = \nz.mem_3748_sv2v_reg ;
  assign \nz.mem [3747] = \nz.mem_3747_sv2v_reg ;
  assign \nz.mem [3746] = \nz.mem_3746_sv2v_reg ;
  assign \nz.mem [3745] = \nz.mem_3745_sv2v_reg ;
  assign \nz.mem [3744] = \nz.mem_3744_sv2v_reg ;
  assign \nz.mem [3743] = \nz.mem_3743_sv2v_reg ;
  assign \nz.mem [3742] = \nz.mem_3742_sv2v_reg ;
  assign \nz.mem [3741] = \nz.mem_3741_sv2v_reg ;
  assign \nz.mem [3740] = \nz.mem_3740_sv2v_reg ;
  assign \nz.mem [3739] = \nz.mem_3739_sv2v_reg ;
  assign \nz.mem [3738] = \nz.mem_3738_sv2v_reg ;
  assign \nz.mem [3737] = \nz.mem_3737_sv2v_reg ;
  assign \nz.mem [3736] = \nz.mem_3736_sv2v_reg ;
  assign \nz.mem [3735] = \nz.mem_3735_sv2v_reg ;
  assign \nz.mem [3734] = \nz.mem_3734_sv2v_reg ;
  assign \nz.mem [3733] = \nz.mem_3733_sv2v_reg ;
  assign \nz.mem [3732] = \nz.mem_3732_sv2v_reg ;
  assign \nz.mem [3731] = \nz.mem_3731_sv2v_reg ;
  assign \nz.mem [3730] = \nz.mem_3730_sv2v_reg ;
  assign \nz.mem [3729] = \nz.mem_3729_sv2v_reg ;
  assign \nz.mem [3728] = \nz.mem_3728_sv2v_reg ;
  assign \nz.mem [3727] = \nz.mem_3727_sv2v_reg ;
  assign \nz.mem [3726] = \nz.mem_3726_sv2v_reg ;
  assign \nz.mem [3725] = \nz.mem_3725_sv2v_reg ;
  assign \nz.mem [3724] = \nz.mem_3724_sv2v_reg ;
  assign \nz.mem [3723] = \nz.mem_3723_sv2v_reg ;
  assign \nz.mem [3722] = \nz.mem_3722_sv2v_reg ;
  assign \nz.mem [3721] = \nz.mem_3721_sv2v_reg ;
  assign \nz.mem [3720] = \nz.mem_3720_sv2v_reg ;
  assign \nz.mem [3719] = \nz.mem_3719_sv2v_reg ;
  assign \nz.mem [3718] = \nz.mem_3718_sv2v_reg ;
  assign \nz.mem [3717] = \nz.mem_3717_sv2v_reg ;
  assign \nz.mem [3716] = \nz.mem_3716_sv2v_reg ;
  assign \nz.mem [3715] = \nz.mem_3715_sv2v_reg ;
  assign \nz.mem [3714] = \nz.mem_3714_sv2v_reg ;
  assign \nz.mem [3713] = \nz.mem_3713_sv2v_reg ;
  assign \nz.mem [3712] = \nz.mem_3712_sv2v_reg ;
  assign \nz.mem [3711] = \nz.mem_3711_sv2v_reg ;
  assign \nz.mem [3710] = \nz.mem_3710_sv2v_reg ;
  assign \nz.mem [3709] = \nz.mem_3709_sv2v_reg ;
  assign \nz.mem [3708] = \nz.mem_3708_sv2v_reg ;
  assign \nz.mem [3707] = \nz.mem_3707_sv2v_reg ;
  assign \nz.mem [3706] = \nz.mem_3706_sv2v_reg ;
  assign \nz.mem [3705] = \nz.mem_3705_sv2v_reg ;
  assign \nz.mem [3704] = \nz.mem_3704_sv2v_reg ;
  assign \nz.mem [3703] = \nz.mem_3703_sv2v_reg ;
  assign \nz.mem [3702] = \nz.mem_3702_sv2v_reg ;
  assign \nz.mem [3701] = \nz.mem_3701_sv2v_reg ;
  assign \nz.mem [3700] = \nz.mem_3700_sv2v_reg ;
  assign \nz.mem [3699] = \nz.mem_3699_sv2v_reg ;
  assign \nz.mem [3698] = \nz.mem_3698_sv2v_reg ;
  assign \nz.mem [3697] = \nz.mem_3697_sv2v_reg ;
  assign \nz.mem [3696] = \nz.mem_3696_sv2v_reg ;
  assign \nz.mem [3695] = \nz.mem_3695_sv2v_reg ;
  assign \nz.mem [3694] = \nz.mem_3694_sv2v_reg ;
  assign \nz.mem [3693] = \nz.mem_3693_sv2v_reg ;
  assign \nz.mem [3692] = \nz.mem_3692_sv2v_reg ;
  assign \nz.mem [3691] = \nz.mem_3691_sv2v_reg ;
  assign \nz.mem [3690] = \nz.mem_3690_sv2v_reg ;
  assign \nz.mem [3689] = \nz.mem_3689_sv2v_reg ;
  assign \nz.mem [3688] = \nz.mem_3688_sv2v_reg ;
  assign \nz.mem [3687] = \nz.mem_3687_sv2v_reg ;
  assign \nz.mem [3686] = \nz.mem_3686_sv2v_reg ;
  assign \nz.mem [3685] = \nz.mem_3685_sv2v_reg ;
  assign \nz.mem [3684] = \nz.mem_3684_sv2v_reg ;
  assign \nz.mem [3683] = \nz.mem_3683_sv2v_reg ;
  assign \nz.mem [3682] = \nz.mem_3682_sv2v_reg ;
  assign \nz.mem [3681] = \nz.mem_3681_sv2v_reg ;
  assign \nz.mem [3680] = \nz.mem_3680_sv2v_reg ;
  assign \nz.mem [3679] = \nz.mem_3679_sv2v_reg ;
  assign \nz.mem [3678] = \nz.mem_3678_sv2v_reg ;
  assign \nz.mem [3677] = \nz.mem_3677_sv2v_reg ;
  assign \nz.mem [3676] = \nz.mem_3676_sv2v_reg ;
  assign \nz.mem [3675] = \nz.mem_3675_sv2v_reg ;
  assign \nz.mem [3674] = \nz.mem_3674_sv2v_reg ;
  assign \nz.mem [3673] = \nz.mem_3673_sv2v_reg ;
  assign \nz.mem [3672] = \nz.mem_3672_sv2v_reg ;
  assign \nz.mem [3671] = \nz.mem_3671_sv2v_reg ;
  assign \nz.mem [3670] = \nz.mem_3670_sv2v_reg ;
  assign \nz.mem [3669] = \nz.mem_3669_sv2v_reg ;
  assign \nz.mem [3668] = \nz.mem_3668_sv2v_reg ;
  assign \nz.mem [3667] = \nz.mem_3667_sv2v_reg ;
  assign \nz.mem [3666] = \nz.mem_3666_sv2v_reg ;
  assign \nz.mem [3665] = \nz.mem_3665_sv2v_reg ;
  assign \nz.mem [3664] = \nz.mem_3664_sv2v_reg ;
  assign \nz.mem [3663] = \nz.mem_3663_sv2v_reg ;
  assign \nz.mem [3662] = \nz.mem_3662_sv2v_reg ;
  assign \nz.mem [3661] = \nz.mem_3661_sv2v_reg ;
  assign \nz.mem [3660] = \nz.mem_3660_sv2v_reg ;
  assign \nz.mem [3659] = \nz.mem_3659_sv2v_reg ;
  assign \nz.mem [3658] = \nz.mem_3658_sv2v_reg ;
  assign \nz.mem [3657] = \nz.mem_3657_sv2v_reg ;
  assign \nz.mem [3656] = \nz.mem_3656_sv2v_reg ;
  assign \nz.mem [3655] = \nz.mem_3655_sv2v_reg ;
  assign \nz.mem [3654] = \nz.mem_3654_sv2v_reg ;
  assign \nz.mem [3653] = \nz.mem_3653_sv2v_reg ;
  assign \nz.mem [3652] = \nz.mem_3652_sv2v_reg ;
  assign \nz.mem [3651] = \nz.mem_3651_sv2v_reg ;
  assign \nz.mem [3650] = \nz.mem_3650_sv2v_reg ;
  assign \nz.mem [3649] = \nz.mem_3649_sv2v_reg ;
  assign \nz.mem [3648] = \nz.mem_3648_sv2v_reg ;
  assign \nz.mem [3647] = \nz.mem_3647_sv2v_reg ;
  assign \nz.mem [3646] = \nz.mem_3646_sv2v_reg ;
  assign \nz.mem [3645] = \nz.mem_3645_sv2v_reg ;
  assign \nz.mem [3644] = \nz.mem_3644_sv2v_reg ;
  assign \nz.mem [3643] = \nz.mem_3643_sv2v_reg ;
  assign \nz.mem [3642] = \nz.mem_3642_sv2v_reg ;
  assign \nz.mem [3641] = \nz.mem_3641_sv2v_reg ;
  assign \nz.mem [3640] = \nz.mem_3640_sv2v_reg ;
  assign \nz.mem [3639] = \nz.mem_3639_sv2v_reg ;
  assign \nz.mem [3638] = \nz.mem_3638_sv2v_reg ;
  assign \nz.mem [3637] = \nz.mem_3637_sv2v_reg ;
  assign \nz.mem [3636] = \nz.mem_3636_sv2v_reg ;
  assign \nz.mem [3635] = \nz.mem_3635_sv2v_reg ;
  assign \nz.mem [3634] = \nz.mem_3634_sv2v_reg ;
  assign \nz.mem [3633] = \nz.mem_3633_sv2v_reg ;
  assign \nz.mem [3632] = \nz.mem_3632_sv2v_reg ;
  assign \nz.mem [3631] = \nz.mem_3631_sv2v_reg ;
  assign \nz.mem [3630] = \nz.mem_3630_sv2v_reg ;
  assign \nz.mem [3629] = \nz.mem_3629_sv2v_reg ;
  assign \nz.mem [3628] = \nz.mem_3628_sv2v_reg ;
  assign \nz.mem [3627] = \nz.mem_3627_sv2v_reg ;
  assign \nz.mem [3626] = \nz.mem_3626_sv2v_reg ;
  assign \nz.mem [3625] = \nz.mem_3625_sv2v_reg ;
  assign \nz.mem [3624] = \nz.mem_3624_sv2v_reg ;
  assign \nz.mem [3623] = \nz.mem_3623_sv2v_reg ;
  assign \nz.mem [3622] = \nz.mem_3622_sv2v_reg ;
  assign \nz.mem [3621] = \nz.mem_3621_sv2v_reg ;
  assign \nz.mem [3620] = \nz.mem_3620_sv2v_reg ;
  assign \nz.mem [3619] = \nz.mem_3619_sv2v_reg ;
  assign \nz.mem [3618] = \nz.mem_3618_sv2v_reg ;
  assign \nz.mem [3617] = \nz.mem_3617_sv2v_reg ;
  assign \nz.mem [3616] = \nz.mem_3616_sv2v_reg ;
  assign \nz.mem [3615] = \nz.mem_3615_sv2v_reg ;
  assign \nz.mem [3614] = \nz.mem_3614_sv2v_reg ;
  assign \nz.mem [3613] = \nz.mem_3613_sv2v_reg ;
  assign \nz.mem [3612] = \nz.mem_3612_sv2v_reg ;
  assign \nz.mem [3611] = \nz.mem_3611_sv2v_reg ;
  assign \nz.mem [3610] = \nz.mem_3610_sv2v_reg ;
  assign \nz.mem [3609] = \nz.mem_3609_sv2v_reg ;
  assign \nz.mem [3608] = \nz.mem_3608_sv2v_reg ;
  assign \nz.mem [3607] = \nz.mem_3607_sv2v_reg ;
  assign \nz.mem [3606] = \nz.mem_3606_sv2v_reg ;
  assign \nz.mem [3605] = \nz.mem_3605_sv2v_reg ;
  assign \nz.mem [3604] = \nz.mem_3604_sv2v_reg ;
  assign \nz.mem [3603] = \nz.mem_3603_sv2v_reg ;
  assign \nz.mem [3602] = \nz.mem_3602_sv2v_reg ;
  assign \nz.mem [3601] = \nz.mem_3601_sv2v_reg ;
  assign \nz.mem [3600] = \nz.mem_3600_sv2v_reg ;
  assign \nz.mem [3599] = \nz.mem_3599_sv2v_reg ;
  assign \nz.mem [3598] = \nz.mem_3598_sv2v_reg ;
  assign \nz.mem [3597] = \nz.mem_3597_sv2v_reg ;
  assign \nz.mem [3596] = \nz.mem_3596_sv2v_reg ;
  assign \nz.mem [3595] = \nz.mem_3595_sv2v_reg ;
  assign \nz.mem [3594] = \nz.mem_3594_sv2v_reg ;
  assign \nz.mem [3593] = \nz.mem_3593_sv2v_reg ;
  assign \nz.mem [3592] = \nz.mem_3592_sv2v_reg ;
  assign \nz.mem [3591] = \nz.mem_3591_sv2v_reg ;
  assign \nz.mem [3590] = \nz.mem_3590_sv2v_reg ;
  assign \nz.mem [3589] = \nz.mem_3589_sv2v_reg ;
  assign \nz.mem [3588] = \nz.mem_3588_sv2v_reg ;
  assign \nz.mem [3587] = \nz.mem_3587_sv2v_reg ;
  assign \nz.mem [3586] = \nz.mem_3586_sv2v_reg ;
  assign \nz.mem [3585] = \nz.mem_3585_sv2v_reg ;
  assign \nz.mem [3584] = \nz.mem_3584_sv2v_reg ;
  assign \nz.mem [3583] = \nz.mem_3583_sv2v_reg ;
  assign \nz.mem [3582] = \nz.mem_3582_sv2v_reg ;
  assign \nz.mem [3581] = \nz.mem_3581_sv2v_reg ;
  assign \nz.mem [3580] = \nz.mem_3580_sv2v_reg ;
  assign \nz.mem [3579] = \nz.mem_3579_sv2v_reg ;
  assign \nz.mem [3578] = \nz.mem_3578_sv2v_reg ;
  assign \nz.mem [3577] = \nz.mem_3577_sv2v_reg ;
  assign \nz.mem [3576] = \nz.mem_3576_sv2v_reg ;
  assign \nz.mem [3575] = \nz.mem_3575_sv2v_reg ;
  assign \nz.mem [3574] = \nz.mem_3574_sv2v_reg ;
  assign \nz.mem [3573] = \nz.mem_3573_sv2v_reg ;
  assign \nz.mem [3572] = \nz.mem_3572_sv2v_reg ;
  assign \nz.mem [3571] = \nz.mem_3571_sv2v_reg ;
  assign \nz.mem [3570] = \nz.mem_3570_sv2v_reg ;
  assign \nz.mem [3569] = \nz.mem_3569_sv2v_reg ;
  assign \nz.mem [3568] = \nz.mem_3568_sv2v_reg ;
  assign \nz.mem [3567] = \nz.mem_3567_sv2v_reg ;
  assign \nz.mem [3566] = \nz.mem_3566_sv2v_reg ;
  assign \nz.mem [3565] = \nz.mem_3565_sv2v_reg ;
  assign \nz.mem [3564] = \nz.mem_3564_sv2v_reg ;
  assign \nz.mem [3563] = \nz.mem_3563_sv2v_reg ;
  assign \nz.mem [3562] = \nz.mem_3562_sv2v_reg ;
  assign \nz.mem [3561] = \nz.mem_3561_sv2v_reg ;
  assign \nz.mem [3560] = \nz.mem_3560_sv2v_reg ;
  assign \nz.mem [3559] = \nz.mem_3559_sv2v_reg ;
  assign \nz.mem [3558] = \nz.mem_3558_sv2v_reg ;
  assign \nz.mem [3557] = \nz.mem_3557_sv2v_reg ;
  assign \nz.mem [3556] = \nz.mem_3556_sv2v_reg ;
  assign \nz.mem [3555] = \nz.mem_3555_sv2v_reg ;
  assign \nz.mem [3554] = \nz.mem_3554_sv2v_reg ;
  assign \nz.mem [3553] = \nz.mem_3553_sv2v_reg ;
  assign \nz.mem [3552] = \nz.mem_3552_sv2v_reg ;
  assign \nz.mem [3551] = \nz.mem_3551_sv2v_reg ;
  assign \nz.mem [3550] = \nz.mem_3550_sv2v_reg ;
  assign \nz.mem [3549] = \nz.mem_3549_sv2v_reg ;
  assign \nz.mem [3548] = \nz.mem_3548_sv2v_reg ;
  assign \nz.mem [3547] = \nz.mem_3547_sv2v_reg ;
  assign \nz.mem [3546] = \nz.mem_3546_sv2v_reg ;
  assign \nz.mem [3545] = \nz.mem_3545_sv2v_reg ;
  assign \nz.mem [3544] = \nz.mem_3544_sv2v_reg ;
  assign \nz.mem [3543] = \nz.mem_3543_sv2v_reg ;
  assign \nz.mem [3542] = \nz.mem_3542_sv2v_reg ;
  assign \nz.mem [3541] = \nz.mem_3541_sv2v_reg ;
  assign \nz.mem [3540] = \nz.mem_3540_sv2v_reg ;
  assign \nz.mem [3539] = \nz.mem_3539_sv2v_reg ;
  assign \nz.mem [3538] = \nz.mem_3538_sv2v_reg ;
  assign \nz.mem [3537] = \nz.mem_3537_sv2v_reg ;
  assign \nz.mem [3536] = \nz.mem_3536_sv2v_reg ;
  assign \nz.mem [3535] = \nz.mem_3535_sv2v_reg ;
  assign \nz.mem [3534] = \nz.mem_3534_sv2v_reg ;
  assign \nz.mem [3533] = \nz.mem_3533_sv2v_reg ;
  assign \nz.mem [3532] = \nz.mem_3532_sv2v_reg ;
  assign \nz.mem [3531] = \nz.mem_3531_sv2v_reg ;
  assign \nz.mem [3530] = \nz.mem_3530_sv2v_reg ;
  assign \nz.mem [3529] = \nz.mem_3529_sv2v_reg ;
  assign \nz.mem [3528] = \nz.mem_3528_sv2v_reg ;
  assign \nz.mem [3527] = \nz.mem_3527_sv2v_reg ;
  assign \nz.mem [3526] = \nz.mem_3526_sv2v_reg ;
  assign \nz.mem [3525] = \nz.mem_3525_sv2v_reg ;
  assign \nz.mem [3524] = \nz.mem_3524_sv2v_reg ;
  assign \nz.mem [3523] = \nz.mem_3523_sv2v_reg ;
  assign \nz.mem [3522] = \nz.mem_3522_sv2v_reg ;
  assign \nz.mem [3521] = \nz.mem_3521_sv2v_reg ;
  assign \nz.mem [3520] = \nz.mem_3520_sv2v_reg ;
  assign \nz.mem [3519] = \nz.mem_3519_sv2v_reg ;
  assign \nz.mem [3518] = \nz.mem_3518_sv2v_reg ;
  assign \nz.mem [3517] = \nz.mem_3517_sv2v_reg ;
  assign \nz.mem [3516] = \nz.mem_3516_sv2v_reg ;
  assign \nz.mem [3515] = \nz.mem_3515_sv2v_reg ;
  assign \nz.mem [3514] = \nz.mem_3514_sv2v_reg ;
  assign \nz.mem [3513] = \nz.mem_3513_sv2v_reg ;
  assign \nz.mem [3512] = \nz.mem_3512_sv2v_reg ;
  assign \nz.mem [3511] = \nz.mem_3511_sv2v_reg ;
  assign \nz.mem [3510] = \nz.mem_3510_sv2v_reg ;
  assign \nz.mem [3509] = \nz.mem_3509_sv2v_reg ;
  assign \nz.mem [3508] = \nz.mem_3508_sv2v_reg ;
  assign \nz.mem [3507] = \nz.mem_3507_sv2v_reg ;
  assign \nz.mem [3506] = \nz.mem_3506_sv2v_reg ;
  assign \nz.mem [3505] = \nz.mem_3505_sv2v_reg ;
  assign \nz.mem [3504] = \nz.mem_3504_sv2v_reg ;
  assign \nz.mem [3503] = \nz.mem_3503_sv2v_reg ;
  assign \nz.mem [3502] = \nz.mem_3502_sv2v_reg ;
  assign \nz.mem [3501] = \nz.mem_3501_sv2v_reg ;
  assign \nz.mem [3500] = \nz.mem_3500_sv2v_reg ;
  assign \nz.mem [3499] = \nz.mem_3499_sv2v_reg ;
  assign \nz.mem [3498] = \nz.mem_3498_sv2v_reg ;
  assign \nz.mem [3497] = \nz.mem_3497_sv2v_reg ;
  assign \nz.mem [3496] = \nz.mem_3496_sv2v_reg ;
  assign \nz.mem [3495] = \nz.mem_3495_sv2v_reg ;
  assign \nz.mem [3494] = \nz.mem_3494_sv2v_reg ;
  assign \nz.mem [3493] = \nz.mem_3493_sv2v_reg ;
  assign \nz.mem [3492] = \nz.mem_3492_sv2v_reg ;
  assign \nz.mem [3491] = \nz.mem_3491_sv2v_reg ;
  assign \nz.mem [3490] = \nz.mem_3490_sv2v_reg ;
  assign \nz.mem [3489] = \nz.mem_3489_sv2v_reg ;
  assign \nz.mem [3488] = \nz.mem_3488_sv2v_reg ;
  assign \nz.mem [3487] = \nz.mem_3487_sv2v_reg ;
  assign \nz.mem [3486] = \nz.mem_3486_sv2v_reg ;
  assign \nz.mem [3485] = \nz.mem_3485_sv2v_reg ;
  assign \nz.mem [3484] = \nz.mem_3484_sv2v_reg ;
  assign \nz.mem [3483] = \nz.mem_3483_sv2v_reg ;
  assign \nz.mem [3482] = \nz.mem_3482_sv2v_reg ;
  assign \nz.mem [3481] = \nz.mem_3481_sv2v_reg ;
  assign \nz.mem [3480] = \nz.mem_3480_sv2v_reg ;
  assign \nz.mem [3479] = \nz.mem_3479_sv2v_reg ;
  assign \nz.mem [3478] = \nz.mem_3478_sv2v_reg ;
  assign \nz.mem [3477] = \nz.mem_3477_sv2v_reg ;
  assign \nz.mem [3476] = \nz.mem_3476_sv2v_reg ;
  assign \nz.mem [3475] = \nz.mem_3475_sv2v_reg ;
  assign \nz.mem [3474] = \nz.mem_3474_sv2v_reg ;
  assign \nz.mem [3473] = \nz.mem_3473_sv2v_reg ;
  assign \nz.mem [3472] = \nz.mem_3472_sv2v_reg ;
  assign \nz.mem [3471] = \nz.mem_3471_sv2v_reg ;
  assign \nz.mem [3470] = \nz.mem_3470_sv2v_reg ;
  assign \nz.mem [3469] = \nz.mem_3469_sv2v_reg ;
  assign \nz.mem [3468] = \nz.mem_3468_sv2v_reg ;
  assign \nz.mem [3467] = \nz.mem_3467_sv2v_reg ;
  assign \nz.mem [3466] = \nz.mem_3466_sv2v_reg ;
  assign \nz.mem [3465] = \nz.mem_3465_sv2v_reg ;
  assign \nz.mem [3464] = \nz.mem_3464_sv2v_reg ;
  assign \nz.mem [3463] = \nz.mem_3463_sv2v_reg ;
  assign \nz.mem [3462] = \nz.mem_3462_sv2v_reg ;
  assign \nz.mem [3461] = \nz.mem_3461_sv2v_reg ;
  assign \nz.mem [3460] = \nz.mem_3460_sv2v_reg ;
  assign \nz.mem [3459] = \nz.mem_3459_sv2v_reg ;
  assign \nz.mem [3458] = \nz.mem_3458_sv2v_reg ;
  assign \nz.mem [3457] = \nz.mem_3457_sv2v_reg ;
  assign \nz.mem [3456] = \nz.mem_3456_sv2v_reg ;
  assign \nz.mem [3455] = \nz.mem_3455_sv2v_reg ;
  assign \nz.mem [3454] = \nz.mem_3454_sv2v_reg ;
  assign \nz.mem [3453] = \nz.mem_3453_sv2v_reg ;
  assign \nz.mem [3452] = \nz.mem_3452_sv2v_reg ;
  assign \nz.mem [3451] = \nz.mem_3451_sv2v_reg ;
  assign \nz.mem [3450] = \nz.mem_3450_sv2v_reg ;
  assign \nz.mem [3449] = \nz.mem_3449_sv2v_reg ;
  assign \nz.mem [3448] = \nz.mem_3448_sv2v_reg ;
  assign \nz.mem [3447] = \nz.mem_3447_sv2v_reg ;
  assign \nz.mem [3446] = \nz.mem_3446_sv2v_reg ;
  assign \nz.mem [3445] = \nz.mem_3445_sv2v_reg ;
  assign \nz.mem [3444] = \nz.mem_3444_sv2v_reg ;
  assign \nz.mem [3443] = \nz.mem_3443_sv2v_reg ;
  assign \nz.mem [3442] = \nz.mem_3442_sv2v_reg ;
  assign \nz.mem [3441] = \nz.mem_3441_sv2v_reg ;
  assign \nz.mem [3440] = \nz.mem_3440_sv2v_reg ;
  assign \nz.mem [3439] = \nz.mem_3439_sv2v_reg ;
  assign \nz.mem [3438] = \nz.mem_3438_sv2v_reg ;
  assign \nz.mem [3437] = \nz.mem_3437_sv2v_reg ;
  assign \nz.mem [3436] = \nz.mem_3436_sv2v_reg ;
  assign \nz.mem [3435] = \nz.mem_3435_sv2v_reg ;
  assign \nz.mem [3434] = \nz.mem_3434_sv2v_reg ;
  assign \nz.mem [3433] = \nz.mem_3433_sv2v_reg ;
  assign \nz.mem [3432] = \nz.mem_3432_sv2v_reg ;
  assign \nz.mem [3431] = \nz.mem_3431_sv2v_reg ;
  assign \nz.mem [3430] = \nz.mem_3430_sv2v_reg ;
  assign \nz.mem [3429] = \nz.mem_3429_sv2v_reg ;
  assign \nz.mem [3428] = \nz.mem_3428_sv2v_reg ;
  assign \nz.mem [3427] = \nz.mem_3427_sv2v_reg ;
  assign \nz.mem [3426] = \nz.mem_3426_sv2v_reg ;
  assign \nz.mem [3425] = \nz.mem_3425_sv2v_reg ;
  assign \nz.mem [3424] = \nz.mem_3424_sv2v_reg ;
  assign \nz.mem [3423] = \nz.mem_3423_sv2v_reg ;
  assign \nz.mem [3422] = \nz.mem_3422_sv2v_reg ;
  assign \nz.mem [3421] = \nz.mem_3421_sv2v_reg ;
  assign \nz.mem [3420] = \nz.mem_3420_sv2v_reg ;
  assign \nz.mem [3419] = \nz.mem_3419_sv2v_reg ;
  assign \nz.mem [3418] = \nz.mem_3418_sv2v_reg ;
  assign \nz.mem [3417] = \nz.mem_3417_sv2v_reg ;
  assign \nz.mem [3416] = \nz.mem_3416_sv2v_reg ;
  assign \nz.mem [3415] = \nz.mem_3415_sv2v_reg ;
  assign \nz.mem [3414] = \nz.mem_3414_sv2v_reg ;
  assign \nz.mem [3413] = \nz.mem_3413_sv2v_reg ;
  assign \nz.mem [3412] = \nz.mem_3412_sv2v_reg ;
  assign \nz.mem [3411] = \nz.mem_3411_sv2v_reg ;
  assign \nz.mem [3410] = \nz.mem_3410_sv2v_reg ;
  assign \nz.mem [3409] = \nz.mem_3409_sv2v_reg ;
  assign \nz.mem [3408] = \nz.mem_3408_sv2v_reg ;
  assign \nz.mem [3407] = \nz.mem_3407_sv2v_reg ;
  assign \nz.mem [3406] = \nz.mem_3406_sv2v_reg ;
  assign \nz.mem [3405] = \nz.mem_3405_sv2v_reg ;
  assign \nz.mem [3404] = \nz.mem_3404_sv2v_reg ;
  assign \nz.mem [3403] = \nz.mem_3403_sv2v_reg ;
  assign \nz.mem [3402] = \nz.mem_3402_sv2v_reg ;
  assign \nz.mem [3401] = \nz.mem_3401_sv2v_reg ;
  assign \nz.mem [3400] = \nz.mem_3400_sv2v_reg ;
  assign \nz.mem [3399] = \nz.mem_3399_sv2v_reg ;
  assign \nz.mem [3398] = \nz.mem_3398_sv2v_reg ;
  assign \nz.mem [3397] = \nz.mem_3397_sv2v_reg ;
  assign \nz.mem [3396] = \nz.mem_3396_sv2v_reg ;
  assign \nz.mem [3395] = \nz.mem_3395_sv2v_reg ;
  assign \nz.mem [3394] = \nz.mem_3394_sv2v_reg ;
  assign \nz.mem [3393] = \nz.mem_3393_sv2v_reg ;
  assign \nz.mem [3392] = \nz.mem_3392_sv2v_reg ;
  assign \nz.mem [3391] = \nz.mem_3391_sv2v_reg ;
  assign \nz.mem [3390] = \nz.mem_3390_sv2v_reg ;
  assign \nz.mem [3389] = \nz.mem_3389_sv2v_reg ;
  assign \nz.mem [3388] = \nz.mem_3388_sv2v_reg ;
  assign \nz.mem [3387] = \nz.mem_3387_sv2v_reg ;
  assign \nz.mem [3386] = \nz.mem_3386_sv2v_reg ;
  assign \nz.mem [3385] = \nz.mem_3385_sv2v_reg ;
  assign \nz.mem [3384] = \nz.mem_3384_sv2v_reg ;
  assign \nz.mem [3383] = \nz.mem_3383_sv2v_reg ;
  assign \nz.mem [3382] = \nz.mem_3382_sv2v_reg ;
  assign \nz.mem [3381] = \nz.mem_3381_sv2v_reg ;
  assign \nz.mem [3380] = \nz.mem_3380_sv2v_reg ;
  assign \nz.mem [3379] = \nz.mem_3379_sv2v_reg ;
  assign \nz.mem [3378] = \nz.mem_3378_sv2v_reg ;
  assign \nz.mem [3377] = \nz.mem_3377_sv2v_reg ;
  assign \nz.mem [3376] = \nz.mem_3376_sv2v_reg ;
  assign \nz.mem [3375] = \nz.mem_3375_sv2v_reg ;
  assign \nz.mem [3374] = \nz.mem_3374_sv2v_reg ;
  assign \nz.mem [3373] = \nz.mem_3373_sv2v_reg ;
  assign \nz.mem [3372] = \nz.mem_3372_sv2v_reg ;
  assign \nz.mem [3371] = \nz.mem_3371_sv2v_reg ;
  assign \nz.mem [3370] = \nz.mem_3370_sv2v_reg ;
  assign \nz.mem [3369] = \nz.mem_3369_sv2v_reg ;
  assign \nz.mem [3368] = \nz.mem_3368_sv2v_reg ;
  assign \nz.mem [3367] = \nz.mem_3367_sv2v_reg ;
  assign \nz.mem [3366] = \nz.mem_3366_sv2v_reg ;
  assign \nz.mem [3365] = \nz.mem_3365_sv2v_reg ;
  assign \nz.mem [3364] = \nz.mem_3364_sv2v_reg ;
  assign \nz.mem [3363] = \nz.mem_3363_sv2v_reg ;
  assign \nz.mem [3362] = \nz.mem_3362_sv2v_reg ;
  assign \nz.mem [3361] = \nz.mem_3361_sv2v_reg ;
  assign \nz.mem [3360] = \nz.mem_3360_sv2v_reg ;
  assign \nz.mem [3359] = \nz.mem_3359_sv2v_reg ;
  assign \nz.mem [3358] = \nz.mem_3358_sv2v_reg ;
  assign \nz.mem [3357] = \nz.mem_3357_sv2v_reg ;
  assign \nz.mem [3356] = \nz.mem_3356_sv2v_reg ;
  assign \nz.mem [3355] = \nz.mem_3355_sv2v_reg ;
  assign \nz.mem [3354] = \nz.mem_3354_sv2v_reg ;
  assign \nz.mem [3353] = \nz.mem_3353_sv2v_reg ;
  assign \nz.mem [3352] = \nz.mem_3352_sv2v_reg ;
  assign \nz.mem [3351] = \nz.mem_3351_sv2v_reg ;
  assign \nz.mem [3350] = \nz.mem_3350_sv2v_reg ;
  assign \nz.mem [3349] = \nz.mem_3349_sv2v_reg ;
  assign \nz.mem [3348] = \nz.mem_3348_sv2v_reg ;
  assign \nz.mem [3347] = \nz.mem_3347_sv2v_reg ;
  assign \nz.mem [3346] = \nz.mem_3346_sv2v_reg ;
  assign \nz.mem [3345] = \nz.mem_3345_sv2v_reg ;
  assign \nz.mem [3344] = \nz.mem_3344_sv2v_reg ;
  assign \nz.mem [3343] = \nz.mem_3343_sv2v_reg ;
  assign \nz.mem [3342] = \nz.mem_3342_sv2v_reg ;
  assign \nz.mem [3341] = \nz.mem_3341_sv2v_reg ;
  assign \nz.mem [3340] = \nz.mem_3340_sv2v_reg ;
  assign \nz.mem [3339] = \nz.mem_3339_sv2v_reg ;
  assign \nz.mem [3338] = \nz.mem_3338_sv2v_reg ;
  assign \nz.mem [3337] = \nz.mem_3337_sv2v_reg ;
  assign \nz.mem [3336] = \nz.mem_3336_sv2v_reg ;
  assign \nz.mem [3335] = \nz.mem_3335_sv2v_reg ;
  assign \nz.mem [3334] = \nz.mem_3334_sv2v_reg ;
  assign \nz.mem [3333] = \nz.mem_3333_sv2v_reg ;
  assign \nz.mem [3332] = \nz.mem_3332_sv2v_reg ;
  assign \nz.mem [3331] = \nz.mem_3331_sv2v_reg ;
  assign \nz.mem [3330] = \nz.mem_3330_sv2v_reg ;
  assign \nz.mem [3329] = \nz.mem_3329_sv2v_reg ;
  assign \nz.mem [3328] = \nz.mem_3328_sv2v_reg ;
  assign \nz.mem [3327] = \nz.mem_3327_sv2v_reg ;
  assign \nz.mem [3326] = \nz.mem_3326_sv2v_reg ;
  assign \nz.mem [3325] = \nz.mem_3325_sv2v_reg ;
  assign \nz.mem [3324] = \nz.mem_3324_sv2v_reg ;
  assign \nz.mem [3323] = \nz.mem_3323_sv2v_reg ;
  assign \nz.mem [3322] = \nz.mem_3322_sv2v_reg ;
  assign \nz.mem [3321] = \nz.mem_3321_sv2v_reg ;
  assign \nz.mem [3320] = \nz.mem_3320_sv2v_reg ;
  assign \nz.mem [3319] = \nz.mem_3319_sv2v_reg ;
  assign \nz.mem [3318] = \nz.mem_3318_sv2v_reg ;
  assign \nz.mem [3317] = \nz.mem_3317_sv2v_reg ;
  assign \nz.mem [3316] = \nz.mem_3316_sv2v_reg ;
  assign \nz.mem [3315] = \nz.mem_3315_sv2v_reg ;
  assign \nz.mem [3314] = \nz.mem_3314_sv2v_reg ;
  assign \nz.mem [3313] = \nz.mem_3313_sv2v_reg ;
  assign \nz.mem [3312] = \nz.mem_3312_sv2v_reg ;
  assign \nz.mem [3311] = \nz.mem_3311_sv2v_reg ;
  assign \nz.mem [3310] = \nz.mem_3310_sv2v_reg ;
  assign \nz.mem [3309] = \nz.mem_3309_sv2v_reg ;
  assign \nz.mem [3308] = \nz.mem_3308_sv2v_reg ;
  assign \nz.mem [3307] = \nz.mem_3307_sv2v_reg ;
  assign \nz.mem [3306] = \nz.mem_3306_sv2v_reg ;
  assign \nz.mem [3305] = \nz.mem_3305_sv2v_reg ;
  assign \nz.mem [3304] = \nz.mem_3304_sv2v_reg ;
  assign \nz.mem [3303] = \nz.mem_3303_sv2v_reg ;
  assign \nz.mem [3302] = \nz.mem_3302_sv2v_reg ;
  assign \nz.mem [3301] = \nz.mem_3301_sv2v_reg ;
  assign \nz.mem [3300] = \nz.mem_3300_sv2v_reg ;
  assign \nz.mem [3299] = \nz.mem_3299_sv2v_reg ;
  assign \nz.mem [3298] = \nz.mem_3298_sv2v_reg ;
  assign \nz.mem [3297] = \nz.mem_3297_sv2v_reg ;
  assign \nz.mem [3296] = \nz.mem_3296_sv2v_reg ;
  assign \nz.mem [3295] = \nz.mem_3295_sv2v_reg ;
  assign \nz.mem [3294] = \nz.mem_3294_sv2v_reg ;
  assign \nz.mem [3293] = \nz.mem_3293_sv2v_reg ;
  assign \nz.mem [3292] = \nz.mem_3292_sv2v_reg ;
  assign \nz.mem [3291] = \nz.mem_3291_sv2v_reg ;
  assign \nz.mem [3290] = \nz.mem_3290_sv2v_reg ;
  assign \nz.mem [3289] = \nz.mem_3289_sv2v_reg ;
  assign \nz.mem [3288] = \nz.mem_3288_sv2v_reg ;
  assign \nz.mem [3287] = \nz.mem_3287_sv2v_reg ;
  assign \nz.mem [3286] = \nz.mem_3286_sv2v_reg ;
  assign \nz.mem [3285] = \nz.mem_3285_sv2v_reg ;
  assign \nz.mem [3284] = \nz.mem_3284_sv2v_reg ;
  assign \nz.mem [3283] = \nz.mem_3283_sv2v_reg ;
  assign \nz.mem [3282] = \nz.mem_3282_sv2v_reg ;
  assign \nz.mem [3281] = \nz.mem_3281_sv2v_reg ;
  assign \nz.mem [3280] = \nz.mem_3280_sv2v_reg ;
  assign \nz.mem [3279] = \nz.mem_3279_sv2v_reg ;
  assign \nz.mem [3278] = \nz.mem_3278_sv2v_reg ;
  assign \nz.mem [3277] = \nz.mem_3277_sv2v_reg ;
  assign \nz.mem [3276] = \nz.mem_3276_sv2v_reg ;
  assign \nz.mem [3275] = \nz.mem_3275_sv2v_reg ;
  assign \nz.mem [3274] = \nz.mem_3274_sv2v_reg ;
  assign \nz.mem [3273] = \nz.mem_3273_sv2v_reg ;
  assign \nz.mem [3272] = \nz.mem_3272_sv2v_reg ;
  assign \nz.mem [3271] = \nz.mem_3271_sv2v_reg ;
  assign \nz.mem [3270] = \nz.mem_3270_sv2v_reg ;
  assign \nz.mem [3269] = \nz.mem_3269_sv2v_reg ;
  assign \nz.mem [3268] = \nz.mem_3268_sv2v_reg ;
  assign \nz.mem [3267] = \nz.mem_3267_sv2v_reg ;
  assign \nz.mem [3266] = \nz.mem_3266_sv2v_reg ;
  assign \nz.mem [3265] = \nz.mem_3265_sv2v_reg ;
  assign \nz.mem [3264] = \nz.mem_3264_sv2v_reg ;
  assign \nz.mem [3263] = \nz.mem_3263_sv2v_reg ;
  assign \nz.mem [3262] = \nz.mem_3262_sv2v_reg ;
  assign \nz.mem [3261] = \nz.mem_3261_sv2v_reg ;
  assign \nz.mem [3260] = \nz.mem_3260_sv2v_reg ;
  assign \nz.mem [3259] = \nz.mem_3259_sv2v_reg ;
  assign \nz.mem [3258] = \nz.mem_3258_sv2v_reg ;
  assign \nz.mem [3257] = \nz.mem_3257_sv2v_reg ;
  assign \nz.mem [3256] = \nz.mem_3256_sv2v_reg ;
  assign \nz.mem [3255] = \nz.mem_3255_sv2v_reg ;
  assign \nz.mem [3254] = \nz.mem_3254_sv2v_reg ;
  assign \nz.mem [3253] = \nz.mem_3253_sv2v_reg ;
  assign \nz.mem [3252] = \nz.mem_3252_sv2v_reg ;
  assign \nz.mem [3251] = \nz.mem_3251_sv2v_reg ;
  assign \nz.mem [3250] = \nz.mem_3250_sv2v_reg ;
  assign \nz.mem [3249] = \nz.mem_3249_sv2v_reg ;
  assign \nz.mem [3248] = \nz.mem_3248_sv2v_reg ;
  assign \nz.mem [3247] = \nz.mem_3247_sv2v_reg ;
  assign \nz.mem [3246] = \nz.mem_3246_sv2v_reg ;
  assign \nz.mem [3245] = \nz.mem_3245_sv2v_reg ;
  assign \nz.mem [3244] = \nz.mem_3244_sv2v_reg ;
  assign \nz.mem [3243] = \nz.mem_3243_sv2v_reg ;
  assign \nz.mem [3242] = \nz.mem_3242_sv2v_reg ;
  assign \nz.mem [3241] = \nz.mem_3241_sv2v_reg ;
  assign \nz.mem [3240] = \nz.mem_3240_sv2v_reg ;
  assign \nz.mem [3239] = \nz.mem_3239_sv2v_reg ;
  assign \nz.mem [3238] = \nz.mem_3238_sv2v_reg ;
  assign \nz.mem [3237] = \nz.mem_3237_sv2v_reg ;
  assign \nz.mem [3236] = \nz.mem_3236_sv2v_reg ;
  assign \nz.mem [3235] = \nz.mem_3235_sv2v_reg ;
  assign \nz.mem [3234] = \nz.mem_3234_sv2v_reg ;
  assign \nz.mem [3233] = \nz.mem_3233_sv2v_reg ;
  assign \nz.mem [3232] = \nz.mem_3232_sv2v_reg ;
  assign \nz.mem [3231] = \nz.mem_3231_sv2v_reg ;
  assign \nz.mem [3230] = \nz.mem_3230_sv2v_reg ;
  assign \nz.mem [3229] = \nz.mem_3229_sv2v_reg ;
  assign \nz.mem [3228] = \nz.mem_3228_sv2v_reg ;
  assign \nz.mem [3227] = \nz.mem_3227_sv2v_reg ;
  assign \nz.mem [3226] = \nz.mem_3226_sv2v_reg ;
  assign \nz.mem [3225] = \nz.mem_3225_sv2v_reg ;
  assign \nz.mem [3224] = \nz.mem_3224_sv2v_reg ;
  assign \nz.mem [3223] = \nz.mem_3223_sv2v_reg ;
  assign \nz.mem [3222] = \nz.mem_3222_sv2v_reg ;
  assign \nz.mem [3221] = \nz.mem_3221_sv2v_reg ;
  assign \nz.mem [3220] = \nz.mem_3220_sv2v_reg ;
  assign \nz.mem [3219] = \nz.mem_3219_sv2v_reg ;
  assign \nz.mem [3218] = \nz.mem_3218_sv2v_reg ;
  assign \nz.mem [3217] = \nz.mem_3217_sv2v_reg ;
  assign \nz.mem [3216] = \nz.mem_3216_sv2v_reg ;
  assign \nz.mem [3215] = \nz.mem_3215_sv2v_reg ;
  assign \nz.mem [3214] = \nz.mem_3214_sv2v_reg ;
  assign \nz.mem [3213] = \nz.mem_3213_sv2v_reg ;
  assign \nz.mem [3212] = \nz.mem_3212_sv2v_reg ;
  assign \nz.mem [3211] = \nz.mem_3211_sv2v_reg ;
  assign \nz.mem [3210] = \nz.mem_3210_sv2v_reg ;
  assign \nz.mem [3209] = \nz.mem_3209_sv2v_reg ;
  assign \nz.mem [3208] = \nz.mem_3208_sv2v_reg ;
  assign \nz.mem [3207] = \nz.mem_3207_sv2v_reg ;
  assign \nz.mem [3206] = \nz.mem_3206_sv2v_reg ;
  assign \nz.mem [3205] = \nz.mem_3205_sv2v_reg ;
  assign \nz.mem [3204] = \nz.mem_3204_sv2v_reg ;
  assign \nz.mem [3203] = \nz.mem_3203_sv2v_reg ;
  assign \nz.mem [3202] = \nz.mem_3202_sv2v_reg ;
  assign \nz.mem [3201] = \nz.mem_3201_sv2v_reg ;
  assign \nz.mem [3200] = \nz.mem_3200_sv2v_reg ;
  assign \nz.mem [3199] = \nz.mem_3199_sv2v_reg ;
  assign \nz.mem [3198] = \nz.mem_3198_sv2v_reg ;
  assign \nz.mem [3197] = \nz.mem_3197_sv2v_reg ;
  assign \nz.mem [3196] = \nz.mem_3196_sv2v_reg ;
  assign \nz.mem [3195] = \nz.mem_3195_sv2v_reg ;
  assign \nz.mem [3194] = \nz.mem_3194_sv2v_reg ;
  assign \nz.mem [3193] = \nz.mem_3193_sv2v_reg ;
  assign \nz.mem [3192] = \nz.mem_3192_sv2v_reg ;
  assign \nz.mem [3191] = \nz.mem_3191_sv2v_reg ;
  assign \nz.mem [3190] = \nz.mem_3190_sv2v_reg ;
  assign \nz.mem [3189] = \nz.mem_3189_sv2v_reg ;
  assign \nz.mem [3188] = \nz.mem_3188_sv2v_reg ;
  assign \nz.mem [3187] = \nz.mem_3187_sv2v_reg ;
  assign \nz.mem [3186] = \nz.mem_3186_sv2v_reg ;
  assign \nz.mem [3185] = \nz.mem_3185_sv2v_reg ;
  assign \nz.mem [3184] = \nz.mem_3184_sv2v_reg ;
  assign \nz.mem [3183] = \nz.mem_3183_sv2v_reg ;
  assign \nz.mem [3182] = \nz.mem_3182_sv2v_reg ;
  assign \nz.mem [3181] = \nz.mem_3181_sv2v_reg ;
  assign \nz.mem [3180] = \nz.mem_3180_sv2v_reg ;
  assign \nz.mem [3179] = \nz.mem_3179_sv2v_reg ;
  assign \nz.mem [3178] = \nz.mem_3178_sv2v_reg ;
  assign \nz.mem [3177] = \nz.mem_3177_sv2v_reg ;
  assign \nz.mem [3176] = \nz.mem_3176_sv2v_reg ;
  assign \nz.mem [3175] = \nz.mem_3175_sv2v_reg ;
  assign \nz.mem [3174] = \nz.mem_3174_sv2v_reg ;
  assign \nz.mem [3173] = \nz.mem_3173_sv2v_reg ;
  assign \nz.mem [3172] = \nz.mem_3172_sv2v_reg ;
  assign \nz.mem [3171] = \nz.mem_3171_sv2v_reg ;
  assign \nz.mem [3170] = \nz.mem_3170_sv2v_reg ;
  assign \nz.mem [3169] = \nz.mem_3169_sv2v_reg ;
  assign \nz.mem [3168] = \nz.mem_3168_sv2v_reg ;
  assign \nz.mem [3167] = \nz.mem_3167_sv2v_reg ;
  assign \nz.mem [3166] = \nz.mem_3166_sv2v_reg ;
  assign \nz.mem [3165] = \nz.mem_3165_sv2v_reg ;
  assign \nz.mem [3164] = \nz.mem_3164_sv2v_reg ;
  assign \nz.mem [3163] = \nz.mem_3163_sv2v_reg ;
  assign \nz.mem [3162] = \nz.mem_3162_sv2v_reg ;
  assign \nz.mem [3161] = \nz.mem_3161_sv2v_reg ;
  assign \nz.mem [3160] = \nz.mem_3160_sv2v_reg ;
  assign \nz.mem [3159] = \nz.mem_3159_sv2v_reg ;
  assign \nz.mem [3158] = \nz.mem_3158_sv2v_reg ;
  assign \nz.mem [3157] = \nz.mem_3157_sv2v_reg ;
  assign \nz.mem [3156] = \nz.mem_3156_sv2v_reg ;
  assign \nz.mem [3155] = \nz.mem_3155_sv2v_reg ;
  assign \nz.mem [3154] = \nz.mem_3154_sv2v_reg ;
  assign \nz.mem [3153] = \nz.mem_3153_sv2v_reg ;
  assign \nz.mem [3152] = \nz.mem_3152_sv2v_reg ;
  assign \nz.mem [3151] = \nz.mem_3151_sv2v_reg ;
  assign \nz.mem [3150] = \nz.mem_3150_sv2v_reg ;
  assign \nz.mem [3149] = \nz.mem_3149_sv2v_reg ;
  assign \nz.mem [3148] = \nz.mem_3148_sv2v_reg ;
  assign \nz.mem [3147] = \nz.mem_3147_sv2v_reg ;
  assign \nz.mem [3146] = \nz.mem_3146_sv2v_reg ;
  assign \nz.mem [3145] = \nz.mem_3145_sv2v_reg ;
  assign \nz.mem [3144] = \nz.mem_3144_sv2v_reg ;
  assign \nz.mem [3143] = \nz.mem_3143_sv2v_reg ;
  assign \nz.mem [3142] = \nz.mem_3142_sv2v_reg ;
  assign \nz.mem [3141] = \nz.mem_3141_sv2v_reg ;
  assign \nz.mem [3140] = \nz.mem_3140_sv2v_reg ;
  assign \nz.mem [3139] = \nz.mem_3139_sv2v_reg ;
  assign \nz.mem [3138] = \nz.mem_3138_sv2v_reg ;
  assign \nz.mem [3137] = \nz.mem_3137_sv2v_reg ;
  assign \nz.mem [3136] = \nz.mem_3136_sv2v_reg ;
  assign \nz.mem [3135] = \nz.mem_3135_sv2v_reg ;
  assign \nz.mem [3134] = \nz.mem_3134_sv2v_reg ;
  assign \nz.mem [3133] = \nz.mem_3133_sv2v_reg ;
  assign \nz.mem [3132] = \nz.mem_3132_sv2v_reg ;
  assign \nz.mem [3131] = \nz.mem_3131_sv2v_reg ;
  assign \nz.mem [3130] = \nz.mem_3130_sv2v_reg ;
  assign \nz.mem [3129] = \nz.mem_3129_sv2v_reg ;
  assign \nz.mem [3128] = \nz.mem_3128_sv2v_reg ;
  assign \nz.mem [3127] = \nz.mem_3127_sv2v_reg ;
  assign \nz.mem [3126] = \nz.mem_3126_sv2v_reg ;
  assign \nz.mem [3125] = \nz.mem_3125_sv2v_reg ;
  assign \nz.mem [3124] = \nz.mem_3124_sv2v_reg ;
  assign \nz.mem [3123] = \nz.mem_3123_sv2v_reg ;
  assign \nz.mem [3122] = \nz.mem_3122_sv2v_reg ;
  assign \nz.mem [3121] = \nz.mem_3121_sv2v_reg ;
  assign \nz.mem [3120] = \nz.mem_3120_sv2v_reg ;
  assign \nz.mem [3119] = \nz.mem_3119_sv2v_reg ;
  assign \nz.mem [3118] = \nz.mem_3118_sv2v_reg ;
  assign \nz.mem [3117] = \nz.mem_3117_sv2v_reg ;
  assign \nz.mem [3116] = \nz.mem_3116_sv2v_reg ;
  assign \nz.mem [3115] = \nz.mem_3115_sv2v_reg ;
  assign \nz.mem [3114] = \nz.mem_3114_sv2v_reg ;
  assign \nz.mem [3113] = \nz.mem_3113_sv2v_reg ;
  assign \nz.mem [3112] = \nz.mem_3112_sv2v_reg ;
  assign \nz.mem [3111] = \nz.mem_3111_sv2v_reg ;
  assign \nz.mem [3110] = \nz.mem_3110_sv2v_reg ;
  assign \nz.mem [3109] = \nz.mem_3109_sv2v_reg ;
  assign \nz.mem [3108] = \nz.mem_3108_sv2v_reg ;
  assign \nz.mem [3107] = \nz.mem_3107_sv2v_reg ;
  assign \nz.mem [3106] = \nz.mem_3106_sv2v_reg ;
  assign \nz.mem [3105] = \nz.mem_3105_sv2v_reg ;
  assign \nz.mem [3104] = \nz.mem_3104_sv2v_reg ;
  assign \nz.mem [3103] = \nz.mem_3103_sv2v_reg ;
  assign \nz.mem [3102] = \nz.mem_3102_sv2v_reg ;
  assign \nz.mem [3101] = \nz.mem_3101_sv2v_reg ;
  assign \nz.mem [3100] = \nz.mem_3100_sv2v_reg ;
  assign \nz.mem [3099] = \nz.mem_3099_sv2v_reg ;
  assign \nz.mem [3098] = \nz.mem_3098_sv2v_reg ;
  assign \nz.mem [3097] = \nz.mem_3097_sv2v_reg ;
  assign \nz.mem [3096] = \nz.mem_3096_sv2v_reg ;
  assign \nz.mem [3095] = \nz.mem_3095_sv2v_reg ;
  assign \nz.mem [3094] = \nz.mem_3094_sv2v_reg ;
  assign \nz.mem [3093] = \nz.mem_3093_sv2v_reg ;
  assign \nz.mem [3092] = \nz.mem_3092_sv2v_reg ;
  assign \nz.mem [3091] = \nz.mem_3091_sv2v_reg ;
  assign \nz.mem [3090] = \nz.mem_3090_sv2v_reg ;
  assign \nz.mem [3089] = \nz.mem_3089_sv2v_reg ;
  assign \nz.mem [3088] = \nz.mem_3088_sv2v_reg ;
  assign \nz.mem [3087] = \nz.mem_3087_sv2v_reg ;
  assign \nz.mem [3086] = \nz.mem_3086_sv2v_reg ;
  assign \nz.mem [3085] = \nz.mem_3085_sv2v_reg ;
  assign \nz.mem [3084] = \nz.mem_3084_sv2v_reg ;
  assign \nz.mem [3083] = \nz.mem_3083_sv2v_reg ;
  assign \nz.mem [3082] = \nz.mem_3082_sv2v_reg ;
  assign \nz.mem [3081] = \nz.mem_3081_sv2v_reg ;
  assign \nz.mem [3080] = \nz.mem_3080_sv2v_reg ;
  assign \nz.mem [3079] = \nz.mem_3079_sv2v_reg ;
  assign \nz.mem [3078] = \nz.mem_3078_sv2v_reg ;
  assign \nz.mem [3077] = \nz.mem_3077_sv2v_reg ;
  assign \nz.mem [3076] = \nz.mem_3076_sv2v_reg ;
  assign \nz.mem [3075] = \nz.mem_3075_sv2v_reg ;
  assign \nz.mem [3074] = \nz.mem_3074_sv2v_reg ;
  assign \nz.mem [3073] = \nz.mem_3073_sv2v_reg ;
  assign \nz.mem [3072] = \nz.mem_3072_sv2v_reg ;
  assign \nz.mem [3071] = \nz.mem_3071_sv2v_reg ;
  assign \nz.mem [3070] = \nz.mem_3070_sv2v_reg ;
  assign \nz.mem [3069] = \nz.mem_3069_sv2v_reg ;
  assign \nz.mem [3068] = \nz.mem_3068_sv2v_reg ;
  assign \nz.mem [3067] = \nz.mem_3067_sv2v_reg ;
  assign \nz.mem [3066] = \nz.mem_3066_sv2v_reg ;
  assign \nz.mem [3065] = \nz.mem_3065_sv2v_reg ;
  assign \nz.mem [3064] = \nz.mem_3064_sv2v_reg ;
  assign \nz.mem [3063] = \nz.mem_3063_sv2v_reg ;
  assign \nz.mem [3062] = \nz.mem_3062_sv2v_reg ;
  assign \nz.mem [3061] = \nz.mem_3061_sv2v_reg ;
  assign \nz.mem [3060] = \nz.mem_3060_sv2v_reg ;
  assign \nz.mem [3059] = \nz.mem_3059_sv2v_reg ;
  assign \nz.mem [3058] = \nz.mem_3058_sv2v_reg ;
  assign \nz.mem [3057] = \nz.mem_3057_sv2v_reg ;
  assign \nz.mem [3056] = \nz.mem_3056_sv2v_reg ;
  assign \nz.mem [3055] = \nz.mem_3055_sv2v_reg ;
  assign \nz.mem [3054] = \nz.mem_3054_sv2v_reg ;
  assign \nz.mem [3053] = \nz.mem_3053_sv2v_reg ;
  assign \nz.mem [3052] = \nz.mem_3052_sv2v_reg ;
  assign \nz.mem [3051] = \nz.mem_3051_sv2v_reg ;
  assign \nz.mem [3050] = \nz.mem_3050_sv2v_reg ;
  assign \nz.mem [3049] = \nz.mem_3049_sv2v_reg ;
  assign \nz.mem [3048] = \nz.mem_3048_sv2v_reg ;
  assign \nz.mem [3047] = \nz.mem_3047_sv2v_reg ;
  assign \nz.mem [3046] = \nz.mem_3046_sv2v_reg ;
  assign \nz.mem [3045] = \nz.mem_3045_sv2v_reg ;
  assign \nz.mem [3044] = \nz.mem_3044_sv2v_reg ;
  assign \nz.mem [3043] = \nz.mem_3043_sv2v_reg ;
  assign \nz.mem [3042] = \nz.mem_3042_sv2v_reg ;
  assign \nz.mem [3041] = \nz.mem_3041_sv2v_reg ;
  assign \nz.mem [3040] = \nz.mem_3040_sv2v_reg ;
  assign \nz.mem [3039] = \nz.mem_3039_sv2v_reg ;
  assign \nz.mem [3038] = \nz.mem_3038_sv2v_reg ;
  assign \nz.mem [3037] = \nz.mem_3037_sv2v_reg ;
  assign \nz.mem [3036] = \nz.mem_3036_sv2v_reg ;
  assign \nz.mem [3035] = \nz.mem_3035_sv2v_reg ;
  assign \nz.mem [3034] = \nz.mem_3034_sv2v_reg ;
  assign \nz.mem [3033] = \nz.mem_3033_sv2v_reg ;
  assign \nz.mem [3032] = \nz.mem_3032_sv2v_reg ;
  assign \nz.mem [3031] = \nz.mem_3031_sv2v_reg ;
  assign \nz.mem [3030] = \nz.mem_3030_sv2v_reg ;
  assign \nz.mem [3029] = \nz.mem_3029_sv2v_reg ;
  assign \nz.mem [3028] = \nz.mem_3028_sv2v_reg ;
  assign \nz.mem [3027] = \nz.mem_3027_sv2v_reg ;
  assign \nz.mem [3026] = \nz.mem_3026_sv2v_reg ;
  assign \nz.mem [3025] = \nz.mem_3025_sv2v_reg ;
  assign \nz.mem [3024] = \nz.mem_3024_sv2v_reg ;
  assign \nz.mem [3023] = \nz.mem_3023_sv2v_reg ;
  assign \nz.mem [3022] = \nz.mem_3022_sv2v_reg ;
  assign \nz.mem [3021] = \nz.mem_3021_sv2v_reg ;
  assign \nz.mem [3020] = \nz.mem_3020_sv2v_reg ;
  assign \nz.mem [3019] = \nz.mem_3019_sv2v_reg ;
  assign \nz.mem [3018] = \nz.mem_3018_sv2v_reg ;
  assign \nz.mem [3017] = \nz.mem_3017_sv2v_reg ;
  assign \nz.mem [3016] = \nz.mem_3016_sv2v_reg ;
  assign \nz.mem [3015] = \nz.mem_3015_sv2v_reg ;
  assign \nz.mem [3014] = \nz.mem_3014_sv2v_reg ;
  assign \nz.mem [3013] = \nz.mem_3013_sv2v_reg ;
  assign \nz.mem [3012] = \nz.mem_3012_sv2v_reg ;
  assign \nz.mem [3011] = \nz.mem_3011_sv2v_reg ;
  assign \nz.mem [3010] = \nz.mem_3010_sv2v_reg ;
  assign \nz.mem [3009] = \nz.mem_3009_sv2v_reg ;
  assign \nz.mem [3008] = \nz.mem_3008_sv2v_reg ;
  assign \nz.mem [3007] = \nz.mem_3007_sv2v_reg ;
  assign \nz.mem [3006] = \nz.mem_3006_sv2v_reg ;
  assign \nz.mem [3005] = \nz.mem_3005_sv2v_reg ;
  assign \nz.mem [3004] = \nz.mem_3004_sv2v_reg ;
  assign \nz.mem [3003] = \nz.mem_3003_sv2v_reg ;
  assign \nz.mem [3002] = \nz.mem_3002_sv2v_reg ;
  assign \nz.mem [3001] = \nz.mem_3001_sv2v_reg ;
  assign \nz.mem [3000] = \nz.mem_3000_sv2v_reg ;
  assign \nz.mem [2999] = \nz.mem_2999_sv2v_reg ;
  assign \nz.mem [2998] = \nz.mem_2998_sv2v_reg ;
  assign \nz.mem [2997] = \nz.mem_2997_sv2v_reg ;
  assign \nz.mem [2996] = \nz.mem_2996_sv2v_reg ;
  assign \nz.mem [2995] = \nz.mem_2995_sv2v_reg ;
  assign \nz.mem [2994] = \nz.mem_2994_sv2v_reg ;
  assign \nz.mem [2993] = \nz.mem_2993_sv2v_reg ;
  assign \nz.mem [2992] = \nz.mem_2992_sv2v_reg ;
  assign \nz.mem [2991] = \nz.mem_2991_sv2v_reg ;
  assign \nz.mem [2990] = \nz.mem_2990_sv2v_reg ;
  assign \nz.mem [2989] = \nz.mem_2989_sv2v_reg ;
  assign \nz.mem [2988] = \nz.mem_2988_sv2v_reg ;
  assign \nz.mem [2987] = \nz.mem_2987_sv2v_reg ;
  assign \nz.mem [2986] = \nz.mem_2986_sv2v_reg ;
  assign \nz.mem [2985] = \nz.mem_2985_sv2v_reg ;
  assign \nz.mem [2984] = \nz.mem_2984_sv2v_reg ;
  assign \nz.mem [2983] = \nz.mem_2983_sv2v_reg ;
  assign \nz.mem [2982] = \nz.mem_2982_sv2v_reg ;
  assign \nz.mem [2981] = \nz.mem_2981_sv2v_reg ;
  assign \nz.mem [2980] = \nz.mem_2980_sv2v_reg ;
  assign \nz.mem [2979] = \nz.mem_2979_sv2v_reg ;
  assign \nz.mem [2978] = \nz.mem_2978_sv2v_reg ;
  assign \nz.mem [2977] = \nz.mem_2977_sv2v_reg ;
  assign \nz.mem [2976] = \nz.mem_2976_sv2v_reg ;
  assign \nz.mem [2975] = \nz.mem_2975_sv2v_reg ;
  assign \nz.mem [2974] = \nz.mem_2974_sv2v_reg ;
  assign \nz.mem [2973] = \nz.mem_2973_sv2v_reg ;
  assign \nz.mem [2972] = \nz.mem_2972_sv2v_reg ;
  assign \nz.mem [2971] = \nz.mem_2971_sv2v_reg ;
  assign \nz.mem [2970] = \nz.mem_2970_sv2v_reg ;
  assign \nz.mem [2969] = \nz.mem_2969_sv2v_reg ;
  assign \nz.mem [2968] = \nz.mem_2968_sv2v_reg ;
  assign \nz.mem [2967] = \nz.mem_2967_sv2v_reg ;
  assign \nz.mem [2966] = \nz.mem_2966_sv2v_reg ;
  assign \nz.mem [2965] = \nz.mem_2965_sv2v_reg ;
  assign \nz.mem [2964] = \nz.mem_2964_sv2v_reg ;
  assign \nz.mem [2963] = \nz.mem_2963_sv2v_reg ;
  assign \nz.mem [2962] = \nz.mem_2962_sv2v_reg ;
  assign \nz.mem [2961] = \nz.mem_2961_sv2v_reg ;
  assign \nz.mem [2960] = \nz.mem_2960_sv2v_reg ;
  assign \nz.mem [2959] = \nz.mem_2959_sv2v_reg ;
  assign \nz.mem [2958] = \nz.mem_2958_sv2v_reg ;
  assign \nz.mem [2957] = \nz.mem_2957_sv2v_reg ;
  assign \nz.mem [2956] = \nz.mem_2956_sv2v_reg ;
  assign \nz.mem [2955] = \nz.mem_2955_sv2v_reg ;
  assign \nz.mem [2954] = \nz.mem_2954_sv2v_reg ;
  assign \nz.mem [2953] = \nz.mem_2953_sv2v_reg ;
  assign \nz.mem [2952] = \nz.mem_2952_sv2v_reg ;
  assign \nz.mem [2951] = \nz.mem_2951_sv2v_reg ;
  assign \nz.mem [2950] = \nz.mem_2950_sv2v_reg ;
  assign \nz.mem [2949] = \nz.mem_2949_sv2v_reg ;
  assign \nz.mem [2948] = \nz.mem_2948_sv2v_reg ;
  assign \nz.mem [2947] = \nz.mem_2947_sv2v_reg ;
  assign \nz.mem [2946] = \nz.mem_2946_sv2v_reg ;
  assign \nz.mem [2945] = \nz.mem_2945_sv2v_reg ;
  assign \nz.mem [2944] = \nz.mem_2944_sv2v_reg ;
  assign \nz.mem [2943] = \nz.mem_2943_sv2v_reg ;
  assign \nz.mem [2942] = \nz.mem_2942_sv2v_reg ;
  assign \nz.mem [2941] = \nz.mem_2941_sv2v_reg ;
  assign \nz.mem [2940] = \nz.mem_2940_sv2v_reg ;
  assign \nz.mem [2939] = \nz.mem_2939_sv2v_reg ;
  assign \nz.mem [2938] = \nz.mem_2938_sv2v_reg ;
  assign \nz.mem [2937] = \nz.mem_2937_sv2v_reg ;
  assign \nz.mem [2936] = \nz.mem_2936_sv2v_reg ;
  assign \nz.mem [2935] = \nz.mem_2935_sv2v_reg ;
  assign \nz.mem [2934] = \nz.mem_2934_sv2v_reg ;
  assign \nz.mem [2933] = \nz.mem_2933_sv2v_reg ;
  assign \nz.mem [2932] = \nz.mem_2932_sv2v_reg ;
  assign \nz.mem [2931] = \nz.mem_2931_sv2v_reg ;
  assign \nz.mem [2930] = \nz.mem_2930_sv2v_reg ;
  assign \nz.mem [2929] = \nz.mem_2929_sv2v_reg ;
  assign \nz.mem [2928] = \nz.mem_2928_sv2v_reg ;
  assign \nz.mem [2927] = \nz.mem_2927_sv2v_reg ;
  assign \nz.mem [2926] = \nz.mem_2926_sv2v_reg ;
  assign \nz.mem [2925] = \nz.mem_2925_sv2v_reg ;
  assign \nz.mem [2924] = \nz.mem_2924_sv2v_reg ;
  assign \nz.mem [2923] = \nz.mem_2923_sv2v_reg ;
  assign \nz.mem [2922] = \nz.mem_2922_sv2v_reg ;
  assign \nz.mem [2921] = \nz.mem_2921_sv2v_reg ;
  assign \nz.mem [2920] = \nz.mem_2920_sv2v_reg ;
  assign \nz.mem [2919] = \nz.mem_2919_sv2v_reg ;
  assign \nz.mem [2918] = \nz.mem_2918_sv2v_reg ;
  assign \nz.mem [2917] = \nz.mem_2917_sv2v_reg ;
  assign \nz.mem [2916] = \nz.mem_2916_sv2v_reg ;
  assign \nz.mem [2915] = \nz.mem_2915_sv2v_reg ;
  assign \nz.mem [2914] = \nz.mem_2914_sv2v_reg ;
  assign \nz.mem [2913] = \nz.mem_2913_sv2v_reg ;
  assign \nz.mem [2912] = \nz.mem_2912_sv2v_reg ;
  assign \nz.mem [2911] = \nz.mem_2911_sv2v_reg ;
  assign \nz.mem [2910] = \nz.mem_2910_sv2v_reg ;
  assign \nz.mem [2909] = \nz.mem_2909_sv2v_reg ;
  assign \nz.mem [2908] = \nz.mem_2908_sv2v_reg ;
  assign \nz.mem [2907] = \nz.mem_2907_sv2v_reg ;
  assign \nz.mem [2906] = \nz.mem_2906_sv2v_reg ;
  assign \nz.mem [2905] = \nz.mem_2905_sv2v_reg ;
  assign \nz.mem [2904] = \nz.mem_2904_sv2v_reg ;
  assign \nz.mem [2903] = \nz.mem_2903_sv2v_reg ;
  assign \nz.mem [2902] = \nz.mem_2902_sv2v_reg ;
  assign \nz.mem [2901] = \nz.mem_2901_sv2v_reg ;
  assign \nz.mem [2900] = \nz.mem_2900_sv2v_reg ;
  assign \nz.mem [2899] = \nz.mem_2899_sv2v_reg ;
  assign \nz.mem [2898] = \nz.mem_2898_sv2v_reg ;
  assign \nz.mem [2897] = \nz.mem_2897_sv2v_reg ;
  assign \nz.mem [2896] = \nz.mem_2896_sv2v_reg ;
  assign \nz.mem [2895] = \nz.mem_2895_sv2v_reg ;
  assign \nz.mem [2894] = \nz.mem_2894_sv2v_reg ;
  assign \nz.mem [2893] = \nz.mem_2893_sv2v_reg ;
  assign \nz.mem [2892] = \nz.mem_2892_sv2v_reg ;
  assign \nz.mem [2891] = \nz.mem_2891_sv2v_reg ;
  assign \nz.mem [2890] = \nz.mem_2890_sv2v_reg ;
  assign \nz.mem [2889] = \nz.mem_2889_sv2v_reg ;
  assign \nz.mem [2888] = \nz.mem_2888_sv2v_reg ;
  assign \nz.mem [2887] = \nz.mem_2887_sv2v_reg ;
  assign \nz.mem [2886] = \nz.mem_2886_sv2v_reg ;
  assign \nz.mem [2885] = \nz.mem_2885_sv2v_reg ;
  assign \nz.mem [2884] = \nz.mem_2884_sv2v_reg ;
  assign \nz.mem [2883] = \nz.mem_2883_sv2v_reg ;
  assign \nz.mem [2882] = \nz.mem_2882_sv2v_reg ;
  assign \nz.mem [2881] = \nz.mem_2881_sv2v_reg ;
  assign \nz.mem [2880] = \nz.mem_2880_sv2v_reg ;
  assign \nz.mem [2879] = \nz.mem_2879_sv2v_reg ;
  assign \nz.mem [2878] = \nz.mem_2878_sv2v_reg ;
  assign \nz.mem [2877] = \nz.mem_2877_sv2v_reg ;
  assign \nz.mem [2876] = \nz.mem_2876_sv2v_reg ;
  assign \nz.mem [2875] = \nz.mem_2875_sv2v_reg ;
  assign \nz.mem [2874] = \nz.mem_2874_sv2v_reg ;
  assign \nz.mem [2873] = \nz.mem_2873_sv2v_reg ;
  assign \nz.mem [2872] = \nz.mem_2872_sv2v_reg ;
  assign \nz.mem [2871] = \nz.mem_2871_sv2v_reg ;
  assign \nz.mem [2870] = \nz.mem_2870_sv2v_reg ;
  assign \nz.mem [2869] = \nz.mem_2869_sv2v_reg ;
  assign \nz.mem [2868] = \nz.mem_2868_sv2v_reg ;
  assign \nz.mem [2867] = \nz.mem_2867_sv2v_reg ;
  assign \nz.mem [2866] = \nz.mem_2866_sv2v_reg ;
  assign \nz.mem [2865] = \nz.mem_2865_sv2v_reg ;
  assign \nz.mem [2864] = \nz.mem_2864_sv2v_reg ;
  assign \nz.mem [2863] = \nz.mem_2863_sv2v_reg ;
  assign \nz.mem [2862] = \nz.mem_2862_sv2v_reg ;
  assign \nz.mem [2861] = \nz.mem_2861_sv2v_reg ;
  assign \nz.mem [2860] = \nz.mem_2860_sv2v_reg ;
  assign \nz.mem [2859] = \nz.mem_2859_sv2v_reg ;
  assign \nz.mem [2858] = \nz.mem_2858_sv2v_reg ;
  assign \nz.mem [2857] = \nz.mem_2857_sv2v_reg ;
  assign \nz.mem [2856] = \nz.mem_2856_sv2v_reg ;
  assign \nz.mem [2855] = \nz.mem_2855_sv2v_reg ;
  assign \nz.mem [2854] = \nz.mem_2854_sv2v_reg ;
  assign \nz.mem [2853] = \nz.mem_2853_sv2v_reg ;
  assign \nz.mem [2852] = \nz.mem_2852_sv2v_reg ;
  assign \nz.mem [2851] = \nz.mem_2851_sv2v_reg ;
  assign \nz.mem [2850] = \nz.mem_2850_sv2v_reg ;
  assign \nz.mem [2849] = \nz.mem_2849_sv2v_reg ;
  assign \nz.mem [2848] = \nz.mem_2848_sv2v_reg ;
  assign \nz.mem [2847] = \nz.mem_2847_sv2v_reg ;
  assign \nz.mem [2846] = \nz.mem_2846_sv2v_reg ;
  assign \nz.mem [2845] = \nz.mem_2845_sv2v_reg ;
  assign \nz.mem [2844] = \nz.mem_2844_sv2v_reg ;
  assign \nz.mem [2843] = \nz.mem_2843_sv2v_reg ;
  assign \nz.mem [2842] = \nz.mem_2842_sv2v_reg ;
  assign \nz.mem [2841] = \nz.mem_2841_sv2v_reg ;
  assign \nz.mem [2840] = \nz.mem_2840_sv2v_reg ;
  assign \nz.mem [2839] = \nz.mem_2839_sv2v_reg ;
  assign \nz.mem [2838] = \nz.mem_2838_sv2v_reg ;
  assign \nz.mem [2837] = \nz.mem_2837_sv2v_reg ;
  assign \nz.mem [2836] = \nz.mem_2836_sv2v_reg ;
  assign \nz.mem [2835] = \nz.mem_2835_sv2v_reg ;
  assign \nz.mem [2834] = \nz.mem_2834_sv2v_reg ;
  assign \nz.mem [2833] = \nz.mem_2833_sv2v_reg ;
  assign \nz.mem [2832] = \nz.mem_2832_sv2v_reg ;
  assign \nz.mem [2831] = \nz.mem_2831_sv2v_reg ;
  assign \nz.mem [2830] = \nz.mem_2830_sv2v_reg ;
  assign \nz.mem [2829] = \nz.mem_2829_sv2v_reg ;
  assign \nz.mem [2828] = \nz.mem_2828_sv2v_reg ;
  assign \nz.mem [2827] = \nz.mem_2827_sv2v_reg ;
  assign \nz.mem [2826] = \nz.mem_2826_sv2v_reg ;
  assign \nz.mem [2825] = \nz.mem_2825_sv2v_reg ;
  assign \nz.mem [2824] = \nz.mem_2824_sv2v_reg ;
  assign \nz.mem [2823] = \nz.mem_2823_sv2v_reg ;
  assign \nz.mem [2822] = \nz.mem_2822_sv2v_reg ;
  assign \nz.mem [2821] = \nz.mem_2821_sv2v_reg ;
  assign \nz.mem [2820] = \nz.mem_2820_sv2v_reg ;
  assign \nz.mem [2819] = \nz.mem_2819_sv2v_reg ;
  assign \nz.mem [2818] = \nz.mem_2818_sv2v_reg ;
  assign \nz.mem [2817] = \nz.mem_2817_sv2v_reg ;
  assign \nz.mem [2816] = \nz.mem_2816_sv2v_reg ;
  assign \nz.mem [2815] = \nz.mem_2815_sv2v_reg ;
  assign \nz.mem [2814] = \nz.mem_2814_sv2v_reg ;
  assign \nz.mem [2813] = \nz.mem_2813_sv2v_reg ;
  assign \nz.mem [2812] = \nz.mem_2812_sv2v_reg ;
  assign \nz.mem [2811] = \nz.mem_2811_sv2v_reg ;
  assign \nz.mem [2810] = \nz.mem_2810_sv2v_reg ;
  assign \nz.mem [2809] = \nz.mem_2809_sv2v_reg ;
  assign \nz.mem [2808] = \nz.mem_2808_sv2v_reg ;
  assign \nz.mem [2807] = \nz.mem_2807_sv2v_reg ;
  assign \nz.mem [2806] = \nz.mem_2806_sv2v_reg ;
  assign \nz.mem [2805] = \nz.mem_2805_sv2v_reg ;
  assign \nz.mem [2804] = \nz.mem_2804_sv2v_reg ;
  assign \nz.mem [2803] = \nz.mem_2803_sv2v_reg ;
  assign \nz.mem [2802] = \nz.mem_2802_sv2v_reg ;
  assign \nz.mem [2801] = \nz.mem_2801_sv2v_reg ;
  assign \nz.mem [2800] = \nz.mem_2800_sv2v_reg ;
  assign \nz.mem [2799] = \nz.mem_2799_sv2v_reg ;
  assign \nz.mem [2798] = \nz.mem_2798_sv2v_reg ;
  assign \nz.mem [2797] = \nz.mem_2797_sv2v_reg ;
  assign \nz.mem [2796] = \nz.mem_2796_sv2v_reg ;
  assign \nz.mem [2795] = \nz.mem_2795_sv2v_reg ;
  assign \nz.mem [2794] = \nz.mem_2794_sv2v_reg ;
  assign \nz.mem [2793] = \nz.mem_2793_sv2v_reg ;
  assign \nz.mem [2792] = \nz.mem_2792_sv2v_reg ;
  assign \nz.mem [2791] = \nz.mem_2791_sv2v_reg ;
  assign \nz.mem [2790] = \nz.mem_2790_sv2v_reg ;
  assign \nz.mem [2789] = \nz.mem_2789_sv2v_reg ;
  assign \nz.mem [2788] = \nz.mem_2788_sv2v_reg ;
  assign \nz.mem [2787] = \nz.mem_2787_sv2v_reg ;
  assign \nz.mem [2786] = \nz.mem_2786_sv2v_reg ;
  assign \nz.mem [2785] = \nz.mem_2785_sv2v_reg ;
  assign \nz.mem [2784] = \nz.mem_2784_sv2v_reg ;
  assign \nz.mem [2783] = \nz.mem_2783_sv2v_reg ;
  assign \nz.mem [2782] = \nz.mem_2782_sv2v_reg ;
  assign \nz.mem [2781] = \nz.mem_2781_sv2v_reg ;
  assign \nz.mem [2780] = \nz.mem_2780_sv2v_reg ;
  assign \nz.mem [2779] = \nz.mem_2779_sv2v_reg ;
  assign \nz.mem [2778] = \nz.mem_2778_sv2v_reg ;
  assign \nz.mem [2777] = \nz.mem_2777_sv2v_reg ;
  assign \nz.mem [2776] = \nz.mem_2776_sv2v_reg ;
  assign \nz.mem [2775] = \nz.mem_2775_sv2v_reg ;
  assign \nz.mem [2774] = \nz.mem_2774_sv2v_reg ;
  assign \nz.mem [2773] = \nz.mem_2773_sv2v_reg ;
  assign \nz.mem [2772] = \nz.mem_2772_sv2v_reg ;
  assign \nz.mem [2771] = \nz.mem_2771_sv2v_reg ;
  assign \nz.mem [2770] = \nz.mem_2770_sv2v_reg ;
  assign \nz.mem [2769] = \nz.mem_2769_sv2v_reg ;
  assign \nz.mem [2768] = \nz.mem_2768_sv2v_reg ;
  assign \nz.mem [2767] = \nz.mem_2767_sv2v_reg ;
  assign \nz.mem [2766] = \nz.mem_2766_sv2v_reg ;
  assign \nz.mem [2765] = \nz.mem_2765_sv2v_reg ;
  assign \nz.mem [2764] = \nz.mem_2764_sv2v_reg ;
  assign \nz.mem [2763] = \nz.mem_2763_sv2v_reg ;
  assign \nz.mem [2762] = \nz.mem_2762_sv2v_reg ;
  assign \nz.mem [2761] = \nz.mem_2761_sv2v_reg ;
  assign \nz.mem [2760] = \nz.mem_2760_sv2v_reg ;
  assign \nz.mem [2759] = \nz.mem_2759_sv2v_reg ;
  assign \nz.mem [2758] = \nz.mem_2758_sv2v_reg ;
  assign \nz.mem [2757] = \nz.mem_2757_sv2v_reg ;
  assign \nz.mem [2756] = \nz.mem_2756_sv2v_reg ;
  assign \nz.mem [2755] = \nz.mem_2755_sv2v_reg ;
  assign \nz.mem [2754] = \nz.mem_2754_sv2v_reg ;
  assign \nz.mem [2753] = \nz.mem_2753_sv2v_reg ;
  assign \nz.mem [2752] = \nz.mem_2752_sv2v_reg ;
  assign \nz.mem [2751] = \nz.mem_2751_sv2v_reg ;
  assign \nz.mem [2750] = \nz.mem_2750_sv2v_reg ;
  assign \nz.mem [2749] = \nz.mem_2749_sv2v_reg ;
  assign \nz.mem [2748] = \nz.mem_2748_sv2v_reg ;
  assign \nz.mem [2747] = \nz.mem_2747_sv2v_reg ;
  assign \nz.mem [2746] = \nz.mem_2746_sv2v_reg ;
  assign \nz.mem [2745] = \nz.mem_2745_sv2v_reg ;
  assign \nz.mem [2744] = \nz.mem_2744_sv2v_reg ;
  assign \nz.mem [2743] = \nz.mem_2743_sv2v_reg ;
  assign \nz.mem [2742] = \nz.mem_2742_sv2v_reg ;
  assign \nz.mem [2741] = \nz.mem_2741_sv2v_reg ;
  assign \nz.mem [2740] = \nz.mem_2740_sv2v_reg ;
  assign \nz.mem [2739] = \nz.mem_2739_sv2v_reg ;
  assign \nz.mem [2738] = \nz.mem_2738_sv2v_reg ;
  assign \nz.mem [2737] = \nz.mem_2737_sv2v_reg ;
  assign \nz.mem [2736] = \nz.mem_2736_sv2v_reg ;
  assign \nz.mem [2735] = \nz.mem_2735_sv2v_reg ;
  assign \nz.mem [2734] = \nz.mem_2734_sv2v_reg ;
  assign \nz.mem [2733] = \nz.mem_2733_sv2v_reg ;
  assign \nz.mem [2732] = \nz.mem_2732_sv2v_reg ;
  assign \nz.mem [2731] = \nz.mem_2731_sv2v_reg ;
  assign \nz.mem [2730] = \nz.mem_2730_sv2v_reg ;
  assign \nz.mem [2729] = \nz.mem_2729_sv2v_reg ;
  assign \nz.mem [2728] = \nz.mem_2728_sv2v_reg ;
  assign \nz.mem [2727] = \nz.mem_2727_sv2v_reg ;
  assign \nz.mem [2726] = \nz.mem_2726_sv2v_reg ;
  assign \nz.mem [2725] = \nz.mem_2725_sv2v_reg ;
  assign \nz.mem [2724] = \nz.mem_2724_sv2v_reg ;
  assign \nz.mem [2723] = \nz.mem_2723_sv2v_reg ;
  assign \nz.mem [2722] = \nz.mem_2722_sv2v_reg ;
  assign \nz.mem [2721] = \nz.mem_2721_sv2v_reg ;
  assign \nz.mem [2720] = \nz.mem_2720_sv2v_reg ;
  assign \nz.mem [2719] = \nz.mem_2719_sv2v_reg ;
  assign \nz.mem [2718] = \nz.mem_2718_sv2v_reg ;
  assign \nz.mem [2717] = \nz.mem_2717_sv2v_reg ;
  assign \nz.mem [2716] = \nz.mem_2716_sv2v_reg ;
  assign \nz.mem [2715] = \nz.mem_2715_sv2v_reg ;
  assign \nz.mem [2714] = \nz.mem_2714_sv2v_reg ;
  assign \nz.mem [2713] = \nz.mem_2713_sv2v_reg ;
  assign \nz.mem [2712] = \nz.mem_2712_sv2v_reg ;
  assign \nz.mem [2711] = \nz.mem_2711_sv2v_reg ;
  assign \nz.mem [2710] = \nz.mem_2710_sv2v_reg ;
  assign \nz.mem [2709] = \nz.mem_2709_sv2v_reg ;
  assign \nz.mem [2708] = \nz.mem_2708_sv2v_reg ;
  assign \nz.mem [2707] = \nz.mem_2707_sv2v_reg ;
  assign \nz.mem [2706] = \nz.mem_2706_sv2v_reg ;
  assign \nz.mem [2705] = \nz.mem_2705_sv2v_reg ;
  assign \nz.mem [2704] = \nz.mem_2704_sv2v_reg ;
  assign \nz.mem [2703] = \nz.mem_2703_sv2v_reg ;
  assign \nz.mem [2702] = \nz.mem_2702_sv2v_reg ;
  assign \nz.mem [2701] = \nz.mem_2701_sv2v_reg ;
  assign \nz.mem [2700] = \nz.mem_2700_sv2v_reg ;
  assign \nz.mem [2699] = \nz.mem_2699_sv2v_reg ;
  assign \nz.mem [2698] = \nz.mem_2698_sv2v_reg ;
  assign \nz.mem [2697] = \nz.mem_2697_sv2v_reg ;
  assign \nz.mem [2696] = \nz.mem_2696_sv2v_reg ;
  assign \nz.mem [2695] = \nz.mem_2695_sv2v_reg ;
  assign \nz.mem [2694] = \nz.mem_2694_sv2v_reg ;
  assign \nz.mem [2693] = \nz.mem_2693_sv2v_reg ;
  assign \nz.mem [2692] = \nz.mem_2692_sv2v_reg ;
  assign \nz.mem [2691] = \nz.mem_2691_sv2v_reg ;
  assign \nz.mem [2690] = \nz.mem_2690_sv2v_reg ;
  assign \nz.mem [2689] = \nz.mem_2689_sv2v_reg ;
  assign \nz.mem [2688] = \nz.mem_2688_sv2v_reg ;
  assign \nz.mem [2687] = \nz.mem_2687_sv2v_reg ;
  assign \nz.mem [2686] = \nz.mem_2686_sv2v_reg ;
  assign \nz.mem [2685] = \nz.mem_2685_sv2v_reg ;
  assign \nz.mem [2684] = \nz.mem_2684_sv2v_reg ;
  assign \nz.mem [2683] = \nz.mem_2683_sv2v_reg ;
  assign \nz.mem [2682] = \nz.mem_2682_sv2v_reg ;
  assign \nz.mem [2681] = \nz.mem_2681_sv2v_reg ;
  assign \nz.mem [2680] = \nz.mem_2680_sv2v_reg ;
  assign \nz.mem [2679] = \nz.mem_2679_sv2v_reg ;
  assign \nz.mem [2678] = \nz.mem_2678_sv2v_reg ;
  assign \nz.mem [2677] = \nz.mem_2677_sv2v_reg ;
  assign \nz.mem [2676] = \nz.mem_2676_sv2v_reg ;
  assign \nz.mem [2675] = \nz.mem_2675_sv2v_reg ;
  assign \nz.mem [2674] = \nz.mem_2674_sv2v_reg ;
  assign \nz.mem [2673] = \nz.mem_2673_sv2v_reg ;
  assign \nz.mem [2672] = \nz.mem_2672_sv2v_reg ;
  assign \nz.mem [2671] = \nz.mem_2671_sv2v_reg ;
  assign \nz.mem [2670] = \nz.mem_2670_sv2v_reg ;
  assign \nz.mem [2669] = \nz.mem_2669_sv2v_reg ;
  assign \nz.mem [2668] = \nz.mem_2668_sv2v_reg ;
  assign \nz.mem [2667] = \nz.mem_2667_sv2v_reg ;
  assign \nz.mem [2666] = \nz.mem_2666_sv2v_reg ;
  assign \nz.mem [2665] = \nz.mem_2665_sv2v_reg ;
  assign \nz.mem [2664] = \nz.mem_2664_sv2v_reg ;
  assign \nz.mem [2663] = \nz.mem_2663_sv2v_reg ;
  assign \nz.mem [2662] = \nz.mem_2662_sv2v_reg ;
  assign \nz.mem [2661] = \nz.mem_2661_sv2v_reg ;
  assign \nz.mem [2660] = \nz.mem_2660_sv2v_reg ;
  assign \nz.mem [2659] = \nz.mem_2659_sv2v_reg ;
  assign \nz.mem [2658] = \nz.mem_2658_sv2v_reg ;
  assign \nz.mem [2657] = \nz.mem_2657_sv2v_reg ;
  assign \nz.mem [2656] = \nz.mem_2656_sv2v_reg ;
  assign \nz.mem [2655] = \nz.mem_2655_sv2v_reg ;
  assign \nz.mem [2654] = \nz.mem_2654_sv2v_reg ;
  assign \nz.mem [2653] = \nz.mem_2653_sv2v_reg ;
  assign \nz.mem [2652] = \nz.mem_2652_sv2v_reg ;
  assign \nz.mem [2651] = \nz.mem_2651_sv2v_reg ;
  assign \nz.mem [2650] = \nz.mem_2650_sv2v_reg ;
  assign \nz.mem [2649] = \nz.mem_2649_sv2v_reg ;
  assign \nz.mem [2648] = \nz.mem_2648_sv2v_reg ;
  assign \nz.mem [2647] = \nz.mem_2647_sv2v_reg ;
  assign \nz.mem [2646] = \nz.mem_2646_sv2v_reg ;
  assign \nz.mem [2645] = \nz.mem_2645_sv2v_reg ;
  assign \nz.mem [2644] = \nz.mem_2644_sv2v_reg ;
  assign \nz.mem [2643] = \nz.mem_2643_sv2v_reg ;
  assign \nz.mem [2642] = \nz.mem_2642_sv2v_reg ;
  assign \nz.mem [2641] = \nz.mem_2641_sv2v_reg ;
  assign \nz.mem [2640] = \nz.mem_2640_sv2v_reg ;
  assign \nz.mem [2639] = \nz.mem_2639_sv2v_reg ;
  assign \nz.mem [2638] = \nz.mem_2638_sv2v_reg ;
  assign \nz.mem [2637] = \nz.mem_2637_sv2v_reg ;
  assign \nz.mem [2636] = \nz.mem_2636_sv2v_reg ;
  assign \nz.mem [2635] = \nz.mem_2635_sv2v_reg ;
  assign \nz.mem [2634] = \nz.mem_2634_sv2v_reg ;
  assign \nz.mem [2633] = \nz.mem_2633_sv2v_reg ;
  assign \nz.mem [2632] = \nz.mem_2632_sv2v_reg ;
  assign \nz.mem [2631] = \nz.mem_2631_sv2v_reg ;
  assign \nz.mem [2630] = \nz.mem_2630_sv2v_reg ;
  assign \nz.mem [2629] = \nz.mem_2629_sv2v_reg ;
  assign \nz.mem [2628] = \nz.mem_2628_sv2v_reg ;
  assign \nz.mem [2627] = \nz.mem_2627_sv2v_reg ;
  assign \nz.mem [2626] = \nz.mem_2626_sv2v_reg ;
  assign \nz.mem [2625] = \nz.mem_2625_sv2v_reg ;
  assign \nz.mem [2624] = \nz.mem_2624_sv2v_reg ;
  assign \nz.mem [2623] = \nz.mem_2623_sv2v_reg ;
  assign \nz.mem [2622] = \nz.mem_2622_sv2v_reg ;
  assign \nz.mem [2621] = \nz.mem_2621_sv2v_reg ;
  assign \nz.mem [2620] = \nz.mem_2620_sv2v_reg ;
  assign \nz.mem [2619] = \nz.mem_2619_sv2v_reg ;
  assign \nz.mem [2618] = \nz.mem_2618_sv2v_reg ;
  assign \nz.mem [2617] = \nz.mem_2617_sv2v_reg ;
  assign \nz.mem [2616] = \nz.mem_2616_sv2v_reg ;
  assign \nz.mem [2615] = \nz.mem_2615_sv2v_reg ;
  assign \nz.mem [2614] = \nz.mem_2614_sv2v_reg ;
  assign \nz.mem [2613] = \nz.mem_2613_sv2v_reg ;
  assign \nz.mem [2612] = \nz.mem_2612_sv2v_reg ;
  assign \nz.mem [2611] = \nz.mem_2611_sv2v_reg ;
  assign \nz.mem [2610] = \nz.mem_2610_sv2v_reg ;
  assign \nz.mem [2609] = \nz.mem_2609_sv2v_reg ;
  assign \nz.mem [2608] = \nz.mem_2608_sv2v_reg ;
  assign \nz.mem [2607] = \nz.mem_2607_sv2v_reg ;
  assign \nz.mem [2606] = \nz.mem_2606_sv2v_reg ;
  assign \nz.mem [2605] = \nz.mem_2605_sv2v_reg ;
  assign \nz.mem [2604] = \nz.mem_2604_sv2v_reg ;
  assign \nz.mem [2603] = \nz.mem_2603_sv2v_reg ;
  assign \nz.mem [2602] = \nz.mem_2602_sv2v_reg ;
  assign \nz.mem [2601] = \nz.mem_2601_sv2v_reg ;
  assign \nz.mem [2600] = \nz.mem_2600_sv2v_reg ;
  assign \nz.mem [2599] = \nz.mem_2599_sv2v_reg ;
  assign \nz.mem [2598] = \nz.mem_2598_sv2v_reg ;
  assign \nz.mem [2597] = \nz.mem_2597_sv2v_reg ;
  assign \nz.mem [2596] = \nz.mem_2596_sv2v_reg ;
  assign \nz.mem [2595] = \nz.mem_2595_sv2v_reg ;
  assign \nz.mem [2594] = \nz.mem_2594_sv2v_reg ;
  assign \nz.mem [2593] = \nz.mem_2593_sv2v_reg ;
  assign \nz.mem [2592] = \nz.mem_2592_sv2v_reg ;
  assign \nz.mem [2591] = \nz.mem_2591_sv2v_reg ;
  assign \nz.mem [2590] = \nz.mem_2590_sv2v_reg ;
  assign \nz.mem [2589] = \nz.mem_2589_sv2v_reg ;
  assign \nz.mem [2588] = \nz.mem_2588_sv2v_reg ;
  assign \nz.mem [2587] = \nz.mem_2587_sv2v_reg ;
  assign \nz.mem [2586] = \nz.mem_2586_sv2v_reg ;
  assign \nz.mem [2585] = \nz.mem_2585_sv2v_reg ;
  assign \nz.mem [2584] = \nz.mem_2584_sv2v_reg ;
  assign \nz.mem [2583] = \nz.mem_2583_sv2v_reg ;
  assign \nz.mem [2582] = \nz.mem_2582_sv2v_reg ;
  assign \nz.mem [2581] = \nz.mem_2581_sv2v_reg ;
  assign \nz.mem [2580] = \nz.mem_2580_sv2v_reg ;
  assign \nz.mem [2579] = \nz.mem_2579_sv2v_reg ;
  assign \nz.mem [2578] = \nz.mem_2578_sv2v_reg ;
  assign \nz.mem [2577] = \nz.mem_2577_sv2v_reg ;
  assign \nz.mem [2576] = \nz.mem_2576_sv2v_reg ;
  assign \nz.mem [2575] = \nz.mem_2575_sv2v_reg ;
  assign \nz.mem [2574] = \nz.mem_2574_sv2v_reg ;
  assign \nz.mem [2573] = \nz.mem_2573_sv2v_reg ;
  assign \nz.mem [2572] = \nz.mem_2572_sv2v_reg ;
  assign \nz.mem [2571] = \nz.mem_2571_sv2v_reg ;
  assign \nz.mem [2570] = \nz.mem_2570_sv2v_reg ;
  assign \nz.mem [2569] = \nz.mem_2569_sv2v_reg ;
  assign \nz.mem [2568] = \nz.mem_2568_sv2v_reg ;
  assign \nz.mem [2567] = \nz.mem_2567_sv2v_reg ;
  assign \nz.mem [2566] = \nz.mem_2566_sv2v_reg ;
  assign \nz.mem [2565] = \nz.mem_2565_sv2v_reg ;
  assign \nz.mem [2564] = \nz.mem_2564_sv2v_reg ;
  assign \nz.mem [2563] = \nz.mem_2563_sv2v_reg ;
  assign \nz.mem [2562] = \nz.mem_2562_sv2v_reg ;
  assign \nz.mem [2561] = \nz.mem_2561_sv2v_reg ;
  assign \nz.mem [2560] = \nz.mem_2560_sv2v_reg ;
  assign \nz.mem [2559] = \nz.mem_2559_sv2v_reg ;
  assign \nz.mem [2558] = \nz.mem_2558_sv2v_reg ;
  assign \nz.mem [2557] = \nz.mem_2557_sv2v_reg ;
  assign \nz.mem [2556] = \nz.mem_2556_sv2v_reg ;
  assign \nz.mem [2555] = \nz.mem_2555_sv2v_reg ;
  assign \nz.mem [2554] = \nz.mem_2554_sv2v_reg ;
  assign \nz.mem [2553] = \nz.mem_2553_sv2v_reg ;
  assign \nz.mem [2552] = \nz.mem_2552_sv2v_reg ;
  assign \nz.mem [2551] = \nz.mem_2551_sv2v_reg ;
  assign \nz.mem [2550] = \nz.mem_2550_sv2v_reg ;
  assign \nz.mem [2549] = \nz.mem_2549_sv2v_reg ;
  assign \nz.mem [2548] = \nz.mem_2548_sv2v_reg ;
  assign \nz.mem [2547] = \nz.mem_2547_sv2v_reg ;
  assign \nz.mem [2546] = \nz.mem_2546_sv2v_reg ;
  assign \nz.mem [2545] = \nz.mem_2545_sv2v_reg ;
  assign \nz.mem [2544] = \nz.mem_2544_sv2v_reg ;
  assign \nz.mem [2543] = \nz.mem_2543_sv2v_reg ;
  assign \nz.mem [2542] = \nz.mem_2542_sv2v_reg ;
  assign \nz.mem [2541] = \nz.mem_2541_sv2v_reg ;
  assign \nz.mem [2540] = \nz.mem_2540_sv2v_reg ;
  assign \nz.mem [2539] = \nz.mem_2539_sv2v_reg ;
  assign \nz.mem [2538] = \nz.mem_2538_sv2v_reg ;
  assign \nz.mem [2537] = \nz.mem_2537_sv2v_reg ;
  assign \nz.mem [2536] = \nz.mem_2536_sv2v_reg ;
  assign \nz.mem [2535] = \nz.mem_2535_sv2v_reg ;
  assign \nz.mem [2534] = \nz.mem_2534_sv2v_reg ;
  assign \nz.mem [2533] = \nz.mem_2533_sv2v_reg ;
  assign \nz.mem [2532] = \nz.mem_2532_sv2v_reg ;
  assign \nz.mem [2531] = \nz.mem_2531_sv2v_reg ;
  assign \nz.mem [2530] = \nz.mem_2530_sv2v_reg ;
  assign \nz.mem [2529] = \nz.mem_2529_sv2v_reg ;
  assign \nz.mem [2528] = \nz.mem_2528_sv2v_reg ;
  assign \nz.mem [2527] = \nz.mem_2527_sv2v_reg ;
  assign \nz.mem [2526] = \nz.mem_2526_sv2v_reg ;
  assign \nz.mem [2525] = \nz.mem_2525_sv2v_reg ;
  assign \nz.mem [2524] = \nz.mem_2524_sv2v_reg ;
  assign \nz.mem [2523] = \nz.mem_2523_sv2v_reg ;
  assign \nz.mem [2522] = \nz.mem_2522_sv2v_reg ;
  assign \nz.mem [2521] = \nz.mem_2521_sv2v_reg ;
  assign \nz.mem [2520] = \nz.mem_2520_sv2v_reg ;
  assign \nz.mem [2519] = \nz.mem_2519_sv2v_reg ;
  assign \nz.mem [2518] = \nz.mem_2518_sv2v_reg ;
  assign \nz.mem [2517] = \nz.mem_2517_sv2v_reg ;
  assign \nz.mem [2516] = \nz.mem_2516_sv2v_reg ;
  assign \nz.mem [2515] = \nz.mem_2515_sv2v_reg ;
  assign \nz.mem [2514] = \nz.mem_2514_sv2v_reg ;
  assign \nz.mem [2513] = \nz.mem_2513_sv2v_reg ;
  assign \nz.mem [2512] = \nz.mem_2512_sv2v_reg ;
  assign \nz.mem [2511] = \nz.mem_2511_sv2v_reg ;
  assign \nz.mem [2510] = \nz.mem_2510_sv2v_reg ;
  assign \nz.mem [2509] = \nz.mem_2509_sv2v_reg ;
  assign \nz.mem [2508] = \nz.mem_2508_sv2v_reg ;
  assign \nz.mem [2507] = \nz.mem_2507_sv2v_reg ;
  assign \nz.mem [2506] = \nz.mem_2506_sv2v_reg ;
  assign \nz.mem [2505] = \nz.mem_2505_sv2v_reg ;
  assign \nz.mem [2504] = \nz.mem_2504_sv2v_reg ;
  assign \nz.mem [2503] = \nz.mem_2503_sv2v_reg ;
  assign \nz.mem [2502] = \nz.mem_2502_sv2v_reg ;
  assign \nz.mem [2501] = \nz.mem_2501_sv2v_reg ;
  assign \nz.mem [2500] = \nz.mem_2500_sv2v_reg ;
  assign \nz.mem [2499] = \nz.mem_2499_sv2v_reg ;
  assign \nz.mem [2498] = \nz.mem_2498_sv2v_reg ;
  assign \nz.mem [2497] = \nz.mem_2497_sv2v_reg ;
  assign \nz.mem [2496] = \nz.mem_2496_sv2v_reg ;
  assign \nz.mem [2495] = \nz.mem_2495_sv2v_reg ;
  assign \nz.mem [2494] = \nz.mem_2494_sv2v_reg ;
  assign \nz.mem [2493] = \nz.mem_2493_sv2v_reg ;
  assign \nz.mem [2492] = \nz.mem_2492_sv2v_reg ;
  assign \nz.mem [2491] = \nz.mem_2491_sv2v_reg ;
  assign \nz.mem [2490] = \nz.mem_2490_sv2v_reg ;
  assign \nz.mem [2489] = \nz.mem_2489_sv2v_reg ;
  assign \nz.mem [2488] = \nz.mem_2488_sv2v_reg ;
  assign \nz.mem [2487] = \nz.mem_2487_sv2v_reg ;
  assign \nz.mem [2486] = \nz.mem_2486_sv2v_reg ;
  assign \nz.mem [2485] = \nz.mem_2485_sv2v_reg ;
  assign \nz.mem [2484] = \nz.mem_2484_sv2v_reg ;
  assign \nz.mem [2483] = \nz.mem_2483_sv2v_reg ;
  assign \nz.mem [2482] = \nz.mem_2482_sv2v_reg ;
  assign \nz.mem [2481] = \nz.mem_2481_sv2v_reg ;
  assign \nz.mem [2480] = \nz.mem_2480_sv2v_reg ;
  assign \nz.mem [2479] = \nz.mem_2479_sv2v_reg ;
  assign \nz.mem [2478] = \nz.mem_2478_sv2v_reg ;
  assign \nz.mem [2477] = \nz.mem_2477_sv2v_reg ;
  assign \nz.mem [2476] = \nz.mem_2476_sv2v_reg ;
  assign \nz.mem [2475] = \nz.mem_2475_sv2v_reg ;
  assign \nz.mem [2474] = \nz.mem_2474_sv2v_reg ;
  assign \nz.mem [2473] = \nz.mem_2473_sv2v_reg ;
  assign \nz.mem [2472] = \nz.mem_2472_sv2v_reg ;
  assign \nz.mem [2471] = \nz.mem_2471_sv2v_reg ;
  assign \nz.mem [2470] = \nz.mem_2470_sv2v_reg ;
  assign \nz.mem [2469] = \nz.mem_2469_sv2v_reg ;
  assign \nz.mem [2468] = \nz.mem_2468_sv2v_reg ;
  assign \nz.mem [2467] = \nz.mem_2467_sv2v_reg ;
  assign \nz.mem [2466] = \nz.mem_2466_sv2v_reg ;
  assign \nz.mem [2465] = \nz.mem_2465_sv2v_reg ;
  assign \nz.mem [2464] = \nz.mem_2464_sv2v_reg ;
  assign \nz.mem [2463] = \nz.mem_2463_sv2v_reg ;
  assign \nz.mem [2462] = \nz.mem_2462_sv2v_reg ;
  assign \nz.mem [2461] = \nz.mem_2461_sv2v_reg ;
  assign \nz.mem [2460] = \nz.mem_2460_sv2v_reg ;
  assign \nz.mem [2459] = \nz.mem_2459_sv2v_reg ;
  assign \nz.mem [2458] = \nz.mem_2458_sv2v_reg ;
  assign \nz.mem [2457] = \nz.mem_2457_sv2v_reg ;
  assign \nz.mem [2456] = \nz.mem_2456_sv2v_reg ;
  assign \nz.mem [2455] = \nz.mem_2455_sv2v_reg ;
  assign \nz.mem [2454] = \nz.mem_2454_sv2v_reg ;
  assign \nz.mem [2453] = \nz.mem_2453_sv2v_reg ;
  assign \nz.mem [2452] = \nz.mem_2452_sv2v_reg ;
  assign \nz.mem [2451] = \nz.mem_2451_sv2v_reg ;
  assign \nz.mem [2450] = \nz.mem_2450_sv2v_reg ;
  assign \nz.mem [2449] = \nz.mem_2449_sv2v_reg ;
  assign \nz.mem [2448] = \nz.mem_2448_sv2v_reg ;
  assign \nz.mem [2447] = \nz.mem_2447_sv2v_reg ;
  assign \nz.mem [2446] = \nz.mem_2446_sv2v_reg ;
  assign \nz.mem [2445] = \nz.mem_2445_sv2v_reg ;
  assign \nz.mem [2444] = \nz.mem_2444_sv2v_reg ;
  assign \nz.mem [2443] = \nz.mem_2443_sv2v_reg ;
  assign \nz.mem [2442] = \nz.mem_2442_sv2v_reg ;
  assign \nz.mem [2441] = \nz.mem_2441_sv2v_reg ;
  assign \nz.mem [2440] = \nz.mem_2440_sv2v_reg ;
  assign \nz.mem [2439] = \nz.mem_2439_sv2v_reg ;
  assign \nz.mem [2438] = \nz.mem_2438_sv2v_reg ;
  assign \nz.mem [2437] = \nz.mem_2437_sv2v_reg ;
  assign \nz.mem [2436] = \nz.mem_2436_sv2v_reg ;
  assign \nz.mem [2435] = \nz.mem_2435_sv2v_reg ;
  assign \nz.mem [2434] = \nz.mem_2434_sv2v_reg ;
  assign \nz.mem [2433] = \nz.mem_2433_sv2v_reg ;
  assign \nz.mem [2432] = \nz.mem_2432_sv2v_reg ;
  assign \nz.mem [2431] = \nz.mem_2431_sv2v_reg ;
  assign \nz.mem [2430] = \nz.mem_2430_sv2v_reg ;
  assign \nz.mem [2429] = \nz.mem_2429_sv2v_reg ;
  assign \nz.mem [2428] = \nz.mem_2428_sv2v_reg ;
  assign \nz.mem [2427] = \nz.mem_2427_sv2v_reg ;
  assign \nz.mem [2426] = \nz.mem_2426_sv2v_reg ;
  assign \nz.mem [2425] = \nz.mem_2425_sv2v_reg ;
  assign \nz.mem [2424] = \nz.mem_2424_sv2v_reg ;
  assign \nz.mem [2423] = \nz.mem_2423_sv2v_reg ;
  assign \nz.mem [2422] = \nz.mem_2422_sv2v_reg ;
  assign \nz.mem [2421] = \nz.mem_2421_sv2v_reg ;
  assign \nz.mem [2420] = \nz.mem_2420_sv2v_reg ;
  assign \nz.mem [2419] = \nz.mem_2419_sv2v_reg ;
  assign \nz.mem [2418] = \nz.mem_2418_sv2v_reg ;
  assign \nz.mem [2417] = \nz.mem_2417_sv2v_reg ;
  assign \nz.mem [2416] = \nz.mem_2416_sv2v_reg ;
  assign \nz.mem [2415] = \nz.mem_2415_sv2v_reg ;
  assign \nz.mem [2414] = \nz.mem_2414_sv2v_reg ;
  assign \nz.mem [2413] = \nz.mem_2413_sv2v_reg ;
  assign \nz.mem [2412] = \nz.mem_2412_sv2v_reg ;
  assign \nz.mem [2411] = \nz.mem_2411_sv2v_reg ;
  assign \nz.mem [2410] = \nz.mem_2410_sv2v_reg ;
  assign \nz.mem [2409] = \nz.mem_2409_sv2v_reg ;
  assign \nz.mem [2408] = \nz.mem_2408_sv2v_reg ;
  assign \nz.mem [2407] = \nz.mem_2407_sv2v_reg ;
  assign \nz.mem [2406] = \nz.mem_2406_sv2v_reg ;
  assign \nz.mem [2405] = \nz.mem_2405_sv2v_reg ;
  assign \nz.mem [2404] = \nz.mem_2404_sv2v_reg ;
  assign \nz.mem [2403] = \nz.mem_2403_sv2v_reg ;
  assign \nz.mem [2402] = \nz.mem_2402_sv2v_reg ;
  assign \nz.mem [2401] = \nz.mem_2401_sv2v_reg ;
  assign \nz.mem [2400] = \nz.mem_2400_sv2v_reg ;
  assign \nz.mem [2399] = \nz.mem_2399_sv2v_reg ;
  assign \nz.mem [2398] = \nz.mem_2398_sv2v_reg ;
  assign \nz.mem [2397] = \nz.mem_2397_sv2v_reg ;
  assign \nz.mem [2396] = \nz.mem_2396_sv2v_reg ;
  assign \nz.mem [2395] = \nz.mem_2395_sv2v_reg ;
  assign \nz.mem [2394] = \nz.mem_2394_sv2v_reg ;
  assign \nz.mem [2393] = \nz.mem_2393_sv2v_reg ;
  assign \nz.mem [2392] = \nz.mem_2392_sv2v_reg ;
  assign \nz.mem [2391] = \nz.mem_2391_sv2v_reg ;
  assign \nz.mem [2390] = \nz.mem_2390_sv2v_reg ;
  assign \nz.mem [2389] = \nz.mem_2389_sv2v_reg ;
  assign \nz.mem [2388] = \nz.mem_2388_sv2v_reg ;
  assign \nz.mem [2387] = \nz.mem_2387_sv2v_reg ;
  assign \nz.mem [2386] = \nz.mem_2386_sv2v_reg ;
  assign \nz.mem [2385] = \nz.mem_2385_sv2v_reg ;
  assign \nz.mem [2384] = \nz.mem_2384_sv2v_reg ;
  assign \nz.mem [2383] = \nz.mem_2383_sv2v_reg ;
  assign \nz.mem [2382] = \nz.mem_2382_sv2v_reg ;
  assign \nz.mem [2381] = \nz.mem_2381_sv2v_reg ;
  assign \nz.mem [2380] = \nz.mem_2380_sv2v_reg ;
  assign \nz.mem [2379] = \nz.mem_2379_sv2v_reg ;
  assign \nz.mem [2378] = \nz.mem_2378_sv2v_reg ;
  assign \nz.mem [2377] = \nz.mem_2377_sv2v_reg ;
  assign \nz.mem [2376] = \nz.mem_2376_sv2v_reg ;
  assign \nz.mem [2375] = \nz.mem_2375_sv2v_reg ;
  assign \nz.mem [2374] = \nz.mem_2374_sv2v_reg ;
  assign \nz.mem [2373] = \nz.mem_2373_sv2v_reg ;
  assign \nz.mem [2372] = \nz.mem_2372_sv2v_reg ;
  assign \nz.mem [2371] = \nz.mem_2371_sv2v_reg ;
  assign \nz.mem [2370] = \nz.mem_2370_sv2v_reg ;
  assign \nz.mem [2369] = \nz.mem_2369_sv2v_reg ;
  assign \nz.mem [2368] = \nz.mem_2368_sv2v_reg ;
  assign \nz.mem [2367] = \nz.mem_2367_sv2v_reg ;
  assign \nz.mem [2366] = \nz.mem_2366_sv2v_reg ;
  assign \nz.mem [2365] = \nz.mem_2365_sv2v_reg ;
  assign \nz.mem [2364] = \nz.mem_2364_sv2v_reg ;
  assign \nz.mem [2363] = \nz.mem_2363_sv2v_reg ;
  assign \nz.mem [2362] = \nz.mem_2362_sv2v_reg ;
  assign \nz.mem [2361] = \nz.mem_2361_sv2v_reg ;
  assign \nz.mem [2360] = \nz.mem_2360_sv2v_reg ;
  assign \nz.mem [2359] = \nz.mem_2359_sv2v_reg ;
  assign \nz.mem [2358] = \nz.mem_2358_sv2v_reg ;
  assign \nz.mem [2357] = \nz.mem_2357_sv2v_reg ;
  assign \nz.mem [2356] = \nz.mem_2356_sv2v_reg ;
  assign \nz.mem [2355] = \nz.mem_2355_sv2v_reg ;
  assign \nz.mem [2354] = \nz.mem_2354_sv2v_reg ;
  assign \nz.mem [2353] = \nz.mem_2353_sv2v_reg ;
  assign \nz.mem [2352] = \nz.mem_2352_sv2v_reg ;
  assign \nz.mem [2351] = \nz.mem_2351_sv2v_reg ;
  assign \nz.mem [2350] = \nz.mem_2350_sv2v_reg ;
  assign \nz.mem [2349] = \nz.mem_2349_sv2v_reg ;
  assign \nz.mem [2348] = \nz.mem_2348_sv2v_reg ;
  assign \nz.mem [2347] = \nz.mem_2347_sv2v_reg ;
  assign \nz.mem [2346] = \nz.mem_2346_sv2v_reg ;
  assign \nz.mem [2345] = \nz.mem_2345_sv2v_reg ;
  assign \nz.mem [2344] = \nz.mem_2344_sv2v_reg ;
  assign \nz.mem [2343] = \nz.mem_2343_sv2v_reg ;
  assign \nz.mem [2342] = \nz.mem_2342_sv2v_reg ;
  assign \nz.mem [2341] = \nz.mem_2341_sv2v_reg ;
  assign \nz.mem [2340] = \nz.mem_2340_sv2v_reg ;
  assign \nz.mem [2339] = \nz.mem_2339_sv2v_reg ;
  assign \nz.mem [2338] = \nz.mem_2338_sv2v_reg ;
  assign \nz.mem [2337] = \nz.mem_2337_sv2v_reg ;
  assign \nz.mem [2336] = \nz.mem_2336_sv2v_reg ;
  assign \nz.mem [2335] = \nz.mem_2335_sv2v_reg ;
  assign \nz.mem [2334] = \nz.mem_2334_sv2v_reg ;
  assign \nz.mem [2333] = \nz.mem_2333_sv2v_reg ;
  assign \nz.mem [2332] = \nz.mem_2332_sv2v_reg ;
  assign \nz.mem [2331] = \nz.mem_2331_sv2v_reg ;
  assign \nz.mem [2330] = \nz.mem_2330_sv2v_reg ;
  assign \nz.mem [2329] = \nz.mem_2329_sv2v_reg ;
  assign \nz.mem [2328] = \nz.mem_2328_sv2v_reg ;
  assign \nz.mem [2327] = \nz.mem_2327_sv2v_reg ;
  assign \nz.mem [2326] = \nz.mem_2326_sv2v_reg ;
  assign \nz.mem [2325] = \nz.mem_2325_sv2v_reg ;
  assign \nz.mem [2324] = \nz.mem_2324_sv2v_reg ;
  assign \nz.mem [2323] = \nz.mem_2323_sv2v_reg ;
  assign \nz.mem [2322] = \nz.mem_2322_sv2v_reg ;
  assign \nz.mem [2321] = \nz.mem_2321_sv2v_reg ;
  assign \nz.mem [2320] = \nz.mem_2320_sv2v_reg ;
  assign \nz.mem [2319] = \nz.mem_2319_sv2v_reg ;
  assign \nz.mem [2318] = \nz.mem_2318_sv2v_reg ;
  assign \nz.mem [2317] = \nz.mem_2317_sv2v_reg ;
  assign \nz.mem [2316] = \nz.mem_2316_sv2v_reg ;
  assign \nz.mem [2315] = \nz.mem_2315_sv2v_reg ;
  assign \nz.mem [2314] = \nz.mem_2314_sv2v_reg ;
  assign \nz.mem [2313] = \nz.mem_2313_sv2v_reg ;
  assign \nz.mem [2312] = \nz.mem_2312_sv2v_reg ;
  assign \nz.mem [2311] = \nz.mem_2311_sv2v_reg ;
  assign \nz.mem [2310] = \nz.mem_2310_sv2v_reg ;
  assign \nz.mem [2309] = \nz.mem_2309_sv2v_reg ;
  assign \nz.mem [2308] = \nz.mem_2308_sv2v_reg ;
  assign \nz.mem [2307] = \nz.mem_2307_sv2v_reg ;
  assign \nz.mem [2306] = \nz.mem_2306_sv2v_reg ;
  assign \nz.mem [2305] = \nz.mem_2305_sv2v_reg ;
  assign \nz.mem [2304] = \nz.mem_2304_sv2v_reg ;
  assign \nz.mem [2303] = \nz.mem_2303_sv2v_reg ;
  assign \nz.mem [2302] = \nz.mem_2302_sv2v_reg ;
  assign \nz.mem [2301] = \nz.mem_2301_sv2v_reg ;
  assign \nz.mem [2300] = \nz.mem_2300_sv2v_reg ;
  assign \nz.mem [2299] = \nz.mem_2299_sv2v_reg ;
  assign \nz.mem [2298] = \nz.mem_2298_sv2v_reg ;
  assign \nz.mem [2297] = \nz.mem_2297_sv2v_reg ;
  assign \nz.mem [2296] = \nz.mem_2296_sv2v_reg ;
  assign \nz.mem [2295] = \nz.mem_2295_sv2v_reg ;
  assign \nz.mem [2294] = \nz.mem_2294_sv2v_reg ;
  assign \nz.mem [2293] = \nz.mem_2293_sv2v_reg ;
  assign \nz.mem [2292] = \nz.mem_2292_sv2v_reg ;
  assign \nz.mem [2291] = \nz.mem_2291_sv2v_reg ;
  assign \nz.mem [2290] = \nz.mem_2290_sv2v_reg ;
  assign \nz.mem [2289] = \nz.mem_2289_sv2v_reg ;
  assign \nz.mem [2288] = \nz.mem_2288_sv2v_reg ;
  assign \nz.mem [2287] = \nz.mem_2287_sv2v_reg ;
  assign \nz.mem [2286] = \nz.mem_2286_sv2v_reg ;
  assign \nz.mem [2285] = \nz.mem_2285_sv2v_reg ;
  assign \nz.mem [2284] = \nz.mem_2284_sv2v_reg ;
  assign \nz.mem [2283] = \nz.mem_2283_sv2v_reg ;
  assign \nz.mem [2282] = \nz.mem_2282_sv2v_reg ;
  assign \nz.mem [2281] = \nz.mem_2281_sv2v_reg ;
  assign \nz.mem [2280] = \nz.mem_2280_sv2v_reg ;
  assign \nz.mem [2279] = \nz.mem_2279_sv2v_reg ;
  assign \nz.mem [2278] = \nz.mem_2278_sv2v_reg ;
  assign \nz.mem [2277] = \nz.mem_2277_sv2v_reg ;
  assign \nz.mem [2276] = \nz.mem_2276_sv2v_reg ;
  assign \nz.mem [2275] = \nz.mem_2275_sv2v_reg ;
  assign \nz.mem [2274] = \nz.mem_2274_sv2v_reg ;
  assign \nz.mem [2273] = \nz.mem_2273_sv2v_reg ;
  assign \nz.mem [2272] = \nz.mem_2272_sv2v_reg ;
  assign \nz.mem [2271] = \nz.mem_2271_sv2v_reg ;
  assign \nz.mem [2270] = \nz.mem_2270_sv2v_reg ;
  assign \nz.mem [2269] = \nz.mem_2269_sv2v_reg ;
  assign \nz.mem [2268] = \nz.mem_2268_sv2v_reg ;
  assign \nz.mem [2267] = \nz.mem_2267_sv2v_reg ;
  assign \nz.mem [2266] = \nz.mem_2266_sv2v_reg ;
  assign \nz.mem [2265] = \nz.mem_2265_sv2v_reg ;
  assign \nz.mem [2264] = \nz.mem_2264_sv2v_reg ;
  assign \nz.mem [2263] = \nz.mem_2263_sv2v_reg ;
  assign \nz.mem [2262] = \nz.mem_2262_sv2v_reg ;
  assign \nz.mem [2261] = \nz.mem_2261_sv2v_reg ;
  assign \nz.mem [2260] = \nz.mem_2260_sv2v_reg ;
  assign \nz.mem [2259] = \nz.mem_2259_sv2v_reg ;
  assign \nz.mem [2258] = \nz.mem_2258_sv2v_reg ;
  assign \nz.mem [2257] = \nz.mem_2257_sv2v_reg ;
  assign \nz.mem [2256] = \nz.mem_2256_sv2v_reg ;
  assign \nz.mem [2255] = \nz.mem_2255_sv2v_reg ;
  assign \nz.mem [2254] = \nz.mem_2254_sv2v_reg ;
  assign \nz.mem [2253] = \nz.mem_2253_sv2v_reg ;
  assign \nz.mem [2252] = \nz.mem_2252_sv2v_reg ;
  assign \nz.mem [2251] = \nz.mem_2251_sv2v_reg ;
  assign \nz.mem [2250] = \nz.mem_2250_sv2v_reg ;
  assign \nz.mem [2249] = \nz.mem_2249_sv2v_reg ;
  assign \nz.mem [2248] = \nz.mem_2248_sv2v_reg ;
  assign \nz.mem [2247] = \nz.mem_2247_sv2v_reg ;
  assign \nz.mem [2246] = \nz.mem_2246_sv2v_reg ;
  assign \nz.mem [2245] = \nz.mem_2245_sv2v_reg ;
  assign \nz.mem [2244] = \nz.mem_2244_sv2v_reg ;
  assign \nz.mem [2243] = \nz.mem_2243_sv2v_reg ;
  assign \nz.mem [2242] = \nz.mem_2242_sv2v_reg ;
  assign \nz.mem [2241] = \nz.mem_2241_sv2v_reg ;
  assign \nz.mem [2240] = \nz.mem_2240_sv2v_reg ;
  assign \nz.mem [2239] = \nz.mem_2239_sv2v_reg ;
  assign \nz.mem [2238] = \nz.mem_2238_sv2v_reg ;
  assign \nz.mem [2237] = \nz.mem_2237_sv2v_reg ;
  assign \nz.mem [2236] = \nz.mem_2236_sv2v_reg ;
  assign \nz.mem [2235] = \nz.mem_2235_sv2v_reg ;
  assign \nz.mem [2234] = \nz.mem_2234_sv2v_reg ;
  assign \nz.mem [2233] = \nz.mem_2233_sv2v_reg ;
  assign \nz.mem [2232] = \nz.mem_2232_sv2v_reg ;
  assign \nz.mem [2231] = \nz.mem_2231_sv2v_reg ;
  assign \nz.mem [2230] = \nz.mem_2230_sv2v_reg ;
  assign \nz.mem [2229] = \nz.mem_2229_sv2v_reg ;
  assign \nz.mem [2228] = \nz.mem_2228_sv2v_reg ;
  assign \nz.mem [2227] = \nz.mem_2227_sv2v_reg ;
  assign \nz.mem [2226] = \nz.mem_2226_sv2v_reg ;
  assign \nz.mem [2225] = \nz.mem_2225_sv2v_reg ;
  assign \nz.mem [2224] = \nz.mem_2224_sv2v_reg ;
  assign \nz.mem [2223] = \nz.mem_2223_sv2v_reg ;
  assign \nz.mem [2222] = \nz.mem_2222_sv2v_reg ;
  assign \nz.mem [2221] = \nz.mem_2221_sv2v_reg ;
  assign \nz.mem [2220] = \nz.mem_2220_sv2v_reg ;
  assign \nz.mem [2219] = \nz.mem_2219_sv2v_reg ;
  assign \nz.mem [2218] = \nz.mem_2218_sv2v_reg ;
  assign \nz.mem [2217] = \nz.mem_2217_sv2v_reg ;
  assign \nz.mem [2216] = \nz.mem_2216_sv2v_reg ;
  assign \nz.mem [2215] = \nz.mem_2215_sv2v_reg ;
  assign \nz.mem [2214] = \nz.mem_2214_sv2v_reg ;
  assign \nz.mem [2213] = \nz.mem_2213_sv2v_reg ;
  assign \nz.mem [2212] = \nz.mem_2212_sv2v_reg ;
  assign \nz.mem [2211] = \nz.mem_2211_sv2v_reg ;
  assign \nz.mem [2210] = \nz.mem_2210_sv2v_reg ;
  assign \nz.mem [2209] = \nz.mem_2209_sv2v_reg ;
  assign \nz.mem [2208] = \nz.mem_2208_sv2v_reg ;
  assign \nz.mem [2207] = \nz.mem_2207_sv2v_reg ;
  assign \nz.mem [2206] = \nz.mem_2206_sv2v_reg ;
  assign \nz.mem [2205] = \nz.mem_2205_sv2v_reg ;
  assign \nz.mem [2204] = \nz.mem_2204_sv2v_reg ;
  assign \nz.mem [2203] = \nz.mem_2203_sv2v_reg ;
  assign \nz.mem [2202] = \nz.mem_2202_sv2v_reg ;
  assign \nz.mem [2201] = \nz.mem_2201_sv2v_reg ;
  assign \nz.mem [2200] = \nz.mem_2200_sv2v_reg ;
  assign \nz.mem [2199] = \nz.mem_2199_sv2v_reg ;
  assign \nz.mem [2198] = \nz.mem_2198_sv2v_reg ;
  assign \nz.mem [2197] = \nz.mem_2197_sv2v_reg ;
  assign \nz.mem [2196] = \nz.mem_2196_sv2v_reg ;
  assign \nz.mem [2195] = \nz.mem_2195_sv2v_reg ;
  assign \nz.mem [2194] = \nz.mem_2194_sv2v_reg ;
  assign \nz.mem [2193] = \nz.mem_2193_sv2v_reg ;
  assign \nz.mem [2192] = \nz.mem_2192_sv2v_reg ;
  assign \nz.mem [2191] = \nz.mem_2191_sv2v_reg ;
  assign \nz.mem [2190] = \nz.mem_2190_sv2v_reg ;
  assign \nz.mem [2189] = \nz.mem_2189_sv2v_reg ;
  assign \nz.mem [2188] = \nz.mem_2188_sv2v_reg ;
  assign \nz.mem [2187] = \nz.mem_2187_sv2v_reg ;
  assign \nz.mem [2186] = \nz.mem_2186_sv2v_reg ;
  assign \nz.mem [2185] = \nz.mem_2185_sv2v_reg ;
  assign \nz.mem [2184] = \nz.mem_2184_sv2v_reg ;
  assign \nz.mem [2183] = \nz.mem_2183_sv2v_reg ;
  assign \nz.mem [2182] = \nz.mem_2182_sv2v_reg ;
  assign \nz.mem [2181] = \nz.mem_2181_sv2v_reg ;
  assign \nz.mem [2180] = \nz.mem_2180_sv2v_reg ;
  assign \nz.mem [2179] = \nz.mem_2179_sv2v_reg ;
  assign \nz.mem [2178] = \nz.mem_2178_sv2v_reg ;
  assign \nz.mem [2177] = \nz.mem_2177_sv2v_reg ;
  assign \nz.mem [2176] = \nz.mem_2176_sv2v_reg ;
  assign \nz.mem [2175] = \nz.mem_2175_sv2v_reg ;
  assign \nz.mem [2174] = \nz.mem_2174_sv2v_reg ;
  assign \nz.mem [2173] = \nz.mem_2173_sv2v_reg ;
  assign \nz.mem [2172] = \nz.mem_2172_sv2v_reg ;
  assign \nz.mem [2171] = \nz.mem_2171_sv2v_reg ;
  assign \nz.mem [2170] = \nz.mem_2170_sv2v_reg ;
  assign \nz.mem [2169] = \nz.mem_2169_sv2v_reg ;
  assign \nz.mem [2168] = \nz.mem_2168_sv2v_reg ;
  assign \nz.mem [2167] = \nz.mem_2167_sv2v_reg ;
  assign \nz.mem [2166] = \nz.mem_2166_sv2v_reg ;
  assign \nz.mem [2165] = \nz.mem_2165_sv2v_reg ;
  assign \nz.mem [2164] = \nz.mem_2164_sv2v_reg ;
  assign \nz.mem [2163] = \nz.mem_2163_sv2v_reg ;
  assign \nz.mem [2162] = \nz.mem_2162_sv2v_reg ;
  assign \nz.mem [2161] = \nz.mem_2161_sv2v_reg ;
  assign \nz.mem [2160] = \nz.mem_2160_sv2v_reg ;
  assign \nz.mem [2159] = \nz.mem_2159_sv2v_reg ;
  assign \nz.mem [2158] = \nz.mem_2158_sv2v_reg ;
  assign \nz.mem [2157] = \nz.mem_2157_sv2v_reg ;
  assign \nz.mem [2156] = \nz.mem_2156_sv2v_reg ;
  assign \nz.mem [2155] = \nz.mem_2155_sv2v_reg ;
  assign \nz.mem [2154] = \nz.mem_2154_sv2v_reg ;
  assign \nz.mem [2153] = \nz.mem_2153_sv2v_reg ;
  assign \nz.mem [2152] = \nz.mem_2152_sv2v_reg ;
  assign \nz.mem [2151] = \nz.mem_2151_sv2v_reg ;
  assign \nz.mem [2150] = \nz.mem_2150_sv2v_reg ;
  assign \nz.mem [2149] = \nz.mem_2149_sv2v_reg ;
  assign \nz.mem [2148] = \nz.mem_2148_sv2v_reg ;
  assign \nz.mem [2147] = \nz.mem_2147_sv2v_reg ;
  assign \nz.mem [2146] = \nz.mem_2146_sv2v_reg ;
  assign \nz.mem [2145] = \nz.mem_2145_sv2v_reg ;
  assign \nz.mem [2144] = \nz.mem_2144_sv2v_reg ;
  assign \nz.mem [2143] = \nz.mem_2143_sv2v_reg ;
  assign \nz.mem [2142] = \nz.mem_2142_sv2v_reg ;
  assign \nz.mem [2141] = \nz.mem_2141_sv2v_reg ;
  assign \nz.mem [2140] = \nz.mem_2140_sv2v_reg ;
  assign \nz.mem [2139] = \nz.mem_2139_sv2v_reg ;
  assign \nz.mem [2138] = \nz.mem_2138_sv2v_reg ;
  assign \nz.mem [2137] = \nz.mem_2137_sv2v_reg ;
  assign \nz.mem [2136] = \nz.mem_2136_sv2v_reg ;
  assign \nz.mem [2135] = \nz.mem_2135_sv2v_reg ;
  assign \nz.mem [2134] = \nz.mem_2134_sv2v_reg ;
  assign \nz.mem [2133] = \nz.mem_2133_sv2v_reg ;
  assign \nz.mem [2132] = \nz.mem_2132_sv2v_reg ;
  assign \nz.mem [2131] = \nz.mem_2131_sv2v_reg ;
  assign \nz.mem [2130] = \nz.mem_2130_sv2v_reg ;
  assign \nz.mem [2129] = \nz.mem_2129_sv2v_reg ;
  assign \nz.mem [2128] = \nz.mem_2128_sv2v_reg ;
  assign \nz.mem [2127] = \nz.mem_2127_sv2v_reg ;
  assign \nz.mem [2126] = \nz.mem_2126_sv2v_reg ;
  assign \nz.mem [2125] = \nz.mem_2125_sv2v_reg ;
  assign \nz.mem [2124] = \nz.mem_2124_sv2v_reg ;
  assign \nz.mem [2123] = \nz.mem_2123_sv2v_reg ;
  assign \nz.mem [2122] = \nz.mem_2122_sv2v_reg ;
  assign \nz.mem [2121] = \nz.mem_2121_sv2v_reg ;
  assign \nz.mem [2120] = \nz.mem_2120_sv2v_reg ;
  assign \nz.mem [2119] = \nz.mem_2119_sv2v_reg ;
  assign \nz.mem [2118] = \nz.mem_2118_sv2v_reg ;
  assign \nz.mem [2117] = \nz.mem_2117_sv2v_reg ;
  assign \nz.mem [2116] = \nz.mem_2116_sv2v_reg ;
  assign \nz.mem [2115] = \nz.mem_2115_sv2v_reg ;
  assign \nz.mem [2114] = \nz.mem_2114_sv2v_reg ;
  assign \nz.mem [2113] = \nz.mem_2113_sv2v_reg ;
  assign \nz.mem [2112] = \nz.mem_2112_sv2v_reg ;
  assign \nz.mem [2111] = \nz.mem_2111_sv2v_reg ;
  assign \nz.mem [2110] = \nz.mem_2110_sv2v_reg ;
  assign \nz.mem [2109] = \nz.mem_2109_sv2v_reg ;
  assign \nz.mem [2108] = \nz.mem_2108_sv2v_reg ;
  assign \nz.mem [2107] = \nz.mem_2107_sv2v_reg ;
  assign \nz.mem [2106] = \nz.mem_2106_sv2v_reg ;
  assign \nz.mem [2105] = \nz.mem_2105_sv2v_reg ;
  assign \nz.mem [2104] = \nz.mem_2104_sv2v_reg ;
  assign \nz.mem [2103] = \nz.mem_2103_sv2v_reg ;
  assign \nz.mem [2102] = \nz.mem_2102_sv2v_reg ;
  assign \nz.mem [2101] = \nz.mem_2101_sv2v_reg ;
  assign \nz.mem [2100] = \nz.mem_2100_sv2v_reg ;
  assign \nz.mem [2099] = \nz.mem_2099_sv2v_reg ;
  assign \nz.mem [2098] = \nz.mem_2098_sv2v_reg ;
  assign \nz.mem [2097] = \nz.mem_2097_sv2v_reg ;
  assign \nz.mem [2096] = \nz.mem_2096_sv2v_reg ;
  assign \nz.mem [2095] = \nz.mem_2095_sv2v_reg ;
  assign \nz.mem [2094] = \nz.mem_2094_sv2v_reg ;
  assign \nz.mem [2093] = \nz.mem_2093_sv2v_reg ;
  assign \nz.mem [2092] = \nz.mem_2092_sv2v_reg ;
  assign \nz.mem [2091] = \nz.mem_2091_sv2v_reg ;
  assign \nz.mem [2090] = \nz.mem_2090_sv2v_reg ;
  assign \nz.mem [2089] = \nz.mem_2089_sv2v_reg ;
  assign \nz.mem [2088] = \nz.mem_2088_sv2v_reg ;
  assign \nz.mem [2087] = \nz.mem_2087_sv2v_reg ;
  assign \nz.mem [2086] = \nz.mem_2086_sv2v_reg ;
  assign \nz.mem [2085] = \nz.mem_2085_sv2v_reg ;
  assign \nz.mem [2084] = \nz.mem_2084_sv2v_reg ;
  assign \nz.mem [2083] = \nz.mem_2083_sv2v_reg ;
  assign \nz.mem [2082] = \nz.mem_2082_sv2v_reg ;
  assign \nz.mem [2081] = \nz.mem_2081_sv2v_reg ;
  assign \nz.mem [2080] = \nz.mem_2080_sv2v_reg ;
  assign \nz.mem [2079] = \nz.mem_2079_sv2v_reg ;
  assign \nz.mem [2078] = \nz.mem_2078_sv2v_reg ;
  assign \nz.mem [2077] = \nz.mem_2077_sv2v_reg ;
  assign \nz.mem [2076] = \nz.mem_2076_sv2v_reg ;
  assign \nz.mem [2075] = \nz.mem_2075_sv2v_reg ;
  assign \nz.mem [2074] = \nz.mem_2074_sv2v_reg ;
  assign \nz.mem [2073] = \nz.mem_2073_sv2v_reg ;
  assign \nz.mem [2072] = \nz.mem_2072_sv2v_reg ;
  assign \nz.mem [2071] = \nz.mem_2071_sv2v_reg ;
  assign \nz.mem [2070] = \nz.mem_2070_sv2v_reg ;
  assign \nz.mem [2069] = \nz.mem_2069_sv2v_reg ;
  assign \nz.mem [2068] = \nz.mem_2068_sv2v_reg ;
  assign \nz.mem [2067] = \nz.mem_2067_sv2v_reg ;
  assign \nz.mem [2066] = \nz.mem_2066_sv2v_reg ;
  assign \nz.mem [2065] = \nz.mem_2065_sv2v_reg ;
  assign \nz.mem [2064] = \nz.mem_2064_sv2v_reg ;
  assign \nz.mem [2063] = \nz.mem_2063_sv2v_reg ;
  assign \nz.mem [2062] = \nz.mem_2062_sv2v_reg ;
  assign \nz.mem [2061] = \nz.mem_2061_sv2v_reg ;
  assign \nz.mem [2060] = \nz.mem_2060_sv2v_reg ;
  assign \nz.mem [2059] = \nz.mem_2059_sv2v_reg ;
  assign \nz.mem [2058] = \nz.mem_2058_sv2v_reg ;
  assign \nz.mem [2057] = \nz.mem_2057_sv2v_reg ;
  assign \nz.mem [2056] = \nz.mem_2056_sv2v_reg ;
  assign \nz.mem [2055] = \nz.mem_2055_sv2v_reg ;
  assign \nz.mem [2054] = \nz.mem_2054_sv2v_reg ;
  assign \nz.mem [2053] = \nz.mem_2053_sv2v_reg ;
  assign \nz.mem [2052] = \nz.mem_2052_sv2v_reg ;
  assign \nz.mem [2051] = \nz.mem_2051_sv2v_reg ;
  assign \nz.mem [2050] = \nz.mem_2050_sv2v_reg ;
  assign \nz.mem [2049] = \nz.mem_2049_sv2v_reg ;
  assign \nz.mem [2048] = \nz.mem_2048_sv2v_reg ;
  assign \nz.mem [2047] = \nz.mem_2047_sv2v_reg ;
  assign \nz.mem [2046] = \nz.mem_2046_sv2v_reg ;
  assign \nz.mem [2045] = \nz.mem_2045_sv2v_reg ;
  assign \nz.mem [2044] = \nz.mem_2044_sv2v_reg ;
  assign \nz.mem [2043] = \nz.mem_2043_sv2v_reg ;
  assign \nz.mem [2042] = \nz.mem_2042_sv2v_reg ;
  assign \nz.mem [2041] = \nz.mem_2041_sv2v_reg ;
  assign \nz.mem [2040] = \nz.mem_2040_sv2v_reg ;
  assign \nz.mem [2039] = \nz.mem_2039_sv2v_reg ;
  assign \nz.mem [2038] = \nz.mem_2038_sv2v_reg ;
  assign \nz.mem [2037] = \nz.mem_2037_sv2v_reg ;
  assign \nz.mem [2036] = \nz.mem_2036_sv2v_reg ;
  assign \nz.mem [2035] = \nz.mem_2035_sv2v_reg ;
  assign \nz.mem [2034] = \nz.mem_2034_sv2v_reg ;
  assign \nz.mem [2033] = \nz.mem_2033_sv2v_reg ;
  assign \nz.mem [2032] = \nz.mem_2032_sv2v_reg ;
  assign \nz.mem [2031] = \nz.mem_2031_sv2v_reg ;
  assign \nz.mem [2030] = \nz.mem_2030_sv2v_reg ;
  assign \nz.mem [2029] = \nz.mem_2029_sv2v_reg ;
  assign \nz.mem [2028] = \nz.mem_2028_sv2v_reg ;
  assign \nz.mem [2027] = \nz.mem_2027_sv2v_reg ;
  assign \nz.mem [2026] = \nz.mem_2026_sv2v_reg ;
  assign \nz.mem [2025] = \nz.mem_2025_sv2v_reg ;
  assign \nz.mem [2024] = \nz.mem_2024_sv2v_reg ;
  assign \nz.mem [2023] = \nz.mem_2023_sv2v_reg ;
  assign \nz.mem [2022] = \nz.mem_2022_sv2v_reg ;
  assign \nz.mem [2021] = \nz.mem_2021_sv2v_reg ;
  assign \nz.mem [2020] = \nz.mem_2020_sv2v_reg ;
  assign \nz.mem [2019] = \nz.mem_2019_sv2v_reg ;
  assign \nz.mem [2018] = \nz.mem_2018_sv2v_reg ;
  assign \nz.mem [2017] = \nz.mem_2017_sv2v_reg ;
  assign \nz.mem [2016] = \nz.mem_2016_sv2v_reg ;
  assign \nz.mem [2015] = \nz.mem_2015_sv2v_reg ;
  assign \nz.mem [2014] = \nz.mem_2014_sv2v_reg ;
  assign \nz.mem [2013] = \nz.mem_2013_sv2v_reg ;
  assign \nz.mem [2012] = \nz.mem_2012_sv2v_reg ;
  assign \nz.mem [2011] = \nz.mem_2011_sv2v_reg ;
  assign \nz.mem [2010] = \nz.mem_2010_sv2v_reg ;
  assign \nz.mem [2009] = \nz.mem_2009_sv2v_reg ;
  assign \nz.mem [2008] = \nz.mem_2008_sv2v_reg ;
  assign \nz.mem [2007] = \nz.mem_2007_sv2v_reg ;
  assign \nz.mem [2006] = \nz.mem_2006_sv2v_reg ;
  assign \nz.mem [2005] = \nz.mem_2005_sv2v_reg ;
  assign \nz.mem [2004] = \nz.mem_2004_sv2v_reg ;
  assign \nz.mem [2003] = \nz.mem_2003_sv2v_reg ;
  assign \nz.mem [2002] = \nz.mem_2002_sv2v_reg ;
  assign \nz.mem [2001] = \nz.mem_2001_sv2v_reg ;
  assign \nz.mem [2000] = \nz.mem_2000_sv2v_reg ;
  assign \nz.mem [1999] = \nz.mem_1999_sv2v_reg ;
  assign \nz.mem [1998] = \nz.mem_1998_sv2v_reg ;
  assign \nz.mem [1997] = \nz.mem_1997_sv2v_reg ;
  assign \nz.mem [1996] = \nz.mem_1996_sv2v_reg ;
  assign \nz.mem [1995] = \nz.mem_1995_sv2v_reg ;
  assign \nz.mem [1994] = \nz.mem_1994_sv2v_reg ;
  assign \nz.mem [1993] = \nz.mem_1993_sv2v_reg ;
  assign \nz.mem [1992] = \nz.mem_1992_sv2v_reg ;
  assign \nz.mem [1991] = \nz.mem_1991_sv2v_reg ;
  assign \nz.mem [1990] = \nz.mem_1990_sv2v_reg ;
  assign \nz.mem [1989] = \nz.mem_1989_sv2v_reg ;
  assign \nz.mem [1988] = \nz.mem_1988_sv2v_reg ;
  assign \nz.mem [1987] = \nz.mem_1987_sv2v_reg ;
  assign \nz.mem [1986] = \nz.mem_1986_sv2v_reg ;
  assign \nz.mem [1985] = \nz.mem_1985_sv2v_reg ;
  assign \nz.mem [1984] = \nz.mem_1984_sv2v_reg ;
  assign \nz.mem [1983] = \nz.mem_1983_sv2v_reg ;
  assign \nz.mem [1982] = \nz.mem_1982_sv2v_reg ;
  assign \nz.mem [1981] = \nz.mem_1981_sv2v_reg ;
  assign \nz.mem [1980] = \nz.mem_1980_sv2v_reg ;
  assign \nz.mem [1979] = \nz.mem_1979_sv2v_reg ;
  assign \nz.mem [1978] = \nz.mem_1978_sv2v_reg ;
  assign \nz.mem [1977] = \nz.mem_1977_sv2v_reg ;
  assign \nz.mem [1976] = \nz.mem_1976_sv2v_reg ;
  assign \nz.mem [1975] = \nz.mem_1975_sv2v_reg ;
  assign \nz.mem [1974] = \nz.mem_1974_sv2v_reg ;
  assign \nz.mem [1973] = \nz.mem_1973_sv2v_reg ;
  assign \nz.mem [1972] = \nz.mem_1972_sv2v_reg ;
  assign \nz.mem [1971] = \nz.mem_1971_sv2v_reg ;
  assign \nz.mem [1970] = \nz.mem_1970_sv2v_reg ;
  assign \nz.mem [1969] = \nz.mem_1969_sv2v_reg ;
  assign \nz.mem [1968] = \nz.mem_1968_sv2v_reg ;
  assign \nz.mem [1967] = \nz.mem_1967_sv2v_reg ;
  assign \nz.mem [1966] = \nz.mem_1966_sv2v_reg ;
  assign \nz.mem [1965] = \nz.mem_1965_sv2v_reg ;
  assign \nz.mem [1964] = \nz.mem_1964_sv2v_reg ;
  assign \nz.mem [1963] = \nz.mem_1963_sv2v_reg ;
  assign \nz.mem [1962] = \nz.mem_1962_sv2v_reg ;
  assign \nz.mem [1961] = \nz.mem_1961_sv2v_reg ;
  assign \nz.mem [1960] = \nz.mem_1960_sv2v_reg ;
  assign \nz.mem [1959] = \nz.mem_1959_sv2v_reg ;
  assign \nz.mem [1958] = \nz.mem_1958_sv2v_reg ;
  assign \nz.mem [1957] = \nz.mem_1957_sv2v_reg ;
  assign \nz.mem [1956] = \nz.mem_1956_sv2v_reg ;
  assign \nz.mem [1955] = \nz.mem_1955_sv2v_reg ;
  assign \nz.mem [1954] = \nz.mem_1954_sv2v_reg ;
  assign \nz.mem [1953] = \nz.mem_1953_sv2v_reg ;
  assign \nz.mem [1952] = \nz.mem_1952_sv2v_reg ;
  assign \nz.mem [1951] = \nz.mem_1951_sv2v_reg ;
  assign \nz.mem [1950] = \nz.mem_1950_sv2v_reg ;
  assign \nz.mem [1949] = \nz.mem_1949_sv2v_reg ;
  assign \nz.mem [1948] = \nz.mem_1948_sv2v_reg ;
  assign \nz.mem [1947] = \nz.mem_1947_sv2v_reg ;
  assign \nz.mem [1946] = \nz.mem_1946_sv2v_reg ;
  assign \nz.mem [1945] = \nz.mem_1945_sv2v_reg ;
  assign \nz.mem [1944] = \nz.mem_1944_sv2v_reg ;
  assign \nz.mem [1943] = \nz.mem_1943_sv2v_reg ;
  assign \nz.mem [1942] = \nz.mem_1942_sv2v_reg ;
  assign \nz.mem [1941] = \nz.mem_1941_sv2v_reg ;
  assign \nz.mem [1940] = \nz.mem_1940_sv2v_reg ;
  assign \nz.mem [1939] = \nz.mem_1939_sv2v_reg ;
  assign \nz.mem [1938] = \nz.mem_1938_sv2v_reg ;
  assign \nz.mem [1937] = \nz.mem_1937_sv2v_reg ;
  assign \nz.mem [1936] = \nz.mem_1936_sv2v_reg ;
  assign \nz.mem [1935] = \nz.mem_1935_sv2v_reg ;
  assign \nz.mem [1934] = \nz.mem_1934_sv2v_reg ;
  assign \nz.mem [1933] = \nz.mem_1933_sv2v_reg ;
  assign \nz.mem [1932] = \nz.mem_1932_sv2v_reg ;
  assign \nz.mem [1931] = \nz.mem_1931_sv2v_reg ;
  assign \nz.mem [1930] = \nz.mem_1930_sv2v_reg ;
  assign \nz.mem [1929] = \nz.mem_1929_sv2v_reg ;
  assign \nz.mem [1928] = \nz.mem_1928_sv2v_reg ;
  assign \nz.mem [1927] = \nz.mem_1927_sv2v_reg ;
  assign \nz.mem [1926] = \nz.mem_1926_sv2v_reg ;
  assign \nz.mem [1925] = \nz.mem_1925_sv2v_reg ;
  assign \nz.mem [1924] = \nz.mem_1924_sv2v_reg ;
  assign \nz.mem [1923] = \nz.mem_1923_sv2v_reg ;
  assign \nz.mem [1922] = \nz.mem_1922_sv2v_reg ;
  assign \nz.mem [1921] = \nz.mem_1921_sv2v_reg ;
  assign \nz.mem [1920] = \nz.mem_1920_sv2v_reg ;
  assign \nz.mem [1919] = \nz.mem_1919_sv2v_reg ;
  assign \nz.mem [1918] = \nz.mem_1918_sv2v_reg ;
  assign \nz.mem [1917] = \nz.mem_1917_sv2v_reg ;
  assign \nz.mem [1916] = \nz.mem_1916_sv2v_reg ;
  assign \nz.mem [1915] = \nz.mem_1915_sv2v_reg ;
  assign \nz.mem [1914] = \nz.mem_1914_sv2v_reg ;
  assign \nz.mem [1913] = \nz.mem_1913_sv2v_reg ;
  assign \nz.mem [1912] = \nz.mem_1912_sv2v_reg ;
  assign \nz.mem [1911] = \nz.mem_1911_sv2v_reg ;
  assign \nz.mem [1910] = \nz.mem_1910_sv2v_reg ;
  assign \nz.mem [1909] = \nz.mem_1909_sv2v_reg ;
  assign \nz.mem [1908] = \nz.mem_1908_sv2v_reg ;
  assign \nz.mem [1907] = \nz.mem_1907_sv2v_reg ;
  assign \nz.mem [1906] = \nz.mem_1906_sv2v_reg ;
  assign \nz.mem [1905] = \nz.mem_1905_sv2v_reg ;
  assign \nz.mem [1904] = \nz.mem_1904_sv2v_reg ;
  assign \nz.mem [1903] = \nz.mem_1903_sv2v_reg ;
  assign \nz.mem [1902] = \nz.mem_1902_sv2v_reg ;
  assign \nz.mem [1901] = \nz.mem_1901_sv2v_reg ;
  assign \nz.mem [1900] = \nz.mem_1900_sv2v_reg ;
  assign \nz.mem [1899] = \nz.mem_1899_sv2v_reg ;
  assign \nz.mem [1898] = \nz.mem_1898_sv2v_reg ;
  assign \nz.mem [1897] = \nz.mem_1897_sv2v_reg ;
  assign \nz.mem [1896] = \nz.mem_1896_sv2v_reg ;
  assign \nz.mem [1895] = \nz.mem_1895_sv2v_reg ;
  assign \nz.mem [1894] = \nz.mem_1894_sv2v_reg ;
  assign \nz.mem [1893] = \nz.mem_1893_sv2v_reg ;
  assign \nz.mem [1892] = \nz.mem_1892_sv2v_reg ;
  assign \nz.mem [1891] = \nz.mem_1891_sv2v_reg ;
  assign \nz.mem [1890] = \nz.mem_1890_sv2v_reg ;
  assign \nz.mem [1889] = \nz.mem_1889_sv2v_reg ;
  assign \nz.mem [1888] = \nz.mem_1888_sv2v_reg ;
  assign \nz.mem [1887] = \nz.mem_1887_sv2v_reg ;
  assign \nz.mem [1886] = \nz.mem_1886_sv2v_reg ;
  assign \nz.mem [1885] = \nz.mem_1885_sv2v_reg ;
  assign \nz.mem [1884] = \nz.mem_1884_sv2v_reg ;
  assign \nz.mem [1883] = \nz.mem_1883_sv2v_reg ;
  assign \nz.mem [1882] = \nz.mem_1882_sv2v_reg ;
  assign \nz.mem [1881] = \nz.mem_1881_sv2v_reg ;
  assign \nz.mem [1880] = \nz.mem_1880_sv2v_reg ;
  assign \nz.mem [1879] = \nz.mem_1879_sv2v_reg ;
  assign \nz.mem [1878] = \nz.mem_1878_sv2v_reg ;
  assign \nz.mem [1877] = \nz.mem_1877_sv2v_reg ;
  assign \nz.mem [1876] = \nz.mem_1876_sv2v_reg ;
  assign \nz.mem [1875] = \nz.mem_1875_sv2v_reg ;
  assign \nz.mem [1874] = \nz.mem_1874_sv2v_reg ;
  assign \nz.mem [1873] = \nz.mem_1873_sv2v_reg ;
  assign \nz.mem [1872] = \nz.mem_1872_sv2v_reg ;
  assign \nz.mem [1871] = \nz.mem_1871_sv2v_reg ;
  assign \nz.mem [1870] = \nz.mem_1870_sv2v_reg ;
  assign \nz.mem [1869] = \nz.mem_1869_sv2v_reg ;
  assign \nz.mem [1868] = \nz.mem_1868_sv2v_reg ;
  assign \nz.mem [1867] = \nz.mem_1867_sv2v_reg ;
  assign \nz.mem [1866] = \nz.mem_1866_sv2v_reg ;
  assign \nz.mem [1865] = \nz.mem_1865_sv2v_reg ;
  assign \nz.mem [1864] = \nz.mem_1864_sv2v_reg ;
  assign \nz.mem [1863] = \nz.mem_1863_sv2v_reg ;
  assign \nz.mem [1862] = \nz.mem_1862_sv2v_reg ;
  assign \nz.mem [1861] = \nz.mem_1861_sv2v_reg ;
  assign \nz.mem [1860] = \nz.mem_1860_sv2v_reg ;
  assign \nz.mem [1859] = \nz.mem_1859_sv2v_reg ;
  assign \nz.mem [1858] = \nz.mem_1858_sv2v_reg ;
  assign \nz.mem [1857] = \nz.mem_1857_sv2v_reg ;
  assign \nz.mem [1856] = \nz.mem_1856_sv2v_reg ;
  assign \nz.mem [1855] = \nz.mem_1855_sv2v_reg ;
  assign \nz.mem [1854] = \nz.mem_1854_sv2v_reg ;
  assign \nz.mem [1853] = \nz.mem_1853_sv2v_reg ;
  assign \nz.mem [1852] = \nz.mem_1852_sv2v_reg ;
  assign \nz.mem [1851] = \nz.mem_1851_sv2v_reg ;
  assign \nz.mem [1850] = \nz.mem_1850_sv2v_reg ;
  assign \nz.mem [1849] = \nz.mem_1849_sv2v_reg ;
  assign \nz.mem [1848] = \nz.mem_1848_sv2v_reg ;
  assign \nz.mem [1847] = \nz.mem_1847_sv2v_reg ;
  assign \nz.mem [1846] = \nz.mem_1846_sv2v_reg ;
  assign \nz.mem [1845] = \nz.mem_1845_sv2v_reg ;
  assign \nz.mem [1844] = \nz.mem_1844_sv2v_reg ;
  assign \nz.mem [1843] = \nz.mem_1843_sv2v_reg ;
  assign \nz.mem [1842] = \nz.mem_1842_sv2v_reg ;
  assign \nz.mem [1841] = \nz.mem_1841_sv2v_reg ;
  assign \nz.mem [1840] = \nz.mem_1840_sv2v_reg ;
  assign \nz.mem [1839] = \nz.mem_1839_sv2v_reg ;
  assign \nz.mem [1838] = \nz.mem_1838_sv2v_reg ;
  assign \nz.mem [1837] = \nz.mem_1837_sv2v_reg ;
  assign \nz.mem [1836] = \nz.mem_1836_sv2v_reg ;
  assign \nz.mem [1835] = \nz.mem_1835_sv2v_reg ;
  assign \nz.mem [1834] = \nz.mem_1834_sv2v_reg ;
  assign \nz.mem [1833] = \nz.mem_1833_sv2v_reg ;
  assign \nz.mem [1832] = \nz.mem_1832_sv2v_reg ;
  assign \nz.mem [1831] = \nz.mem_1831_sv2v_reg ;
  assign \nz.mem [1830] = \nz.mem_1830_sv2v_reg ;
  assign \nz.mem [1829] = \nz.mem_1829_sv2v_reg ;
  assign \nz.mem [1828] = \nz.mem_1828_sv2v_reg ;
  assign \nz.mem [1827] = \nz.mem_1827_sv2v_reg ;
  assign \nz.mem [1826] = \nz.mem_1826_sv2v_reg ;
  assign \nz.mem [1825] = \nz.mem_1825_sv2v_reg ;
  assign \nz.mem [1824] = \nz.mem_1824_sv2v_reg ;
  assign \nz.mem [1823] = \nz.mem_1823_sv2v_reg ;
  assign \nz.mem [1822] = \nz.mem_1822_sv2v_reg ;
  assign \nz.mem [1821] = \nz.mem_1821_sv2v_reg ;
  assign \nz.mem [1820] = \nz.mem_1820_sv2v_reg ;
  assign \nz.mem [1819] = \nz.mem_1819_sv2v_reg ;
  assign \nz.mem [1818] = \nz.mem_1818_sv2v_reg ;
  assign \nz.mem [1817] = \nz.mem_1817_sv2v_reg ;
  assign \nz.mem [1816] = \nz.mem_1816_sv2v_reg ;
  assign \nz.mem [1815] = \nz.mem_1815_sv2v_reg ;
  assign \nz.mem [1814] = \nz.mem_1814_sv2v_reg ;
  assign \nz.mem [1813] = \nz.mem_1813_sv2v_reg ;
  assign \nz.mem [1812] = \nz.mem_1812_sv2v_reg ;
  assign \nz.mem [1811] = \nz.mem_1811_sv2v_reg ;
  assign \nz.mem [1810] = \nz.mem_1810_sv2v_reg ;
  assign \nz.mem [1809] = \nz.mem_1809_sv2v_reg ;
  assign \nz.mem [1808] = \nz.mem_1808_sv2v_reg ;
  assign \nz.mem [1807] = \nz.mem_1807_sv2v_reg ;
  assign \nz.mem [1806] = \nz.mem_1806_sv2v_reg ;
  assign \nz.mem [1805] = \nz.mem_1805_sv2v_reg ;
  assign \nz.mem [1804] = \nz.mem_1804_sv2v_reg ;
  assign \nz.mem [1803] = \nz.mem_1803_sv2v_reg ;
  assign \nz.mem [1802] = \nz.mem_1802_sv2v_reg ;
  assign \nz.mem [1801] = \nz.mem_1801_sv2v_reg ;
  assign \nz.mem [1800] = \nz.mem_1800_sv2v_reg ;
  assign \nz.mem [1799] = \nz.mem_1799_sv2v_reg ;
  assign \nz.mem [1798] = \nz.mem_1798_sv2v_reg ;
  assign \nz.mem [1797] = \nz.mem_1797_sv2v_reg ;
  assign \nz.mem [1796] = \nz.mem_1796_sv2v_reg ;
  assign \nz.mem [1795] = \nz.mem_1795_sv2v_reg ;
  assign \nz.mem [1794] = \nz.mem_1794_sv2v_reg ;
  assign \nz.mem [1793] = \nz.mem_1793_sv2v_reg ;
  assign \nz.mem [1792] = \nz.mem_1792_sv2v_reg ;
  assign \nz.mem [1791] = \nz.mem_1791_sv2v_reg ;
  assign \nz.mem [1790] = \nz.mem_1790_sv2v_reg ;
  assign \nz.mem [1789] = \nz.mem_1789_sv2v_reg ;
  assign \nz.mem [1788] = \nz.mem_1788_sv2v_reg ;
  assign \nz.mem [1787] = \nz.mem_1787_sv2v_reg ;
  assign \nz.mem [1786] = \nz.mem_1786_sv2v_reg ;
  assign \nz.mem [1785] = \nz.mem_1785_sv2v_reg ;
  assign \nz.mem [1784] = \nz.mem_1784_sv2v_reg ;
  assign \nz.mem [1783] = \nz.mem_1783_sv2v_reg ;
  assign \nz.mem [1782] = \nz.mem_1782_sv2v_reg ;
  assign \nz.mem [1781] = \nz.mem_1781_sv2v_reg ;
  assign \nz.mem [1780] = \nz.mem_1780_sv2v_reg ;
  assign \nz.mem [1779] = \nz.mem_1779_sv2v_reg ;
  assign \nz.mem [1778] = \nz.mem_1778_sv2v_reg ;
  assign \nz.mem [1777] = \nz.mem_1777_sv2v_reg ;
  assign \nz.mem [1776] = \nz.mem_1776_sv2v_reg ;
  assign \nz.mem [1775] = \nz.mem_1775_sv2v_reg ;
  assign \nz.mem [1774] = \nz.mem_1774_sv2v_reg ;
  assign \nz.mem [1773] = \nz.mem_1773_sv2v_reg ;
  assign \nz.mem [1772] = \nz.mem_1772_sv2v_reg ;
  assign \nz.mem [1771] = \nz.mem_1771_sv2v_reg ;
  assign \nz.mem [1770] = \nz.mem_1770_sv2v_reg ;
  assign \nz.mem [1769] = \nz.mem_1769_sv2v_reg ;
  assign \nz.mem [1768] = \nz.mem_1768_sv2v_reg ;
  assign \nz.mem [1767] = \nz.mem_1767_sv2v_reg ;
  assign \nz.mem [1766] = \nz.mem_1766_sv2v_reg ;
  assign \nz.mem [1765] = \nz.mem_1765_sv2v_reg ;
  assign \nz.mem [1764] = \nz.mem_1764_sv2v_reg ;
  assign \nz.mem [1763] = \nz.mem_1763_sv2v_reg ;
  assign \nz.mem [1762] = \nz.mem_1762_sv2v_reg ;
  assign \nz.mem [1761] = \nz.mem_1761_sv2v_reg ;
  assign \nz.mem [1760] = \nz.mem_1760_sv2v_reg ;
  assign \nz.mem [1759] = \nz.mem_1759_sv2v_reg ;
  assign \nz.mem [1758] = \nz.mem_1758_sv2v_reg ;
  assign \nz.mem [1757] = \nz.mem_1757_sv2v_reg ;
  assign \nz.mem [1756] = \nz.mem_1756_sv2v_reg ;
  assign \nz.mem [1755] = \nz.mem_1755_sv2v_reg ;
  assign \nz.mem [1754] = \nz.mem_1754_sv2v_reg ;
  assign \nz.mem [1753] = \nz.mem_1753_sv2v_reg ;
  assign \nz.mem [1752] = \nz.mem_1752_sv2v_reg ;
  assign \nz.mem [1751] = \nz.mem_1751_sv2v_reg ;
  assign \nz.mem [1750] = \nz.mem_1750_sv2v_reg ;
  assign \nz.mem [1749] = \nz.mem_1749_sv2v_reg ;
  assign \nz.mem [1748] = \nz.mem_1748_sv2v_reg ;
  assign \nz.mem [1747] = \nz.mem_1747_sv2v_reg ;
  assign \nz.mem [1746] = \nz.mem_1746_sv2v_reg ;
  assign \nz.mem [1745] = \nz.mem_1745_sv2v_reg ;
  assign \nz.mem [1744] = \nz.mem_1744_sv2v_reg ;
  assign \nz.mem [1743] = \nz.mem_1743_sv2v_reg ;
  assign \nz.mem [1742] = \nz.mem_1742_sv2v_reg ;
  assign \nz.mem [1741] = \nz.mem_1741_sv2v_reg ;
  assign \nz.mem [1740] = \nz.mem_1740_sv2v_reg ;
  assign \nz.mem [1739] = \nz.mem_1739_sv2v_reg ;
  assign \nz.mem [1738] = \nz.mem_1738_sv2v_reg ;
  assign \nz.mem [1737] = \nz.mem_1737_sv2v_reg ;
  assign \nz.mem [1736] = \nz.mem_1736_sv2v_reg ;
  assign \nz.mem [1735] = \nz.mem_1735_sv2v_reg ;
  assign \nz.mem [1734] = \nz.mem_1734_sv2v_reg ;
  assign \nz.mem [1733] = \nz.mem_1733_sv2v_reg ;
  assign \nz.mem [1732] = \nz.mem_1732_sv2v_reg ;
  assign \nz.mem [1731] = \nz.mem_1731_sv2v_reg ;
  assign \nz.mem [1730] = \nz.mem_1730_sv2v_reg ;
  assign \nz.mem [1729] = \nz.mem_1729_sv2v_reg ;
  assign \nz.mem [1728] = \nz.mem_1728_sv2v_reg ;
  assign \nz.mem [1727] = \nz.mem_1727_sv2v_reg ;
  assign \nz.mem [1726] = \nz.mem_1726_sv2v_reg ;
  assign \nz.mem [1725] = \nz.mem_1725_sv2v_reg ;
  assign \nz.mem [1724] = \nz.mem_1724_sv2v_reg ;
  assign \nz.mem [1723] = \nz.mem_1723_sv2v_reg ;
  assign \nz.mem [1722] = \nz.mem_1722_sv2v_reg ;
  assign \nz.mem [1721] = \nz.mem_1721_sv2v_reg ;
  assign \nz.mem [1720] = \nz.mem_1720_sv2v_reg ;
  assign \nz.mem [1719] = \nz.mem_1719_sv2v_reg ;
  assign \nz.mem [1718] = \nz.mem_1718_sv2v_reg ;
  assign \nz.mem [1717] = \nz.mem_1717_sv2v_reg ;
  assign \nz.mem [1716] = \nz.mem_1716_sv2v_reg ;
  assign \nz.mem [1715] = \nz.mem_1715_sv2v_reg ;
  assign \nz.mem [1714] = \nz.mem_1714_sv2v_reg ;
  assign \nz.mem [1713] = \nz.mem_1713_sv2v_reg ;
  assign \nz.mem [1712] = \nz.mem_1712_sv2v_reg ;
  assign \nz.mem [1711] = \nz.mem_1711_sv2v_reg ;
  assign \nz.mem [1710] = \nz.mem_1710_sv2v_reg ;
  assign \nz.mem [1709] = \nz.mem_1709_sv2v_reg ;
  assign \nz.mem [1708] = \nz.mem_1708_sv2v_reg ;
  assign \nz.mem [1707] = \nz.mem_1707_sv2v_reg ;
  assign \nz.mem [1706] = \nz.mem_1706_sv2v_reg ;
  assign \nz.mem [1705] = \nz.mem_1705_sv2v_reg ;
  assign \nz.mem [1704] = \nz.mem_1704_sv2v_reg ;
  assign \nz.mem [1703] = \nz.mem_1703_sv2v_reg ;
  assign \nz.mem [1702] = \nz.mem_1702_sv2v_reg ;
  assign \nz.mem [1701] = \nz.mem_1701_sv2v_reg ;
  assign \nz.mem [1700] = \nz.mem_1700_sv2v_reg ;
  assign \nz.mem [1699] = \nz.mem_1699_sv2v_reg ;
  assign \nz.mem [1698] = \nz.mem_1698_sv2v_reg ;
  assign \nz.mem [1697] = \nz.mem_1697_sv2v_reg ;
  assign \nz.mem [1696] = \nz.mem_1696_sv2v_reg ;
  assign \nz.mem [1695] = \nz.mem_1695_sv2v_reg ;
  assign \nz.mem [1694] = \nz.mem_1694_sv2v_reg ;
  assign \nz.mem [1693] = \nz.mem_1693_sv2v_reg ;
  assign \nz.mem [1692] = \nz.mem_1692_sv2v_reg ;
  assign \nz.mem [1691] = \nz.mem_1691_sv2v_reg ;
  assign \nz.mem [1690] = \nz.mem_1690_sv2v_reg ;
  assign \nz.mem [1689] = \nz.mem_1689_sv2v_reg ;
  assign \nz.mem [1688] = \nz.mem_1688_sv2v_reg ;
  assign \nz.mem [1687] = \nz.mem_1687_sv2v_reg ;
  assign \nz.mem [1686] = \nz.mem_1686_sv2v_reg ;
  assign \nz.mem [1685] = \nz.mem_1685_sv2v_reg ;
  assign \nz.mem [1684] = \nz.mem_1684_sv2v_reg ;
  assign \nz.mem [1683] = \nz.mem_1683_sv2v_reg ;
  assign \nz.mem [1682] = \nz.mem_1682_sv2v_reg ;
  assign \nz.mem [1681] = \nz.mem_1681_sv2v_reg ;
  assign \nz.mem [1680] = \nz.mem_1680_sv2v_reg ;
  assign \nz.mem [1679] = \nz.mem_1679_sv2v_reg ;
  assign \nz.mem [1678] = \nz.mem_1678_sv2v_reg ;
  assign \nz.mem [1677] = \nz.mem_1677_sv2v_reg ;
  assign \nz.mem [1676] = \nz.mem_1676_sv2v_reg ;
  assign \nz.mem [1675] = \nz.mem_1675_sv2v_reg ;
  assign \nz.mem [1674] = \nz.mem_1674_sv2v_reg ;
  assign \nz.mem [1673] = \nz.mem_1673_sv2v_reg ;
  assign \nz.mem [1672] = \nz.mem_1672_sv2v_reg ;
  assign \nz.mem [1671] = \nz.mem_1671_sv2v_reg ;
  assign \nz.mem [1670] = \nz.mem_1670_sv2v_reg ;
  assign \nz.mem [1669] = \nz.mem_1669_sv2v_reg ;
  assign \nz.mem [1668] = \nz.mem_1668_sv2v_reg ;
  assign \nz.mem [1667] = \nz.mem_1667_sv2v_reg ;
  assign \nz.mem [1666] = \nz.mem_1666_sv2v_reg ;
  assign \nz.mem [1665] = \nz.mem_1665_sv2v_reg ;
  assign \nz.mem [1664] = \nz.mem_1664_sv2v_reg ;
  assign \nz.mem [1663] = \nz.mem_1663_sv2v_reg ;
  assign \nz.mem [1662] = \nz.mem_1662_sv2v_reg ;
  assign \nz.mem [1661] = \nz.mem_1661_sv2v_reg ;
  assign \nz.mem [1660] = \nz.mem_1660_sv2v_reg ;
  assign \nz.mem [1659] = \nz.mem_1659_sv2v_reg ;
  assign \nz.mem [1658] = \nz.mem_1658_sv2v_reg ;
  assign \nz.mem [1657] = \nz.mem_1657_sv2v_reg ;
  assign \nz.mem [1656] = \nz.mem_1656_sv2v_reg ;
  assign \nz.mem [1655] = \nz.mem_1655_sv2v_reg ;
  assign \nz.mem [1654] = \nz.mem_1654_sv2v_reg ;
  assign \nz.mem [1653] = \nz.mem_1653_sv2v_reg ;
  assign \nz.mem [1652] = \nz.mem_1652_sv2v_reg ;
  assign \nz.mem [1651] = \nz.mem_1651_sv2v_reg ;
  assign \nz.mem [1650] = \nz.mem_1650_sv2v_reg ;
  assign \nz.mem [1649] = \nz.mem_1649_sv2v_reg ;
  assign \nz.mem [1648] = \nz.mem_1648_sv2v_reg ;
  assign \nz.mem [1647] = \nz.mem_1647_sv2v_reg ;
  assign \nz.mem [1646] = \nz.mem_1646_sv2v_reg ;
  assign \nz.mem [1645] = \nz.mem_1645_sv2v_reg ;
  assign \nz.mem [1644] = \nz.mem_1644_sv2v_reg ;
  assign \nz.mem [1643] = \nz.mem_1643_sv2v_reg ;
  assign \nz.mem [1642] = \nz.mem_1642_sv2v_reg ;
  assign \nz.mem [1641] = \nz.mem_1641_sv2v_reg ;
  assign \nz.mem [1640] = \nz.mem_1640_sv2v_reg ;
  assign \nz.mem [1639] = \nz.mem_1639_sv2v_reg ;
  assign \nz.mem [1638] = \nz.mem_1638_sv2v_reg ;
  assign \nz.mem [1637] = \nz.mem_1637_sv2v_reg ;
  assign \nz.mem [1636] = \nz.mem_1636_sv2v_reg ;
  assign \nz.mem [1635] = \nz.mem_1635_sv2v_reg ;
  assign \nz.mem [1634] = \nz.mem_1634_sv2v_reg ;
  assign \nz.mem [1633] = \nz.mem_1633_sv2v_reg ;
  assign \nz.mem [1632] = \nz.mem_1632_sv2v_reg ;
  assign \nz.mem [1631] = \nz.mem_1631_sv2v_reg ;
  assign \nz.mem [1630] = \nz.mem_1630_sv2v_reg ;
  assign \nz.mem [1629] = \nz.mem_1629_sv2v_reg ;
  assign \nz.mem [1628] = \nz.mem_1628_sv2v_reg ;
  assign \nz.mem [1627] = \nz.mem_1627_sv2v_reg ;
  assign \nz.mem [1626] = \nz.mem_1626_sv2v_reg ;
  assign \nz.mem [1625] = \nz.mem_1625_sv2v_reg ;
  assign \nz.mem [1624] = \nz.mem_1624_sv2v_reg ;
  assign \nz.mem [1623] = \nz.mem_1623_sv2v_reg ;
  assign \nz.mem [1622] = \nz.mem_1622_sv2v_reg ;
  assign \nz.mem [1621] = \nz.mem_1621_sv2v_reg ;
  assign \nz.mem [1620] = \nz.mem_1620_sv2v_reg ;
  assign \nz.mem [1619] = \nz.mem_1619_sv2v_reg ;
  assign \nz.mem [1618] = \nz.mem_1618_sv2v_reg ;
  assign \nz.mem [1617] = \nz.mem_1617_sv2v_reg ;
  assign \nz.mem [1616] = \nz.mem_1616_sv2v_reg ;
  assign \nz.mem [1615] = \nz.mem_1615_sv2v_reg ;
  assign \nz.mem [1614] = \nz.mem_1614_sv2v_reg ;
  assign \nz.mem [1613] = \nz.mem_1613_sv2v_reg ;
  assign \nz.mem [1612] = \nz.mem_1612_sv2v_reg ;
  assign \nz.mem [1611] = \nz.mem_1611_sv2v_reg ;
  assign \nz.mem [1610] = \nz.mem_1610_sv2v_reg ;
  assign \nz.mem [1609] = \nz.mem_1609_sv2v_reg ;
  assign \nz.mem [1608] = \nz.mem_1608_sv2v_reg ;
  assign \nz.mem [1607] = \nz.mem_1607_sv2v_reg ;
  assign \nz.mem [1606] = \nz.mem_1606_sv2v_reg ;
  assign \nz.mem [1605] = \nz.mem_1605_sv2v_reg ;
  assign \nz.mem [1604] = \nz.mem_1604_sv2v_reg ;
  assign \nz.mem [1603] = \nz.mem_1603_sv2v_reg ;
  assign \nz.mem [1602] = \nz.mem_1602_sv2v_reg ;
  assign \nz.mem [1601] = \nz.mem_1601_sv2v_reg ;
  assign \nz.mem [1600] = \nz.mem_1600_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [79] = (N163)? \nz.mem [79] : 
                             (N165)? \nz.mem [159] : 
                             (N167)? \nz.mem [239] : 
                             (N169)? \nz.mem [319] : 
                             (N171)? \nz.mem [399] : 
                             (N173)? \nz.mem [479] : 
                             (N175)? \nz.mem [559] : 
                             (N177)? \nz.mem [639] : 
                             (N179)? \nz.mem [719] : 
                             (N181)? \nz.mem [799] : 
                             (N183)? \nz.mem [879] : 
                             (N185)? \nz.mem [959] : 
                             (N187)? \nz.mem [1039] : 
                             (N189)? \nz.mem [1119] : 
                             (N191)? \nz.mem [1199] : 
                             (N193)? \nz.mem [1279] : 
                             (N195)? \nz.mem [1359] : 
                             (N197)? \nz.mem [1439] : 
                             (N199)? \nz.mem [1519] : 
                             (N201)? \nz.mem [1599] : 
                             (N203)? \nz.mem [1679] : 
                             (N205)? \nz.mem [1759] : 
                             (N207)? \nz.mem [1839] : 
                             (N209)? \nz.mem [1919] : 
                             (N211)? \nz.mem [1999] : 
                             (N213)? \nz.mem [2079] : 
                             (N215)? \nz.mem [2159] : 
                             (N217)? \nz.mem [2239] : 
                             (N219)? \nz.mem [2319] : 
                             (N221)? \nz.mem [2399] : 
                             (N223)? \nz.mem [2479] : 
                             (N225)? \nz.mem [2559] : 
                             (N164)? \nz.mem [2639] : 
                             (N166)? \nz.mem [2719] : 
                             (N168)? \nz.mem [2799] : 
                             (N170)? \nz.mem [2879] : 
                             (N172)? \nz.mem [2959] : 
                             (N174)? \nz.mem [3039] : 
                             (N176)? \nz.mem [3119] : 
                             (N178)? \nz.mem [3199] : 
                             (N180)? \nz.mem [3279] : 
                             (N182)? \nz.mem [3359] : 
                             (N184)? \nz.mem [3439] : 
                             (N186)? \nz.mem [3519] : 
                             (N188)? \nz.mem [3599] : 
                             (N190)? \nz.mem [3679] : 
                             (N192)? \nz.mem [3759] : 
                             (N194)? \nz.mem [3839] : 
                             (N196)? \nz.mem [3919] : 
                             (N198)? \nz.mem [3999] : 
                             (N200)? \nz.mem [4079] : 
                             (N202)? \nz.mem [4159] : 
                             (N204)? \nz.mem [4239] : 
                             (N206)? \nz.mem [4319] : 
                             (N208)? \nz.mem [4399] : 
                             (N210)? \nz.mem [4479] : 
                             (N212)? \nz.mem [4559] : 
                             (N214)? \nz.mem [4639] : 
                             (N216)? \nz.mem [4719] : 
                             (N218)? \nz.mem [4799] : 
                             (N220)? \nz.mem [4879] : 
                             (N222)? \nz.mem [4959] : 
                             (N224)? \nz.mem [5039] : 
                             (N226)? \nz.mem [5119] : 1'b0;
  assign \nz.data_out [78] = (N163)? \nz.mem [78] : 
                             (N165)? \nz.mem [158] : 
                             (N167)? \nz.mem [238] : 
                             (N169)? \nz.mem [318] : 
                             (N171)? \nz.mem [398] : 
                             (N173)? \nz.mem [478] : 
                             (N175)? \nz.mem [558] : 
                             (N177)? \nz.mem [638] : 
                             (N179)? \nz.mem [718] : 
                             (N181)? \nz.mem [798] : 
                             (N183)? \nz.mem [878] : 
                             (N185)? \nz.mem [958] : 
                             (N187)? \nz.mem [1038] : 
                             (N189)? \nz.mem [1118] : 
                             (N191)? \nz.mem [1198] : 
                             (N193)? \nz.mem [1278] : 
                             (N195)? \nz.mem [1358] : 
                             (N197)? \nz.mem [1438] : 
                             (N199)? \nz.mem [1518] : 
                             (N201)? \nz.mem [1598] : 
                             (N203)? \nz.mem [1678] : 
                             (N205)? \nz.mem [1758] : 
                             (N207)? \nz.mem [1838] : 
                             (N209)? \nz.mem [1918] : 
                             (N211)? \nz.mem [1998] : 
                             (N213)? \nz.mem [2078] : 
                             (N215)? \nz.mem [2158] : 
                             (N217)? \nz.mem [2238] : 
                             (N219)? \nz.mem [2318] : 
                             (N221)? \nz.mem [2398] : 
                             (N223)? \nz.mem [2478] : 
                             (N225)? \nz.mem [2558] : 
                             (N164)? \nz.mem [2638] : 
                             (N166)? \nz.mem [2718] : 
                             (N168)? \nz.mem [2798] : 
                             (N170)? \nz.mem [2878] : 
                             (N172)? \nz.mem [2958] : 
                             (N174)? \nz.mem [3038] : 
                             (N176)? \nz.mem [3118] : 
                             (N178)? \nz.mem [3198] : 
                             (N180)? \nz.mem [3278] : 
                             (N182)? \nz.mem [3358] : 
                             (N184)? \nz.mem [3438] : 
                             (N186)? \nz.mem [3518] : 
                             (N188)? \nz.mem [3598] : 
                             (N190)? \nz.mem [3678] : 
                             (N192)? \nz.mem [3758] : 
                             (N194)? \nz.mem [3838] : 
                             (N196)? \nz.mem [3918] : 
                             (N198)? \nz.mem [3998] : 
                             (N200)? \nz.mem [4078] : 
                             (N202)? \nz.mem [4158] : 
                             (N204)? \nz.mem [4238] : 
                             (N206)? \nz.mem [4318] : 
                             (N208)? \nz.mem [4398] : 
                             (N210)? \nz.mem [4478] : 
                             (N212)? \nz.mem [4558] : 
                             (N214)? \nz.mem [4638] : 
                             (N216)? \nz.mem [4718] : 
                             (N218)? \nz.mem [4798] : 
                             (N220)? \nz.mem [4878] : 
                             (N222)? \nz.mem [4958] : 
                             (N224)? \nz.mem [5038] : 
                             (N226)? \nz.mem [5118] : 1'b0;
  assign \nz.data_out [77] = (N163)? \nz.mem [77] : 
                             (N165)? \nz.mem [157] : 
                             (N167)? \nz.mem [237] : 
                             (N169)? \nz.mem [317] : 
                             (N171)? \nz.mem [397] : 
                             (N173)? \nz.mem [477] : 
                             (N175)? \nz.mem [557] : 
                             (N177)? \nz.mem [637] : 
                             (N179)? \nz.mem [717] : 
                             (N181)? \nz.mem [797] : 
                             (N183)? \nz.mem [877] : 
                             (N185)? \nz.mem [957] : 
                             (N187)? \nz.mem [1037] : 
                             (N189)? \nz.mem [1117] : 
                             (N191)? \nz.mem [1197] : 
                             (N193)? \nz.mem [1277] : 
                             (N195)? \nz.mem [1357] : 
                             (N197)? \nz.mem [1437] : 
                             (N199)? \nz.mem [1517] : 
                             (N201)? \nz.mem [1597] : 
                             (N203)? \nz.mem [1677] : 
                             (N205)? \nz.mem [1757] : 
                             (N207)? \nz.mem [1837] : 
                             (N209)? \nz.mem [1917] : 
                             (N211)? \nz.mem [1997] : 
                             (N213)? \nz.mem [2077] : 
                             (N215)? \nz.mem [2157] : 
                             (N217)? \nz.mem [2237] : 
                             (N219)? \nz.mem [2317] : 
                             (N221)? \nz.mem [2397] : 
                             (N223)? \nz.mem [2477] : 
                             (N225)? \nz.mem [2557] : 
                             (N164)? \nz.mem [2637] : 
                             (N166)? \nz.mem [2717] : 
                             (N168)? \nz.mem [2797] : 
                             (N170)? \nz.mem [2877] : 
                             (N172)? \nz.mem [2957] : 
                             (N174)? \nz.mem [3037] : 
                             (N176)? \nz.mem [3117] : 
                             (N178)? \nz.mem [3197] : 
                             (N180)? \nz.mem [3277] : 
                             (N182)? \nz.mem [3357] : 
                             (N184)? \nz.mem [3437] : 
                             (N186)? \nz.mem [3517] : 
                             (N188)? \nz.mem [3597] : 
                             (N190)? \nz.mem [3677] : 
                             (N192)? \nz.mem [3757] : 
                             (N194)? \nz.mem [3837] : 
                             (N196)? \nz.mem [3917] : 
                             (N198)? \nz.mem [3997] : 
                             (N200)? \nz.mem [4077] : 
                             (N202)? \nz.mem [4157] : 
                             (N204)? \nz.mem [4237] : 
                             (N206)? \nz.mem [4317] : 
                             (N208)? \nz.mem [4397] : 
                             (N210)? \nz.mem [4477] : 
                             (N212)? \nz.mem [4557] : 
                             (N214)? \nz.mem [4637] : 
                             (N216)? \nz.mem [4717] : 
                             (N218)? \nz.mem [4797] : 
                             (N220)? \nz.mem [4877] : 
                             (N222)? \nz.mem [4957] : 
                             (N224)? \nz.mem [5037] : 
                             (N226)? \nz.mem [5117] : 1'b0;
  assign \nz.data_out [76] = (N163)? \nz.mem [76] : 
                             (N165)? \nz.mem [156] : 
                             (N167)? \nz.mem [236] : 
                             (N169)? \nz.mem [316] : 
                             (N171)? \nz.mem [396] : 
                             (N173)? \nz.mem [476] : 
                             (N175)? \nz.mem [556] : 
                             (N177)? \nz.mem [636] : 
                             (N179)? \nz.mem [716] : 
                             (N181)? \nz.mem [796] : 
                             (N183)? \nz.mem [876] : 
                             (N185)? \nz.mem [956] : 
                             (N187)? \nz.mem [1036] : 
                             (N189)? \nz.mem [1116] : 
                             (N191)? \nz.mem [1196] : 
                             (N193)? \nz.mem [1276] : 
                             (N195)? \nz.mem [1356] : 
                             (N197)? \nz.mem [1436] : 
                             (N199)? \nz.mem [1516] : 
                             (N201)? \nz.mem [1596] : 
                             (N203)? \nz.mem [1676] : 
                             (N205)? \nz.mem [1756] : 
                             (N207)? \nz.mem [1836] : 
                             (N209)? \nz.mem [1916] : 
                             (N211)? \nz.mem [1996] : 
                             (N213)? \nz.mem [2076] : 
                             (N215)? \nz.mem [2156] : 
                             (N217)? \nz.mem [2236] : 
                             (N219)? \nz.mem [2316] : 
                             (N221)? \nz.mem [2396] : 
                             (N223)? \nz.mem [2476] : 
                             (N225)? \nz.mem [2556] : 
                             (N164)? \nz.mem [2636] : 
                             (N166)? \nz.mem [2716] : 
                             (N168)? \nz.mem [2796] : 
                             (N170)? \nz.mem [2876] : 
                             (N172)? \nz.mem [2956] : 
                             (N174)? \nz.mem [3036] : 
                             (N176)? \nz.mem [3116] : 
                             (N178)? \nz.mem [3196] : 
                             (N180)? \nz.mem [3276] : 
                             (N182)? \nz.mem [3356] : 
                             (N184)? \nz.mem [3436] : 
                             (N186)? \nz.mem [3516] : 
                             (N188)? \nz.mem [3596] : 
                             (N190)? \nz.mem [3676] : 
                             (N192)? \nz.mem [3756] : 
                             (N194)? \nz.mem [3836] : 
                             (N196)? \nz.mem [3916] : 
                             (N198)? \nz.mem [3996] : 
                             (N200)? \nz.mem [4076] : 
                             (N202)? \nz.mem [4156] : 
                             (N204)? \nz.mem [4236] : 
                             (N206)? \nz.mem [4316] : 
                             (N208)? \nz.mem [4396] : 
                             (N210)? \nz.mem [4476] : 
                             (N212)? \nz.mem [4556] : 
                             (N214)? \nz.mem [4636] : 
                             (N216)? \nz.mem [4716] : 
                             (N218)? \nz.mem [4796] : 
                             (N220)? \nz.mem [4876] : 
                             (N222)? \nz.mem [4956] : 
                             (N224)? \nz.mem [5036] : 
                             (N226)? \nz.mem [5116] : 1'b0;
  assign \nz.data_out [75] = (N163)? \nz.mem [75] : 
                             (N165)? \nz.mem [155] : 
                             (N167)? \nz.mem [235] : 
                             (N169)? \nz.mem [315] : 
                             (N171)? \nz.mem [395] : 
                             (N173)? \nz.mem [475] : 
                             (N175)? \nz.mem [555] : 
                             (N177)? \nz.mem [635] : 
                             (N179)? \nz.mem [715] : 
                             (N181)? \nz.mem [795] : 
                             (N183)? \nz.mem [875] : 
                             (N185)? \nz.mem [955] : 
                             (N187)? \nz.mem [1035] : 
                             (N189)? \nz.mem [1115] : 
                             (N191)? \nz.mem [1195] : 
                             (N193)? \nz.mem [1275] : 
                             (N195)? \nz.mem [1355] : 
                             (N197)? \nz.mem [1435] : 
                             (N199)? \nz.mem [1515] : 
                             (N201)? \nz.mem [1595] : 
                             (N203)? \nz.mem [1675] : 
                             (N205)? \nz.mem [1755] : 
                             (N207)? \nz.mem [1835] : 
                             (N209)? \nz.mem [1915] : 
                             (N211)? \nz.mem [1995] : 
                             (N213)? \nz.mem [2075] : 
                             (N215)? \nz.mem [2155] : 
                             (N217)? \nz.mem [2235] : 
                             (N219)? \nz.mem [2315] : 
                             (N221)? \nz.mem [2395] : 
                             (N223)? \nz.mem [2475] : 
                             (N225)? \nz.mem [2555] : 
                             (N164)? \nz.mem [2635] : 
                             (N166)? \nz.mem [2715] : 
                             (N168)? \nz.mem [2795] : 
                             (N170)? \nz.mem [2875] : 
                             (N172)? \nz.mem [2955] : 
                             (N174)? \nz.mem [3035] : 
                             (N176)? \nz.mem [3115] : 
                             (N178)? \nz.mem [3195] : 
                             (N180)? \nz.mem [3275] : 
                             (N182)? \nz.mem [3355] : 
                             (N184)? \nz.mem [3435] : 
                             (N186)? \nz.mem [3515] : 
                             (N188)? \nz.mem [3595] : 
                             (N190)? \nz.mem [3675] : 
                             (N192)? \nz.mem [3755] : 
                             (N194)? \nz.mem [3835] : 
                             (N196)? \nz.mem [3915] : 
                             (N198)? \nz.mem [3995] : 
                             (N200)? \nz.mem [4075] : 
                             (N202)? \nz.mem [4155] : 
                             (N204)? \nz.mem [4235] : 
                             (N206)? \nz.mem [4315] : 
                             (N208)? \nz.mem [4395] : 
                             (N210)? \nz.mem [4475] : 
                             (N212)? \nz.mem [4555] : 
                             (N214)? \nz.mem [4635] : 
                             (N216)? \nz.mem [4715] : 
                             (N218)? \nz.mem [4795] : 
                             (N220)? \nz.mem [4875] : 
                             (N222)? \nz.mem [4955] : 
                             (N224)? \nz.mem [5035] : 
                             (N226)? \nz.mem [5115] : 1'b0;
  assign \nz.data_out [74] = (N163)? \nz.mem [74] : 
                             (N165)? \nz.mem [154] : 
                             (N167)? \nz.mem [234] : 
                             (N169)? \nz.mem [314] : 
                             (N171)? \nz.mem [394] : 
                             (N173)? \nz.mem [474] : 
                             (N175)? \nz.mem [554] : 
                             (N177)? \nz.mem [634] : 
                             (N179)? \nz.mem [714] : 
                             (N181)? \nz.mem [794] : 
                             (N183)? \nz.mem [874] : 
                             (N185)? \nz.mem [954] : 
                             (N187)? \nz.mem [1034] : 
                             (N189)? \nz.mem [1114] : 
                             (N191)? \nz.mem [1194] : 
                             (N193)? \nz.mem [1274] : 
                             (N195)? \nz.mem [1354] : 
                             (N197)? \nz.mem [1434] : 
                             (N199)? \nz.mem [1514] : 
                             (N201)? \nz.mem [1594] : 
                             (N203)? \nz.mem [1674] : 
                             (N205)? \nz.mem [1754] : 
                             (N207)? \nz.mem [1834] : 
                             (N209)? \nz.mem [1914] : 
                             (N211)? \nz.mem [1994] : 
                             (N213)? \nz.mem [2074] : 
                             (N215)? \nz.mem [2154] : 
                             (N217)? \nz.mem [2234] : 
                             (N219)? \nz.mem [2314] : 
                             (N221)? \nz.mem [2394] : 
                             (N223)? \nz.mem [2474] : 
                             (N225)? \nz.mem [2554] : 
                             (N164)? \nz.mem [2634] : 
                             (N166)? \nz.mem [2714] : 
                             (N168)? \nz.mem [2794] : 
                             (N170)? \nz.mem [2874] : 
                             (N172)? \nz.mem [2954] : 
                             (N174)? \nz.mem [3034] : 
                             (N176)? \nz.mem [3114] : 
                             (N178)? \nz.mem [3194] : 
                             (N180)? \nz.mem [3274] : 
                             (N182)? \nz.mem [3354] : 
                             (N184)? \nz.mem [3434] : 
                             (N186)? \nz.mem [3514] : 
                             (N188)? \nz.mem [3594] : 
                             (N190)? \nz.mem [3674] : 
                             (N192)? \nz.mem [3754] : 
                             (N194)? \nz.mem [3834] : 
                             (N196)? \nz.mem [3914] : 
                             (N198)? \nz.mem [3994] : 
                             (N200)? \nz.mem [4074] : 
                             (N202)? \nz.mem [4154] : 
                             (N204)? \nz.mem [4234] : 
                             (N206)? \nz.mem [4314] : 
                             (N208)? \nz.mem [4394] : 
                             (N210)? \nz.mem [4474] : 
                             (N212)? \nz.mem [4554] : 
                             (N214)? \nz.mem [4634] : 
                             (N216)? \nz.mem [4714] : 
                             (N218)? \nz.mem [4794] : 
                             (N220)? \nz.mem [4874] : 
                             (N222)? \nz.mem [4954] : 
                             (N224)? \nz.mem [5034] : 
                             (N226)? \nz.mem [5114] : 1'b0;
  assign \nz.data_out [73] = (N163)? \nz.mem [73] : 
                             (N165)? \nz.mem [153] : 
                             (N167)? \nz.mem [233] : 
                             (N169)? \nz.mem [313] : 
                             (N171)? \nz.mem [393] : 
                             (N173)? \nz.mem [473] : 
                             (N175)? \nz.mem [553] : 
                             (N177)? \nz.mem [633] : 
                             (N179)? \nz.mem [713] : 
                             (N181)? \nz.mem [793] : 
                             (N183)? \nz.mem [873] : 
                             (N185)? \nz.mem [953] : 
                             (N187)? \nz.mem [1033] : 
                             (N189)? \nz.mem [1113] : 
                             (N191)? \nz.mem [1193] : 
                             (N193)? \nz.mem [1273] : 
                             (N195)? \nz.mem [1353] : 
                             (N197)? \nz.mem [1433] : 
                             (N199)? \nz.mem [1513] : 
                             (N201)? \nz.mem [1593] : 
                             (N203)? \nz.mem [1673] : 
                             (N205)? \nz.mem [1753] : 
                             (N207)? \nz.mem [1833] : 
                             (N209)? \nz.mem [1913] : 
                             (N211)? \nz.mem [1993] : 
                             (N213)? \nz.mem [2073] : 
                             (N215)? \nz.mem [2153] : 
                             (N217)? \nz.mem [2233] : 
                             (N219)? \nz.mem [2313] : 
                             (N221)? \nz.mem [2393] : 
                             (N223)? \nz.mem [2473] : 
                             (N225)? \nz.mem [2553] : 
                             (N164)? \nz.mem [2633] : 
                             (N166)? \nz.mem [2713] : 
                             (N168)? \nz.mem [2793] : 
                             (N170)? \nz.mem [2873] : 
                             (N172)? \nz.mem [2953] : 
                             (N174)? \nz.mem [3033] : 
                             (N176)? \nz.mem [3113] : 
                             (N178)? \nz.mem [3193] : 
                             (N180)? \nz.mem [3273] : 
                             (N182)? \nz.mem [3353] : 
                             (N184)? \nz.mem [3433] : 
                             (N186)? \nz.mem [3513] : 
                             (N188)? \nz.mem [3593] : 
                             (N190)? \nz.mem [3673] : 
                             (N192)? \nz.mem [3753] : 
                             (N194)? \nz.mem [3833] : 
                             (N196)? \nz.mem [3913] : 
                             (N198)? \nz.mem [3993] : 
                             (N200)? \nz.mem [4073] : 
                             (N202)? \nz.mem [4153] : 
                             (N204)? \nz.mem [4233] : 
                             (N206)? \nz.mem [4313] : 
                             (N208)? \nz.mem [4393] : 
                             (N210)? \nz.mem [4473] : 
                             (N212)? \nz.mem [4553] : 
                             (N214)? \nz.mem [4633] : 
                             (N216)? \nz.mem [4713] : 
                             (N218)? \nz.mem [4793] : 
                             (N220)? \nz.mem [4873] : 
                             (N222)? \nz.mem [4953] : 
                             (N224)? \nz.mem [5033] : 
                             (N226)? \nz.mem [5113] : 1'b0;
  assign \nz.data_out [72] = (N163)? \nz.mem [72] : 
                             (N165)? \nz.mem [152] : 
                             (N167)? \nz.mem [232] : 
                             (N169)? \nz.mem [312] : 
                             (N171)? \nz.mem [392] : 
                             (N173)? \nz.mem [472] : 
                             (N175)? \nz.mem [552] : 
                             (N177)? \nz.mem [632] : 
                             (N179)? \nz.mem [712] : 
                             (N181)? \nz.mem [792] : 
                             (N183)? \nz.mem [872] : 
                             (N185)? \nz.mem [952] : 
                             (N187)? \nz.mem [1032] : 
                             (N189)? \nz.mem [1112] : 
                             (N191)? \nz.mem [1192] : 
                             (N193)? \nz.mem [1272] : 
                             (N195)? \nz.mem [1352] : 
                             (N197)? \nz.mem [1432] : 
                             (N199)? \nz.mem [1512] : 
                             (N201)? \nz.mem [1592] : 
                             (N203)? \nz.mem [1672] : 
                             (N205)? \nz.mem [1752] : 
                             (N207)? \nz.mem [1832] : 
                             (N209)? \nz.mem [1912] : 
                             (N211)? \nz.mem [1992] : 
                             (N213)? \nz.mem [2072] : 
                             (N215)? \nz.mem [2152] : 
                             (N217)? \nz.mem [2232] : 
                             (N219)? \nz.mem [2312] : 
                             (N221)? \nz.mem [2392] : 
                             (N223)? \nz.mem [2472] : 
                             (N225)? \nz.mem [2552] : 
                             (N164)? \nz.mem [2632] : 
                             (N166)? \nz.mem [2712] : 
                             (N168)? \nz.mem [2792] : 
                             (N170)? \nz.mem [2872] : 
                             (N172)? \nz.mem [2952] : 
                             (N174)? \nz.mem [3032] : 
                             (N176)? \nz.mem [3112] : 
                             (N178)? \nz.mem [3192] : 
                             (N180)? \nz.mem [3272] : 
                             (N182)? \nz.mem [3352] : 
                             (N184)? \nz.mem [3432] : 
                             (N186)? \nz.mem [3512] : 
                             (N188)? \nz.mem [3592] : 
                             (N190)? \nz.mem [3672] : 
                             (N192)? \nz.mem [3752] : 
                             (N194)? \nz.mem [3832] : 
                             (N196)? \nz.mem [3912] : 
                             (N198)? \nz.mem [3992] : 
                             (N200)? \nz.mem [4072] : 
                             (N202)? \nz.mem [4152] : 
                             (N204)? \nz.mem [4232] : 
                             (N206)? \nz.mem [4312] : 
                             (N208)? \nz.mem [4392] : 
                             (N210)? \nz.mem [4472] : 
                             (N212)? \nz.mem [4552] : 
                             (N214)? \nz.mem [4632] : 
                             (N216)? \nz.mem [4712] : 
                             (N218)? \nz.mem [4792] : 
                             (N220)? \nz.mem [4872] : 
                             (N222)? \nz.mem [4952] : 
                             (N224)? \nz.mem [5032] : 
                             (N226)? \nz.mem [5112] : 1'b0;
  assign \nz.data_out [71] = (N163)? \nz.mem [71] : 
                             (N165)? \nz.mem [151] : 
                             (N167)? \nz.mem [231] : 
                             (N169)? \nz.mem [311] : 
                             (N171)? \nz.mem [391] : 
                             (N173)? \nz.mem [471] : 
                             (N175)? \nz.mem [551] : 
                             (N177)? \nz.mem [631] : 
                             (N179)? \nz.mem [711] : 
                             (N181)? \nz.mem [791] : 
                             (N183)? \nz.mem [871] : 
                             (N185)? \nz.mem [951] : 
                             (N187)? \nz.mem [1031] : 
                             (N189)? \nz.mem [1111] : 
                             (N191)? \nz.mem [1191] : 
                             (N193)? \nz.mem [1271] : 
                             (N195)? \nz.mem [1351] : 
                             (N197)? \nz.mem [1431] : 
                             (N199)? \nz.mem [1511] : 
                             (N201)? \nz.mem [1591] : 
                             (N203)? \nz.mem [1671] : 
                             (N205)? \nz.mem [1751] : 
                             (N207)? \nz.mem [1831] : 
                             (N209)? \nz.mem [1911] : 
                             (N211)? \nz.mem [1991] : 
                             (N213)? \nz.mem [2071] : 
                             (N215)? \nz.mem [2151] : 
                             (N217)? \nz.mem [2231] : 
                             (N219)? \nz.mem [2311] : 
                             (N221)? \nz.mem [2391] : 
                             (N223)? \nz.mem [2471] : 
                             (N225)? \nz.mem [2551] : 
                             (N164)? \nz.mem [2631] : 
                             (N166)? \nz.mem [2711] : 
                             (N168)? \nz.mem [2791] : 
                             (N170)? \nz.mem [2871] : 
                             (N172)? \nz.mem [2951] : 
                             (N174)? \nz.mem [3031] : 
                             (N176)? \nz.mem [3111] : 
                             (N178)? \nz.mem [3191] : 
                             (N180)? \nz.mem [3271] : 
                             (N182)? \nz.mem [3351] : 
                             (N184)? \nz.mem [3431] : 
                             (N186)? \nz.mem [3511] : 
                             (N188)? \nz.mem [3591] : 
                             (N190)? \nz.mem [3671] : 
                             (N192)? \nz.mem [3751] : 
                             (N194)? \nz.mem [3831] : 
                             (N196)? \nz.mem [3911] : 
                             (N198)? \nz.mem [3991] : 
                             (N200)? \nz.mem [4071] : 
                             (N202)? \nz.mem [4151] : 
                             (N204)? \nz.mem [4231] : 
                             (N206)? \nz.mem [4311] : 
                             (N208)? \nz.mem [4391] : 
                             (N210)? \nz.mem [4471] : 
                             (N212)? \nz.mem [4551] : 
                             (N214)? \nz.mem [4631] : 
                             (N216)? \nz.mem [4711] : 
                             (N218)? \nz.mem [4791] : 
                             (N220)? \nz.mem [4871] : 
                             (N222)? \nz.mem [4951] : 
                             (N224)? \nz.mem [5031] : 
                             (N226)? \nz.mem [5111] : 1'b0;
  assign \nz.data_out [70] = (N163)? \nz.mem [70] : 
                             (N165)? \nz.mem [150] : 
                             (N167)? \nz.mem [230] : 
                             (N169)? \nz.mem [310] : 
                             (N171)? \nz.mem [390] : 
                             (N173)? \nz.mem [470] : 
                             (N175)? \nz.mem [550] : 
                             (N177)? \nz.mem [630] : 
                             (N179)? \nz.mem [710] : 
                             (N181)? \nz.mem [790] : 
                             (N183)? \nz.mem [870] : 
                             (N185)? \nz.mem [950] : 
                             (N187)? \nz.mem [1030] : 
                             (N189)? \nz.mem [1110] : 
                             (N191)? \nz.mem [1190] : 
                             (N193)? \nz.mem [1270] : 
                             (N195)? \nz.mem [1350] : 
                             (N197)? \nz.mem [1430] : 
                             (N199)? \nz.mem [1510] : 
                             (N201)? \nz.mem [1590] : 
                             (N203)? \nz.mem [1670] : 
                             (N205)? \nz.mem [1750] : 
                             (N207)? \nz.mem [1830] : 
                             (N209)? \nz.mem [1910] : 
                             (N211)? \nz.mem [1990] : 
                             (N213)? \nz.mem [2070] : 
                             (N215)? \nz.mem [2150] : 
                             (N217)? \nz.mem [2230] : 
                             (N219)? \nz.mem [2310] : 
                             (N221)? \nz.mem [2390] : 
                             (N223)? \nz.mem [2470] : 
                             (N225)? \nz.mem [2550] : 
                             (N164)? \nz.mem [2630] : 
                             (N166)? \nz.mem [2710] : 
                             (N168)? \nz.mem [2790] : 
                             (N170)? \nz.mem [2870] : 
                             (N172)? \nz.mem [2950] : 
                             (N174)? \nz.mem [3030] : 
                             (N176)? \nz.mem [3110] : 
                             (N178)? \nz.mem [3190] : 
                             (N180)? \nz.mem [3270] : 
                             (N182)? \nz.mem [3350] : 
                             (N184)? \nz.mem [3430] : 
                             (N186)? \nz.mem [3510] : 
                             (N188)? \nz.mem [3590] : 
                             (N190)? \nz.mem [3670] : 
                             (N192)? \nz.mem [3750] : 
                             (N194)? \nz.mem [3830] : 
                             (N196)? \nz.mem [3910] : 
                             (N198)? \nz.mem [3990] : 
                             (N200)? \nz.mem [4070] : 
                             (N202)? \nz.mem [4150] : 
                             (N204)? \nz.mem [4230] : 
                             (N206)? \nz.mem [4310] : 
                             (N208)? \nz.mem [4390] : 
                             (N210)? \nz.mem [4470] : 
                             (N212)? \nz.mem [4550] : 
                             (N214)? \nz.mem [4630] : 
                             (N216)? \nz.mem [4710] : 
                             (N218)? \nz.mem [4790] : 
                             (N220)? \nz.mem [4870] : 
                             (N222)? \nz.mem [4950] : 
                             (N224)? \nz.mem [5030] : 
                             (N226)? \nz.mem [5110] : 1'b0;
  assign \nz.data_out [69] = (N163)? \nz.mem [69] : 
                             (N165)? \nz.mem [149] : 
                             (N167)? \nz.mem [229] : 
                             (N169)? \nz.mem [309] : 
                             (N171)? \nz.mem [389] : 
                             (N173)? \nz.mem [469] : 
                             (N175)? \nz.mem [549] : 
                             (N177)? \nz.mem [629] : 
                             (N179)? \nz.mem [709] : 
                             (N181)? \nz.mem [789] : 
                             (N183)? \nz.mem [869] : 
                             (N185)? \nz.mem [949] : 
                             (N187)? \nz.mem [1029] : 
                             (N189)? \nz.mem [1109] : 
                             (N191)? \nz.mem [1189] : 
                             (N193)? \nz.mem [1269] : 
                             (N195)? \nz.mem [1349] : 
                             (N197)? \nz.mem [1429] : 
                             (N199)? \nz.mem [1509] : 
                             (N201)? \nz.mem [1589] : 
                             (N203)? \nz.mem [1669] : 
                             (N205)? \nz.mem [1749] : 
                             (N207)? \nz.mem [1829] : 
                             (N209)? \nz.mem [1909] : 
                             (N211)? \nz.mem [1989] : 
                             (N213)? \nz.mem [2069] : 
                             (N215)? \nz.mem [2149] : 
                             (N217)? \nz.mem [2229] : 
                             (N219)? \nz.mem [2309] : 
                             (N221)? \nz.mem [2389] : 
                             (N223)? \nz.mem [2469] : 
                             (N225)? \nz.mem [2549] : 
                             (N164)? \nz.mem [2629] : 
                             (N166)? \nz.mem [2709] : 
                             (N168)? \nz.mem [2789] : 
                             (N170)? \nz.mem [2869] : 
                             (N172)? \nz.mem [2949] : 
                             (N174)? \nz.mem [3029] : 
                             (N176)? \nz.mem [3109] : 
                             (N178)? \nz.mem [3189] : 
                             (N180)? \nz.mem [3269] : 
                             (N182)? \nz.mem [3349] : 
                             (N184)? \nz.mem [3429] : 
                             (N186)? \nz.mem [3509] : 
                             (N188)? \nz.mem [3589] : 
                             (N190)? \nz.mem [3669] : 
                             (N192)? \nz.mem [3749] : 
                             (N194)? \nz.mem [3829] : 
                             (N196)? \nz.mem [3909] : 
                             (N198)? \nz.mem [3989] : 
                             (N200)? \nz.mem [4069] : 
                             (N202)? \nz.mem [4149] : 
                             (N204)? \nz.mem [4229] : 
                             (N206)? \nz.mem [4309] : 
                             (N208)? \nz.mem [4389] : 
                             (N210)? \nz.mem [4469] : 
                             (N212)? \nz.mem [4549] : 
                             (N214)? \nz.mem [4629] : 
                             (N216)? \nz.mem [4709] : 
                             (N218)? \nz.mem [4789] : 
                             (N220)? \nz.mem [4869] : 
                             (N222)? \nz.mem [4949] : 
                             (N224)? \nz.mem [5029] : 
                             (N226)? \nz.mem [5109] : 1'b0;
  assign \nz.data_out [68] = (N163)? \nz.mem [68] : 
                             (N165)? \nz.mem [148] : 
                             (N167)? \nz.mem [228] : 
                             (N169)? \nz.mem [308] : 
                             (N171)? \nz.mem [388] : 
                             (N173)? \nz.mem [468] : 
                             (N175)? \nz.mem [548] : 
                             (N177)? \nz.mem [628] : 
                             (N179)? \nz.mem [708] : 
                             (N181)? \nz.mem [788] : 
                             (N183)? \nz.mem [868] : 
                             (N185)? \nz.mem [948] : 
                             (N187)? \nz.mem [1028] : 
                             (N189)? \nz.mem [1108] : 
                             (N191)? \nz.mem [1188] : 
                             (N193)? \nz.mem [1268] : 
                             (N195)? \nz.mem [1348] : 
                             (N197)? \nz.mem [1428] : 
                             (N199)? \nz.mem [1508] : 
                             (N201)? \nz.mem [1588] : 
                             (N203)? \nz.mem [1668] : 
                             (N205)? \nz.mem [1748] : 
                             (N207)? \nz.mem [1828] : 
                             (N209)? \nz.mem [1908] : 
                             (N211)? \nz.mem [1988] : 
                             (N213)? \nz.mem [2068] : 
                             (N215)? \nz.mem [2148] : 
                             (N217)? \nz.mem [2228] : 
                             (N219)? \nz.mem [2308] : 
                             (N221)? \nz.mem [2388] : 
                             (N223)? \nz.mem [2468] : 
                             (N225)? \nz.mem [2548] : 
                             (N164)? \nz.mem [2628] : 
                             (N166)? \nz.mem [2708] : 
                             (N168)? \nz.mem [2788] : 
                             (N170)? \nz.mem [2868] : 
                             (N172)? \nz.mem [2948] : 
                             (N174)? \nz.mem [3028] : 
                             (N176)? \nz.mem [3108] : 
                             (N178)? \nz.mem [3188] : 
                             (N180)? \nz.mem [3268] : 
                             (N182)? \nz.mem [3348] : 
                             (N184)? \nz.mem [3428] : 
                             (N186)? \nz.mem [3508] : 
                             (N188)? \nz.mem [3588] : 
                             (N190)? \nz.mem [3668] : 
                             (N192)? \nz.mem [3748] : 
                             (N194)? \nz.mem [3828] : 
                             (N196)? \nz.mem [3908] : 
                             (N198)? \nz.mem [3988] : 
                             (N200)? \nz.mem [4068] : 
                             (N202)? \nz.mem [4148] : 
                             (N204)? \nz.mem [4228] : 
                             (N206)? \nz.mem [4308] : 
                             (N208)? \nz.mem [4388] : 
                             (N210)? \nz.mem [4468] : 
                             (N212)? \nz.mem [4548] : 
                             (N214)? \nz.mem [4628] : 
                             (N216)? \nz.mem [4708] : 
                             (N218)? \nz.mem [4788] : 
                             (N220)? \nz.mem [4868] : 
                             (N222)? \nz.mem [4948] : 
                             (N224)? \nz.mem [5028] : 
                             (N226)? \nz.mem [5108] : 1'b0;
  assign \nz.data_out [67] = (N163)? \nz.mem [67] : 
                             (N165)? \nz.mem [147] : 
                             (N167)? \nz.mem [227] : 
                             (N169)? \nz.mem [307] : 
                             (N171)? \nz.mem [387] : 
                             (N173)? \nz.mem [467] : 
                             (N175)? \nz.mem [547] : 
                             (N177)? \nz.mem [627] : 
                             (N179)? \nz.mem [707] : 
                             (N181)? \nz.mem [787] : 
                             (N183)? \nz.mem [867] : 
                             (N185)? \nz.mem [947] : 
                             (N187)? \nz.mem [1027] : 
                             (N189)? \nz.mem [1107] : 
                             (N191)? \nz.mem [1187] : 
                             (N193)? \nz.mem [1267] : 
                             (N195)? \nz.mem [1347] : 
                             (N197)? \nz.mem [1427] : 
                             (N199)? \nz.mem [1507] : 
                             (N201)? \nz.mem [1587] : 
                             (N203)? \nz.mem [1667] : 
                             (N205)? \nz.mem [1747] : 
                             (N207)? \nz.mem [1827] : 
                             (N209)? \nz.mem [1907] : 
                             (N211)? \nz.mem [1987] : 
                             (N213)? \nz.mem [2067] : 
                             (N215)? \nz.mem [2147] : 
                             (N217)? \nz.mem [2227] : 
                             (N219)? \nz.mem [2307] : 
                             (N221)? \nz.mem [2387] : 
                             (N223)? \nz.mem [2467] : 
                             (N225)? \nz.mem [2547] : 
                             (N164)? \nz.mem [2627] : 
                             (N166)? \nz.mem [2707] : 
                             (N168)? \nz.mem [2787] : 
                             (N170)? \nz.mem [2867] : 
                             (N172)? \nz.mem [2947] : 
                             (N174)? \nz.mem [3027] : 
                             (N176)? \nz.mem [3107] : 
                             (N178)? \nz.mem [3187] : 
                             (N180)? \nz.mem [3267] : 
                             (N182)? \nz.mem [3347] : 
                             (N184)? \nz.mem [3427] : 
                             (N186)? \nz.mem [3507] : 
                             (N188)? \nz.mem [3587] : 
                             (N190)? \nz.mem [3667] : 
                             (N192)? \nz.mem [3747] : 
                             (N194)? \nz.mem [3827] : 
                             (N196)? \nz.mem [3907] : 
                             (N198)? \nz.mem [3987] : 
                             (N200)? \nz.mem [4067] : 
                             (N202)? \nz.mem [4147] : 
                             (N204)? \nz.mem [4227] : 
                             (N206)? \nz.mem [4307] : 
                             (N208)? \nz.mem [4387] : 
                             (N210)? \nz.mem [4467] : 
                             (N212)? \nz.mem [4547] : 
                             (N214)? \nz.mem [4627] : 
                             (N216)? \nz.mem [4707] : 
                             (N218)? \nz.mem [4787] : 
                             (N220)? \nz.mem [4867] : 
                             (N222)? \nz.mem [4947] : 
                             (N224)? \nz.mem [5027] : 
                             (N226)? \nz.mem [5107] : 1'b0;
  assign \nz.data_out [66] = (N163)? \nz.mem [66] : 
                             (N165)? \nz.mem [146] : 
                             (N167)? \nz.mem [226] : 
                             (N169)? \nz.mem [306] : 
                             (N171)? \nz.mem [386] : 
                             (N173)? \nz.mem [466] : 
                             (N175)? \nz.mem [546] : 
                             (N177)? \nz.mem [626] : 
                             (N179)? \nz.mem [706] : 
                             (N181)? \nz.mem [786] : 
                             (N183)? \nz.mem [866] : 
                             (N185)? \nz.mem [946] : 
                             (N187)? \nz.mem [1026] : 
                             (N189)? \nz.mem [1106] : 
                             (N191)? \nz.mem [1186] : 
                             (N193)? \nz.mem [1266] : 
                             (N195)? \nz.mem [1346] : 
                             (N197)? \nz.mem [1426] : 
                             (N199)? \nz.mem [1506] : 
                             (N201)? \nz.mem [1586] : 
                             (N203)? \nz.mem [1666] : 
                             (N205)? \nz.mem [1746] : 
                             (N207)? \nz.mem [1826] : 
                             (N209)? \nz.mem [1906] : 
                             (N211)? \nz.mem [1986] : 
                             (N213)? \nz.mem [2066] : 
                             (N215)? \nz.mem [2146] : 
                             (N217)? \nz.mem [2226] : 
                             (N219)? \nz.mem [2306] : 
                             (N221)? \nz.mem [2386] : 
                             (N223)? \nz.mem [2466] : 
                             (N225)? \nz.mem [2546] : 
                             (N164)? \nz.mem [2626] : 
                             (N166)? \nz.mem [2706] : 
                             (N168)? \nz.mem [2786] : 
                             (N170)? \nz.mem [2866] : 
                             (N172)? \nz.mem [2946] : 
                             (N174)? \nz.mem [3026] : 
                             (N176)? \nz.mem [3106] : 
                             (N178)? \nz.mem [3186] : 
                             (N180)? \nz.mem [3266] : 
                             (N182)? \nz.mem [3346] : 
                             (N184)? \nz.mem [3426] : 
                             (N186)? \nz.mem [3506] : 
                             (N188)? \nz.mem [3586] : 
                             (N190)? \nz.mem [3666] : 
                             (N192)? \nz.mem [3746] : 
                             (N194)? \nz.mem [3826] : 
                             (N196)? \nz.mem [3906] : 
                             (N198)? \nz.mem [3986] : 
                             (N200)? \nz.mem [4066] : 
                             (N202)? \nz.mem [4146] : 
                             (N204)? \nz.mem [4226] : 
                             (N206)? \nz.mem [4306] : 
                             (N208)? \nz.mem [4386] : 
                             (N210)? \nz.mem [4466] : 
                             (N212)? \nz.mem [4546] : 
                             (N214)? \nz.mem [4626] : 
                             (N216)? \nz.mem [4706] : 
                             (N218)? \nz.mem [4786] : 
                             (N220)? \nz.mem [4866] : 
                             (N222)? \nz.mem [4946] : 
                             (N224)? \nz.mem [5026] : 
                             (N226)? \nz.mem [5106] : 1'b0;
  assign \nz.data_out [65] = (N163)? \nz.mem [65] : 
                             (N165)? \nz.mem [145] : 
                             (N167)? \nz.mem [225] : 
                             (N169)? \nz.mem [305] : 
                             (N171)? \nz.mem [385] : 
                             (N173)? \nz.mem [465] : 
                             (N175)? \nz.mem [545] : 
                             (N177)? \nz.mem [625] : 
                             (N179)? \nz.mem [705] : 
                             (N181)? \nz.mem [785] : 
                             (N183)? \nz.mem [865] : 
                             (N185)? \nz.mem [945] : 
                             (N187)? \nz.mem [1025] : 
                             (N189)? \nz.mem [1105] : 
                             (N191)? \nz.mem [1185] : 
                             (N193)? \nz.mem [1265] : 
                             (N195)? \nz.mem [1345] : 
                             (N197)? \nz.mem [1425] : 
                             (N199)? \nz.mem [1505] : 
                             (N201)? \nz.mem [1585] : 
                             (N203)? \nz.mem [1665] : 
                             (N205)? \nz.mem [1745] : 
                             (N207)? \nz.mem [1825] : 
                             (N209)? \nz.mem [1905] : 
                             (N211)? \nz.mem [1985] : 
                             (N213)? \nz.mem [2065] : 
                             (N215)? \nz.mem [2145] : 
                             (N217)? \nz.mem [2225] : 
                             (N219)? \nz.mem [2305] : 
                             (N221)? \nz.mem [2385] : 
                             (N223)? \nz.mem [2465] : 
                             (N225)? \nz.mem [2545] : 
                             (N164)? \nz.mem [2625] : 
                             (N166)? \nz.mem [2705] : 
                             (N168)? \nz.mem [2785] : 
                             (N170)? \nz.mem [2865] : 
                             (N172)? \nz.mem [2945] : 
                             (N174)? \nz.mem [3025] : 
                             (N176)? \nz.mem [3105] : 
                             (N178)? \nz.mem [3185] : 
                             (N180)? \nz.mem [3265] : 
                             (N182)? \nz.mem [3345] : 
                             (N184)? \nz.mem [3425] : 
                             (N186)? \nz.mem [3505] : 
                             (N188)? \nz.mem [3585] : 
                             (N190)? \nz.mem [3665] : 
                             (N192)? \nz.mem [3745] : 
                             (N194)? \nz.mem [3825] : 
                             (N196)? \nz.mem [3905] : 
                             (N198)? \nz.mem [3985] : 
                             (N200)? \nz.mem [4065] : 
                             (N202)? \nz.mem [4145] : 
                             (N204)? \nz.mem [4225] : 
                             (N206)? \nz.mem [4305] : 
                             (N208)? \nz.mem [4385] : 
                             (N210)? \nz.mem [4465] : 
                             (N212)? \nz.mem [4545] : 
                             (N214)? \nz.mem [4625] : 
                             (N216)? \nz.mem [4705] : 
                             (N218)? \nz.mem [4785] : 
                             (N220)? \nz.mem [4865] : 
                             (N222)? \nz.mem [4945] : 
                             (N224)? \nz.mem [5025] : 
                             (N226)? \nz.mem [5105] : 1'b0;
  assign \nz.data_out [64] = (N163)? \nz.mem [64] : 
                             (N165)? \nz.mem [144] : 
                             (N167)? \nz.mem [224] : 
                             (N169)? \nz.mem [304] : 
                             (N171)? \nz.mem [384] : 
                             (N173)? \nz.mem [464] : 
                             (N175)? \nz.mem [544] : 
                             (N177)? \nz.mem [624] : 
                             (N179)? \nz.mem [704] : 
                             (N181)? \nz.mem [784] : 
                             (N183)? \nz.mem [864] : 
                             (N185)? \nz.mem [944] : 
                             (N187)? \nz.mem [1024] : 
                             (N189)? \nz.mem [1104] : 
                             (N191)? \nz.mem [1184] : 
                             (N193)? \nz.mem [1264] : 
                             (N195)? \nz.mem [1344] : 
                             (N197)? \nz.mem [1424] : 
                             (N199)? \nz.mem [1504] : 
                             (N201)? \nz.mem [1584] : 
                             (N203)? \nz.mem [1664] : 
                             (N205)? \nz.mem [1744] : 
                             (N207)? \nz.mem [1824] : 
                             (N209)? \nz.mem [1904] : 
                             (N211)? \nz.mem [1984] : 
                             (N213)? \nz.mem [2064] : 
                             (N215)? \nz.mem [2144] : 
                             (N217)? \nz.mem [2224] : 
                             (N219)? \nz.mem [2304] : 
                             (N221)? \nz.mem [2384] : 
                             (N223)? \nz.mem [2464] : 
                             (N225)? \nz.mem [2544] : 
                             (N164)? \nz.mem [2624] : 
                             (N166)? \nz.mem [2704] : 
                             (N168)? \nz.mem [2784] : 
                             (N170)? \nz.mem [2864] : 
                             (N172)? \nz.mem [2944] : 
                             (N174)? \nz.mem [3024] : 
                             (N176)? \nz.mem [3104] : 
                             (N178)? \nz.mem [3184] : 
                             (N180)? \nz.mem [3264] : 
                             (N182)? \nz.mem [3344] : 
                             (N184)? \nz.mem [3424] : 
                             (N186)? \nz.mem [3504] : 
                             (N188)? \nz.mem [3584] : 
                             (N190)? \nz.mem [3664] : 
                             (N192)? \nz.mem [3744] : 
                             (N194)? \nz.mem [3824] : 
                             (N196)? \nz.mem [3904] : 
                             (N198)? \nz.mem [3984] : 
                             (N200)? \nz.mem [4064] : 
                             (N202)? \nz.mem [4144] : 
                             (N204)? \nz.mem [4224] : 
                             (N206)? \nz.mem [4304] : 
                             (N208)? \nz.mem [4384] : 
                             (N210)? \nz.mem [4464] : 
                             (N212)? \nz.mem [4544] : 
                             (N214)? \nz.mem [4624] : 
                             (N216)? \nz.mem [4704] : 
                             (N218)? \nz.mem [4784] : 
                             (N220)? \nz.mem [4864] : 
                             (N222)? \nz.mem [4944] : 
                             (N224)? \nz.mem [5024] : 
                             (N226)? \nz.mem [5104] : 1'b0;
  assign \nz.data_out [63] = (N163)? \nz.mem [63] : 
                             (N165)? \nz.mem [143] : 
                             (N167)? \nz.mem [223] : 
                             (N169)? \nz.mem [303] : 
                             (N171)? \nz.mem [383] : 
                             (N173)? \nz.mem [463] : 
                             (N175)? \nz.mem [543] : 
                             (N177)? \nz.mem [623] : 
                             (N179)? \nz.mem [703] : 
                             (N181)? \nz.mem [783] : 
                             (N183)? \nz.mem [863] : 
                             (N185)? \nz.mem [943] : 
                             (N187)? \nz.mem [1023] : 
                             (N189)? \nz.mem [1103] : 
                             (N191)? \nz.mem [1183] : 
                             (N193)? \nz.mem [1263] : 
                             (N195)? \nz.mem [1343] : 
                             (N197)? \nz.mem [1423] : 
                             (N199)? \nz.mem [1503] : 
                             (N201)? \nz.mem [1583] : 
                             (N203)? \nz.mem [1663] : 
                             (N205)? \nz.mem [1743] : 
                             (N207)? \nz.mem [1823] : 
                             (N209)? \nz.mem [1903] : 
                             (N211)? \nz.mem [1983] : 
                             (N213)? \nz.mem [2063] : 
                             (N215)? \nz.mem [2143] : 
                             (N217)? \nz.mem [2223] : 
                             (N219)? \nz.mem [2303] : 
                             (N221)? \nz.mem [2383] : 
                             (N223)? \nz.mem [2463] : 
                             (N225)? \nz.mem [2543] : 
                             (N164)? \nz.mem [2623] : 
                             (N166)? \nz.mem [2703] : 
                             (N168)? \nz.mem [2783] : 
                             (N170)? \nz.mem [2863] : 
                             (N172)? \nz.mem [2943] : 
                             (N174)? \nz.mem [3023] : 
                             (N176)? \nz.mem [3103] : 
                             (N178)? \nz.mem [3183] : 
                             (N180)? \nz.mem [3263] : 
                             (N182)? \nz.mem [3343] : 
                             (N184)? \nz.mem [3423] : 
                             (N186)? \nz.mem [3503] : 
                             (N188)? \nz.mem [3583] : 
                             (N190)? \nz.mem [3663] : 
                             (N192)? \nz.mem [3743] : 
                             (N194)? \nz.mem [3823] : 
                             (N196)? \nz.mem [3903] : 
                             (N198)? \nz.mem [3983] : 
                             (N200)? \nz.mem [4063] : 
                             (N202)? \nz.mem [4143] : 
                             (N204)? \nz.mem [4223] : 
                             (N206)? \nz.mem [4303] : 
                             (N208)? \nz.mem [4383] : 
                             (N210)? \nz.mem [4463] : 
                             (N212)? \nz.mem [4543] : 
                             (N214)? \nz.mem [4623] : 
                             (N216)? \nz.mem [4703] : 
                             (N218)? \nz.mem [4783] : 
                             (N220)? \nz.mem [4863] : 
                             (N222)? \nz.mem [4943] : 
                             (N224)? \nz.mem [5023] : 
                             (N226)? \nz.mem [5103] : 1'b0;
  assign \nz.data_out [62] = (N163)? \nz.mem [62] : 
                             (N165)? \nz.mem [142] : 
                             (N167)? \nz.mem [222] : 
                             (N169)? \nz.mem [302] : 
                             (N171)? \nz.mem [382] : 
                             (N173)? \nz.mem [462] : 
                             (N175)? \nz.mem [542] : 
                             (N177)? \nz.mem [622] : 
                             (N179)? \nz.mem [702] : 
                             (N181)? \nz.mem [782] : 
                             (N183)? \nz.mem [862] : 
                             (N185)? \nz.mem [942] : 
                             (N187)? \nz.mem [1022] : 
                             (N189)? \nz.mem [1102] : 
                             (N191)? \nz.mem [1182] : 
                             (N193)? \nz.mem [1262] : 
                             (N195)? \nz.mem [1342] : 
                             (N197)? \nz.mem [1422] : 
                             (N199)? \nz.mem [1502] : 
                             (N201)? \nz.mem [1582] : 
                             (N203)? \nz.mem [1662] : 
                             (N205)? \nz.mem [1742] : 
                             (N207)? \nz.mem [1822] : 
                             (N209)? \nz.mem [1902] : 
                             (N211)? \nz.mem [1982] : 
                             (N213)? \nz.mem [2062] : 
                             (N215)? \nz.mem [2142] : 
                             (N217)? \nz.mem [2222] : 
                             (N219)? \nz.mem [2302] : 
                             (N221)? \nz.mem [2382] : 
                             (N223)? \nz.mem [2462] : 
                             (N225)? \nz.mem [2542] : 
                             (N164)? \nz.mem [2622] : 
                             (N166)? \nz.mem [2702] : 
                             (N168)? \nz.mem [2782] : 
                             (N170)? \nz.mem [2862] : 
                             (N172)? \nz.mem [2942] : 
                             (N174)? \nz.mem [3022] : 
                             (N176)? \nz.mem [3102] : 
                             (N178)? \nz.mem [3182] : 
                             (N180)? \nz.mem [3262] : 
                             (N182)? \nz.mem [3342] : 
                             (N184)? \nz.mem [3422] : 
                             (N186)? \nz.mem [3502] : 
                             (N188)? \nz.mem [3582] : 
                             (N190)? \nz.mem [3662] : 
                             (N192)? \nz.mem [3742] : 
                             (N194)? \nz.mem [3822] : 
                             (N196)? \nz.mem [3902] : 
                             (N198)? \nz.mem [3982] : 
                             (N200)? \nz.mem [4062] : 
                             (N202)? \nz.mem [4142] : 
                             (N204)? \nz.mem [4222] : 
                             (N206)? \nz.mem [4302] : 
                             (N208)? \nz.mem [4382] : 
                             (N210)? \nz.mem [4462] : 
                             (N212)? \nz.mem [4542] : 
                             (N214)? \nz.mem [4622] : 
                             (N216)? \nz.mem [4702] : 
                             (N218)? \nz.mem [4782] : 
                             (N220)? \nz.mem [4862] : 
                             (N222)? \nz.mem [4942] : 
                             (N224)? \nz.mem [5022] : 
                             (N226)? \nz.mem [5102] : 1'b0;
  assign \nz.data_out [61] = (N163)? \nz.mem [61] : 
                             (N165)? \nz.mem [141] : 
                             (N167)? \nz.mem [221] : 
                             (N169)? \nz.mem [301] : 
                             (N171)? \nz.mem [381] : 
                             (N173)? \nz.mem [461] : 
                             (N175)? \nz.mem [541] : 
                             (N177)? \nz.mem [621] : 
                             (N179)? \nz.mem [701] : 
                             (N181)? \nz.mem [781] : 
                             (N183)? \nz.mem [861] : 
                             (N185)? \nz.mem [941] : 
                             (N187)? \nz.mem [1021] : 
                             (N189)? \nz.mem [1101] : 
                             (N191)? \nz.mem [1181] : 
                             (N193)? \nz.mem [1261] : 
                             (N195)? \nz.mem [1341] : 
                             (N197)? \nz.mem [1421] : 
                             (N199)? \nz.mem [1501] : 
                             (N201)? \nz.mem [1581] : 
                             (N203)? \nz.mem [1661] : 
                             (N205)? \nz.mem [1741] : 
                             (N207)? \nz.mem [1821] : 
                             (N209)? \nz.mem [1901] : 
                             (N211)? \nz.mem [1981] : 
                             (N213)? \nz.mem [2061] : 
                             (N215)? \nz.mem [2141] : 
                             (N217)? \nz.mem [2221] : 
                             (N219)? \nz.mem [2301] : 
                             (N221)? \nz.mem [2381] : 
                             (N223)? \nz.mem [2461] : 
                             (N225)? \nz.mem [2541] : 
                             (N164)? \nz.mem [2621] : 
                             (N166)? \nz.mem [2701] : 
                             (N168)? \nz.mem [2781] : 
                             (N170)? \nz.mem [2861] : 
                             (N172)? \nz.mem [2941] : 
                             (N174)? \nz.mem [3021] : 
                             (N176)? \nz.mem [3101] : 
                             (N178)? \nz.mem [3181] : 
                             (N180)? \nz.mem [3261] : 
                             (N182)? \nz.mem [3341] : 
                             (N184)? \nz.mem [3421] : 
                             (N186)? \nz.mem [3501] : 
                             (N188)? \nz.mem [3581] : 
                             (N190)? \nz.mem [3661] : 
                             (N192)? \nz.mem [3741] : 
                             (N194)? \nz.mem [3821] : 
                             (N196)? \nz.mem [3901] : 
                             (N198)? \nz.mem [3981] : 
                             (N200)? \nz.mem [4061] : 
                             (N202)? \nz.mem [4141] : 
                             (N204)? \nz.mem [4221] : 
                             (N206)? \nz.mem [4301] : 
                             (N208)? \nz.mem [4381] : 
                             (N210)? \nz.mem [4461] : 
                             (N212)? \nz.mem [4541] : 
                             (N214)? \nz.mem [4621] : 
                             (N216)? \nz.mem [4701] : 
                             (N218)? \nz.mem [4781] : 
                             (N220)? \nz.mem [4861] : 
                             (N222)? \nz.mem [4941] : 
                             (N224)? \nz.mem [5021] : 
                             (N226)? \nz.mem [5101] : 1'b0;
  assign \nz.data_out [60] = (N163)? \nz.mem [60] : 
                             (N165)? \nz.mem [140] : 
                             (N167)? \nz.mem [220] : 
                             (N169)? \nz.mem [300] : 
                             (N171)? \nz.mem [380] : 
                             (N173)? \nz.mem [460] : 
                             (N175)? \nz.mem [540] : 
                             (N177)? \nz.mem [620] : 
                             (N179)? \nz.mem [700] : 
                             (N181)? \nz.mem [780] : 
                             (N183)? \nz.mem [860] : 
                             (N185)? \nz.mem [940] : 
                             (N187)? \nz.mem [1020] : 
                             (N189)? \nz.mem [1100] : 
                             (N191)? \nz.mem [1180] : 
                             (N193)? \nz.mem [1260] : 
                             (N195)? \nz.mem [1340] : 
                             (N197)? \nz.mem [1420] : 
                             (N199)? \nz.mem [1500] : 
                             (N201)? \nz.mem [1580] : 
                             (N203)? \nz.mem [1660] : 
                             (N205)? \nz.mem [1740] : 
                             (N207)? \nz.mem [1820] : 
                             (N209)? \nz.mem [1900] : 
                             (N211)? \nz.mem [1980] : 
                             (N213)? \nz.mem [2060] : 
                             (N215)? \nz.mem [2140] : 
                             (N217)? \nz.mem [2220] : 
                             (N219)? \nz.mem [2300] : 
                             (N221)? \nz.mem [2380] : 
                             (N223)? \nz.mem [2460] : 
                             (N225)? \nz.mem [2540] : 
                             (N164)? \nz.mem [2620] : 
                             (N166)? \nz.mem [2700] : 
                             (N168)? \nz.mem [2780] : 
                             (N170)? \nz.mem [2860] : 
                             (N172)? \nz.mem [2940] : 
                             (N174)? \nz.mem [3020] : 
                             (N176)? \nz.mem [3100] : 
                             (N178)? \nz.mem [3180] : 
                             (N180)? \nz.mem [3260] : 
                             (N182)? \nz.mem [3340] : 
                             (N184)? \nz.mem [3420] : 
                             (N186)? \nz.mem [3500] : 
                             (N188)? \nz.mem [3580] : 
                             (N190)? \nz.mem [3660] : 
                             (N192)? \nz.mem [3740] : 
                             (N194)? \nz.mem [3820] : 
                             (N196)? \nz.mem [3900] : 
                             (N198)? \nz.mem [3980] : 
                             (N200)? \nz.mem [4060] : 
                             (N202)? \nz.mem [4140] : 
                             (N204)? \nz.mem [4220] : 
                             (N206)? \nz.mem [4300] : 
                             (N208)? \nz.mem [4380] : 
                             (N210)? \nz.mem [4460] : 
                             (N212)? \nz.mem [4540] : 
                             (N214)? \nz.mem [4620] : 
                             (N216)? \nz.mem [4700] : 
                             (N218)? \nz.mem [4780] : 
                             (N220)? \nz.mem [4860] : 
                             (N222)? \nz.mem [4940] : 
                             (N224)? \nz.mem [5020] : 
                             (N226)? \nz.mem [5100] : 1'b0;
  assign \nz.data_out [59] = (N163)? \nz.mem [59] : 
                             (N165)? \nz.mem [139] : 
                             (N167)? \nz.mem [219] : 
                             (N169)? \nz.mem [299] : 
                             (N171)? \nz.mem [379] : 
                             (N173)? \nz.mem [459] : 
                             (N175)? \nz.mem [539] : 
                             (N177)? \nz.mem [619] : 
                             (N179)? \nz.mem [699] : 
                             (N181)? \nz.mem [779] : 
                             (N183)? \nz.mem [859] : 
                             (N185)? \nz.mem [939] : 
                             (N187)? \nz.mem [1019] : 
                             (N189)? \nz.mem [1099] : 
                             (N191)? \nz.mem [1179] : 
                             (N193)? \nz.mem [1259] : 
                             (N195)? \nz.mem [1339] : 
                             (N197)? \nz.mem [1419] : 
                             (N199)? \nz.mem [1499] : 
                             (N201)? \nz.mem [1579] : 
                             (N203)? \nz.mem [1659] : 
                             (N205)? \nz.mem [1739] : 
                             (N207)? \nz.mem [1819] : 
                             (N209)? \nz.mem [1899] : 
                             (N211)? \nz.mem [1979] : 
                             (N213)? \nz.mem [2059] : 
                             (N215)? \nz.mem [2139] : 
                             (N217)? \nz.mem [2219] : 
                             (N219)? \nz.mem [2299] : 
                             (N221)? \nz.mem [2379] : 
                             (N223)? \nz.mem [2459] : 
                             (N225)? \nz.mem [2539] : 
                             (N164)? \nz.mem [2619] : 
                             (N166)? \nz.mem [2699] : 
                             (N168)? \nz.mem [2779] : 
                             (N170)? \nz.mem [2859] : 
                             (N172)? \nz.mem [2939] : 
                             (N174)? \nz.mem [3019] : 
                             (N176)? \nz.mem [3099] : 
                             (N178)? \nz.mem [3179] : 
                             (N180)? \nz.mem [3259] : 
                             (N182)? \nz.mem [3339] : 
                             (N184)? \nz.mem [3419] : 
                             (N186)? \nz.mem [3499] : 
                             (N188)? \nz.mem [3579] : 
                             (N190)? \nz.mem [3659] : 
                             (N192)? \nz.mem [3739] : 
                             (N194)? \nz.mem [3819] : 
                             (N196)? \nz.mem [3899] : 
                             (N198)? \nz.mem [3979] : 
                             (N200)? \nz.mem [4059] : 
                             (N202)? \nz.mem [4139] : 
                             (N204)? \nz.mem [4219] : 
                             (N206)? \nz.mem [4299] : 
                             (N208)? \nz.mem [4379] : 
                             (N210)? \nz.mem [4459] : 
                             (N212)? \nz.mem [4539] : 
                             (N214)? \nz.mem [4619] : 
                             (N216)? \nz.mem [4699] : 
                             (N218)? \nz.mem [4779] : 
                             (N220)? \nz.mem [4859] : 
                             (N222)? \nz.mem [4939] : 
                             (N224)? \nz.mem [5019] : 
                             (N226)? \nz.mem [5099] : 1'b0;
  assign \nz.data_out [58] = (N163)? \nz.mem [58] : 
                             (N165)? \nz.mem [138] : 
                             (N167)? \nz.mem [218] : 
                             (N169)? \nz.mem [298] : 
                             (N171)? \nz.mem [378] : 
                             (N173)? \nz.mem [458] : 
                             (N175)? \nz.mem [538] : 
                             (N177)? \nz.mem [618] : 
                             (N179)? \nz.mem [698] : 
                             (N181)? \nz.mem [778] : 
                             (N183)? \nz.mem [858] : 
                             (N185)? \nz.mem [938] : 
                             (N187)? \nz.mem [1018] : 
                             (N189)? \nz.mem [1098] : 
                             (N191)? \nz.mem [1178] : 
                             (N193)? \nz.mem [1258] : 
                             (N195)? \nz.mem [1338] : 
                             (N197)? \nz.mem [1418] : 
                             (N199)? \nz.mem [1498] : 
                             (N201)? \nz.mem [1578] : 
                             (N203)? \nz.mem [1658] : 
                             (N205)? \nz.mem [1738] : 
                             (N207)? \nz.mem [1818] : 
                             (N209)? \nz.mem [1898] : 
                             (N211)? \nz.mem [1978] : 
                             (N213)? \nz.mem [2058] : 
                             (N215)? \nz.mem [2138] : 
                             (N217)? \nz.mem [2218] : 
                             (N219)? \nz.mem [2298] : 
                             (N221)? \nz.mem [2378] : 
                             (N223)? \nz.mem [2458] : 
                             (N225)? \nz.mem [2538] : 
                             (N164)? \nz.mem [2618] : 
                             (N166)? \nz.mem [2698] : 
                             (N168)? \nz.mem [2778] : 
                             (N170)? \nz.mem [2858] : 
                             (N172)? \nz.mem [2938] : 
                             (N174)? \nz.mem [3018] : 
                             (N176)? \nz.mem [3098] : 
                             (N178)? \nz.mem [3178] : 
                             (N180)? \nz.mem [3258] : 
                             (N182)? \nz.mem [3338] : 
                             (N184)? \nz.mem [3418] : 
                             (N186)? \nz.mem [3498] : 
                             (N188)? \nz.mem [3578] : 
                             (N190)? \nz.mem [3658] : 
                             (N192)? \nz.mem [3738] : 
                             (N194)? \nz.mem [3818] : 
                             (N196)? \nz.mem [3898] : 
                             (N198)? \nz.mem [3978] : 
                             (N200)? \nz.mem [4058] : 
                             (N202)? \nz.mem [4138] : 
                             (N204)? \nz.mem [4218] : 
                             (N206)? \nz.mem [4298] : 
                             (N208)? \nz.mem [4378] : 
                             (N210)? \nz.mem [4458] : 
                             (N212)? \nz.mem [4538] : 
                             (N214)? \nz.mem [4618] : 
                             (N216)? \nz.mem [4698] : 
                             (N218)? \nz.mem [4778] : 
                             (N220)? \nz.mem [4858] : 
                             (N222)? \nz.mem [4938] : 
                             (N224)? \nz.mem [5018] : 
                             (N226)? \nz.mem [5098] : 1'b0;
  assign \nz.data_out [57] = (N163)? \nz.mem [57] : 
                             (N165)? \nz.mem [137] : 
                             (N167)? \nz.mem [217] : 
                             (N169)? \nz.mem [297] : 
                             (N171)? \nz.mem [377] : 
                             (N173)? \nz.mem [457] : 
                             (N175)? \nz.mem [537] : 
                             (N177)? \nz.mem [617] : 
                             (N179)? \nz.mem [697] : 
                             (N181)? \nz.mem [777] : 
                             (N183)? \nz.mem [857] : 
                             (N185)? \nz.mem [937] : 
                             (N187)? \nz.mem [1017] : 
                             (N189)? \nz.mem [1097] : 
                             (N191)? \nz.mem [1177] : 
                             (N193)? \nz.mem [1257] : 
                             (N195)? \nz.mem [1337] : 
                             (N197)? \nz.mem [1417] : 
                             (N199)? \nz.mem [1497] : 
                             (N201)? \nz.mem [1577] : 
                             (N203)? \nz.mem [1657] : 
                             (N205)? \nz.mem [1737] : 
                             (N207)? \nz.mem [1817] : 
                             (N209)? \nz.mem [1897] : 
                             (N211)? \nz.mem [1977] : 
                             (N213)? \nz.mem [2057] : 
                             (N215)? \nz.mem [2137] : 
                             (N217)? \nz.mem [2217] : 
                             (N219)? \nz.mem [2297] : 
                             (N221)? \nz.mem [2377] : 
                             (N223)? \nz.mem [2457] : 
                             (N225)? \nz.mem [2537] : 
                             (N164)? \nz.mem [2617] : 
                             (N166)? \nz.mem [2697] : 
                             (N168)? \nz.mem [2777] : 
                             (N170)? \nz.mem [2857] : 
                             (N172)? \nz.mem [2937] : 
                             (N174)? \nz.mem [3017] : 
                             (N176)? \nz.mem [3097] : 
                             (N178)? \nz.mem [3177] : 
                             (N180)? \nz.mem [3257] : 
                             (N182)? \nz.mem [3337] : 
                             (N184)? \nz.mem [3417] : 
                             (N186)? \nz.mem [3497] : 
                             (N188)? \nz.mem [3577] : 
                             (N190)? \nz.mem [3657] : 
                             (N192)? \nz.mem [3737] : 
                             (N194)? \nz.mem [3817] : 
                             (N196)? \nz.mem [3897] : 
                             (N198)? \nz.mem [3977] : 
                             (N200)? \nz.mem [4057] : 
                             (N202)? \nz.mem [4137] : 
                             (N204)? \nz.mem [4217] : 
                             (N206)? \nz.mem [4297] : 
                             (N208)? \nz.mem [4377] : 
                             (N210)? \nz.mem [4457] : 
                             (N212)? \nz.mem [4537] : 
                             (N214)? \nz.mem [4617] : 
                             (N216)? \nz.mem [4697] : 
                             (N218)? \nz.mem [4777] : 
                             (N220)? \nz.mem [4857] : 
                             (N222)? \nz.mem [4937] : 
                             (N224)? \nz.mem [5017] : 
                             (N226)? \nz.mem [5097] : 1'b0;
  assign \nz.data_out [56] = (N163)? \nz.mem [56] : 
                             (N165)? \nz.mem [136] : 
                             (N167)? \nz.mem [216] : 
                             (N169)? \nz.mem [296] : 
                             (N171)? \nz.mem [376] : 
                             (N173)? \nz.mem [456] : 
                             (N175)? \nz.mem [536] : 
                             (N177)? \nz.mem [616] : 
                             (N179)? \nz.mem [696] : 
                             (N181)? \nz.mem [776] : 
                             (N183)? \nz.mem [856] : 
                             (N185)? \nz.mem [936] : 
                             (N187)? \nz.mem [1016] : 
                             (N189)? \nz.mem [1096] : 
                             (N191)? \nz.mem [1176] : 
                             (N193)? \nz.mem [1256] : 
                             (N195)? \nz.mem [1336] : 
                             (N197)? \nz.mem [1416] : 
                             (N199)? \nz.mem [1496] : 
                             (N201)? \nz.mem [1576] : 
                             (N203)? \nz.mem [1656] : 
                             (N205)? \nz.mem [1736] : 
                             (N207)? \nz.mem [1816] : 
                             (N209)? \nz.mem [1896] : 
                             (N211)? \nz.mem [1976] : 
                             (N213)? \nz.mem [2056] : 
                             (N215)? \nz.mem [2136] : 
                             (N217)? \nz.mem [2216] : 
                             (N219)? \nz.mem [2296] : 
                             (N221)? \nz.mem [2376] : 
                             (N223)? \nz.mem [2456] : 
                             (N225)? \nz.mem [2536] : 
                             (N164)? \nz.mem [2616] : 
                             (N166)? \nz.mem [2696] : 
                             (N168)? \nz.mem [2776] : 
                             (N170)? \nz.mem [2856] : 
                             (N172)? \nz.mem [2936] : 
                             (N174)? \nz.mem [3016] : 
                             (N176)? \nz.mem [3096] : 
                             (N178)? \nz.mem [3176] : 
                             (N180)? \nz.mem [3256] : 
                             (N182)? \nz.mem [3336] : 
                             (N184)? \nz.mem [3416] : 
                             (N186)? \nz.mem [3496] : 
                             (N188)? \nz.mem [3576] : 
                             (N190)? \nz.mem [3656] : 
                             (N192)? \nz.mem [3736] : 
                             (N194)? \nz.mem [3816] : 
                             (N196)? \nz.mem [3896] : 
                             (N198)? \nz.mem [3976] : 
                             (N200)? \nz.mem [4056] : 
                             (N202)? \nz.mem [4136] : 
                             (N204)? \nz.mem [4216] : 
                             (N206)? \nz.mem [4296] : 
                             (N208)? \nz.mem [4376] : 
                             (N210)? \nz.mem [4456] : 
                             (N212)? \nz.mem [4536] : 
                             (N214)? \nz.mem [4616] : 
                             (N216)? \nz.mem [4696] : 
                             (N218)? \nz.mem [4776] : 
                             (N220)? \nz.mem [4856] : 
                             (N222)? \nz.mem [4936] : 
                             (N224)? \nz.mem [5016] : 
                             (N226)? \nz.mem [5096] : 1'b0;
  assign \nz.data_out [55] = (N163)? \nz.mem [55] : 
                             (N165)? \nz.mem [135] : 
                             (N167)? \nz.mem [215] : 
                             (N169)? \nz.mem [295] : 
                             (N171)? \nz.mem [375] : 
                             (N173)? \nz.mem [455] : 
                             (N175)? \nz.mem [535] : 
                             (N177)? \nz.mem [615] : 
                             (N179)? \nz.mem [695] : 
                             (N181)? \nz.mem [775] : 
                             (N183)? \nz.mem [855] : 
                             (N185)? \nz.mem [935] : 
                             (N187)? \nz.mem [1015] : 
                             (N189)? \nz.mem [1095] : 
                             (N191)? \nz.mem [1175] : 
                             (N193)? \nz.mem [1255] : 
                             (N195)? \nz.mem [1335] : 
                             (N197)? \nz.mem [1415] : 
                             (N199)? \nz.mem [1495] : 
                             (N201)? \nz.mem [1575] : 
                             (N203)? \nz.mem [1655] : 
                             (N205)? \nz.mem [1735] : 
                             (N207)? \nz.mem [1815] : 
                             (N209)? \nz.mem [1895] : 
                             (N211)? \nz.mem [1975] : 
                             (N213)? \nz.mem [2055] : 
                             (N215)? \nz.mem [2135] : 
                             (N217)? \nz.mem [2215] : 
                             (N219)? \nz.mem [2295] : 
                             (N221)? \nz.mem [2375] : 
                             (N223)? \nz.mem [2455] : 
                             (N225)? \nz.mem [2535] : 
                             (N164)? \nz.mem [2615] : 
                             (N166)? \nz.mem [2695] : 
                             (N168)? \nz.mem [2775] : 
                             (N170)? \nz.mem [2855] : 
                             (N172)? \nz.mem [2935] : 
                             (N174)? \nz.mem [3015] : 
                             (N176)? \nz.mem [3095] : 
                             (N178)? \nz.mem [3175] : 
                             (N180)? \nz.mem [3255] : 
                             (N182)? \nz.mem [3335] : 
                             (N184)? \nz.mem [3415] : 
                             (N186)? \nz.mem [3495] : 
                             (N188)? \nz.mem [3575] : 
                             (N190)? \nz.mem [3655] : 
                             (N192)? \nz.mem [3735] : 
                             (N194)? \nz.mem [3815] : 
                             (N196)? \nz.mem [3895] : 
                             (N198)? \nz.mem [3975] : 
                             (N200)? \nz.mem [4055] : 
                             (N202)? \nz.mem [4135] : 
                             (N204)? \nz.mem [4215] : 
                             (N206)? \nz.mem [4295] : 
                             (N208)? \nz.mem [4375] : 
                             (N210)? \nz.mem [4455] : 
                             (N212)? \nz.mem [4535] : 
                             (N214)? \nz.mem [4615] : 
                             (N216)? \nz.mem [4695] : 
                             (N218)? \nz.mem [4775] : 
                             (N220)? \nz.mem [4855] : 
                             (N222)? \nz.mem [4935] : 
                             (N224)? \nz.mem [5015] : 
                             (N226)? \nz.mem [5095] : 1'b0;
  assign \nz.data_out [54] = (N163)? \nz.mem [54] : 
                             (N165)? \nz.mem [134] : 
                             (N167)? \nz.mem [214] : 
                             (N169)? \nz.mem [294] : 
                             (N171)? \nz.mem [374] : 
                             (N173)? \nz.mem [454] : 
                             (N175)? \nz.mem [534] : 
                             (N177)? \nz.mem [614] : 
                             (N179)? \nz.mem [694] : 
                             (N181)? \nz.mem [774] : 
                             (N183)? \nz.mem [854] : 
                             (N185)? \nz.mem [934] : 
                             (N187)? \nz.mem [1014] : 
                             (N189)? \nz.mem [1094] : 
                             (N191)? \nz.mem [1174] : 
                             (N193)? \nz.mem [1254] : 
                             (N195)? \nz.mem [1334] : 
                             (N197)? \nz.mem [1414] : 
                             (N199)? \nz.mem [1494] : 
                             (N201)? \nz.mem [1574] : 
                             (N203)? \nz.mem [1654] : 
                             (N205)? \nz.mem [1734] : 
                             (N207)? \nz.mem [1814] : 
                             (N209)? \nz.mem [1894] : 
                             (N211)? \nz.mem [1974] : 
                             (N213)? \nz.mem [2054] : 
                             (N215)? \nz.mem [2134] : 
                             (N217)? \nz.mem [2214] : 
                             (N219)? \nz.mem [2294] : 
                             (N221)? \nz.mem [2374] : 
                             (N223)? \nz.mem [2454] : 
                             (N225)? \nz.mem [2534] : 
                             (N164)? \nz.mem [2614] : 
                             (N166)? \nz.mem [2694] : 
                             (N168)? \nz.mem [2774] : 
                             (N170)? \nz.mem [2854] : 
                             (N172)? \nz.mem [2934] : 
                             (N174)? \nz.mem [3014] : 
                             (N176)? \nz.mem [3094] : 
                             (N178)? \nz.mem [3174] : 
                             (N180)? \nz.mem [3254] : 
                             (N182)? \nz.mem [3334] : 
                             (N184)? \nz.mem [3414] : 
                             (N186)? \nz.mem [3494] : 
                             (N188)? \nz.mem [3574] : 
                             (N190)? \nz.mem [3654] : 
                             (N192)? \nz.mem [3734] : 
                             (N194)? \nz.mem [3814] : 
                             (N196)? \nz.mem [3894] : 
                             (N198)? \nz.mem [3974] : 
                             (N200)? \nz.mem [4054] : 
                             (N202)? \nz.mem [4134] : 
                             (N204)? \nz.mem [4214] : 
                             (N206)? \nz.mem [4294] : 
                             (N208)? \nz.mem [4374] : 
                             (N210)? \nz.mem [4454] : 
                             (N212)? \nz.mem [4534] : 
                             (N214)? \nz.mem [4614] : 
                             (N216)? \nz.mem [4694] : 
                             (N218)? \nz.mem [4774] : 
                             (N220)? \nz.mem [4854] : 
                             (N222)? \nz.mem [4934] : 
                             (N224)? \nz.mem [5014] : 
                             (N226)? \nz.mem [5094] : 1'b0;
  assign \nz.data_out [53] = (N163)? \nz.mem [53] : 
                             (N165)? \nz.mem [133] : 
                             (N167)? \nz.mem [213] : 
                             (N169)? \nz.mem [293] : 
                             (N171)? \nz.mem [373] : 
                             (N173)? \nz.mem [453] : 
                             (N175)? \nz.mem [533] : 
                             (N177)? \nz.mem [613] : 
                             (N179)? \nz.mem [693] : 
                             (N181)? \nz.mem [773] : 
                             (N183)? \nz.mem [853] : 
                             (N185)? \nz.mem [933] : 
                             (N187)? \nz.mem [1013] : 
                             (N189)? \nz.mem [1093] : 
                             (N191)? \nz.mem [1173] : 
                             (N193)? \nz.mem [1253] : 
                             (N195)? \nz.mem [1333] : 
                             (N197)? \nz.mem [1413] : 
                             (N199)? \nz.mem [1493] : 
                             (N201)? \nz.mem [1573] : 
                             (N203)? \nz.mem [1653] : 
                             (N205)? \nz.mem [1733] : 
                             (N207)? \nz.mem [1813] : 
                             (N209)? \nz.mem [1893] : 
                             (N211)? \nz.mem [1973] : 
                             (N213)? \nz.mem [2053] : 
                             (N215)? \nz.mem [2133] : 
                             (N217)? \nz.mem [2213] : 
                             (N219)? \nz.mem [2293] : 
                             (N221)? \nz.mem [2373] : 
                             (N223)? \nz.mem [2453] : 
                             (N225)? \nz.mem [2533] : 
                             (N164)? \nz.mem [2613] : 
                             (N166)? \nz.mem [2693] : 
                             (N168)? \nz.mem [2773] : 
                             (N170)? \nz.mem [2853] : 
                             (N172)? \nz.mem [2933] : 
                             (N174)? \nz.mem [3013] : 
                             (N176)? \nz.mem [3093] : 
                             (N178)? \nz.mem [3173] : 
                             (N180)? \nz.mem [3253] : 
                             (N182)? \nz.mem [3333] : 
                             (N184)? \nz.mem [3413] : 
                             (N186)? \nz.mem [3493] : 
                             (N188)? \nz.mem [3573] : 
                             (N190)? \nz.mem [3653] : 
                             (N192)? \nz.mem [3733] : 
                             (N194)? \nz.mem [3813] : 
                             (N196)? \nz.mem [3893] : 
                             (N198)? \nz.mem [3973] : 
                             (N200)? \nz.mem [4053] : 
                             (N202)? \nz.mem [4133] : 
                             (N204)? \nz.mem [4213] : 
                             (N206)? \nz.mem [4293] : 
                             (N208)? \nz.mem [4373] : 
                             (N210)? \nz.mem [4453] : 
                             (N212)? \nz.mem [4533] : 
                             (N214)? \nz.mem [4613] : 
                             (N216)? \nz.mem [4693] : 
                             (N218)? \nz.mem [4773] : 
                             (N220)? \nz.mem [4853] : 
                             (N222)? \nz.mem [4933] : 
                             (N224)? \nz.mem [5013] : 
                             (N226)? \nz.mem [5093] : 1'b0;
  assign \nz.data_out [52] = (N163)? \nz.mem [52] : 
                             (N165)? \nz.mem [132] : 
                             (N167)? \nz.mem [212] : 
                             (N169)? \nz.mem [292] : 
                             (N171)? \nz.mem [372] : 
                             (N173)? \nz.mem [452] : 
                             (N175)? \nz.mem [532] : 
                             (N177)? \nz.mem [612] : 
                             (N179)? \nz.mem [692] : 
                             (N181)? \nz.mem [772] : 
                             (N183)? \nz.mem [852] : 
                             (N185)? \nz.mem [932] : 
                             (N187)? \nz.mem [1012] : 
                             (N189)? \nz.mem [1092] : 
                             (N191)? \nz.mem [1172] : 
                             (N193)? \nz.mem [1252] : 
                             (N195)? \nz.mem [1332] : 
                             (N197)? \nz.mem [1412] : 
                             (N199)? \nz.mem [1492] : 
                             (N201)? \nz.mem [1572] : 
                             (N203)? \nz.mem [1652] : 
                             (N205)? \nz.mem [1732] : 
                             (N207)? \nz.mem [1812] : 
                             (N209)? \nz.mem [1892] : 
                             (N211)? \nz.mem [1972] : 
                             (N213)? \nz.mem [2052] : 
                             (N215)? \nz.mem [2132] : 
                             (N217)? \nz.mem [2212] : 
                             (N219)? \nz.mem [2292] : 
                             (N221)? \nz.mem [2372] : 
                             (N223)? \nz.mem [2452] : 
                             (N225)? \nz.mem [2532] : 
                             (N164)? \nz.mem [2612] : 
                             (N166)? \nz.mem [2692] : 
                             (N168)? \nz.mem [2772] : 
                             (N170)? \nz.mem [2852] : 
                             (N172)? \nz.mem [2932] : 
                             (N174)? \nz.mem [3012] : 
                             (N176)? \nz.mem [3092] : 
                             (N178)? \nz.mem [3172] : 
                             (N180)? \nz.mem [3252] : 
                             (N182)? \nz.mem [3332] : 
                             (N184)? \nz.mem [3412] : 
                             (N186)? \nz.mem [3492] : 
                             (N188)? \nz.mem [3572] : 
                             (N190)? \nz.mem [3652] : 
                             (N192)? \nz.mem [3732] : 
                             (N194)? \nz.mem [3812] : 
                             (N196)? \nz.mem [3892] : 
                             (N198)? \nz.mem [3972] : 
                             (N200)? \nz.mem [4052] : 
                             (N202)? \nz.mem [4132] : 
                             (N204)? \nz.mem [4212] : 
                             (N206)? \nz.mem [4292] : 
                             (N208)? \nz.mem [4372] : 
                             (N210)? \nz.mem [4452] : 
                             (N212)? \nz.mem [4532] : 
                             (N214)? \nz.mem [4612] : 
                             (N216)? \nz.mem [4692] : 
                             (N218)? \nz.mem [4772] : 
                             (N220)? \nz.mem [4852] : 
                             (N222)? \nz.mem [4932] : 
                             (N224)? \nz.mem [5012] : 
                             (N226)? \nz.mem [5092] : 1'b0;
  assign \nz.data_out [51] = (N163)? \nz.mem [51] : 
                             (N165)? \nz.mem [131] : 
                             (N167)? \nz.mem [211] : 
                             (N169)? \nz.mem [291] : 
                             (N171)? \nz.mem [371] : 
                             (N173)? \nz.mem [451] : 
                             (N175)? \nz.mem [531] : 
                             (N177)? \nz.mem [611] : 
                             (N179)? \nz.mem [691] : 
                             (N181)? \nz.mem [771] : 
                             (N183)? \nz.mem [851] : 
                             (N185)? \nz.mem [931] : 
                             (N187)? \nz.mem [1011] : 
                             (N189)? \nz.mem [1091] : 
                             (N191)? \nz.mem [1171] : 
                             (N193)? \nz.mem [1251] : 
                             (N195)? \nz.mem [1331] : 
                             (N197)? \nz.mem [1411] : 
                             (N199)? \nz.mem [1491] : 
                             (N201)? \nz.mem [1571] : 
                             (N203)? \nz.mem [1651] : 
                             (N205)? \nz.mem [1731] : 
                             (N207)? \nz.mem [1811] : 
                             (N209)? \nz.mem [1891] : 
                             (N211)? \nz.mem [1971] : 
                             (N213)? \nz.mem [2051] : 
                             (N215)? \nz.mem [2131] : 
                             (N217)? \nz.mem [2211] : 
                             (N219)? \nz.mem [2291] : 
                             (N221)? \nz.mem [2371] : 
                             (N223)? \nz.mem [2451] : 
                             (N225)? \nz.mem [2531] : 
                             (N164)? \nz.mem [2611] : 
                             (N166)? \nz.mem [2691] : 
                             (N168)? \nz.mem [2771] : 
                             (N170)? \nz.mem [2851] : 
                             (N172)? \nz.mem [2931] : 
                             (N174)? \nz.mem [3011] : 
                             (N176)? \nz.mem [3091] : 
                             (N178)? \nz.mem [3171] : 
                             (N180)? \nz.mem [3251] : 
                             (N182)? \nz.mem [3331] : 
                             (N184)? \nz.mem [3411] : 
                             (N186)? \nz.mem [3491] : 
                             (N188)? \nz.mem [3571] : 
                             (N190)? \nz.mem [3651] : 
                             (N192)? \nz.mem [3731] : 
                             (N194)? \nz.mem [3811] : 
                             (N196)? \nz.mem [3891] : 
                             (N198)? \nz.mem [3971] : 
                             (N200)? \nz.mem [4051] : 
                             (N202)? \nz.mem [4131] : 
                             (N204)? \nz.mem [4211] : 
                             (N206)? \nz.mem [4291] : 
                             (N208)? \nz.mem [4371] : 
                             (N210)? \nz.mem [4451] : 
                             (N212)? \nz.mem [4531] : 
                             (N214)? \nz.mem [4611] : 
                             (N216)? \nz.mem [4691] : 
                             (N218)? \nz.mem [4771] : 
                             (N220)? \nz.mem [4851] : 
                             (N222)? \nz.mem [4931] : 
                             (N224)? \nz.mem [5011] : 
                             (N226)? \nz.mem [5091] : 1'b0;
  assign \nz.data_out [50] = (N163)? \nz.mem [50] : 
                             (N165)? \nz.mem [130] : 
                             (N167)? \nz.mem [210] : 
                             (N169)? \nz.mem [290] : 
                             (N171)? \nz.mem [370] : 
                             (N173)? \nz.mem [450] : 
                             (N175)? \nz.mem [530] : 
                             (N177)? \nz.mem [610] : 
                             (N179)? \nz.mem [690] : 
                             (N181)? \nz.mem [770] : 
                             (N183)? \nz.mem [850] : 
                             (N185)? \nz.mem [930] : 
                             (N187)? \nz.mem [1010] : 
                             (N189)? \nz.mem [1090] : 
                             (N191)? \nz.mem [1170] : 
                             (N193)? \nz.mem [1250] : 
                             (N195)? \nz.mem [1330] : 
                             (N197)? \nz.mem [1410] : 
                             (N199)? \nz.mem [1490] : 
                             (N201)? \nz.mem [1570] : 
                             (N203)? \nz.mem [1650] : 
                             (N205)? \nz.mem [1730] : 
                             (N207)? \nz.mem [1810] : 
                             (N209)? \nz.mem [1890] : 
                             (N211)? \nz.mem [1970] : 
                             (N213)? \nz.mem [2050] : 
                             (N215)? \nz.mem [2130] : 
                             (N217)? \nz.mem [2210] : 
                             (N219)? \nz.mem [2290] : 
                             (N221)? \nz.mem [2370] : 
                             (N223)? \nz.mem [2450] : 
                             (N225)? \nz.mem [2530] : 
                             (N164)? \nz.mem [2610] : 
                             (N166)? \nz.mem [2690] : 
                             (N168)? \nz.mem [2770] : 
                             (N170)? \nz.mem [2850] : 
                             (N172)? \nz.mem [2930] : 
                             (N174)? \nz.mem [3010] : 
                             (N176)? \nz.mem [3090] : 
                             (N178)? \nz.mem [3170] : 
                             (N180)? \nz.mem [3250] : 
                             (N182)? \nz.mem [3330] : 
                             (N184)? \nz.mem [3410] : 
                             (N186)? \nz.mem [3490] : 
                             (N188)? \nz.mem [3570] : 
                             (N190)? \nz.mem [3650] : 
                             (N192)? \nz.mem [3730] : 
                             (N194)? \nz.mem [3810] : 
                             (N196)? \nz.mem [3890] : 
                             (N198)? \nz.mem [3970] : 
                             (N200)? \nz.mem [4050] : 
                             (N202)? \nz.mem [4130] : 
                             (N204)? \nz.mem [4210] : 
                             (N206)? \nz.mem [4290] : 
                             (N208)? \nz.mem [4370] : 
                             (N210)? \nz.mem [4450] : 
                             (N212)? \nz.mem [4530] : 
                             (N214)? \nz.mem [4610] : 
                             (N216)? \nz.mem [4690] : 
                             (N218)? \nz.mem [4770] : 
                             (N220)? \nz.mem [4850] : 
                             (N222)? \nz.mem [4930] : 
                             (N224)? \nz.mem [5010] : 
                             (N226)? \nz.mem [5090] : 1'b0;
  assign \nz.data_out [49] = (N163)? \nz.mem [49] : 
                             (N165)? \nz.mem [129] : 
                             (N167)? \nz.mem [209] : 
                             (N169)? \nz.mem [289] : 
                             (N171)? \nz.mem [369] : 
                             (N173)? \nz.mem [449] : 
                             (N175)? \nz.mem [529] : 
                             (N177)? \nz.mem [609] : 
                             (N179)? \nz.mem [689] : 
                             (N181)? \nz.mem [769] : 
                             (N183)? \nz.mem [849] : 
                             (N185)? \nz.mem [929] : 
                             (N187)? \nz.mem [1009] : 
                             (N189)? \nz.mem [1089] : 
                             (N191)? \nz.mem [1169] : 
                             (N193)? \nz.mem [1249] : 
                             (N195)? \nz.mem [1329] : 
                             (N197)? \nz.mem [1409] : 
                             (N199)? \nz.mem [1489] : 
                             (N201)? \nz.mem [1569] : 
                             (N203)? \nz.mem [1649] : 
                             (N205)? \nz.mem [1729] : 
                             (N207)? \nz.mem [1809] : 
                             (N209)? \nz.mem [1889] : 
                             (N211)? \nz.mem [1969] : 
                             (N213)? \nz.mem [2049] : 
                             (N215)? \nz.mem [2129] : 
                             (N217)? \nz.mem [2209] : 
                             (N219)? \nz.mem [2289] : 
                             (N221)? \nz.mem [2369] : 
                             (N223)? \nz.mem [2449] : 
                             (N225)? \nz.mem [2529] : 
                             (N164)? \nz.mem [2609] : 
                             (N166)? \nz.mem [2689] : 
                             (N168)? \nz.mem [2769] : 
                             (N170)? \nz.mem [2849] : 
                             (N172)? \nz.mem [2929] : 
                             (N174)? \nz.mem [3009] : 
                             (N176)? \nz.mem [3089] : 
                             (N178)? \nz.mem [3169] : 
                             (N180)? \nz.mem [3249] : 
                             (N182)? \nz.mem [3329] : 
                             (N184)? \nz.mem [3409] : 
                             (N186)? \nz.mem [3489] : 
                             (N188)? \nz.mem [3569] : 
                             (N190)? \nz.mem [3649] : 
                             (N192)? \nz.mem [3729] : 
                             (N194)? \nz.mem [3809] : 
                             (N196)? \nz.mem [3889] : 
                             (N198)? \nz.mem [3969] : 
                             (N200)? \nz.mem [4049] : 
                             (N202)? \nz.mem [4129] : 
                             (N204)? \nz.mem [4209] : 
                             (N206)? \nz.mem [4289] : 
                             (N208)? \nz.mem [4369] : 
                             (N210)? \nz.mem [4449] : 
                             (N212)? \nz.mem [4529] : 
                             (N214)? \nz.mem [4609] : 
                             (N216)? \nz.mem [4689] : 
                             (N218)? \nz.mem [4769] : 
                             (N220)? \nz.mem [4849] : 
                             (N222)? \nz.mem [4929] : 
                             (N224)? \nz.mem [5009] : 
                             (N226)? \nz.mem [5089] : 1'b0;
  assign \nz.data_out [48] = (N163)? \nz.mem [48] : 
                             (N165)? \nz.mem [128] : 
                             (N167)? \nz.mem [208] : 
                             (N169)? \nz.mem [288] : 
                             (N171)? \nz.mem [368] : 
                             (N173)? \nz.mem [448] : 
                             (N175)? \nz.mem [528] : 
                             (N177)? \nz.mem [608] : 
                             (N179)? \nz.mem [688] : 
                             (N181)? \nz.mem [768] : 
                             (N183)? \nz.mem [848] : 
                             (N185)? \nz.mem [928] : 
                             (N187)? \nz.mem [1008] : 
                             (N189)? \nz.mem [1088] : 
                             (N191)? \nz.mem [1168] : 
                             (N193)? \nz.mem [1248] : 
                             (N195)? \nz.mem [1328] : 
                             (N197)? \nz.mem [1408] : 
                             (N199)? \nz.mem [1488] : 
                             (N201)? \nz.mem [1568] : 
                             (N203)? \nz.mem [1648] : 
                             (N205)? \nz.mem [1728] : 
                             (N207)? \nz.mem [1808] : 
                             (N209)? \nz.mem [1888] : 
                             (N211)? \nz.mem [1968] : 
                             (N213)? \nz.mem [2048] : 
                             (N215)? \nz.mem [2128] : 
                             (N217)? \nz.mem [2208] : 
                             (N219)? \nz.mem [2288] : 
                             (N221)? \nz.mem [2368] : 
                             (N223)? \nz.mem [2448] : 
                             (N225)? \nz.mem [2528] : 
                             (N164)? \nz.mem [2608] : 
                             (N166)? \nz.mem [2688] : 
                             (N168)? \nz.mem [2768] : 
                             (N170)? \nz.mem [2848] : 
                             (N172)? \nz.mem [2928] : 
                             (N174)? \nz.mem [3008] : 
                             (N176)? \nz.mem [3088] : 
                             (N178)? \nz.mem [3168] : 
                             (N180)? \nz.mem [3248] : 
                             (N182)? \nz.mem [3328] : 
                             (N184)? \nz.mem [3408] : 
                             (N186)? \nz.mem [3488] : 
                             (N188)? \nz.mem [3568] : 
                             (N190)? \nz.mem [3648] : 
                             (N192)? \nz.mem [3728] : 
                             (N194)? \nz.mem [3808] : 
                             (N196)? \nz.mem [3888] : 
                             (N198)? \nz.mem [3968] : 
                             (N200)? \nz.mem [4048] : 
                             (N202)? \nz.mem [4128] : 
                             (N204)? \nz.mem [4208] : 
                             (N206)? \nz.mem [4288] : 
                             (N208)? \nz.mem [4368] : 
                             (N210)? \nz.mem [4448] : 
                             (N212)? \nz.mem [4528] : 
                             (N214)? \nz.mem [4608] : 
                             (N216)? \nz.mem [4688] : 
                             (N218)? \nz.mem [4768] : 
                             (N220)? \nz.mem [4848] : 
                             (N222)? \nz.mem [4928] : 
                             (N224)? \nz.mem [5008] : 
                             (N226)? \nz.mem [5088] : 1'b0;
  assign \nz.data_out [47] = (N163)? \nz.mem [47] : 
                             (N165)? \nz.mem [127] : 
                             (N167)? \nz.mem [207] : 
                             (N169)? \nz.mem [287] : 
                             (N171)? \nz.mem [367] : 
                             (N173)? \nz.mem [447] : 
                             (N175)? \nz.mem [527] : 
                             (N177)? \nz.mem [607] : 
                             (N179)? \nz.mem [687] : 
                             (N181)? \nz.mem [767] : 
                             (N183)? \nz.mem [847] : 
                             (N185)? \nz.mem [927] : 
                             (N187)? \nz.mem [1007] : 
                             (N189)? \nz.mem [1087] : 
                             (N191)? \nz.mem [1167] : 
                             (N193)? \nz.mem [1247] : 
                             (N195)? \nz.mem [1327] : 
                             (N197)? \nz.mem [1407] : 
                             (N199)? \nz.mem [1487] : 
                             (N201)? \nz.mem [1567] : 
                             (N203)? \nz.mem [1647] : 
                             (N205)? \nz.mem [1727] : 
                             (N207)? \nz.mem [1807] : 
                             (N209)? \nz.mem [1887] : 
                             (N211)? \nz.mem [1967] : 
                             (N213)? \nz.mem [2047] : 
                             (N215)? \nz.mem [2127] : 
                             (N217)? \nz.mem [2207] : 
                             (N219)? \nz.mem [2287] : 
                             (N221)? \nz.mem [2367] : 
                             (N223)? \nz.mem [2447] : 
                             (N225)? \nz.mem [2527] : 
                             (N164)? \nz.mem [2607] : 
                             (N166)? \nz.mem [2687] : 
                             (N168)? \nz.mem [2767] : 
                             (N170)? \nz.mem [2847] : 
                             (N172)? \nz.mem [2927] : 
                             (N174)? \nz.mem [3007] : 
                             (N176)? \nz.mem [3087] : 
                             (N178)? \nz.mem [3167] : 
                             (N180)? \nz.mem [3247] : 
                             (N182)? \nz.mem [3327] : 
                             (N184)? \nz.mem [3407] : 
                             (N186)? \nz.mem [3487] : 
                             (N188)? \nz.mem [3567] : 
                             (N190)? \nz.mem [3647] : 
                             (N192)? \nz.mem [3727] : 
                             (N194)? \nz.mem [3807] : 
                             (N196)? \nz.mem [3887] : 
                             (N198)? \nz.mem [3967] : 
                             (N200)? \nz.mem [4047] : 
                             (N202)? \nz.mem [4127] : 
                             (N204)? \nz.mem [4207] : 
                             (N206)? \nz.mem [4287] : 
                             (N208)? \nz.mem [4367] : 
                             (N210)? \nz.mem [4447] : 
                             (N212)? \nz.mem [4527] : 
                             (N214)? \nz.mem [4607] : 
                             (N216)? \nz.mem [4687] : 
                             (N218)? \nz.mem [4767] : 
                             (N220)? \nz.mem [4847] : 
                             (N222)? \nz.mem [4927] : 
                             (N224)? \nz.mem [5007] : 
                             (N226)? \nz.mem [5087] : 1'b0;
  assign \nz.data_out [46] = (N163)? \nz.mem [46] : 
                             (N165)? \nz.mem [126] : 
                             (N167)? \nz.mem [206] : 
                             (N169)? \nz.mem [286] : 
                             (N171)? \nz.mem [366] : 
                             (N173)? \nz.mem [446] : 
                             (N175)? \nz.mem [526] : 
                             (N177)? \nz.mem [606] : 
                             (N179)? \nz.mem [686] : 
                             (N181)? \nz.mem [766] : 
                             (N183)? \nz.mem [846] : 
                             (N185)? \nz.mem [926] : 
                             (N187)? \nz.mem [1006] : 
                             (N189)? \nz.mem [1086] : 
                             (N191)? \nz.mem [1166] : 
                             (N193)? \nz.mem [1246] : 
                             (N195)? \nz.mem [1326] : 
                             (N197)? \nz.mem [1406] : 
                             (N199)? \nz.mem [1486] : 
                             (N201)? \nz.mem [1566] : 
                             (N203)? \nz.mem [1646] : 
                             (N205)? \nz.mem [1726] : 
                             (N207)? \nz.mem [1806] : 
                             (N209)? \nz.mem [1886] : 
                             (N211)? \nz.mem [1966] : 
                             (N213)? \nz.mem [2046] : 
                             (N215)? \nz.mem [2126] : 
                             (N217)? \nz.mem [2206] : 
                             (N219)? \nz.mem [2286] : 
                             (N221)? \nz.mem [2366] : 
                             (N223)? \nz.mem [2446] : 
                             (N225)? \nz.mem [2526] : 
                             (N164)? \nz.mem [2606] : 
                             (N166)? \nz.mem [2686] : 
                             (N168)? \nz.mem [2766] : 
                             (N170)? \nz.mem [2846] : 
                             (N172)? \nz.mem [2926] : 
                             (N174)? \nz.mem [3006] : 
                             (N176)? \nz.mem [3086] : 
                             (N178)? \nz.mem [3166] : 
                             (N180)? \nz.mem [3246] : 
                             (N182)? \nz.mem [3326] : 
                             (N184)? \nz.mem [3406] : 
                             (N186)? \nz.mem [3486] : 
                             (N188)? \nz.mem [3566] : 
                             (N190)? \nz.mem [3646] : 
                             (N192)? \nz.mem [3726] : 
                             (N194)? \nz.mem [3806] : 
                             (N196)? \nz.mem [3886] : 
                             (N198)? \nz.mem [3966] : 
                             (N200)? \nz.mem [4046] : 
                             (N202)? \nz.mem [4126] : 
                             (N204)? \nz.mem [4206] : 
                             (N206)? \nz.mem [4286] : 
                             (N208)? \nz.mem [4366] : 
                             (N210)? \nz.mem [4446] : 
                             (N212)? \nz.mem [4526] : 
                             (N214)? \nz.mem [4606] : 
                             (N216)? \nz.mem [4686] : 
                             (N218)? \nz.mem [4766] : 
                             (N220)? \nz.mem [4846] : 
                             (N222)? \nz.mem [4926] : 
                             (N224)? \nz.mem [5006] : 
                             (N226)? \nz.mem [5086] : 1'b0;
  assign \nz.data_out [45] = (N163)? \nz.mem [45] : 
                             (N165)? \nz.mem [125] : 
                             (N167)? \nz.mem [205] : 
                             (N169)? \nz.mem [285] : 
                             (N171)? \nz.mem [365] : 
                             (N173)? \nz.mem [445] : 
                             (N175)? \nz.mem [525] : 
                             (N177)? \nz.mem [605] : 
                             (N179)? \nz.mem [685] : 
                             (N181)? \nz.mem [765] : 
                             (N183)? \nz.mem [845] : 
                             (N185)? \nz.mem [925] : 
                             (N187)? \nz.mem [1005] : 
                             (N189)? \nz.mem [1085] : 
                             (N191)? \nz.mem [1165] : 
                             (N193)? \nz.mem [1245] : 
                             (N195)? \nz.mem [1325] : 
                             (N197)? \nz.mem [1405] : 
                             (N199)? \nz.mem [1485] : 
                             (N201)? \nz.mem [1565] : 
                             (N203)? \nz.mem [1645] : 
                             (N205)? \nz.mem [1725] : 
                             (N207)? \nz.mem [1805] : 
                             (N209)? \nz.mem [1885] : 
                             (N211)? \nz.mem [1965] : 
                             (N213)? \nz.mem [2045] : 
                             (N215)? \nz.mem [2125] : 
                             (N217)? \nz.mem [2205] : 
                             (N219)? \nz.mem [2285] : 
                             (N221)? \nz.mem [2365] : 
                             (N223)? \nz.mem [2445] : 
                             (N225)? \nz.mem [2525] : 
                             (N164)? \nz.mem [2605] : 
                             (N166)? \nz.mem [2685] : 
                             (N168)? \nz.mem [2765] : 
                             (N170)? \nz.mem [2845] : 
                             (N172)? \nz.mem [2925] : 
                             (N174)? \nz.mem [3005] : 
                             (N176)? \nz.mem [3085] : 
                             (N178)? \nz.mem [3165] : 
                             (N180)? \nz.mem [3245] : 
                             (N182)? \nz.mem [3325] : 
                             (N184)? \nz.mem [3405] : 
                             (N186)? \nz.mem [3485] : 
                             (N188)? \nz.mem [3565] : 
                             (N190)? \nz.mem [3645] : 
                             (N192)? \nz.mem [3725] : 
                             (N194)? \nz.mem [3805] : 
                             (N196)? \nz.mem [3885] : 
                             (N198)? \nz.mem [3965] : 
                             (N200)? \nz.mem [4045] : 
                             (N202)? \nz.mem [4125] : 
                             (N204)? \nz.mem [4205] : 
                             (N206)? \nz.mem [4285] : 
                             (N208)? \nz.mem [4365] : 
                             (N210)? \nz.mem [4445] : 
                             (N212)? \nz.mem [4525] : 
                             (N214)? \nz.mem [4605] : 
                             (N216)? \nz.mem [4685] : 
                             (N218)? \nz.mem [4765] : 
                             (N220)? \nz.mem [4845] : 
                             (N222)? \nz.mem [4925] : 
                             (N224)? \nz.mem [5005] : 
                             (N226)? \nz.mem [5085] : 1'b0;
  assign \nz.data_out [44] = (N163)? \nz.mem [44] : 
                             (N165)? \nz.mem [124] : 
                             (N167)? \nz.mem [204] : 
                             (N169)? \nz.mem [284] : 
                             (N171)? \nz.mem [364] : 
                             (N173)? \nz.mem [444] : 
                             (N175)? \nz.mem [524] : 
                             (N177)? \nz.mem [604] : 
                             (N179)? \nz.mem [684] : 
                             (N181)? \nz.mem [764] : 
                             (N183)? \nz.mem [844] : 
                             (N185)? \nz.mem [924] : 
                             (N187)? \nz.mem [1004] : 
                             (N189)? \nz.mem [1084] : 
                             (N191)? \nz.mem [1164] : 
                             (N193)? \nz.mem [1244] : 
                             (N195)? \nz.mem [1324] : 
                             (N197)? \nz.mem [1404] : 
                             (N199)? \nz.mem [1484] : 
                             (N201)? \nz.mem [1564] : 
                             (N203)? \nz.mem [1644] : 
                             (N205)? \nz.mem [1724] : 
                             (N207)? \nz.mem [1804] : 
                             (N209)? \nz.mem [1884] : 
                             (N211)? \nz.mem [1964] : 
                             (N213)? \nz.mem [2044] : 
                             (N215)? \nz.mem [2124] : 
                             (N217)? \nz.mem [2204] : 
                             (N219)? \nz.mem [2284] : 
                             (N221)? \nz.mem [2364] : 
                             (N223)? \nz.mem [2444] : 
                             (N225)? \nz.mem [2524] : 
                             (N164)? \nz.mem [2604] : 
                             (N166)? \nz.mem [2684] : 
                             (N168)? \nz.mem [2764] : 
                             (N170)? \nz.mem [2844] : 
                             (N172)? \nz.mem [2924] : 
                             (N174)? \nz.mem [3004] : 
                             (N176)? \nz.mem [3084] : 
                             (N178)? \nz.mem [3164] : 
                             (N180)? \nz.mem [3244] : 
                             (N182)? \nz.mem [3324] : 
                             (N184)? \nz.mem [3404] : 
                             (N186)? \nz.mem [3484] : 
                             (N188)? \nz.mem [3564] : 
                             (N190)? \nz.mem [3644] : 
                             (N192)? \nz.mem [3724] : 
                             (N194)? \nz.mem [3804] : 
                             (N196)? \nz.mem [3884] : 
                             (N198)? \nz.mem [3964] : 
                             (N200)? \nz.mem [4044] : 
                             (N202)? \nz.mem [4124] : 
                             (N204)? \nz.mem [4204] : 
                             (N206)? \nz.mem [4284] : 
                             (N208)? \nz.mem [4364] : 
                             (N210)? \nz.mem [4444] : 
                             (N212)? \nz.mem [4524] : 
                             (N214)? \nz.mem [4604] : 
                             (N216)? \nz.mem [4684] : 
                             (N218)? \nz.mem [4764] : 
                             (N220)? \nz.mem [4844] : 
                             (N222)? \nz.mem [4924] : 
                             (N224)? \nz.mem [5004] : 
                             (N226)? \nz.mem [5084] : 1'b0;
  assign \nz.data_out [43] = (N163)? \nz.mem [43] : 
                             (N165)? \nz.mem [123] : 
                             (N167)? \nz.mem [203] : 
                             (N169)? \nz.mem [283] : 
                             (N171)? \nz.mem [363] : 
                             (N173)? \nz.mem [443] : 
                             (N175)? \nz.mem [523] : 
                             (N177)? \nz.mem [603] : 
                             (N179)? \nz.mem [683] : 
                             (N181)? \nz.mem [763] : 
                             (N183)? \nz.mem [843] : 
                             (N185)? \nz.mem [923] : 
                             (N187)? \nz.mem [1003] : 
                             (N189)? \nz.mem [1083] : 
                             (N191)? \nz.mem [1163] : 
                             (N193)? \nz.mem [1243] : 
                             (N195)? \nz.mem [1323] : 
                             (N197)? \nz.mem [1403] : 
                             (N199)? \nz.mem [1483] : 
                             (N201)? \nz.mem [1563] : 
                             (N203)? \nz.mem [1643] : 
                             (N205)? \nz.mem [1723] : 
                             (N207)? \nz.mem [1803] : 
                             (N209)? \nz.mem [1883] : 
                             (N211)? \nz.mem [1963] : 
                             (N213)? \nz.mem [2043] : 
                             (N215)? \nz.mem [2123] : 
                             (N217)? \nz.mem [2203] : 
                             (N219)? \nz.mem [2283] : 
                             (N221)? \nz.mem [2363] : 
                             (N223)? \nz.mem [2443] : 
                             (N225)? \nz.mem [2523] : 
                             (N164)? \nz.mem [2603] : 
                             (N166)? \nz.mem [2683] : 
                             (N168)? \nz.mem [2763] : 
                             (N170)? \nz.mem [2843] : 
                             (N172)? \nz.mem [2923] : 
                             (N174)? \nz.mem [3003] : 
                             (N176)? \nz.mem [3083] : 
                             (N178)? \nz.mem [3163] : 
                             (N180)? \nz.mem [3243] : 
                             (N182)? \nz.mem [3323] : 
                             (N184)? \nz.mem [3403] : 
                             (N186)? \nz.mem [3483] : 
                             (N188)? \nz.mem [3563] : 
                             (N190)? \nz.mem [3643] : 
                             (N192)? \nz.mem [3723] : 
                             (N194)? \nz.mem [3803] : 
                             (N196)? \nz.mem [3883] : 
                             (N198)? \nz.mem [3963] : 
                             (N200)? \nz.mem [4043] : 
                             (N202)? \nz.mem [4123] : 
                             (N204)? \nz.mem [4203] : 
                             (N206)? \nz.mem [4283] : 
                             (N208)? \nz.mem [4363] : 
                             (N210)? \nz.mem [4443] : 
                             (N212)? \nz.mem [4523] : 
                             (N214)? \nz.mem [4603] : 
                             (N216)? \nz.mem [4683] : 
                             (N218)? \nz.mem [4763] : 
                             (N220)? \nz.mem [4843] : 
                             (N222)? \nz.mem [4923] : 
                             (N224)? \nz.mem [5003] : 
                             (N226)? \nz.mem [5083] : 1'b0;
  assign \nz.data_out [42] = (N163)? \nz.mem [42] : 
                             (N165)? \nz.mem [122] : 
                             (N167)? \nz.mem [202] : 
                             (N169)? \nz.mem [282] : 
                             (N171)? \nz.mem [362] : 
                             (N173)? \nz.mem [442] : 
                             (N175)? \nz.mem [522] : 
                             (N177)? \nz.mem [602] : 
                             (N179)? \nz.mem [682] : 
                             (N181)? \nz.mem [762] : 
                             (N183)? \nz.mem [842] : 
                             (N185)? \nz.mem [922] : 
                             (N187)? \nz.mem [1002] : 
                             (N189)? \nz.mem [1082] : 
                             (N191)? \nz.mem [1162] : 
                             (N193)? \nz.mem [1242] : 
                             (N195)? \nz.mem [1322] : 
                             (N197)? \nz.mem [1402] : 
                             (N199)? \nz.mem [1482] : 
                             (N201)? \nz.mem [1562] : 
                             (N203)? \nz.mem [1642] : 
                             (N205)? \nz.mem [1722] : 
                             (N207)? \nz.mem [1802] : 
                             (N209)? \nz.mem [1882] : 
                             (N211)? \nz.mem [1962] : 
                             (N213)? \nz.mem [2042] : 
                             (N215)? \nz.mem [2122] : 
                             (N217)? \nz.mem [2202] : 
                             (N219)? \nz.mem [2282] : 
                             (N221)? \nz.mem [2362] : 
                             (N223)? \nz.mem [2442] : 
                             (N225)? \nz.mem [2522] : 
                             (N164)? \nz.mem [2602] : 
                             (N166)? \nz.mem [2682] : 
                             (N168)? \nz.mem [2762] : 
                             (N170)? \nz.mem [2842] : 
                             (N172)? \nz.mem [2922] : 
                             (N174)? \nz.mem [3002] : 
                             (N176)? \nz.mem [3082] : 
                             (N178)? \nz.mem [3162] : 
                             (N180)? \nz.mem [3242] : 
                             (N182)? \nz.mem [3322] : 
                             (N184)? \nz.mem [3402] : 
                             (N186)? \nz.mem [3482] : 
                             (N188)? \nz.mem [3562] : 
                             (N190)? \nz.mem [3642] : 
                             (N192)? \nz.mem [3722] : 
                             (N194)? \nz.mem [3802] : 
                             (N196)? \nz.mem [3882] : 
                             (N198)? \nz.mem [3962] : 
                             (N200)? \nz.mem [4042] : 
                             (N202)? \nz.mem [4122] : 
                             (N204)? \nz.mem [4202] : 
                             (N206)? \nz.mem [4282] : 
                             (N208)? \nz.mem [4362] : 
                             (N210)? \nz.mem [4442] : 
                             (N212)? \nz.mem [4522] : 
                             (N214)? \nz.mem [4602] : 
                             (N216)? \nz.mem [4682] : 
                             (N218)? \nz.mem [4762] : 
                             (N220)? \nz.mem [4842] : 
                             (N222)? \nz.mem [4922] : 
                             (N224)? \nz.mem [5002] : 
                             (N226)? \nz.mem [5082] : 1'b0;
  assign \nz.data_out [41] = (N163)? \nz.mem [41] : 
                             (N165)? \nz.mem [121] : 
                             (N167)? \nz.mem [201] : 
                             (N169)? \nz.mem [281] : 
                             (N171)? \nz.mem [361] : 
                             (N173)? \nz.mem [441] : 
                             (N175)? \nz.mem [521] : 
                             (N177)? \nz.mem [601] : 
                             (N179)? \nz.mem [681] : 
                             (N181)? \nz.mem [761] : 
                             (N183)? \nz.mem [841] : 
                             (N185)? \nz.mem [921] : 
                             (N187)? \nz.mem [1001] : 
                             (N189)? \nz.mem [1081] : 
                             (N191)? \nz.mem [1161] : 
                             (N193)? \nz.mem [1241] : 
                             (N195)? \nz.mem [1321] : 
                             (N197)? \nz.mem [1401] : 
                             (N199)? \nz.mem [1481] : 
                             (N201)? \nz.mem [1561] : 
                             (N203)? \nz.mem [1641] : 
                             (N205)? \nz.mem [1721] : 
                             (N207)? \nz.mem [1801] : 
                             (N209)? \nz.mem [1881] : 
                             (N211)? \nz.mem [1961] : 
                             (N213)? \nz.mem [2041] : 
                             (N215)? \nz.mem [2121] : 
                             (N217)? \nz.mem [2201] : 
                             (N219)? \nz.mem [2281] : 
                             (N221)? \nz.mem [2361] : 
                             (N223)? \nz.mem [2441] : 
                             (N225)? \nz.mem [2521] : 
                             (N164)? \nz.mem [2601] : 
                             (N166)? \nz.mem [2681] : 
                             (N168)? \nz.mem [2761] : 
                             (N170)? \nz.mem [2841] : 
                             (N172)? \nz.mem [2921] : 
                             (N174)? \nz.mem [3001] : 
                             (N176)? \nz.mem [3081] : 
                             (N178)? \nz.mem [3161] : 
                             (N180)? \nz.mem [3241] : 
                             (N182)? \nz.mem [3321] : 
                             (N184)? \nz.mem [3401] : 
                             (N186)? \nz.mem [3481] : 
                             (N188)? \nz.mem [3561] : 
                             (N190)? \nz.mem [3641] : 
                             (N192)? \nz.mem [3721] : 
                             (N194)? \nz.mem [3801] : 
                             (N196)? \nz.mem [3881] : 
                             (N198)? \nz.mem [3961] : 
                             (N200)? \nz.mem [4041] : 
                             (N202)? \nz.mem [4121] : 
                             (N204)? \nz.mem [4201] : 
                             (N206)? \nz.mem [4281] : 
                             (N208)? \nz.mem [4361] : 
                             (N210)? \nz.mem [4441] : 
                             (N212)? \nz.mem [4521] : 
                             (N214)? \nz.mem [4601] : 
                             (N216)? \nz.mem [4681] : 
                             (N218)? \nz.mem [4761] : 
                             (N220)? \nz.mem [4841] : 
                             (N222)? \nz.mem [4921] : 
                             (N224)? \nz.mem [5001] : 
                             (N226)? \nz.mem [5081] : 1'b0;
  assign \nz.data_out [40] = (N163)? \nz.mem [40] : 
                             (N165)? \nz.mem [120] : 
                             (N167)? \nz.mem [200] : 
                             (N169)? \nz.mem [280] : 
                             (N171)? \nz.mem [360] : 
                             (N173)? \nz.mem [440] : 
                             (N175)? \nz.mem [520] : 
                             (N177)? \nz.mem [600] : 
                             (N179)? \nz.mem [680] : 
                             (N181)? \nz.mem [760] : 
                             (N183)? \nz.mem [840] : 
                             (N185)? \nz.mem [920] : 
                             (N187)? \nz.mem [1000] : 
                             (N189)? \nz.mem [1080] : 
                             (N191)? \nz.mem [1160] : 
                             (N193)? \nz.mem [1240] : 
                             (N195)? \nz.mem [1320] : 
                             (N197)? \nz.mem [1400] : 
                             (N199)? \nz.mem [1480] : 
                             (N201)? \nz.mem [1560] : 
                             (N203)? \nz.mem [1640] : 
                             (N205)? \nz.mem [1720] : 
                             (N207)? \nz.mem [1800] : 
                             (N209)? \nz.mem [1880] : 
                             (N211)? \nz.mem [1960] : 
                             (N213)? \nz.mem [2040] : 
                             (N215)? \nz.mem [2120] : 
                             (N217)? \nz.mem [2200] : 
                             (N219)? \nz.mem [2280] : 
                             (N221)? \nz.mem [2360] : 
                             (N223)? \nz.mem [2440] : 
                             (N225)? \nz.mem [2520] : 
                             (N164)? \nz.mem [2600] : 
                             (N166)? \nz.mem [2680] : 
                             (N168)? \nz.mem [2760] : 
                             (N170)? \nz.mem [2840] : 
                             (N172)? \nz.mem [2920] : 
                             (N174)? \nz.mem [3000] : 
                             (N176)? \nz.mem [3080] : 
                             (N178)? \nz.mem [3160] : 
                             (N180)? \nz.mem [3240] : 
                             (N182)? \nz.mem [3320] : 
                             (N184)? \nz.mem [3400] : 
                             (N186)? \nz.mem [3480] : 
                             (N188)? \nz.mem [3560] : 
                             (N190)? \nz.mem [3640] : 
                             (N192)? \nz.mem [3720] : 
                             (N194)? \nz.mem [3800] : 
                             (N196)? \nz.mem [3880] : 
                             (N198)? \nz.mem [3960] : 
                             (N200)? \nz.mem [4040] : 
                             (N202)? \nz.mem [4120] : 
                             (N204)? \nz.mem [4200] : 
                             (N206)? \nz.mem [4280] : 
                             (N208)? \nz.mem [4360] : 
                             (N210)? \nz.mem [4440] : 
                             (N212)? \nz.mem [4520] : 
                             (N214)? \nz.mem [4600] : 
                             (N216)? \nz.mem [4680] : 
                             (N218)? \nz.mem [4760] : 
                             (N220)? \nz.mem [4840] : 
                             (N222)? \nz.mem [4920] : 
                             (N224)? \nz.mem [5000] : 
                             (N226)? \nz.mem [5080] : 1'b0;
  assign \nz.data_out [39] = (N163)? \nz.mem [39] : 
                             (N165)? \nz.mem [119] : 
                             (N167)? \nz.mem [199] : 
                             (N169)? \nz.mem [279] : 
                             (N171)? \nz.mem [359] : 
                             (N173)? \nz.mem [439] : 
                             (N175)? \nz.mem [519] : 
                             (N177)? \nz.mem [599] : 
                             (N179)? \nz.mem [679] : 
                             (N181)? \nz.mem [759] : 
                             (N183)? \nz.mem [839] : 
                             (N185)? \nz.mem [919] : 
                             (N187)? \nz.mem [999] : 
                             (N189)? \nz.mem [1079] : 
                             (N191)? \nz.mem [1159] : 
                             (N193)? \nz.mem [1239] : 
                             (N195)? \nz.mem [1319] : 
                             (N197)? \nz.mem [1399] : 
                             (N199)? \nz.mem [1479] : 
                             (N201)? \nz.mem [1559] : 
                             (N203)? \nz.mem [1639] : 
                             (N205)? \nz.mem [1719] : 
                             (N207)? \nz.mem [1799] : 
                             (N209)? \nz.mem [1879] : 
                             (N211)? \nz.mem [1959] : 
                             (N213)? \nz.mem [2039] : 
                             (N215)? \nz.mem [2119] : 
                             (N217)? \nz.mem [2199] : 
                             (N219)? \nz.mem [2279] : 
                             (N221)? \nz.mem [2359] : 
                             (N223)? \nz.mem [2439] : 
                             (N225)? \nz.mem [2519] : 
                             (N164)? \nz.mem [2599] : 
                             (N166)? \nz.mem [2679] : 
                             (N168)? \nz.mem [2759] : 
                             (N170)? \nz.mem [2839] : 
                             (N172)? \nz.mem [2919] : 
                             (N174)? \nz.mem [2999] : 
                             (N176)? \nz.mem [3079] : 
                             (N178)? \nz.mem [3159] : 
                             (N180)? \nz.mem [3239] : 
                             (N182)? \nz.mem [3319] : 
                             (N184)? \nz.mem [3399] : 
                             (N186)? \nz.mem [3479] : 
                             (N188)? \nz.mem [3559] : 
                             (N190)? \nz.mem [3639] : 
                             (N192)? \nz.mem [3719] : 
                             (N194)? \nz.mem [3799] : 
                             (N196)? \nz.mem [3879] : 
                             (N198)? \nz.mem [3959] : 
                             (N200)? \nz.mem [4039] : 
                             (N202)? \nz.mem [4119] : 
                             (N204)? \nz.mem [4199] : 
                             (N206)? \nz.mem [4279] : 
                             (N208)? \nz.mem [4359] : 
                             (N210)? \nz.mem [4439] : 
                             (N212)? \nz.mem [4519] : 
                             (N214)? \nz.mem [4599] : 
                             (N216)? \nz.mem [4679] : 
                             (N218)? \nz.mem [4759] : 
                             (N220)? \nz.mem [4839] : 
                             (N222)? \nz.mem [4919] : 
                             (N224)? \nz.mem [4999] : 
                             (N226)? \nz.mem [5079] : 1'b0;
  assign \nz.data_out [38] = (N163)? \nz.mem [38] : 
                             (N165)? \nz.mem [118] : 
                             (N167)? \nz.mem [198] : 
                             (N169)? \nz.mem [278] : 
                             (N171)? \nz.mem [358] : 
                             (N173)? \nz.mem [438] : 
                             (N175)? \nz.mem [518] : 
                             (N177)? \nz.mem [598] : 
                             (N179)? \nz.mem [678] : 
                             (N181)? \nz.mem [758] : 
                             (N183)? \nz.mem [838] : 
                             (N185)? \nz.mem [918] : 
                             (N187)? \nz.mem [998] : 
                             (N189)? \nz.mem [1078] : 
                             (N191)? \nz.mem [1158] : 
                             (N193)? \nz.mem [1238] : 
                             (N195)? \nz.mem [1318] : 
                             (N197)? \nz.mem [1398] : 
                             (N199)? \nz.mem [1478] : 
                             (N201)? \nz.mem [1558] : 
                             (N203)? \nz.mem [1638] : 
                             (N205)? \nz.mem [1718] : 
                             (N207)? \nz.mem [1798] : 
                             (N209)? \nz.mem [1878] : 
                             (N211)? \nz.mem [1958] : 
                             (N213)? \nz.mem [2038] : 
                             (N215)? \nz.mem [2118] : 
                             (N217)? \nz.mem [2198] : 
                             (N219)? \nz.mem [2278] : 
                             (N221)? \nz.mem [2358] : 
                             (N223)? \nz.mem [2438] : 
                             (N225)? \nz.mem [2518] : 
                             (N164)? \nz.mem [2598] : 
                             (N166)? \nz.mem [2678] : 
                             (N168)? \nz.mem [2758] : 
                             (N170)? \nz.mem [2838] : 
                             (N172)? \nz.mem [2918] : 
                             (N174)? \nz.mem [2998] : 
                             (N176)? \nz.mem [3078] : 
                             (N178)? \nz.mem [3158] : 
                             (N180)? \nz.mem [3238] : 
                             (N182)? \nz.mem [3318] : 
                             (N184)? \nz.mem [3398] : 
                             (N186)? \nz.mem [3478] : 
                             (N188)? \nz.mem [3558] : 
                             (N190)? \nz.mem [3638] : 
                             (N192)? \nz.mem [3718] : 
                             (N194)? \nz.mem [3798] : 
                             (N196)? \nz.mem [3878] : 
                             (N198)? \nz.mem [3958] : 
                             (N200)? \nz.mem [4038] : 
                             (N202)? \nz.mem [4118] : 
                             (N204)? \nz.mem [4198] : 
                             (N206)? \nz.mem [4278] : 
                             (N208)? \nz.mem [4358] : 
                             (N210)? \nz.mem [4438] : 
                             (N212)? \nz.mem [4518] : 
                             (N214)? \nz.mem [4598] : 
                             (N216)? \nz.mem [4678] : 
                             (N218)? \nz.mem [4758] : 
                             (N220)? \nz.mem [4838] : 
                             (N222)? \nz.mem [4918] : 
                             (N224)? \nz.mem [4998] : 
                             (N226)? \nz.mem [5078] : 1'b0;
  assign \nz.data_out [37] = (N163)? \nz.mem [37] : 
                             (N165)? \nz.mem [117] : 
                             (N167)? \nz.mem [197] : 
                             (N169)? \nz.mem [277] : 
                             (N171)? \nz.mem [357] : 
                             (N173)? \nz.mem [437] : 
                             (N175)? \nz.mem [517] : 
                             (N177)? \nz.mem [597] : 
                             (N179)? \nz.mem [677] : 
                             (N181)? \nz.mem [757] : 
                             (N183)? \nz.mem [837] : 
                             (N185)? \nz.mem [917] : 
                             (N187)? \nz.mem [997] : 
                             (N189)? \nz.mem [1077] : 
                             (N191)? \nz.mem [1157] : 
                             (N193)? \nz.mem [1237] : 
                             (N195)? \nz.mem [1317] : 
                             (N197)? \nz.mem [1397] : 
                             (N199)? \nz.mem [1477] : 
                             (N201)? \nz.mem [1557] : 
                             (N203)? \nz.mem [1637] : 
                             (N205)? \nz.mem [1717] : 
                             (N207)? \nz.mem [1797] : 
                             (N209)? \nz.mem [1877] : 
                             (N211)? \nz.mem [1957] : 
                             (N213)? \nz.mem [2037] : 
                             (N215)? \nz.mem [2117] : 
                             (N217)? \nz.mem [2197] : 
                             (N219)? \nz.mem [2277] : 
                             (N221)? \nz.mem [2357] : 
                             (N223)? \nz.mem [2437] : 
                             (N225)? \nz.mem [2517] : 
                             (N164)? \nz.mem [2597] : 
                             (N166)? \nz.mem [2677] : 
                             (N168)? \nz.mem [2757] : 
                             (N170)? \nz.mem [2837] : 
                             (N172)? \nz.mem [2917] : 
                             (N174)? \nz.mem [2997] : 
                             (N176)? \nz.mem [3077] : 
                             (N178)? \nz.mem [3157] : 
                             (N180)? \nz.mem [3237] : 
                             (N182)? \nz.mem [3317] : 
                             (N184)? \nz.mem [3397] : 
                             (N186)? \nz.mem [3477] : 
                             (N188)? \nz.mem [3557] : 
                             (N190)? \nz.mem [3637] : 
                             (N192)? \nz.mem [3717] : 
                             (N194)? \nz.mem [3797] : 
                             (N196)? \nz.mem [3877] : 
                             (N198)? \nz.mem [3957] : 
                             (N200)? \nz.mem [4037] : 
                             (N202)? \nz.mem [4117] : 
                             (N204)? \nz.mem [4197] : 
                             (N206)? \nz.mem [4277] : 
                             (N208)? \nz.mem [4357] : 
                             (N210)? \nz.mem [4437] : 
                             (N212)? \nz.mem [4517] : 
                             (N214)? \nz.mem [4597] : 
                             (N216)? \nz.mem [4677] : 
                             (N218)? \nz.mem [4757] : 
                             (N220)? \nz.mem [4837] : 
                             (N222)? \nz.mem [4917] : 
                             (N224)? \nz.mem [4997] : 
                             (N226)? \nz.mem [5077] : 1'b0;
  assign \nz.data_out [36] = (N163)? \nz.mem [36] : 
                             (N165)? \nz.mem [116] : 
                             (N167)? \nz.mem [196] : 
                             (N169)? \nz.mem [276] : 
                             (N171)? \nz.mem [356] : 
                             (N173)? \nz.mem [436] : 
                             (N175)? \nz.mem [516] : 
                             (N177)? \nz.mem [596] : 
                             (N179)? \nz.mem [676] : 
                             (N181)? \nz.mem [756] : 
                             (N183)? \nz.mem [836] : 
                             (N185)? \nz.mem [916] : 
                             (N187)? \nz.mem [996] : 
                             (N189)? \nz.mem [1076] : 
                             (N191)? \nz.mem [1156] : 
                             (N193)? \nz.mem [1236] : 
                             (N195)? \nz.mem [1316] : 
                             (N197)? \nz.mem [1396] : 
                             (N199)? \nz.mem [1476] : 
                             (N201)? \nz.mem [1556] : 
                             (N203)? \nz.mem [1636] : 
                             (N205)? \nz.mem [1716] : 
                             (N207)? \nz.mem [1796] : 
                             (N209)? \nz.mem [1876] : 
                             (N211)? \nz.mem [1956] : 
                             (N213)? \nz.mem [2036] : 
                             (N215)? \nz.mem [2116] : 
                             (N217)? \nz.mem [2196] : 
                             (N219)? \nz.mem [2276] : 
                             (N221)? \nz.mem [2356] : 
                             (N223)? \nz.mem [2436] : 
                             (N225)? \nz.mem [2516] : 
                             (N164)? \nz.mem [2596] : 
                             (N166)? \nz.mem [2676] : 
                             (N168)? \nz.mem [2756] : 
                             (N170)? \nz.mem [2836] : 
                             (N172)? \nz.mem [2916] : 
                             (N174)? \nz.mem [2996] : 
                             (N176)? \nz.mem [3076] : 
                             (N178)? \nz.mem [3156] : 
                             (N180)? \nz.mem [3236] : 
                             (N182)? \nz.mem [3316] : 
                             (N184)? \nz.mem [3396] : 
                             (N186)? \nz.mem [3476] : 
                             (N188)? \nz.mem [3556] : 
                             (N190)? \nz.mem [3636] : 
                             (N192)? \nz.mem [3716] : 
                             (N194)? \nz.mem [3796] : 
                             (N196)? \nz.mem [3876] : 
                             (N198)? \nz.mem [3956] : 
                             (N200)? \nz.mem [4036] : 
                             (N202)? \nz.mem [4116] : 
                             (N204)? \nz.mem [4196] : 
                             (N206)? \nz.mem [4276] : 
                             (N208)? \nz.mem [4356] : 
                             (N210)? \nz.mem [4436] : 
                             (N212)? \nz.mem [4516] : 
                             (N214)? \nz.mem [4596] : 
                             (N216)? \nz.mem [4676] : 
                             (N218)? \nz.mem [4756] : 
                             (N220)? \nz.mem [4836] : 
                             (N222)? \nz.mem [4916] : 
                             (N224)? \nz.mem [4996] : 
                             (N226)? \nz.mem [5076] : 1'b0;
  assign \nz.data_out [35] = (N163)? \nz.mem [35] : 
                             (N165)? \nz.mem [115] : 
                             (N167)? \nz.mem [195] : 
                             (N169)? \nz.mem [275] : 
                             (N171)? \nz.mem [355] : 
                             (N173)? \nz.mem [435] : 
                             (N175)? \nz.mem [515] : 
                             (N177)? \nz.mem [595] : 
                             (N179)? \nz.mem [675] : 
                             (N181)? \nz.mem [755] : 
                             (N183)? \nz.mem [835] : 
                             (N185)? \nz.mem [915] : 
                             (N187)? \nz.mem [995] : 
                             (N189)? \nz.mem [1075] : 
                             (N191)? \nz.mem [1155] : 
                             (N193)? \nz.mem [1235] : 
                             (N195)? \nz.mem [1315] : 
                             (N197)? \nz.mem [1395] : 
                             (N199)? \nz.mem [1475] : 
                             (N201)? \nz.mem [1555] : 
                             (N203)? \nz.mem [1635] : 
                             (N205)? \nz.mem [1715] : 
                             (N207)? \nz.mem [1795] : 
                             (N209)? \nz.mem [1875] : 
                             (N211)? \nz.mem [1955] : 
                             (N213)? \nz.mem [2035] : 
                             (N215)? \nz.mem [2115] : 
                             (N217)? \nz.mem [2195] : 
                             (N219)? \nz.mem [2275] : 
                             (N221)? \nz.mem [2355] : 
                             (N223)? \nz.mem [2435] : 
                             (N225)? \nz.mem [2515] : 
                             (N164)? \nz.mem [2595] : 
                             (N166)? \nz.mem [2675] : 
                             (N168)? \nz.mem [2755] : 
                             (N170)? \nz.mem [2835] : 
                             (N172)? \nz.mem [2915] : 
                             (N174)? \nz.mem [2995] : 
                             (N176)? \nz.mem [3075] : 
                             (N178)? \nz.mem [3155] : 
                             (N180)? \nz.mem [3235] : 
                             (N182)? \nz.mem [3315] : 
                             (N184)? \nz.mem [3395] : 
                             (N186)? \nz.mem [3475] : 
                             (N188)? \nz.mem [3555] : 
                             (N190)? \nz.mem [3635] : 
                             (N192)? \nz.mem [3715] : 
                             (N194)? \nz.mem [3795] : 
                             (N196)? \nz.mem [3875] : 
                             (N198)? \nz.mem [3955] : 
                             (N200)? \nz.mem [4035] : 
                             (N202)? \nz.mem [4115] : 
                             (N204)? \nz.mem [4195] : 
                             (N206)? \nz.mem [4275] : 
                             (N208)? \nz.mem [4355] : 
                             (N210)? \nz.mem [4435] : 
                             (N212)? \nz.mem [4515] : 
                             (N214)? \nz.mem [4595] : 
                             (N216)? \nz.mem [4675] : 
                             (N218)? \nz.mem [4755] : 
                             (N220)? \nz.mem [4835] : 
                             (N222)? \nz.mem [4915] : 
                             (N224)? \nz.mem [4995] : 
                             (N226)? \nz.mem [5075] : 1'b0;
  assign \nz.data_out [34] = (N163)? \nz.mem [34] : 
                             (N165)? \nz.mem [114] : 
                             (N167)? \nz.mem [194] : 
                             (N169)? \nz.mem [274] : 
                             (N171)? \nz.mem [354] : 
                             (N173)? \nz.mem [434] : 
                             (N175)? \nz.mem [514] : 
                             (N177)? \nz.mem [594] : 
                             (N179)? \nz.mem [674] : 
                             (N181)? \nz.mem [754] : 
                             (N183)? \nz.mem [834] : 
                             (N185)? \nz.mem [914] : 
                             (N187)? \nz.mem [994] : 
                             (N189)? \nz.mem [1074] : 
                             (N191)? \nz.mem [1154] : 
                             (N193)? \nz.mem [1234] : 
                             (N195)? \nz.mem [1314] : 
                             (N197)? \nz.mem [1394] : 
                             (N199)? \nz.mem [1474] : 
                             (N201)? \nz.mem [1554] : 
                             (N203)? \nz.mem [1634] : 
                             (N205)? \nz.mem [1714] : 
                             (N207)? \nz.mem [1794] : 
                             (N209)? \nz.mem [1874] : 
                             (N211)? \nz.mem [1954] : 
                             (N213)? \nz.mem [2034] : 
                             (N215)? \nz.mem [2114] : 
                             (N217)? \nz.mem [2194] : 
                             (N219)? \nz.mem [2274] : 
                             (N221)? \nz.mem [2354] : 
                             (N223)? \nz.mem [2434] : 
                             (N225)? \nz.mem [2514] : 
                             (N164)? \nz.mem [2594] : 
                             (N166)? \nz.mem [2674] : 
                             (N168)? \nz.mem [2754] : 
                             (N170)? \nz.mem [2834] : 
                             (N172)? \nz.mem [2914] : 
                             (N174)? \nz.mem [2994] : 
                             (N176)? \nz.mem [3074] : 
                             (N178)? \nz.mem [3154] : 
                             (N180)? \nz.mem [3234] : 
                             (N182)? \nz.mem [3314] : 
                             (N184)? \nz.mem [3394] : 
                             (N186)? \nz.mem [3474] : 
                             (N188)? \nz.mem [3554] : 
                             (N190)? \nz.mem [3634] : 
                             (N192)? \nz.mem [3714] : 
                             (N194)? \nz.mem [3794] : 
                             (N196)? \nz.mem [3874] : 
                             (N198)? \nz.mem [3954] : 
                             (N200)? \nz.mem [4034] : 
                             (N202)? \nz.mem [4114] : 
                             (N204)? \nz.mem [4194] : 
                             (N206)? \nz.mem [4274] : 
                             (N208)? \nz.mem [4354] : 
                             (N210)? \nz.mem [4434] : 
                             (N212)? \nz.mem [4514] : 
                             (N214)? \nz.mem [4594] : 
                             (N216)? \nz.mem [4674] : 
                             (N218)? \nz.mem [4754] : 
                             (N220)? \nz.mem [4834] : 
                             (N222)? \nz.mem [4914] : 
                             (N224)? \nz.mem [4994] : 
                             (N226)? \nz.mem [5074] : 1'b0;
  assign \nz.data_out [33] = (N163)? \nz.mem [33] : 
                             (N165)? \nz.mem [113] : 
                             (N167)? \nz.mem [193] : 
                             (N169)? \nz.mem [273] : 
                             (N171)? \nz.mem [353] : 
                             (N173)? \nz.mem [433] : 
                             (N175)? \nz.mem [513] : 
                             (N177)? \nz.mem [593] : 
                             (N179)? \nz.mem [673] : 
                             (N181)? \nz.mem [753] : 
                             (N183)? \nz.mem [833] : 
                             (N185)? \nz.mem [913] : 
                             (N187)? \nz.mem [993] : 
                             (N189)? \nz.mem [1073] : 
                             (N191)? \nz.mem [1153] : 
                             (N193)? \nz.mem [1233] : 
                             (N195)? \nz.mem [1313] : 
                             (N197)? \nz.mem [1393] : 
                             (N199)? \nz.mem [1473] : 
                             (N201)? \nz.mem [1553] : 
                             (N203)? \nz.mem [1633] : 
                             (N205)? \nz.mem [1713] : 
                             (N207)? \nz.mem [1793] : 
                             (N209)? \nz.mem [1873] : 
                             (N211)? \nz.mem [1953] : 
                             (N213)? \nz.mem [2033] : 
                             (N215)? \nz.mem [2113] : 
                             (N217)? \nz.mem [2193] : 
                             (N219)? \nz.mem [2273] : 
                             (N221)? \nz.mem [2353] : 
                             (N223)? \nz.mem [2433] : 
                             (N225)? \nz.mem [2513] : 
                             (N164)? \nz.mem [2593] : 
                             (N166)? \nz.mem [2673] : 
                             (N168)? \nz.mem [2753] : 
                             (N170)? \nz.mem [2833] : 
                             (N172)? \nz.mem [2913] : 
                             (N174)? \nz.mem [2993] : 
                             (N176)? \nz.mem [3073] : 
                             (N178)? \nz.mem [3153] : 
                             (N180)? \nz.mem [3233] : 
                             (N182)? \nz.mem [3313] : 
                             (N184)? \nz.mem [3393] : 
                             (N186)? \nz.mem [3473] : 
                             (N188)? \nz.mem [3553] : 
                             (N190)? \nz.mem [3633] : 
                             (N192)? \nz.mem [3713] : 
                             (N194)? \nz.mem [3793] : 
                             (N196)? \nz.mem [3873] : 
                             (N198)? \nz.mem [3953] : 
                             (N200)? \nz.mem [4033] : 
                             (N202)? \nz.mem [4113] : 
                             (N204)? \nz.mem [4193] : 
                             (N206)? \nz.mem [4273] : 
                             (N208)? \nz.mem [4353] : 
                             (N210)? \nz.mem [4433] : 
                             (N212)? \nz.mem [4513] : 
                             (N214)? \nz.mem [4593] : 
                             (N216)? \nz.mem [4673] : 
                             (N218)? \nz.mem [4753] : 
                             (N220)? \nz.mem [4833] : 
                             (N222)? \nz.mem [4913] : 
                             (N224)? \nz.mem [4993] : 
                             (N226)? \nz.mem [5073] : 1'b0;
  assign \nz.data_out [32] = (N163)? \nz.mem [32] : 
                             (N165)? \nz.mem [112] : 
                             (N167)? \nz.mem [192] : 
                             (N169)? \nz.mem [272] : 
                             (N171)? \nz.mem [352] : 
                             (N173)? \nz.mem [432] : 
                             (N175)? \nz.mem [512] : 
                             (N177)? \nz.mem [592] : 
                             (N179)? \nz.mem [672] : 
                             (N181)? \nz.mem [752] : 
                             (N183)? \nz.mem [832] : 
                             (N185)? \nz.mem [912] : 
                             (N187)? \nz.mem [992] : 
                             (N189)? \nz.mem [1072] : 
                             (N191)? \nz.mem [1152] : 
                             (N193)? \nz.mem [1232] : 
                             (N195)? \nz.mem [1312] : 
                             (N197)? \nz.mem [1392] : 
                             (N199)? \nz.mem [1472] : 
                             (N201)? \nz.mem [1552] : 
                             (N203)? \nz.mem [1632] : 
                             (N205)? \nz.mem [1712] : 
                             (N207)? \nz.mem [1792] : 
                             (N209)? \nz.mem [1872] : 
                             (N211)? \nz.mem [1952] : 
                             (N213)? \nz.mem [2032] : 
                             (N215)? \nz.mem [2112] : 
                             (N217)? \nz.mem [2192] : 
                             (N219)? \nz.mem [2272] : 
                             (N221)? \nz.mem [2352] : 
                             (N223)? \nz.mem [2432] : 
                             (N225)? \nz.mem [2512] : 
                             (N164)? \nz.mem [2592] : 
                             (N166)? \nz.mem [2672] : 
                             (N168)? \nz.mem [2752] : 
                             (N170)? \nz.mem [2832] : 
                             (N172)? \nz.mem [2912] : 
                             (N174)? \nz.mem [2992] : 
                             (N176)? \nz.mem [3072] : 
                             (N178)? \nz.mem [3152] : 
                             (N180)? \nz.mem [3232] : 
                             (N182)? \nz.mem [3312] : 
                             (N184)? \nz.mem [3392] : 
                             (N186)? \nz.mem [3472] : 
                             (N188)? \nz.mem [3552] : 
                             (N190)? \nz.mem [3632] : 
                             (N192)? \nz.mem [3712] : 
                             (N194)? \nz.mem [3792] : 
                             (N196)? \nz.mem [3872] : 
                             (N198)? \nz.mem [3952] : 
                             (N200)? \nz.mem [4032] : 
                             (N202)? \nz.mem [4112] : 
                             (N204)? \nz.mem [4192] : 
                             (N206)? \nz.mem [4272] : 
                             (N208)? \nz.mem [4352] : 
                             (N210)? \nz.mem [4432] : 
                             (N212)? \nz.mem [4512] : 
                             (N214)? \nz.mem [4592] : 
                             (N216)? \nz.mem [4672] : 
                             (N218)? \nz.mem [4752] : 
                             (N220)? \nz.mem [4832] : 
                             (N222)? \nz.mem [4912] : 
                             (N224)? \nz.mem [4992] : 
                             (N226)? \nz.mem [5072] : 1'b0;
  assign \nz.data_out [31] = (N163)? \nz.mem [31] : 
                             (N165)? \nz.mem [111] : 
                             (N167)? \nz.mem [191] : 
                             (N169)? \nz.mem [271] : 
                             (N171)? \nz.mem [351] : 
                             (N173)? \nz.mem [431] : 
                             (N175)? \nz.mem [511] : 
                             (N177)? \nz.mem [591] : 
                             (N179)? \nz.mem [671] : 
                             (N181)? \nz.mem [751] : 
                             (N183)? \nz.mem [831] : 
                             (N185)? \nz.mem [911] : 
                             (N187)? \nz.mem [991] : 
                             (N189)? \nz.mem [1071] : 
                             (N191)? \nz.mem [1151] : 
                             (N193)? \nz.mem [1231] : 
                             (N195)? \nz.mem [1311] : 
                             (N197)? \nz.mem [1391] : 
                             (N199)? \nz.mem [1471] : 
                             (N201)? \nz.mem [1551] : 
                             (N203)? \nz.mem [1631] : 
                             (N205)? \nz.mem [1711] : 
                             (N207)? \nz.mem [1791] : 
                             (N209)? \nz.mem [1871] : 
                             (N211)? \nz.mem [1951] : 
                             (N213)? \nz.mem [2031] : 
                             (N215)? \nz.mem [2111] : 
                             (N217)? \nz.mem [2191] : 
                             (N219)? \nz.mem [2271] : 
                             (N221)? \nz.mem [2351] : 
                             (N223)? \nz.mem [2431] : 
                             (N225)? \nz.mem [2511] : 
                             (N164)? \nz.mem [2591] : 
                             (N166)? \nz.mem [2671] : 
                             (N168)? \nz.mem [2751] : 
                             (N170)? \nz.mem [2831] : 
                             (N172)? \nz.mem [2911] : 
                             (N174)? \nz.mem [2991] : 
                             (N176)? \nz.mem [3071] : 
                             (N178)? \nz.mem [3151] : 
                             (N180)? \nz.mem [3231] : 
                             (N182)? \nz.mem [3311] : 
                             (N184)? \nz.mem [3391] : 
                             (N186)? \nz.mem [3471] : 
                             (N188)? \nz.mem [3551] : 
                             (N190)? \nz.mem [3631] : 
                             (N192)? \nz.mem [3711] : 
                             (N194)? \nz.mem [3791] : 
                             (N196)? \nz.mem [3871] : 
                             (N198)? \nz.mem [3951] : 
                             (N200)? \nz.mem [4031] : 
                             (N202)? \nz.mem [4111] : 
                             (N204)? \nz.mem [4191] : 
                             (N206)? \nz.mem [4271] : 
                             (N208)? \nz.mem [4351] : 
                             (N210)? \nz.mem [4431] : 
                             (N212)? \nz.mem [4511] : 
                             (N214)? \nz.mem [4591] : 
                             (N216)? \nz.mem [4671] : 
                             (N218)? \nz.mem [4751] : 
                             (N220)? \nz.mem [4831] : 
                             (N222)? \nz.mem [4911] : 
                             (N224)? \nz.mem [4991] : 
                             (N226)? \nz.mem [5071] : 1'b0;
  assign \nz.data_out [30] = (N163)? \nz.mem [30] : 
                             (N165)? \nz.mem [110] : 
                             (N167)? \nz.mem [190] : 
                             (N169)? \nz.mem [270] : 
                             (N171)? \nz.mem [350] : 
                             (N173)? \nz.mem [430] : 
                             (N175)? \nz.mem [510] : 
                             (N177)? \nz.mem [590] : 
                             (N179)? \nz.mem [670] : 
                             (N181)? \nz.mem [750] : 
                             (N183)? \nz.mem [830] : 
                             (N185)? \nz.mem [910] : 
                             (N187)? \nz.mem [990] : 
                             (N189)? \nz.mem [1070] : 
                             (N191)? \nz.mem [1150] : 
                             (N193)? \nz.mem [1230] : 
                             (N195)? \nz.mem [1310] : 
                             (N197)? \nz.mem [1390] : 
                             (N199)? \nz.mem [1470] : 
                             (N201)? \nz.mem [1550] : 
                             (N203)? \nz.mem [1630] : 
                             (N205)? \nz.mem [1710] : 
                             (N207)? \nz.mem [1790] : 
                             (N209)? \nz.mem [1870] : 
                             (N211)? \nz.mem [1950] : 
                             (N213)? \nz.mem [2030] : 
                             (N215)? \nz.mem [2110] : 
                             (N217)? \nz.mem [2190] : 
                             (N219)? \nz.mem [2270] : 
                             (N221)? \nz.mem [2350] : 
                             (N223)? \nz.mem [2430] : 
                             (N225)? \nz.mem [2510] : 
                             (N164)? \nz.mem [2590] : 
                             (N166)? \nz.mem [2670] : 
                             (N168)? \nz.mem [2750] : 
                             (N170)? \nz.mem [2830] : 
                             (N172)? \nz.mem [2910] : 
                             (N174)? \nz.mem [2990] : 
                             (N176)? \nz.mem [3070] : 
                             (N178)? \nz.mem [3150] : 
                             (N180)? \nz.mem [3230] : 
                             (N182)? \nz.mem [3310] : 
                             (N184)? \nz.mem [3390] : 
                             (N186)? \nz.mem [3470] : 
                             (N188)? \nz.mem [3550] : 
                             (N190)? \nz.mem [3630] : 
                             (N192)? \nz.mem [3710] : 
                             (N194)? \nz.mem [3790] : 
                             (N196)? \nz.mem [3870] : 
                             (N198)? \nz.mem [3950] : 
                             (N200)? \nz.mem [4030] : 
                             (N202)? \nz.mem [4110] : 
                             (N204)? \nz.mem [4190] : 
                             (N206)? \nz.mem [4270] : 
                             (N208)? \nz.mem [4350] : 
                             (N210)? \nz.mem [4430] : 
                             (N212)? \nz.mem [4510] : 
                             (N214)? \nz.mem [4590] : 
                             (N216)? \nz.mem [4670] : 
                             (N218)? \nz.mem [4750] : 
                             (N220)? \nz.mem [4830] : 
                             (N222)? \nz.mem [4910] : 
                             (N224)? \nz.mem [4990] : 
                             (N226)? \nz.mem [5070] : 1'b0;
  assign \nz.data_out [29] = (N163)? \nz.mem [29] : 
                             (N165)? \nz.mem [109] : 
                             (N167)? \nz.mem [189] : 
                             (N169)? \nz.mem [269] : 
                             (N171)? \nz.mem [349] : 
                             (N173)? \nz.mem [429] : 
                             (N175)? \nz.mem [509] : 
                             (N177)? \nz.mem [589] : 
                             (N179)? \nz.mem [669] : 
                             (N181)? \nz.mem [749] : 
                             (N183)? \nz.mem [829] : 
                             (N185)? \nz.mem [909] : 
                             (N187)? \nz.mem [989] : 
                             (N189)? \nz.mem [1069] : 
                             (N191)? \nz.mem [1149] : 
                             (N193)? \nz.mem [1229] : 
                             (N195)? \nz.mem [1309] : 
                             (N197)? \nz.mem [1389] : 
                             (N199)? \nz.mem [1469] : 
                             (N201)? \nz.mem [1549] : 
                             (N203)? \nz.mem [1629] : 
                             (N205)? \nz.mem [1709] : 
                             (N207)? \nz.mem [1789] : 
                             (N209)? \nz.mem [1869] : 
                             (N211)? \nz.mem [1949] : 
                             (N213)? \nz.mem [2029] : 
                             (N215)? \nz.mem [2109] : 
                             (N217)? \nz.mem [2189] : 
                             (N219)? \nz.mem [2269] : 
                             (N221)? \nz.mem [2349] : 
                             (N223)? \nz.mem [2429] : 
                             (N225)? \nz.mem [2509] : 
                             (N164)? \nz.mem [2589] : 
                             (N166)? \nz.mem [2669] : 
                             (N168)? \nz.mem [2749] : 
                             (N170)? \nz.mem [2829] : 
                             (N172)? \nz.mem [2909] : 
                             (N174)? \nz.mem [2989] : 
                             (N176)? \nz.mem [3069] : 
                             (N178)? \nz.mem [3149] : 
                             (N180)? \nz.mem [3229] : 
                             (N182)? \nz.mem [3309] : 
                             (N184)? \nz.mem [3389] : 
                             (N186)? \nz.mem [3469] : 
                             (N188)? \nz.mem [3549] : 
                             (N190)? \nz.mem [3629] : 
                             (N192)? \nz.mem [3709] : 
                             (N194)? \nz.mem [3789] : 
                             (N196)? \nz.mem [3869] : 
                             (N198)? \nz.mem [3949] : 
                             (N200)? \nz.mem [4029] : 
                             (N202)? \nz.mem [4109] : 
                             (N204)? \nz.mem [4189] : 
                             (N206)? \nz.mem [4269] : 
                             (N208)? \nz.mem [4349] : 
                             (N210)? \nz.mem [4429] : 
                             (N212)? \nz.mem [4509] : 
                             (N214)? \nz.mem [4589] : 
                             (N216)? \nz.mem [4669] : 
                             (N218)? \nz.mem [4749] : 
                             (N220)? \nz.mem [4829] : 
                             (N222)? \nz.mem [4909] : 
                             (N224)? \nz.mem [4989] : 
                             (N226)? \nz.mem [5069] : 1'b0;
  assign \nz.data_out [28] = (N163)? \nz.mem [28] : 
                             (N165)? \nz.mem [108] : 
                             (N167)? \nz.mem [188] : 
                             (N169)? \nz.mem [268] : 
                             (N171)? \nz.mem [348] : 
                             (N173)? \nz.mem [428] : 
                             (N175)? \nz.mem [508] : 
                             (N177)? \nz.mem [588] : 
                             (N179)? \nz.mem [668] : 
                             (N181)? \nz.mem [748] : 
                             (N183)? \nz.mem [828] : 
                             (N185)? \nz.mem [908] : 
                             (N187)? \nz.mem [988] : 
                             (N189)? \nz.mem [1068] : 
                             (N191)? \nz.mem [1148] : 
                             (N193)? \nz.mem [1228] : 
                             (N195)? \nz.mem [1308] : 
                             (N197)? \nz.mem [1388] : 
                             (N199)? \nz.mem [1468] : 
                             (N201)? \nz.mem [1548] : 
                             (N203)? \nz.mem [1628] : 
                             (N205)? \nz.mem [1708] : 
                             (N207)? \nz.mem [1788] : 
                             (N209)? \nz.mem [1868] : 
                             (N211)? \nz.mem [1948] : 
                             (N213)? \nz.mem [2028] : 
                             (N215)? \nz.mem [2108] : 
                             (N217)? \nz.mem [2188] : 
                             (N219)? \nz.mem [2268] : 
                             (N221)? \nz.mem [2348] : 
                             (N223)? \nz.mem [2428] : 
                             (N225)? \nz.mem [2508] : 
                             (N164)? \nz.mem [2588] : 
                             (N166)? \nz.mem [2668] : 
                             (N168)? \nz.mem [2748] : 
                             (N170)? \nz.mem [2828] : 
                             (N172)? \nz.mem [2908] : 
                             (N174)? \nz.mem [2988] : 
                             (N176)? \nz.mem [3068] : 
                             (N178)? \nz.mem [3148] : 
                             (N180)? \nz.mem [3228] : 
                             (N182)? \nz.mem [3308] : 
                             (N184)? \nz.mem [3388] : 
                             (N186)? \nz.mem [3468] : 
                             (N188)? \nz.mem [3548] : 
                             (N190)? \nz.mem [3628] : 
                             (N192)? \nz.mem [3708] : 
                             (N194)? \nz.mem [3788] : 
                             (N196)? \nz.mem [3868] : 
                             (N198)? \nz.mem [3948] : 
                             (N200)? \nz.mem [4028] : 
                             (N202)? \nz.mem [4108] : 
                             (N204)? \nz.mem [4188] : 
                             (N206)? \nz.mem [4268] : 
                             (N208)? \nz.mem [4348] : 
                             (N210)? \nz.mem [4428] : 
                             (N212)? \nz.mem [4508] : 
                             (N214)? \nz.mem [4588] : 
                             (N216)? \nz.mem [4668] : 
                             (N218)? \nz.mem [4748] : 
                             (N220)? \nz.mem [4828] : 
                             (N222)? \nz.mem [4908] : 
                             (N224)? \nz.mem [4988] : 
                             (N226)? \nz.mem [5068] : 1'b0;
  assign \nz.data_out [27] = (N163)? \nz.mem [27] : 
                             (N165)? \nz.mem [107] : 
                             (N167)? \nz.mem [187] : 
                             (N169)? \nz.mem [267] : 
                             (N171)? \nz.mem [347] : 
                             (N173)? \nz.mem [427] : 
                             (N175)? \nz.mem [507] : 
                             (N177)? \nz.mem [587] : 
                             (N179)? \nz.mem [667] : 
                             (N181)? \nz.mem [747] : 
                             (N183)? \nz.mem [827] : 
                             (N185)? \nz.mem [907] : 
                             (N187)? \nz.mem [987] : 
                             (N189)? \nz.mem [1067] : 
                             (N191)? \nz.mem [1147] : 
                             (N193)? \nz.mem [1227] : 
                             (N195)? \nz.mem [1307] : 
                             (N197)? \nz.mem [1387] : 
                             (N199)? \nz.mem [1467] : 
                             (N201)? \nz.mem [1547] : 
                             (N203)? \nz.mem [1627] : 
                             (N205)? \nz.mem [1707] : 
                             (N207)? \nz.mem [1787] : 
                             (N209)? \nz.mem [1867] : 
                             (N211)? \nz.mem [1947] : 
                             (N213)? \nz.mem [2027] : 
                             (N215)? \nz.mem [2107] : 
                             (N217)? \nz.mem [2187] : 
                             (N219)? \nz.mem [2267] : 
                             (N221)? \nz.mem [2347] : 
                             (N223)? \nz.mem [2427] : 
                             (N225)? \nz.mem [2507] : 
                             (N164)? \nz.mem [2587] : 
                             (N166)? \nz.mem [2667] : 
                             (N168)? \nz.mem [2747] : 
                             (N170)? \nz.mem [2827] : 
                             (N172)? \nz.mem [2907] : 
                             (N174)? \nz.mem [2987] : 
                             (N176)? \nz.mem [3067] : 
                             (N178)? \nz.mem [3147] : 
                             (N180)? \nz.mem [3227] : 
                             (N182)? \nz.mem [3307] : 
                             (N184)? \nz.mem [3387] : 
                             (N186)? \nz.mem [3467] : 
                             (N188)? \nz.mem [3547] : 
                             (N190)? \nz.mem [3627] : 
                             (N192)? \nz.mem [3707] : 
                             (N194)? \nz.mem [3787] : 
                             (N196)? \nz.mem [3867] : 
                             (N198)? \nz.mem [3947] : 
                             (N200)? \nz.mem [4027] : 
                             (N202)? \nz.mem [4107] : 
                             (N204)? \nz.mem [4187] : 
                             (N206)? \nz.mem [4267] : 
                             (N208)? \nz.mem [4347] : 
                             (N210)? \nz.mem [4427] : 
                             (N212)? \nz.mem [4507] : 
                             (N214)? \nz.mem [4587] : 
                             (N216)? \nz.mem [4667] : 
                             (N218)? \nz.mem [4747] : 
                             (N220)? \nz.mem [4827] : 
                             (N222)? \nz.mem [4907] : 
                             (N224)? \nz.mem [4987] : 
                             (N226)? \nz.mem [5067] : 1'b0;
  assign \nz.data_out [26] = (N163)? \nz.mem [26] : 
                             (N165)? \nz.mem [106] : 
                             (N167)? \nz.mem [186] : 
                             (N169)? \nz.mem [266] : 
                             (N171)? \nz.mem [346] : 
                             (N173)? \nz.mem [426] : 
                             (N175)? \nz.mem [506] : 
                             (N177)? \nz.mem [586] : 
                             (N179)? \nz.mem [666] : 
                             (N181)? \nz.mem [746] : 
                             (N183)? \nz.mem [826] : 
                             (N185)? \nz.mem [906] : 
                             (N187)? \nz.mem [986] : 
                             (N189)? \nz.mem [1066] : 
                             (N191)? \nz.mem [1146] : 
                             (N193)? \nz.mem [1226] : 
                             (N195)? \nz.mem [1306] : 
                             (N197)? \nz.mem [1386] : 
                             (N199)? \nz.mem [1466] : 
                             (N201)? \nz.mem [1546] : 
                             (N203)? \nz.mem [1626] : 
                             (N205)? \nz.mem [1706] : 
                             (N207)? \nz.mem [1786] : 
                             (N209)? \nz.mem [1866] : 
                             (N211)? \nz.mem [1946] : 
                             (N213)? \nz.mem [2026] : 
                             (N215)? \nz.mem [2106] : 
                             (N217)? \nz.mem [2186] : 
                             (N219)? \nz.mem [2266] : 
                             (N221)? \nz.mem [2346] : 
                             (N223)? \nz.mem [2426] : 
                             (N225)? \nz.mem [2506] : 
                             (N164)? \nz.mem [2586] : 
                             (N166)? \nz.mem [2666] : 
                             (N168)? \nz.mem [2746] : 
                             (N170)? \nz.mem [2826] : 
                             (N172)? \nz.mem [2906] : 
                             (N174)? \nz.mem [2986] : 
                             (N176)? \nz.mem [3066] : 
                             (N178)? \nz.mem [3146] : 
                             (N180)? \nz.mem [3226] : 
                             (N182)? \nz.mem [3306] : 
                             (N184)? \nz.mem [3386] : 
                             (N186)? \nz.mem [3466] : 
                             (N188)? \nz.mem [3546] : 
                             (N190)? \nz.mem [3626] : 
                             (N192)? \nz.mem [3706] : 
                             (N194)? \nz.mem [3786] : 
                             (N196)? \nz.mem [3866] : 
                             (N198)? \nz.mem [3946] : 
                             (N200)? \nz.mem [4026] : 
                             (N202)? \nz.mem [4106] : 
                             (N204)? \nz.mem [4186] : 
                             (N206)? \nz.mem [4266] : 
                             (N208)? \nz.mem [4346] : 
                             (N210)? \nz.mem [4426] : 
                             (N212)? \nz.mem [4506] : 
                             (N214)? \nz.mem [4586] : 
                             (N216)? \nz.mem [4666] : 
                             (N218)? \nz.mem [4746] : 
                             (N220)? \nz.mem [4826] : 
                             (N222)? \nz.mem [4906] : 
                             (N224)? \nz.mem [4986] : 
                             (N226)? \nz.mem [5066] : 1'b0;
  assign \nz.data_out [25] = (N163)? \nz.mem [25] : 
                             (N165)? \nz.mem [105] : 
                             (N167)? \nz.mem [185] : 
                             (N169)? \nz.mem [265] : 
                             (N171)? \nz.mem [345] : 
                             (N173)? \nz.mem [425] : 
                             (N175)? \nz.mem [505] : 
                             (N177)? \nz.mem [585] : 
                             (N179)? \nz.mem [665] : 
                             (N181)? \nz.mem [745] : 
                             (N183)? \nz.mem [825] : 
                             (N185)? \nz.mem [905] : 
                             (N187)? \nz.mem [985] : 
                             (N189)? \nz.mem [1065] : 
                             (N191)? \nz.mem [1145] : 
                             (N193)? \nz.mem [1225] : 
                             (N195)? \nz.mem [1305] : 
                             (N197)? \nz.mem [1385] : 
                             (N199)? \nz.mem [1465] : 
                             (N201)? \nz.mem [1545] : 
                             (N203)? \nz.mem [1625] : 
                             (N205)? \nz.mem [1705] : 
                             (N207)? \nz.mem [1785] : 
                             (N209)? \nz.mem [1865] : 
                             (N211)? \nz.mem [1945] : 
                             (N213)? \nz.mem [2025] : 
                             (N215)? \nz.mem [2105] : 
                             (N217)? \nz.mem [2185] : 
                             (N219)? \nz.mem [2265] : 
                             (N221)? \nz.mem [2345] : 
                             (N223)? \nz.mem [2425] : 
                             (N225)? \nz.mem [2505] : 
                             (N164)? \nz.mem [2585] : 
                             (N166)? \nz.mem [2665] : 
                             (N168)? \nz.mem [2745] : 
                             (N170)? \nz.mem [2825] : 
                             (N172)? \nz.mem [2905] : 
                             (N174)? \nz.mem [2985] : 
                             (N176)? \nz.mem [3065] : 
                             (N178)? \nz.mem [3145] : 
                             (N180)? \nz.mem [3225] : 
                             (N182)? \nz.mem [3305] : 
                             (N184)? \nz.mem [3385] : 
                             (N186)? \nz.mem [3465] : 
                             (N188)? \nz.mem [3545] : 
                             (N190)? \nz.mem [3625] : 
                             (N192)? \nz.mem [3705] : 
                             (N194)? \nz.mem [3785] : 
                             (N196)? \nz.mem [3865] : 
                             (N198)? \nz.mem [3945] : 
                             (N200)? \nz.mem [4025] : 
                             (N202)? \nz.mem [4105] : 
                             (N204)? \nz.mem [4185] : 
                             (N206)? \nz.mem [4265] : 
                             (N208)? \nz.mem [4345] : 
                             (N210)? \nz.mem [4425] : 
                             (N212)? \nz.mem [4505] : 
                             (N214)? \nz.mem [4585] : 
                             (N216)? \nz.mem [4665] : 
                             (N218)? \nz.mem [4745] : 
                             (N220)? \nz.mem [4825] : 
                             (N222)? \nz.mem [4905] : 
                             (N224)? \nz.mem [4985] : 
                             (N226)? \nz.mem [5065] : 1'b0;
  assign \nz.data_out [24] = (N163)? \nz.mem [24] : 
                             (N165)? \nz.mem [104] : 
                             (N167)? \nz.mem [184] : 
                             (N169)? \nz.mem [264] : 
                             (N171)? \nz.mem [344] : 
                             (N173)? \nz.mem [424] : 
                             (N175)? \nz.mem [504] : 
                             (N177)? \nz.mem [584] : 
                             (N179)? \nz.mem [664] : 
                             (N181)? \nz.mem [744] : 
                             (N183)? \nz.mem [824] : 
                             (N185)? \nz.mem [904] : 
                             (N187)? \nz.mem [984] : 
                             (N189)? \nz.mem [1064] : 
                             (N191)? \nz.mem [1144] : 
                             (N193)? \nz.mem [1224] : 
                             (N195)? \nz.mem [1304] : 
                             (N197)? \nz.mem [1384] : 
                             (N199)? \nz.mem [1464] : 
                             (N201)? \nz.mem [1544] : 
                             (N203)? \nz.mem [1624] : 
                             (N205)? \nz.mem [1704] : 
                             (N207)? \nz.mem [1784] : 
                             (N209)? \nz.mem [1864] : 
                             (N211)? \nz.mem [1944] : 
                             (N213)? \nz.mem [2024] : 
                             (N215)? \nz.mem [2104] : 
                             (N217)? \nz.mem [2184] : 
                             (N219)? \nz.mem [2264] : 
                             (N221)? \nz.mem [2344] : 
                             (N223)? \nz.mem [2424] : 
                             (N225)? \nz.mem [2504] : 
                             (N164)? \nz.mem [2584] : 
                             (N166)? \nz.mem [2664] : 
                             (N168)? \nz.mem [2744] : 
                             (N170)? \nz.mem [2824] : 
                             (N172)? \nz.mem [2904] : 
                             (N174)? \nz.mem [2984] : 
                             (N176)? \nz.mem [3064] : 
                             (N178)? \nz.mem [3144] : 
                             (N180)? \nz.mem [3224] : 
                             (N182)? \nz.mem [3304] : 
                             (N184)? \nz.mem [3384] : 
                             (N186)? \nz.mem [3464] : 
                             (N188)? \nz.mem [3544] : 
                             (N190)? \nz.mem [3624] : 
                             (N192)? \nz.mem [3704] : 
                             (N194)? \nz.mem [3784] : 
                             (N196)? \nz.mem [3864] : 
                             (N198)? \nz.mem [3944] : 
                             (N200)? \nz.mem [4024] : 
                             (N202)? \nz.mem [4104] : 
                             (N204)? \nz.mem [4184] : 
                             (N206)? \nz.mem [4264] : 
                             (N208)? \nz.mem [4344] : 
                             (N210)? \nz.mem [4424] : 
                             (N212)? \nz.mem [4504] : 
                             (N214)? \nz.mem [4584] : 
                             (N216)? \nz.mem [4664] : 
                             (N218)? \nz.mem [4744] : 
                             (N220)? \nz.mem [4824] : 
                             (N222)? \nz.mem [4904] : 
                             (N224)? \nz.mem [4984] : 
                             (N226)? \nz.mem [5064] : 1'b0;
  assign \nz.data_out [23] = (N163)? \nz.mem [23] : 
                             (N165)? \nz.mem [103] : 
                             (N167)? \nz.mem [183] : 
                             (N169)? \nz.mem [263] : 
                             (N171)? \nz.mem [343] : 
                             (N173)? \nz.mem [423] : 
                             (N175)? \nz.mem [503] : 
                             (N177)? \nz.mem [583] : 
                             (N179)? \nz.mem [663] : 
                             (N181)? \nz.mem [743] : 
                             (N183)? \nz.mem [823] : 
                             (N185)? \nz.mem [903] : 
                             (N187)? \nz.mem [983] : 
                             (N189)? \nz.mem [1063] : 
                             (N191)? \nz.mem [1143] : 
                             (N193)? \nz.mem [1223] : 
                             (N195)? \nz.mem [1303] : 
                             (N197)? \nz.mem [1383] : 
                             (N199)? \nz.mem [1463] : 
                             (N201)? \nz.mem [1543] : 
                             (N203)? \nz.mem [1623] : 
                             (N205)? \nz.mem [1703] : 
                             (N207)? \nz.mem [1783] : 
                             (N209)? \nz.mem [1863] : 
                             (N211)? \nz.mem [1943] : 
                             (N213)? \nz.mem [2023] : 
                             (N215)? \nz.mem [2103] : 
                             (N217)? \nz.mem [2183] : 
                             (N219)? \nz.mem [2263] : 
                             (N221)? \nz.mem [2343] : 
                             (N223)? \nz.mem [2423] : 
                             (N225)? \nz.mem [2503] : 
                             (N164)? \nz.mem [2583] : 
                             (N166)? \nz.mem [2663] : 
                             (N168)? \nz.mem [2743] : 
                             (N170)? \nz.mem [2823] : 
                             (N172)? \nz.mem [2903] : 
                             (N174)? \nz.mem [2983] : 
                             (N176)? \nz.mem [3063] : 
                             (N178)? \nz.mem [3143] : 
                             (N180)? \nz.mem [3223] : 
                             (N182)? \nz.mem [3303] : 
                             (N184)? \nz.mem [3383] : 
                             (N186)? \nz.mem [3463] : 
                             (N188)? \nz.mem [3543] : 
                             (N190)? \nz.mem [3623] : 
                             (N192)? \nz.mem [3703] : 
                             (N194)? \nz.mem [3783] : 
                             (N196)? \nz.mem [3863] : 
                             (N198)? \nz.mem [3943] : 
                             (N200)? \nz.mem [4023] : 
                             (N202)? \nz.mem [4103] : 
                             (N204)? \nz.mem [4183] : 
                             (N206)? \nz.mem [4263] : 
                             (N208)? \nz.mem [4343] : 
                             (N210)? \nz.mem [4423] : 
                             (N212)? \nz.mem [4503] : 
                             (N214)? \nz.mem [4583] : 
                             (N216)? \nz.mem [4663] : 
                             (N218)? \nz.mem [4743] : 
                             (N220)? \nz.mem [4823] : 
                             (N222)? \nz.mem [4903] : 
                             (N224)? \nz.mem [4983] : 
                             (N226)? \nz.mem [5063] : 1'b0;
  assign \nz.data_out [22] = (N163)? \nz.mem [22] : 
                             (N165)? \nz.mem [102] : 
                             (N167)? \nz.mem [182] : 
                             (N169)? \nz.mem [262] : 
                             (N171)? \nz.mem [342] : 
                             (N173)? \nz.mem [422] : 
                             (N175)? \nz.mem [502] : 
                             (N177)? \nz.mem [582] : 
                             (N179)? \nz.mem [662] : 
                             (N181)? \nz.mem [742] : 
                             (N183)? \nz.mem [822] : 
                             (N185)? \nz.mem [902] : 
                             (N187)? \nz.mem [982] : 
                             (N189)? \nz.mem [1062] : 
                             (N191)? \nz.mem [1142] : 
                             (N193)? \nz.mem [1222] : 
                             (N195)? \nz.mem [1302] : 
                             (N197)? \nz.mem [1382] : 
                             (N199)? \nz.mem [1462] : 
                             (N201)? \nz.mem [1542] : 
                             (N203)? \nz.mem [1622] : 
                             (N205)? \nz.mem [1702] : 
                             (N207)? \nz.mem [1782] : 
                             (N209)? \nz.mem [1862] : 
                             (N211)? \nz.mem [1942] : 
                             (N213)? \nz.mem [2022] : 
                             (N215)? \nz.mem [2102] : 
                             (N217)? \nz.mem [2182] : 
                             (N219)? \nz.mem [2262] : 
                             (N221)? \nz.mem [2342] : 
                             (N223)? \nz.mem [2422] : 
                             (N225)? \nz.mem [2502] : 
                             (N164)? \nz.mem [2582] : 
                             (N166)? \nz.mem [2662] : 
                             (N168)? \nz.mem [2742] : 
                             (N170)? \nz.mem [2822] : 
                             (N172)? \nz.mem [2902] : 
                             (N174)? \nz.mem [2982] : 
                             (N176)? \nz.mem [3062] : 
                             (N178)? \nz.mem [3142] : 
                             (N180)? \nz.mem [3222] : 
                             (N182)? \nz.mem [3302] : 
                             (N184)? \nz.mem [3382] : 
                             (N186)? \nz.mem [3462] : 
                             (N188)? \nz.mem [3542] : 
                             (N190)? \nz.mem [3622] : 
                             (N192)? \nz.mem [3702] : 
                             (N194)? \nz.mem [3782] : 
                             (N196)? \nz.mem [3862] : 
                             (N198)? \nz.mem [3942] : 
                             (N200)? \nz.mem [4022] : 
                             (N202)? \nz.mem [4102] : 
                             (N204)? \nz.mem [4182] : 
                             (N206)? \nz.mem [4262] : 
                             (N208)? \nz.mem [4342] : 
                             (N210)? \nz.mem [4422] : 
                             (N212)? \nz.mem [4502] : 
                             (N214)? \nz.mem [4582] : 
                             (N216)? \nz.mem [4662] : 
                             (N218)? \nz.mem [4742] : 
                             (N220)? \nz.mem [4822] : 
                             (N222)? \nz.mem [4902] : 
                             (N224)? \nz.mem [4982] : 
                             (N226)? \nz.mem [5062] : 1'b0;
  assign \nz.data_out [21] = (N163)? \nz.mem [21] : 
                             (N165)? \nz.mem [101] : 
                             (N167)? \nz.mem [181] : 
                             (N169)? \nz.mem [261] : 
                             (N171)? \nz.mem [341] : 
                             (N173)? \nz.mem [421] : 
                             (N175)? \nz.mem [501] : 
                             (N177)? \nz.mem [581] : 
                             (N179)? \nz.mem [661] : 
                             (N181)? \nz.mem [741] : 
                             (N183)? \nz.mem [821] : 
                             (N185)? \nz.mem [901] : 
                             (N187)? \nz.mem [981] : 
                             (N189)? \nz.mem [1061] : 
                             (N191)? \nz.mem [1141] : 
                             (N193)? \nz.mem [1221] : 
                             (N195)? \nz.mem [1301] : 
                             (N197)? \nz.mem [1381] : 
                             (N199)? \nz.mem [1461] : 
                             (N201)? \nz.mem [1541] : 
                             (N203)? \nz.mem [1621] : 
                             (N205)? \nz.mem [1701] : 
                             (N207)? \nz.mem [1781] : 
                             (N209)? \nz.mem [1861] : 
                             (N211)? \nz.mem [1941] : 
                             (N213)? \nz.mem [2021] : 
                             (N215)? \nz.mem [2101] : 
                             (N217)? \nz.mem [2181] : 
                             (N219)? \nz.mem [2261] : 
                             (N221)? \nz.mem [2341] : 
                             (N223)? \nz.mem [2421] : 
                             (N225)? \nz.mem [2501] : 
                             (N164)? \nz.mem [2581] : 
                             (N166)? \nz.mem [2661] : 
                             (N168)? \nz.mem [2741] : 
                             (N170)? \nz.mem [2821] : 
                             (N172)? \nz.mem [2901] : 
                             (N174)? \nz.mem [2981] : 
                             (N176)? \nz.mem [3061] : 
                             (N178)? \nz.mem [3141] : 
                             (N180)? \nz.mem [3221] : 
                             (N182)? \nz.mem [3301] : 
                             (N184)? \nz.mem [3381] : 
                             (N186)? \nz.mem [3461] : 
                             (N188)? \nz.mem [3541] : 
                             (N190)? \nz.mem [3621] : 
                             (N192)? \nz.mem [3701] : 
                             (N194)? \nz.mem [3781] : 
                             (N196)? \nz.mem [3861] : 
                             (N198)? \nz.mem [3941] : 
                             (N200)? \nz.mem [4021] : 
                             (N202)? \nz.mem [4101] : 
                             (N204)? \nz.mem [4181] : 
                             (N206)? \nz.mem [4261] : 
                             (N208)? \nz.mem [4341] : 
                             (N210)? \nz.mem [4421] : 
                             (N212)? \nz.mem [4501] : 
                             (N214)? \nz.mem [4581] : 
                             (N216)? \nz.mem [4661] : 
                             (N218)? \nz.mem [4741] : 
                             (N220)? \nz.mem [4821] : 
                             (N222)? \nz.mem [4901] : 
                             (N224)? \nz.mem [4981] : 
                             (N226)? \nz.mem [5061] : 1'b0;
  assign \nz.data_out [20] = (N163)? \nz.mem [20] : 
                             (N165)? \nz.mem [100] : 
                             (N167)? \nz.mem [180] : 
                             (N169)? \nz.mem [260] : 
                             (N171)? \nz.mem [340] : 
                             (N173)? \nz.mem [420] : 
                             (N175)? \nz.mem [500] : 
                             (N177)? \nz.mem [580] : 
                             (N179)? \nz.mem [660] : 
                             (N181)? \nz.mem [740] : 
                             (N183)? \nz.mem [820] : 
                             (N185)? \nz.mem [900] : 
                             (N187)? \nz.mem [980] : 
                             (N189)? \nz.mem [1060] : 
                             (N191)? \nz.mem [1140] : 
                             (N193)? \nz.mem [1220] : 
                             (N195)? \nz.mem [1300] : 
                             (N197)? \nz.mem [1380] : 
                             (N199)? \nz.mem [1460] : 
                             (N201)? \nz.mem [1540] : 
                             (N203)? \nz.mem [1620] : 
                             (N205)? \nz.mem [1700] : 
                             (N207)? \nz.mem [1780] : 
                             (N209)? \nz.mem [1860] : 
                             (N211)? \nz.mem [1940] : 
                             (N213)? \nz.mem [2020] : 
                             (N215)? \nz.mem [2100] : 
                             (N217)? \nz.mem [2180] : 
                             (N219)? \nz.mem [2260] : 
                             (N221)? \nz.mem [2340] : 
                             (N223)? \nz.mem [2420] : 
                             (N225)? \nz.mem [2500] : 
                             (N164)? \nz.mem [2580] : 
                             (N166)? \nz.mem [2660] : 
                             (N168)? \nz.mem [2740] : 
                             (N170)? \nz.mem [2820] : 
                             (N172)? \nz.mem [2900] : 
                             (N174)? \nz.mem [2980] : 
                             (N176)? \nz.mem [3060] : 
                             (N178)? \nz.mem [3140] : 
                             (N180)? \nz.mem [3220] : 
                             (N182)? \nz.mem [3300] : 
                             (N184)? \nz.mem [3380] : 
                             (N186)? \nz.mem [3460] : 
                             (N188)? \nz.mem [3540] : 
                             (N190)? \nz.mem [3620] : 
                             (N192)? \nz.mem [3700] : 
                             (N194)? \nz.mem [3780] : 
                             (N196)? \nz.mem [3860] : 
                             (N198)? \nz.mem [3940] : 
                             (N200)? \nz.mem [4020] : 
                             (N202)? \nz.mem [4100] : 
                             (N204)? \nz.mem [4180] : 
                             (N206)? \nz.mem [4260] : 
                             (N208)? \nz.mem [4340] : 
                             (N210)? \nz.mem [4420] : 
                             (N212)? \nz.mem [4500] : 
                             (N214)? \nz.mem [4580] : 
                             (N216)? \nz.mem [4660] : 
                             (N218)? \nz.mem [4740] : 
                             (N220)? \nz.mem [4820] : 
                             (N222)? \nz.mem [4900] : 
                             (N224)? \nz.mem [4980] : 
                             (N226)? \nz.mem [5060] : 1'b0;
  assign \nz.data_out [19] = (N163)? \nz.mem [19] : 
                             (N165)? \nz.mem [99] : 
                             (N167)? \nz.mem [179] : 
                             (N169)? \nz.mem [259] : 
                             (N171)? \nz.mem [339] : 
                             (N173)? \nz.mem [419] : 
                             (N175)? \nz.mem [499] : 
                             (N177)? \nz.mem [579] : 
                             (N179)? \nz.mem [659] : 
                             (N181)? \nz.mem [739] : 
                             (N183)? \nz.mem [819] : 
                             (N185)? \nz.mem [899] : 
                             (N187)? \nz.mem [979] : 
                             (N189)? \nz.mem [1059] : 
                             (N191)? \nz.mem [1139] : 
                             (N193)? \nz.mem [1219] : 
                             (N195)? \nz.mem [1299] : 
                             (N197)? \nz.mem [1379] : 
                             (N199)? \nz.mem [1459] : 
                             (N201)? \nz.mem [1539] : 
                             (N203)? \nz.mem [1619] : 
                             (N205)? \nz.mem [1699] : 
                             (N207)? \nz.mem [1779] : 
                             (N209)? \nz.mem [1859] : 
                             (N211)? \nz.mem [1939] : 
                             (N213)? \nz.mem [2019] : 
                             (N215)? \nz.mem [2099] : 
                             (N217)? \nz.mem [2179] : 
                             (N219)? \nz.mem [2259] : 
                             (N221)? \nz.mem [2339] : 
                             (N223)? \nz.mem [2419] : 
                             (N225)? \nz.mem [2499] : 
                             (N164)? \nz.mem [2579] : 
                             (N166)? \nz.mem [2659] : 
                             (N168)? \nz.mem [2739] : 
                             (N170)? \nz.mem [2819] : 
                             (N172)? \nz.mem [2899] : 
                             (N174)? \nz.mem [2979] : 
                             (N176)? \nz.mem [3059] : 
                             (N178)? \nz.mem [3139] : 
                             (N180)? \nz.mem [3219] : 
                             (N182)? \nz.mem [3299] : 
                             (N184)? \nz.mem [3379] : 
                             (N186)? \nz.mem [3459] : 
                             (N188)? \nz.mem [3539] : 
                             (N190)? \nz.mem [3619] : 
                             (N192)? \nz.mem [3699] : 
                             (N194)? \nz.mem [3779] : 
                             (N196)? \nz.mem [3859] : 
                             (N198)? \nz.mem [3939] : 
                             (N200)? \nz.mem [4019] : 
                             (N202)? \nz.mem [4099] : 
                             (N204)? \nz.mem [4179] : 
                             (N206)? \nz.mem [4259] : 
                             (N208)? \nz.mem [4339] : 
                             (N210)? \nz.mem [4419] : 
                             (N212)? \nz.mem [4499] : 
                             (N214)? \nz.mem [4579] : 
                             (N216)? \nz.mem [4659] : 
                             (N218)? \nz.mem [4739] : 
                             (N220)? \nz.mem [4819] : 
                             (N222)? \nz.mem [4899] : 
                             (N224)? \nz.mem [4979] : 
                             (N226)? \nz.mem [5059] : 1'b0;
  assign \nz.data_out [18] = (N163)? \nz.mem [18] : 
                             (N165)? \nz.mem [98] : 
                             (N167)? \nz.mem [178] : 
                             (N169)? \nz.mem [258] : 
                             (N171)? \nz.mem [338] : 
                             (N173)? \nz.mem [418] : 
                             (N175)? \nz.mem [498] : 
                             (N177)? \nz.mem [578] : 
                             (N179)? \nz.mem [658] : 
                             (N181)? \nz.mem [738] : 
                             (N183)? \nz.mem [818] : 
                             (N185)? \nz.mem [898] : 
                             (N187)? \nz.mem [978] : 
                             (N189)? \nz.mem [1058] : 
                             (N191)? \nz.mem [1138] : 
                             (N193)? \nz.mem [1218] : 
                             (N195)? \nz.mem [1298] : 
                             (N197)? \nz.mem [1378] : 
                             (N199)? \nz.mem [1458] : 
                             (N201)? \nz.mem [1538] : 
                             (N203)? \nz.mem [1618] : 
                             (N205)? \nz.mem [1698] : 
                             (N207)? \nz.mem [1778] : 
                             (N209)? \nz.mem [1858] : 
                             (N211)? \nz.mem [1938] : 
                             (N213)? \nz.mem [2018] : 
                             (N215)? \nz.mem [2098] : 
                             (N217)? \nz.mem [2178] : 
                             (N219)? \nz.mem [2258] : 
                             (N221)? \nz.mem [2338] : 
                             (N223)? \nz.mem [2418] : 
                             (N225)? \nz.mem [2498] : 
                             (N164)? \nz.mem [2578] : 
                             (N166)? \nz.mem [2658] : 
                             (N168)? \nz.mem [2738] : 
                             (N170)? \nz.mem [2818] : 
                             (N172)? \nz.mem [2898] : 
                             (N174)? \nz.mem [2978] : 
                             (N176)? \nz.mem [3058] : 
                             (N178)? \nz.mem [3138] : 
                             (N180)? \nz.mem [3218] : 
                             (N182)? \nz.mem [3298] : 
                             (N184)? \nz.mem [3378] : 
                             (N186)? \nz.mem [3458] : 
                             (N188)? \nz.mem [3538] : 
                             (N190)? \nz.mem [3618] : 
                             (N192)? \nz.mem [3698] : 
                             (N194)? \nz.mem [3778] : 
                             (N196)? \nz.mem [3858] : 
                             (N198)? \nz.mem [3938] : 
                             (N200)? \nz.mem [4018] : 
                             (N202)? \nz.mem [4098] : 
                             (N204)? \nz.mem [4178] : 
                             (N206)? \nz.mem [4258] : 
                             (N208)? \nz.mem [4338] : 
                             (N210)? \nz.mem [4418] : 
                             (N212)? \nz.mem [4498] : 
                             (N214)? \nz.mem [4578] : 
                             (N216)? \nz.mem [4658] : 
                             (N218)? \nz.mem [4738] : 
                             (N220)? \nz.mem [4818] : 
                             (N222)? \nz.mem [4898] : 
                             (N224)? \nz.mem [4978] : 
                             (N226)? \nz.mem [5058] : 1'b0;
  assign \nz.data_out [17] = (N163)? \nz.mem [17] : 
                             (N165)? \nz.mem [97] : 
                             (N167)? \nz.mem [177] : 
                             (N169)? \nz.mem [257] : 
                             (N171)? \nz.mem [337] : 
                             (N173)? \nz.mem [417] : 
                             (N175)? \nz.mem [497] : 
                             (N177)? \nz.mem [577] : 
                             (N179)? \nz.mem [657] : 
                             (N181)? \nz.mem [737] : 
                             (N183)? \nz.mem [817] : 
                             (N185)? \nz.mem [897] : 
                             (N187)? \nz.mem [977] : 
                             (N189)? \nz.mem [1057] : 
                             (N191)? \nz.mem [1137] : 
                             (N193)? \nz.mem [1217] : 
                             (N195)? \nz.mem [1297] : 
                             (N197)? \nz.mem [1377] : 
                             (N199)? \nz.mem [1457] : 
                             (N201)? \nz.mem [1537] : 
                             (N203)? \nz.mem [1617] : 
                             (N205)? \nz.mem [1697] : 
                             (N207)? \nz.mem [1777] : 
                             (N209)? \nz.mem [1857] : 
                             (N211)? \nz.mem [1937] : 
                             (N213)? \nz.mem [2017] : 
                             (N215)? \nz.mem [2097] : 
                             (N217)? \nz.mem [2177] : 
                             (N219)? \nz.mem [2257] : 
                             (N221)? \nz.mem [2337] : 
                             (N223)? \nz.mem [2417] : 
                             (N225)? \nz.mem [2497] : 
                             (N164)? \nz.mem [2577] : 
                             (N166)? \nz.mem [2657] : 
                             (N168)? \nz.mem [2737] : 
                             (N170)? \nz.mem [2817] : 
                             (N172)? \nz.mem [2897] : 
                             (N174)? \nz.mem [2977] : 
                             (N176)? \nz.mem [3057] : 
                             (N178)? \nz.mem [3137] : 
                             (N180)? \nz.mem [3217] : 
                             (N182)? \nz.mem [3297] : 
                             (N184)? \nz.mem [3377] : 
                             (N186)? \nz.mem [3457] : 
                             (N188)? \nz.mem [3537] : 
                             (N190)? \nz.mem [3617] : 
                             (N192)? \nz.mem [3697] : 
                             (N194)? \nz.mem [3777] : 
                             (N196)? \nz.mem [3857] : 
                             (N198)? \nz.mem [3937] : 
                             (N200)? \nz.mem [4017] : 
                             (N202)? \nz.mem [4097] : 
                             (N204)? \nz.mem [4177] : 
                             (N206)? \nz.mem [4257] : 
                             (N208)? \nz.mem [4337] : 
                             (N210)? \nz.mem [4417] : 
                             (N212)? \nz.mem [4497] : 
                             (N214)? \nz.mem [4577] : 
                             (N216)? \nz.mem [4657] : 
                             (N218)? \nz.mem [4737] : 
                             (N220)? \nz.mem [4817] : 
                             (N222)? \nz.mem [4897] : 
                             (N224)? \nz.mem [4977] : 
                             (N226)? \nz.mem [5057] : 1'b0;
  assign \nz.data_out [16] = (N163)? \nz.mem [16] : 
                             (N165)? \nz.mem [96] : 
                             (N167)? \nz.mem [176] : 
                             (N169)? \nz.mem [256] : 
                             (N171)? \nz.mem [336] : 
                             (N173)? \nz.mem [416] : 
                             (N175)? \nz.mem [496] : 
                             (N177)? \nz.mem [576] : 
                             (N179)? \nz.mem [656] : 
                             (N181)? \nz.mem [736] : 
                             (N183)? \nz.mem [816] : 
                             (N185)? \nz.mem [896] : 
                             (N187)? \nz.mem [976] : 
                             (N189)? \nz.mem [1056] : 
                             (N191)? \nz.mem [1136] : 
                             (N193)? \nz.mem [1216] : 
                             (N195)? \nz.mem [1296] : 
                             (N197)? \nz.mem [1376] : 
                             (N199)? \nz.mem [1456] : 
                             (N201)? \nz.mem [1536] : 
                             (N203)? \nz.mem [1616] : 
                             (N205)? \nz.mem [1696] : 
                             (N207)? \nz.mem [1776] : 
                             (N209)? \nz.mem [1856] : 
                             (N211)? \nz.mem [1936] : 
                             (N213)? \nz.mem [2016] : 
                             (N215)? \nz.mem [2096] : 
                             (N217)? \nz.mem [2176] : 
                             (N219)? \nz.mem [2256] : 
                             (N221)? \nz.mem [2336] : 
                             (N223)? \nz.mem [2416] : 
                             (N225)? \nz.mem [2496] : 
                             (N164)? \nz.mem [2576] : 
                             (N166)? \nz.mem [2656] : 
                             (N168)? \nz.mem [2736] : 
                             (N170)? \nz.mem [2816] : 
                             (N172)? \nz.mem [2896] : 
                             (N174)? \nz.mem [2976] : 
                             (N176)? \nz.mem [3056] : 
                             (N178)? \nz.mem [3136] : 
                             (N180)? \nz.mem [3216] : 
                             (N182)? \nz.mem [3296] : 
                             (N184)? \nz.mem [3376] : 
                             (N186)? \nz.mem [3456] : 
                             (N188)? \nz.mem [3536] : 
                             (N190)? \nz.mem [3616] : 
                             (N192)? \nz.mem [3696] : 
                             (N194)? \nz.mem [3776] : 
                             (N196)? \nz.mem [3856] : 
                             (N198)? \nz.mem [3936] : 
                             (N200)? \nz.mem [4016] : 
                             (N202)? \nz.mem [4096] : 
                             (N204)? \nz.mem [4176] : 
                             (N206)? \nz.mem [4256] : 
                             (N208)? \nz.mem [4336] : 
                             (N210)? \nz.mem [4416] : 
                             (N212)? \nz.mem [4496] : 
                             (N214)? \nz.mem [4576] : 
                             (N216)? \nz.mem [4656] : 
                             (N218)? \nz.mem [4736] : 
                             (N220)? \nz.mem [4816] : 
                             (N222)? \nz.mem [4896] : 
                             (N224)? \nz.mem [4976] : 
                             (N226)? \nz.mem [5056] : 1'b0;
  assign \nz.data_out [15] = (N163)? \nz.mem [15] : 
                             (N165)? \nz.mem [95] : 
                             (N167)? \nz.mem [175] : 
                             (N169)? \nz.mem [255] : 
                             (N171)? \nz.mem [335] : 
                             (N173)? \nz.mem [415] : 
                             (N175)? \nz.mem [495] : 
                             (N177)? \nz.mem [575] : 
                             (N179)? \nz.mem [655] : 
                             (N181)? \nz.mem [735] : 
                             (N183)? \nz.mem [815] : 
                             (N185)? \nz.mem [895] : 
                             (N187)? \nz.mem [975] : 
                             (N189)? \nz.mem [1055] : 
                             (N191)? \nz.mem [1135] : 
                             (N193)? \nz.mem [1215] : 
                             (N195)? \nz.mem [1295] : 
                             (N197)? \nz.mem [1375] : 
                             (N199)? \nz.mem [1455] : 
                             (N201)? \nz.mem [1535] : 
                             (N203)? \nz.mem [1615] : 
                             (N205)? \nz.mem [1695] : 
                             (N207)? \nz.mem [1775] : 
                             (N209)? \nz.mem [1855] : 
                             (N211)? \nz.mem [1935] : 
                             (N213)? \nz.mem [2015] : 
                             (N215)? \nz.mem [2095] : 
                             (N217)? \nz.mem [2175] : 
                             (N219)? \nz.mem [2255] : 
                             (N221)? \nz.mem [2335] : 
                             (N223)? \nz.mem [2415] : 
                             (N225)? \nz.mem [2495] : 
                             (N164)? \nz.mem [2575] : 
                             (N166)? \nz.mem [2655] : 
                             (N168)? \nz.mem [2735] : 
                             (N170)? \nz.mem [2815] : 
                             (N172)? \nz.mem [2895] : 
                             (N174)? \nz.mem [2975] : 
                             (N176)? \nz.mem [3055] : 
                             (N178)? \nz.mem [3135] : 
                             (N180)? \nz.mem [3215] : 
                             (N182)? \nz.mem [3295] : 
                             (N184)? \nz.mem [3375] : 
                             (N186)? \nz.mem [3455] : 
                             (N188)? \nz.mem [3535] : 
                             (N190)? \nz.mem [3615] : 
                             (N192)? \nz.mem [3695] : 
                             (N194)? \nz.mem [3775] : 
                             (N196)? \nz.mem [3855] : 
                             (N198)? \nz.mem [3935] : 
                             (N200)? \nz.mem [4015] : 
                             (N202)? \nz.mem [4095] : 
                             (N204)? \nz.mem [4175] : 
                             (N206)? \nz.mem [4255] : 
                             (N208)? \nz.mem [4335] : 
                             (N210)? \nz.mem [4415] : 
                             (N212)? \nz.mem [4495] : 
                             (N214)? \nz.mem [4575] : 
                             (N216)? \nz.mem [4655] : 
                             (N218)? \nz.mem [4735] : 
                             (N220)? \nz.mem [4815] : 
                             (N222)? \nz.mem [4895] : 
                             (N224)? \nz.mem [4975] : 
                             (N226)? \nz.mem [5055] : 1'b0;
  assign \nz.data_out [14] = (N163)? \nz.mem [14] : 
                             (N165)? \nz.mem [94] : 
                             (N167)? \nz.mem [174] : 
                             (N169)? \nz.mem [254] : 
                             (N171)? \nz.mem [334] : 
                             (N173)? \nz.mem [414] : 
                             (N175)? \nz.mem [494] : 
                             (N177)? \nz.mem [574] : 
                             (N179)? \nz.mem [654] : 
                             (N181)? \nz.mem [734] : 
                             (N183)? \nz.mem [814] : 
                             (N185)? \nz.mem [894] : 
                             (N187)? \nz.mem [974] : 
                             (N189)? \nz.mem [1054] : 
                             (N191)? \nz.mem [1134] : 
                             (N193)? \nz.mem [1214] : 
                             (N195)? \nz.mem [1294] : 
                             (N197)? \nz.mem [1374] : 
                             (N199)? \nz.mem [1454] : 
                             (N201)? \nz.mem [1534] : 
                             (N203)? \nz.mem [1614] : 
                             (N205)? \nz.mem [1694] : 
                             (N207)? \nz.mem [1774] : 
                             (N209)? \nz.mem [1854] : 
                             (N211)? \nz.mem [1934] : 
                             (N213)? \nz.mem [2014] : 
                             (N215)? \nz.mem [2094] : 
                             (N217)? \nz.mem [2174] : 
                             (N219)? \nz.mem [2254] : 
                             (N221)? \nz.mem [2334] : 
                             (N223)? \nz.mem [2414] : 
                             (N225)? \nz.mem [2494] : 
                             (N164)? \nz.mem [2574] : 
                             (N166)? \nz.mem [2654] : 
                             (N168)? \nz.mem [2734] : 
                             (N170)? \nz.mem [2814] : 
                             (N172)? \nz.mem [2894] : 
                             (N174)? \nz.mem [2974] : 
                             (N176)? \nz.mem [3054] : 
                             (N178)? \nz.mem [3134] : 
                             (N180)? \nz.mem [3214] : 
                             (N182)? \nz.mem [3294] : 
                             (N184)? \nz.mem [3374] : 
                             (N186)? \nz.mem [3454] : 
                             (N188)? \nz.mem [3534] : 
                             (N190)? \nz.mem [3614] : 
                             (N192)? \nz.mem [3694] : 
                             (N194)? \nz.mem [3774] : 
                             (N196)? \nz.mem [3854] : 
                             (N198)? \nz.mem [3934] : 
                             (N200)? \nz.mem [4014] : 
                             (N202)? \nz.mem [4094] : 
                             (N204)? \nz.mem [4174] : 
                             (N206)? \nz.mem [4254] : 
                             (N208)? \nz.mem [4334] : 
                             (N210)? \nz.mem [4414] : 
                             (N212)? \nz.mem [4494] : 
                             (N214)? \nz.mem [4574] : 
                             (N216)? \nz.mem [4654] : 
                             (N218)? \nz.mem [4734] : 
                             (N220)? \nz.mem [4814] : 
                             (N222)? \nz.mem [4894] : 
                             (N224)? \nz.mem [4974] : 
                             (N226)? \nz.mem [5054] : 1'b0;
  assign \nz.data_out [13] = (N163)? \nz.mem [13] : 
                             (N165)? \nz.mem [93] : 
                             (N167)? \nz.mem [173] : 
                             (N169)? \nz.mem [253] : 
                             (N171)? \nz.mem [333] : 
                             (N173)? \nz.mem [413] : 
                             (N175)? \nz.mem [493] : 
                             (N177)? \nz.mem [573] : 
                             (N179)? \nz.mem [653] : 
                             (N181)? \nz.mem [733] : 
                             (N183)? \nz.mem [813] : 
                             (N185)? \nz.mem [893] : 
                             (N187)? \nz.mem [973] : 
                             (N189)? \nz.mem [1053] : 
                             (N191)? \nz.mem [1133] : 
                             (N193)? \nz.mem [1213] : 
                             (N195)? \nz.mem [1293] : 
                             (N197)? \nz.mem [1373] : 
                             (N199)? \nz.mem [1453] : 
                             (N201)? \nz.mem [1533] : 
                             (N203)? \nz.mem [1613] : 
                             (N205)? \nz.mem [1693] : 
                             (N207)? \nz.mem [1773] : 
                             (N209)? \nz.mem [1853] : 
                             (N211)? \nz.mem [1933] : 
                             (N213)? \nz.mem [2013] : 
                             (N215)? \nz.mem [2093] : 
                             (N217)? \nz.mem [2173] : 
                             (N219)? \nz.mem [2253] : 
                             (N221)? \nz.mem [2333] : 
                             (N223)? \nz.mem [2413] : 
                             (N225)? \nz.mem [2493] : 
                             (N164)? \nz.mem [2573] : 
                             (N166)? \nz.mem [2653] : 
                             (N168)? \nz.mem [2733] : 
                             (N170)? \nz.mem [2813] : 
                             (N172)? \nz.mem [2893] : 
                             (N174)? \nz.mem [2973] : 
                             (N176)? \nz.mem [3053] : 
                             (N178)? \nz.mem [3133] : 
                             (N180)? \nz.mem [3213] : 
                             (N182)? \nz.mem [3293] : 
                             (N184)? \nz.mem [3373] : 
                             (N186)? \nz.mem [3453] : 
                             (N188)? \nz.mem [3533] : 
                             (N190)? \nz.mem [3613] : 
                             (N192)? \nz.mem [3693] : 
                             (N194)? \nz.mem [3773] : 
                             (N196)? \nz.mem [3853] : 
                             (N198)? \nz.mem [3933] : 
                             (N200)? \nz.mem [4013] : 
                             (N202)? \nz.mem [4093] : 
                             (N204)? \nz.mem [4173] : 
                             (N206)? \nz.mem [4253] : 
                             (N208)? \nz.mem [4333] : 
                             (N210)? \nz.mem [4413] : 
                             (N212)? \nz.mem [4493] : 
                             (N214)? \nz.mem [4573] : 
                             (N216)? \nz.mem [4653] : 
                             (N218)? \nz.mem [4733] : 
                             (N220)? \nz.mem [4813] : 
                             (N222)? \nz.mem [4893] : 
                             (N224)? \nz.mem [4973] : 
                             (N226)? \nz.mem [5053] : 1'b0;
  assign \nz.data_out [12] = (N163)? \nz.mem [12] : 
                             (N165)? \nz.mem [92] : 
                             (N167)? \nz.mem [172] : 
                             (N169)? \nz.mem [252] : 
                             (N171)? \nz.mem [332] : 
                             (N173)? \nz.mem [412] : 
                             (N175)? \nz.mem [492] : 
                             (N177)? \nz.mem [572] : 
                             (N179)? \nz.mem [652] : 
                             (N181)? \nz.mem [732] : 
                             (N183)? \nz.mem [812] : 
                             (N185)? \nz.mem [892] : 
                             (N187)? \nz.mem [972] : 
                             (N189)? \nz.mem [1052] : 
                             (N191)? \nz.mem [1132] : 
                             (N193)? \nz.mem [1212] : 
                             (N195)? \nz.mem [1292] : 
                             (N197)? \nz.mem [1372] : 
                             (N199)? \nz.mem [1452] : 
                             (N201)? \nz.mem [1532] : 
                             (N203)? \nz.mem [1612] : 
                             (N205)? \nz.mem [1692] : 
                             (N207)? \nz.mem [1772] : 
                             (N209)? \nz.mem [1852] : 
                             (N211)? \nz.mem [1932] : 
                             (N213)? \nz.mem [2012] : 
                             (N215)? \nz.mem [2092] : 
                             (N217)? \nz.mem [2172] : 
                             (N219)? \nz.mem [2252] : 
                             (N221)? \nz.mem [2332] : 
                             (N223)? \nz.mem [2412] : 
                             (N225)? \nz.mem [2492] : 
                             (N164)? \nz.mem [2572] : 
                             (N166)? \nz.mem [2652] : 
                             (N168)? \nz.mem [2732] : 
                             (N170)? \nz.mem [2812] : 
                             (N172)? \nz.mem [2892] : 
                             (N174)? \nz.mem [2972] : 
                             (N176)? \nz.mem [3052] : 
                             (N178)? \nz.mem [3132] : 
                             (N180)? \nz.mem [3212] : 
                             (N182)? \nz.mem [3292] : 
                             (N184)? \nz.mem [3372] : 
                             (N186)? \nz.mem [3452] : 
                             (N188)? \nz.mem [3532] : 
                             (N190)? \nz.mem [3612] : 
                             (N192)? \nz.mem [3692] : 
                             (N194)? \nz.mem [3772] : 
                             (N196)? \nz.mem [3852] : 
                             (N198)? \nz.mem [3932] : 
                             (N200)? \nz.mem [4012] : 
                             (N202)? \nz.mem [4092] : 
                             (N204)? \nz.mem [4172] : 
                             (N206)? \nz.mem [4252] : 
                             (N208)? \nz.mem [4332] : 
                             (N210)? \nz.mem [4412] : 
                             (N212)? \nz.mem [4492] : 
                             (N214)? \nz.mem [4572] : 
                             (N216)? \nz.mem [4652] : 
                             (N218)? \nz.mem [4732] : 
                             (N220)? \nz.mem [4812] : 
                             (N222)? \nz.mem [4892] : 
                             (N224)? \nz.mem [4972] : 
                             (N226)? \nz.mem [5052] : 1'b0;
  assign \nz.data_out [11] = (N163)? \nz.mem [11] : 
                             (N165)? \nz.mem [91] : 
                             (N167)? \nz.mem [171] : 
                             (N169)? \nz.mem [251] : 
                             (N171)? \nz.mem [331] : 
                             (N173)? \nz.mem [411] : 
                             (N175)? \nz.mem [491] : 
                             (N177)? \nz.mem [571] : 
                             (N179)? \nz.mem [651] : 
                             (N181)? \nz.mem [731] : 
                             (N183)? \nz.mem [811] : 
                             (N185)? \nz.mem [891] : 
                             (N187)? \nz.mem [971] : 
                             (N189)? \nz.mem [1051] : 
                             (N191)? \nz.mem [1131] : 
                             (N193)? \nz.mem [1211] : 
                             (N195)? \nz.mem [1291] : 
                             (N197)? \nz.mem [1371] : 
                             (N199)? \nz.mem [1451] : 
                             (N201)? \nz.mem [1531] : 
                             (N203)? \nz.mem [1611] : 
                             (N205)? \nz.mem [1691] : 
                             (N207)? \nz.mem [1771] : 
                             (N209)? \nz.mem [1851] : 
                             (N211)? \nz.mem [1931] : 
                             (N213)? \nz.mem [2011] : 
                             (N215)? \nz.mem [2091] : 
                             (N217)? \nz.mem [2171] : 
                             (N219)? \nz.mem [2251] : 
                             (N221)? \nz.mem [2331] : 
                             (N223)? \nz.mem [2411] : 
                             (N225)? \nz.mem [2491] : 
                             (N164)? \nz.mem [2571] : 
                             (N166)? \nz.mem [2651] : 
                             (N168)? \nz.mem [2731] : 
                             (N170)? \nz.mem [2811] : 
                             (N172)? \nz.mem [2891] : 
                             (N174)? \nz.mem [2971] : 
                             (N176)? \nz.mem [3051] : 
                             (N178)? \nz.mem [3131] : 
                             (N180)? \nz.mem [3211] : 
                             (N182)? \nz.mem [3291] : 
                             (N184)? \nz.mem [3371] : 
                             (N186)? \nz.mem [3451] : 
                             (N188)? \nz.mem [3531] : 
                             (N190)? \nz.mem [3611] : 
                             (N192)? \nz.mem [3691] : 
                             (N194)? \nz.mem [3771] : 
                             (N196)? \nz.mem [3851] : 
                             (N198)? \nz.mem [3931] : 
                             (N200)? \nz.mem [4011] : 
                             (N202)? \nz.mem [4091] : 
                             (N204)? \nz.mem [4171] : 
                             (N206)? \nz.mem [4251] : 
                             (N208)? \nz.mem [4331] : 
                             (N210)? \nz.mem [4411] : 
                             (N212)? \nz.mem [4491] : 
                             (N214)? \nz.mem [4571] : 
                             (N216)? \nz.mem [4651] : 
                             (N218)? \nz.mem [4731] : 
                             (N220)? \nz.mem [4811] : 
                             (N222)? \nz.mem [4891] : 
                             (N224)? \nz.mem [4971] : 
                             (N226)? \nz.mem [5051] : 1'b0;
  assign \nz.data_out [10] = (N163)? \nz.mem [10] : 
                             (N165)? \nz.mem [90] : 
                             (N167)? \nz.mem [170] : 
                             (N169)? \nz.mem [250] : 
                             (N171)? \nz.mem [330] : 
                             (N173)? \nz.mem [410] : 
                             (N175)? \nz.mem [490] : 
                             (N177)? \nz.mem [570] : 
                             (N179)? \nz.mem [650] : 
                             (N181)? \nz.mem [730] : 
                             (N183)? \nz.mem [810] : 
                             (N185)? \nz.mem [890] : 
                             (N187)? \nz.mem [970] : 
                             (N189)? \nz.mem [1050] : 
                             (N191)? \nz.mem [1130] : 
                             (N193)? \nz.mem [1210] : 
                             (N195)? \nz.mem [1290] : 
                             (N197)? \nz.mem [1370] : 
                             (N199)? \nz.mem [1450] : 
                             (N201)? \nz.mem [1530] : 
                             (N203)? \nz.mem [1610] : 
                             (N205)? \nz.mem [1690] : 
                             (N207)? \nz.mem [1770] : 
                             (N209)? \nz.mem [1850] : 
                             (N211)? \nz.mem [1930] : 
                             (N213)? \nz.mem [2010] : 
                             (N215)? \nz.mem [2090] : 
                             (N217)? \nz.mem [2170] : 
                             (N219)? \nz.mem [2250] : 
                             (N221)? \nz.mem [2330] : 
                             (N223)? \nz.mem [2410] : 
                             (N225)? \nz.mem [2490] : 
                             (N164)? \nz.mem [2570] : 
                             (N166)? \nz.mem [2650] : 
                             (N168)? \nz.mem [2730] : 
                             (N170)? \nz.mem [2810] : 
                             (N172)? \nz.mem [2890] : 
                             (N174)? \nz.mem [2970] : 
                             (N176)? \nz.mem [3050] : 
                             (N178)? \nz.mem [3130] : 
                             (N180)? \nz.mem [3210] : 
                             (N182)? \nz.mem [3290] : 
                             (N184)? \nz.mem [3370] : 
                             (N186)? \nz.mem [3450] : 
                             (N188)? \nz.mem [3530] : 
                             (N190)? \nz.mem [3610] : 
                             (N192)? \nz.mem [3690] : 
                             (N194)? \nz.mem [3770] : 
                             (N196)? \nz.mem [3850] : 
                             (N198)? \nz.mem [3930] : 
                             (N200)? \nz.mem [4010] : 
                             (N202)? \nz.mem [4090] : 
                             (N204)? \nz.mem [4170] : 
                             (N206)? \nz.mem [4250] : 
                             (N208)? \nz.mem [4330] : 
                             (N210)? \nz.mem [4410] : 
                             (N212)? \nz.mem [4490] : 
                             (N214)? \nz.mem [4570] : 
                             (N216)? \nz.mem [4650] : 
                             (N218)? \nz.mem [4730] : 
                             (N220)? \nz.mem [4810] : 
                             (N222)? \nz.mem [4890] : 
                             (N224)? \nz.mem [4970] : 
                             (N226)? \nz.mem [5050] : 1'b0;
  assign \nz.data_out [9] = (N163)? \nz.mem [9] : 
                            (N165)? \nz.mem [89] : 
                            (N167)? \nz.mem [169] : 
                            (N169)? \nz.mem [249] : 
                            (N171)? \nz.mem [329] : 
                            (N173)? \nz.mem [409] : 
                            (N175)? \nz.mem [489] : 
                            (N177)? \nz.mem [569] : 
                            (N179)? \nz.mem [649] : 
                            (N181)? \nz.mem [729] : 
                            (N183)? \nz.mem [809] : 
                            (N185)? \nz.mem [889] : 
                            (N187)? \nz.mem [969] : 
                            (N189)? \nz.mem [1049] : 
                            (N191)? \nz.mem [1129] : 
                            (N193)? \nz.mem [1209] : 
                            (N195)? \nz.mem [1289] : 
                            (N197)? \nz.mem [1369] : 
                            (N199)? \nz.mem [1449] : 
                            (N201)? \nz.mem [1529] : 
                            (N203)? \nz.mem [1609] : 
                            (N205)? \nz.mem [1689] : 
                            (N207)? \nz.mem [1769] : 
                            (N209)? \nz.mem [1849] : 
                            (N211)? \nz.mem [1929] : 
                            (N213)? \nz.mem [2009] : 
                            (N215)? \nz.mem [2089] : 
                            (N217)? \nz.mem [2169] : 
                            (N219)? \nz.mem [2249] : 
                            (N221)? \nz.mem [2329] : 
                            (N223)? \nz.mem [2409] : 
                            (N225)? \nz.mem [2489] : 
                            (N164)? \nz.mem [2569] : 
                            (N166)? \nz.mem [2649] : 
                            (N168)? \nz.mem [2729] : 
                            (N170)? \nz.mem [2809] : 
                            (N172)? \nz.mem [2889] : 
                            (N174)? \nz.mem [2969] : 
                            (N176)? \nz.mem [3049] : 
                            (N178)? \nz.mem [3129] : 
                            (N180)? \nz.mem [3209] : 
                            (N182)? \nz.mem [3289] : 
                            (N184)? \nz.mem [3369] : 
                            (N186)? \nz.mem [3449] : 
                            (N188)? \nz.mem [3529] : 
                            (N190)? \nz.mem [3609] : 
                            (N192)? \nz.mem [3689] : 
                            (N194)? \nz.mem [3769] : 
                            (N196)? \nz.mem [3849] : 
                            (N198)? \nz.mem [3929] : 
                            (N200)? \nz.mem [4009] : 
                            (N202)? \nz.mem [4089] : 
                            (N204)? \nz.mem [4169] : 
                            (N206)? \nz.mem [4249] : 
                            (N208)? \nz.mem [4329] : 
                            (N210)? \nz.mem [4409] : 
                            (N212)? \nz.mem [4489] : 
                            (N214)? \nz.mem [4569] : 
                            (N216)? \nz.mem [4649] : 
                            (N218)? \nz.mem [4729] : 
                            (N220)? \nz.mem [4809] : 
                            (N222)? \nz.mem [4889] : 
                            (N224)? \nz.mem [4969] : 
                            (N226)? \nz.mem [5049] : 1'b0;
  assign \nz.data_out [8] = (N163)? \nz.mem [8] : 
                            (N165)? \nz.mem [88] : 
                            (N167)? \nz.mem [168] : 
                            (N169)? \nz.mem [248] : 
                            (N171)? \nz.mem [328] : 
                            (N173)? \nz.mem [408] : 
                            (N175)? \nz.mem [488] : 
                            (N177)? \nz.mem [568] : 
                            (N179)? \nz.mem [648] : 
                            (N181)? \nz.mem [728] : 
                            (N183)? \nz.mem [808] : 
                            (N185)? \nz.mem [888] : 
                            (N187)? \nz.mem [968] : 
                            (N189)? \nz.mem [1048] : 
                            (N191)? \nz.mem [1128] : 
                            (N193)? \nz.mem [1208] : 
                            (N195)? \nz.mem [1288] : 
                            (N197)? \nz.mem [1368] : 
                            (N199)? \nz.mem [1448] : 
                            (N201)? \nz.mem [1528] : 
                            (N203)? \nz.mem [1608] : 
                            (N205)? \nz.mem [1688] : 
                            (N207)? \nz.mem [1768] : 
                            (N209)? \nz.mem [1848] : 
                            (N211)? \nz.mem [1928] : 
                            (N213)? \nz.mem [2008] : 
                            (N215)? \nz.mem [2088] : 
                            (N217)? \nz.mem [2168] : 
                            (N219)? \nz.mem [2248] : 
                            (N221)? \nz.mem [2328] : 
                            (N223)? \nz.mem [2408] : 
                            (N225)? \nz.mem [2488] : 
                            (N164)? \nz.mem [2568] : 
                            (N166)? \nz.mem [2648] : 
                            (N168)? \nz.mem [2728] : 
                            (N170)? \nz.mem [2808] : 
                            (N172)? \nz.mem [2888] : 
                            (N174)? \nz.mem [2968] : 
                            (N176)? \nz.mem [3048] : 
                            (N178)? \nz.mem [3128] : 
                            (N180)? \nz.mem [3208] : 
                            (N182)? \nz.mem [3288] : 
                            (N184)? \nz.mem [3368] : 
                            (N186)? \nz.mem [3448] : 
                            (N188)? \nz.mem [3528] : 
                            (N190)? \nz.mem [3608] : 
                            (N192)? \nz.mem [3688] : 
                            (N194)? \nz.mem [3768] : 
                            (N196)? \nz.mem [3848] : 
                            (N198)? \nz.mem [3928] : 
                            (N200)? \nz.mem [4008] : 
                            (N202)? \nz.mem [4088] : 
                            (N204)? \nz.mem [4168] : 
                            (N206)? \nz.mem [4248] : 
                            (N208)? \nz.mem [4328] : 
                            (N210)? \nz.mem [4408] : 
                            (N212)? \nz.mem [4488] : 
                            (N214)? \nz.mem [4568] : 
                            (N216)? \nz.mem [4648] : 
                            (N218)? \nz.mem [4728] : 
                            (N220)? \nz.mem [4808] : 
                            (N222)? \nz.mem [4888] : 
                            (N224)? \nz.mem [4968] : 
                            (N226)? \nz.mem [5048] : 1'b0;
  assign \nz.data_out [7] = (N163)? \nz.mem [7] : 
                            (N165)? \nz.mem [87] : 
                            (N167)? \nz.mem [167] : 
                            (N169)? \nz.mem [247] : 
                            (N171)? \nz.mem [327] : 
                            (N173)? \nz.mem [407] : 
                            (N175)? \nz.mem [487] : 
                            (N177)? \nz.mem [567] : 
                            (N179)? \nz.mem [647] : 
                            (N181)? \nz.mem [727] : 
                            (N183)? \nz.mem [807] : 
                            (N185)? \nz.mem [887] : 
                            (N187)? \nz.mem [967] : 
                            (N189)? \nz.mem [1047] : 
                            (N191)? \nz.mem [1127] : 
                            (N193)? \nz.mem [1207] : 
                            (N195)? \nz.mem [1287] : 
                            (N197)? \nz.mem [1367] : 
                            (N199)? \nz.mem [1447] : 
                            (N201)? \nz.mem [1527] : 
                            (N203)? \nz.mem [1607] : 
                            (N205)? \nz.mem [1687] : 
                            (N207)? \nz.mem [1767] : 
                            (N209)? \nz.mem [1847] : 
                            (N211)? \nz.mem [1927] : 
                            (N213)? \nz.mem [2007] : 
                            (N215)? \nz.mem [2087] : 
                            (N217)? \nz.mem [2167] : 
                            (N219)? \nz.mem [2247] : 
                            (N221)? \nz.mem [2327] : 
                            (N223)? \nz.mem [2407] : 
                            (N225)? \nz.mem [2487] : 
                            (N164)? \nz.mem [2567] : 
                            (N166)? \nz.mem [2647] : 
                            (N168)? \nz.mem [2727] : 
                            (N170)? \nz.mem [2807] : 
                            (N172)? \nz.mem [2887] : 
                            (N174)? \nz.mem [2967] : 
                            (N176)? \nz.mem [3047] : 
                            (N178)? \nz.mem [3127] : 
                            (N180)? \nz.mem [3207] : 
                            (N182)? \nz.mem [3287] : 
                            (N184)? \nz.mem [3367] : 
                            (N186)? \nz.mem [3447] : 
                            (N188)? \nz.mem [3527] : 
                            (N190)? \nz.mem [3607] : 
                            (N192)? \nz.mem [3687] : 
                            (N194)? \nz.mem [3767] : 
                            (N196)? \nz.mem [3847] : 
                            (N198)? \nz.mem [3927] : 
                            (N200)? \nz.mem [4007] : 
                            (N202)? \nz.mem [4087] : 
                            (N204)? \nz.mem [4167] : 
                            (N206)? \nz.mem [4247] : 
                            (N208)? \nz.mem [4327] : 
                            (N210)? \nz.mem [4407] : 
                            (N212)? \nz.mem [4487] : 
                            (N214)? \nz.mem [4567] : 
                            (N216)? \nz.mem [4647] : 
                            (N218)? \nz.mem [4727] : 
                            (N220)? \nz.mem [4807] : 
                            (N222)? \nz.mem [4887] : 
                            (N224)? \nz.mem [4967] : 
                            (N226)? \nz.mem [5047] : 1'b0;
  assign \nz.data_out [6] = (N163)? \nz.mem [6] : 
                            (N165)? \nz.mem [86] : 
                            (N167)? \nz.mem [166] : 
                            (N169)? \nz.mem [246] : 
                            (N171)? \nz.mem [326] : 
                            (N173)? \nz.mem [406] : 
                            (N175)? \nz.mem [486] : 
                            (N177)? \nz.mem [566] : 
                            (N179)? \nz.mem [646] : 
                            (N181)? \nz.mem [726] : 
                            (N183)? \nz.mem [806] : 
                            (N185)? \nz.mem [886] : 
                            (N187)? \nz.mem [966] : 
                            (N189)? \nz.mem [1046] : 
                            (N191)? \nz.mem [1126] : 
                            (N193)? \nz.mem [1206] : 
                            (N195)? \nz.mem [1286] : 
                            (N197)? \nz.mem [1366] : 
                            (N199)? \nz.mem [1446] : 
                            (N201)? \nz.mem [1526] : 
                            (N203)? \nz.mem [1606] : 
                            (N205)? \nz.mem [1686] : 
                            (N207)? \nz.mem [1766] : 
                            (N209)? \nz.mem [1846] : 
                            (N211)? \nz.mem [1926] : 
                            (N213)? \nz.mem [2006] : 
                            (N215)? \nz.mem [2086] : 
                            (N217)? \nz.mem [2166] : 
                            (N219)? \nz.mem [2246] : 
                            (N221)? \nz.mem [2326] : 
                            (N223)? \nz.mem [2406] : 
                            (N225)? \nz.mem [2486] : 
                            (N164)? \nz.mem [2566] : 
                            (N166)? \nz.mem [2646] : 
                            (N168)? \nz.mem [2726] : 
                            (N170)? \nz.mem [2806] : 
                            (N172)? \nz.mem [2886] : 
                            (N174)? \nz.mem [2966] : 
                            (N176)? \nz.mem [3046] : 
                            (N178)? \nz.mem [3126] : 
                            (N180)? \nz.mem [3206] : 
                            (N182)? \nz.mem [3286] : 
                            (N184)? \nz.mem [3366] : 
                            (N186)? \nz.mem [3446] : 
                            (N188)? \nz.mem [3526] : 
                            (N190)? \nz.mem [3606] : 
                            (N192)? \nz.mem [3686] : 
                            (N194)? \nz.mem [3766] : 
                            (N196)? \nz.mem [3846] : 
                            (N198)? \nz.mem [3926] : 
                            (N200)? \nz.mem [4006] : 
                            (N202)? \nz.mem [4086] : 
                            (N204)? \nz.mem [4166] : 
                            (N206)? \nz.mem [4246] : 
                            (N208)? \nz.mem [4326] : 
                            (N210)? \nz.mem [4406] : 
                            (N212)? \nz.mem [4486] : 
                            (N214)? \nz.mem [4566] : 
                            (N216)? \nz.mem [4646] : 
                            (N218)? \nz.mem [4726] : 
                            (N220)? \nz.mem [4806] : 
                            (N222)? \nz.mem [4886] : 
                            (N224)? \nz.mem [4966] : 
                            (N226)? \nz.mem [5046] : 1'b0;
  assign \nz.data_out [5] = (N163)? \nz.mem [5] : 
                            (N165)? \nz.mem [85] : 
                            (N167)? \nz.mem [165] : 
                            (N169)? \nz.mem [245] : 
                            (N171)? \nz.mem [325] : 
                            (N173)? \nz.mem [405] : 
                            (N175)? \nz.mem [485] : 
                            (N177)? \nz.mem [565] : 
                            (N179)? \nz.mem [645] : 
                            (N181)? \nz.mem [725] : 
                            (N183)? \nz.mem [805] : 
                            (N185)? \nz.mem [885] : 
                            (N187)? \nz.mem [965] : 
                            (N189)? \nz.mem [1045] : 
                            (N191)? \nz.mem [1125] : 
                            (N193)? \nz.mem [1205] : 
                            (N195)? \nz.mem [1285] : 
                            (N197)? \nz.mem [1365] : 
                            (N199)? \nz.mem [1445] : 
                            (N201)? \nz.mem [1525] : 
                            (N203)? \nz.mem [1605] : 
                            (N205)? \nz.mem [1685] : 
                            (N207)? \nz.mem [1765] : 
                            (N209)? \nz.mem [1845] : 
                            (N211)? \nz.mem [1925] : 
                            (N213)? \nz.mem [2005] : 
                            (N215)? \nz.mem [2085] : 
                            (N217)? \nz.mem [2165] : 
                            (N219)? \nz.mem [2245] : 
                            (N221)? \nz.mem [2325] : 
                            (N223)? \nz.mem [2405] : 
                            (N225)? \nz.mem [2485] : 
                            (N164)? \nz.mem [2565] : 
                            (N166)? \nz.mem [2645] : 
                            (N168)? \nz.mem [2725] : 
                            (N170)? \nz.mem [2805] : 
                            (N172)? \nz.mem [2885] : 
                            (N174)? \nz.mem [2965] : 
                            (N176)? \nz.mem [3045] : 
                            (N178)? \nz.mem [3125] : 
                            (N180)? \nz.mem [3205] : 
                            (N182)? \nz.mem [3285] : 
                            (N184)? \nz.mem [3365] : 
                            (N186)? \nz.mem [3445] : 
                            (N188)? \nz.mem [3525] : 
                            (N190)? \nz.mem [3605] : 
                            (N192)? \nz.mem [3685] : 
                            (N194)? \nz.mem [3765] : 
                            (N196)? \nz.mem [3845] : 
                            (N198)? \nz.mem [3925] : 
                            (N200)? \nz.mem [4005] : 
                            (N202)? \nz.mem [4085] : 
                            (N204)? \nz.mem [4165] : 
                            (N206)? \nz.mem [4245] : 
                            (N208)? \nz.mem [4325] : 
                            (N210)? \nz.mem [4405] : 
                            (N212)? \nz.mem [4485] : 
                            (N214)? \nz.mem [4565] : 
                            (N216)? \nz.mem [4645] : 
                            (N218)? \nz.mem [4725] : 
                            (N220)? \nz.mem [4805] : 
                            (N222)? \nz.mem [4885] : 
                            (N224)? \nz.mem [4965] : 
                            (N226)? \nz.mem [5045] : 1'b0;
  assign \nz.data_out [4] = (N163)? \nz.mem [4] : 
                            (N165)? \nz.mem [84] : 
                            (N167)? \nz.mem [164] : 
                            (N169)? \nz.mem [244] : 
                            (N171)? \nz.mem [324] : 
                            (N173)? \nz.mem [404] : 
                            (N175)? \nz.mem [484] : 
                            (N177)? \nz.mem [564] : 
                            (N179)? \nz.mem [644] : 
                            (N181)? \nz.mem [724] : 
                            (N183)? \nz.mem [804] : 
                            (N185)? \nz.mem [884] : 
                            (N187)? \nz.mem [964] : 
                            (N189)? \nz.mem [1044] : 
                            (N191)? \nz.mem [1124] : 
                            (N193)? \nz.mem [1204] : 
                            (N195)? \nz.mem [1284] : 
                            (N197)? \nz.mem [1364] : 
                            (N199)? \nz.mem [1444] : 
                            (N201)? \nz.mem [1524] : 
                            (N203)? \nz.mem [1604] : 
                            (N205)? \nz.mem [1684] : 
                            (N207)? \nz.mem [1764] : 
                            (N209)? \nz.mem [1844] : 
                            (N211)? \nz.mem [1924] : 
                            (N213)? \nz.mem [2004] : 
                            (N215)? \nz.mem [2084] : 
                            (N217)? \nz.mem [2164] : 
                            (N219)? \nz.mem [2244] : 
                            (N221)? \nz.mem [2324] : 
                            (N223)? \nz.mem [2404] : 
                            (N225)? \nz.mem [2484] : 
                            (N164)? \nz.mem [2564] : 
                            (N166)? \nz.mem [2644] : 
                            (N168)? \nz.mem [2724] : 
                            (N170)? \nz.mem [2804] : 
                            (N172)? \nz.mem [2884] : 
                            (N174)? \nz.mem [2964] : 
                            (N176)? \nz.mem [3044] : 
                            (N178)? \nz.mem [3124] : 
                            (N180)? \nz.mem [3204] : 
                            (N182)? \nz.mem [3284] : 
                            (N184)? \nz.mem [3364] : 
                            (N186)? \nz.mem [3444] : 
                            (N188)? \nz.mem [3524] : 
                            (N190)? \nz.mem [3604] : 
                            (N192)? \nz.mem [3684] : 
                            (N194)? \nz.mem [3764] : 
                            (N196)? \nz.mem [3844] : 
                            (N198)? \nz.mem [3924] : 
                            (N200)? \nz.mem [4004] : 
                            (N202)? \nz.mem [4084] : 
                            (N204)? \nz.mem [4164] : 
                            (N206)? \nz.mem [4244] : 
                            (N208)? \nz.mem [4324] : 
                            (N210)? \nz.mem [4404] : 
                            (N212)? \nz.mem [4484] : 
                            (N214)? \nz.mem [4564] : 
                            (N216)? \nz.mem [4644] : 
                            (N218)? \nz.mem [4724] : 
                            (N220)? \nz.mem [4804] : 
                            (N222)? \nz.mem [4884] : 
                            (N224)? \nz.mem [4964] : 
                            (N226)? \nz.mem [5044] : 1'b0;
  assign \nz.data_out [3] = (N163)? \nz.mem [3] : 
                            (N165)? \nz.mem [83] : 
                            (N167)? \nz.mem [163] : 
                            (N169)? \nz.mem [243] : 
                            (N171)? \nz.mem [323] : 
                            (N173)? \nz.mem [403] : 
                            (N175)? \nz.mem [483] : 
                            (N177)? \nz.mem [563] : 
                            (N179)? \nz.mem [643] : 
                            (N181)? \nz.mem [723] : 
                            (N183)? \nz.mem [803] : 
                            (N185)? \nz.mem [883] : 
                            (N187)? \nz.mem [963] : 
                            (N189)? \nz.mem [1043] : 
                            (N191)? \nz.mem [1123] : 
                            (N193)? \nz.mem [1203] : 
                            (N195)? \nz.mem [1283] : 
                            (N197)? \nz.mem [1363] : 
                            (N199)? \nz.mem [1443] : 
                            (N201)? \nz.mem [1523] : 
                            (N203)? \nz.mem [1603] : 
                            (N205)? \nz.mem [1683] : 
                            (N207)? \nz.mem [1763] : 
                            (N209)? \nz.mem [1843] : 
                            (N211)? \nz.mem [1923] : 
                            (N213)? \nz.mem [2003] : 
                            (N215)? \nz.mem [2083] : 
                            (N217)? \nz.mem [2163] : 
                            (N219)? \nz.mem [2243] : 
                            (N221)? \nz.mem [2323] : 
                            (N223)? \nz.mem [2403] : 
                            (N225)? \nz.mem [2483] : 
                            (N164)? \nz.mem [2563] : 
                            (N166)? \nz.mem [2643] : 
                            (N168)? \nz.mem [2723] : 
                            (N170)? \nz.mem [2803] : 
                            (N172)? \nz.mem [2883] : 
                            (N174)? \nz.mem [2963] : 
                            (N176)? \nz.mem [3043] : 
                            (N178)? \nz.mem [3123] : 
                            (N180)? \nz.mem [3203] : 
                            (N182)? \nz.mem [3283] : 
                            (N184)? \nz.mem [3363] : 
                            (N186)? \nz.mem [3443] : 
                            (N188)? \nz.mem [3523] : 
                            (N190)? \nz.mem [3603] : 
                            (N192)? \nz.mem [3683] : 
                            (N194)? \nz.mem [3763] : 
                            (N196)? \nz.mem [3843] : 
                            (N198)? \nz.mem [3923] : 
                            (N200)? \nz.mem [4003] : 
                            (N202)? \nz.mem [4083] : 
                            (N204)? \nz.mem [4163] : 
                            (N206)? \nz.mem [4243] : 
                            (N208)? \nz.mem [4323] : 
                            (N210)? \nz.mem [4403] : 
                            (N212)? \nz.mem [4483] : 
                            (N214)? \nz.mem [4563] : 
                            (N216)? \nz.mem [4643] : 
                            (N218)? \nz.mem [4723] : 
                            (N220)? \nz.mem [4803] : 
                            (N222)? \nz.mem [4883] : 
                            (N224)? \nz.mem [4963] : 
                            (N226)? \nz.mem [5043] : 1'b0;
  assign \nz.data_out [2] = (N163)? \nz.mem [2] : 
                            (N165)? \nz.mem [82] : 
                            (N167)? \nz.mem [162] : 
                            (N169)? \nz.mem [242] : 
                            (N171)? \nz.mem [322] : 
                            (N173)? \nz.mem [402] : 
                            (N175)? \nz.mem [482] : 
                            (N177)? \nz.mem [562] : 
                            (N179)? \nz.mem [642] : 
                            (N181)? \nz.mem [722] : 
                            (N183)? \nz.mem [802] : 
                            (N185)? \nz.mem [882] : 
                            (N187)? \nz.mem [962] : 
                            (N189)? \nz.mem [1042] : 
                            (N191)? \nz.mem [1122] : 
                            (N193)? \nz.mem [1202] : 
                            (N195)? \nz.mem [1282] : 
                            (N197)? \nz.mem [1362] : 
                            (N199)? \nz.mem [1442] : 
                            (N201)? \nz.mem [1522] : 
                            (N203)? \nz.mem [1602] : 
                            (N205)? \nz.mem [1682] : 
                            (N207)? \nz.mem [1762] : 
                            (N209)? \nz.mem [1842] : 
                            (N211)? \nz.mem [1922] : 
                            (N213)? \nz.mem [2002] : 
                            (N215)? \nz.mem [2082] : 
                            (N217)? \nz.mem [2162] : 
                            (N219)? \nz.mem [2242] : 
                            (N221)? \nz.mem [2322] : 
                            (N223)? \nz.mem [2402] : 
                            (N225)? \nz.mem [2482] : 
                            (N164)? \nz.mem [2562] : 
                            (N166)? \nz.mem [2642] : 
                            (N168)? \nz.mem [2722] : 
                            (N170)? \nz.mem [2802] : 
                            (N172)? \nz.mem [2882] : 
                            (N174)? \nz.mem [2962] : 
                            (N176)? \nz.mem [3042] : 
                            (N178)? \nz.mem [3122] : 
                            (N180)? \nz.mem [3202] : 
                            (N182)? \nz.mem [3282] : 
                            (N184)? \nz.mem [3362] : 
                            (N186)? \nz.mem [3442] : 
                            (N188)? \nz.mem [3522] : 
                            (N190)? \nz.mem [3602] : 
                            (N192)? \nz.mem [3682] : 
                            (N194)? \nz.mem [3762] : 
                            (N196)? \nz.mem [3842] : 
                            (N198)? \nz.mem [3922] : 
                            (N200)? \nz.mem [4002] : 
                            (N202)? \nz.mem [4082] : 
                            (N204)? \nz.mem [4162] : 
                            (N206)? \nz.mem [4242] : 
                            (N208)? \nz.mem [4322] : 
                            (N210)? \nz.mem [4402] : 
                            (N212)? \nz.mem [4482] : 
                            (N214)? \nz.mem [4562] : 
                            (N216)? \nz.mem [4642] : 
                            (N218)? \nz.mem [4722] : 
                            (N220)? \nz.mem [4802] : 
                            (N222)? \nz.mem [4882] : 
                            (N224)? \nz.mem [4962] : 
                            (N226)? \nz.mem [5042] : 1'b0;
  assign \nz.data_out [1] = (N163)? \nz.mem [1] : 
                            (N165)? \nz.mem [81] : 
                            (N167)? \nz.mem [161] : 
                            (N169)? \nz.mem [241] : 
                            (N171)? \nz.mem [321] : 
                            (N173)? \nz.mem [401] : 
                            (N175)? \nz.mem [481] : 
                            (N177)? \nz.mem [561] : 
                            (N179)? \nz.mem [641] : 
                            (N181)? \nz.mem [721] : 
                            (N183)? \nz.mem [801] : 
                            (N185)? \nz.mem [881] : 
                            (N187)? \nz.mem [961] : 
                            (N189)? \nz.mem [1041] : 
                            (N191)? \nz.mem [1121] : 
                            (N193)? \nz.mem [1201] : 
                            (N195)? \nz.mem [1281] : 
                            (N197)? \nz.mem [1361] : 
                            (N199)? \nz.mem [1441] : 
                            (N201)? \nz.mem [1521] : 
                            (N203)? \nz.mem [1601] : 
                            (N205)? \nz.mem [1681] : 
                            (N207)? \nz.mem [1761] : 
                            (N209)? \nz.mem [1841] : 
                            (N211)? \nz.mem [1921] : 
                            (N213)? \nz.mem [2001] : 
                            (N215)? \nz.mem [2081] : 
                            (N217)? \nz.mem [2161] : 
                            (N219)? \nz.mem [2241] : 
                            (N221)? \nz.mem [2321] : 
                            (N223)? \nz.mem [2401] : 
                            (N225)? \nz.mem [2481] : 
                            (N164)? \nz.mem [2561] : 
                            (N166)? \nz.mem [2641] : 
                            (N168)? \nz.mem [2721] : 
                            (N170)? \nz.mem [2801] : 
                            (N172)? \nz.mem [2881] : 
                            (N174)? \nz.mem [2961] : 
                            (N176)? \nz.mem [3041] : 
                            (N178)? \nz.mem [3121] : 
                            (N180)? \nz.mem [3201] : 
                            (N182)? \nz.mem [3281] : 
                            (N184)? \nz.mem [3361] : 
                            (N186)? \nz.mem [3441] : 
                            (N188)? \nz.mem [3521] : 
                            (N190)? \nz.mem [3601] : 
                            (N192)? \nz.mem [3681] : 
                            (N194)? \nz.mem [3761] : 
                            (N196)? \nz.mem [3841] : 
                            (N198)? \nz.mem [3921] : 
                            (N200)? \nz.mem [4001] : 
                            (N202)? \nz.mem [4081] : 
                            (N204)? \nz.mem [4161] : 
                            (N206)? \nz.mem [4241] : 
                            (N208)? \nz.mem [4321] : 
                            (N210)? \nz.mem [4401] : 
                            (N212)? \nz.mem [4481] : 
                            (N214)? \nz.mem [4561] : 
                            (N216)? \nz.mem [4641] : 
                            (N218)? \nz.mem [4721] : 
                            (N220)? \nz.mem [4801] : 
                            (N222)? \nz.mem [4881] : 
                            (N224)? \nz.mem [4961] : 
                            (N226)? \nz.mem [5041] : 1'b0;
  assign \nz.data_out [0] = (N163)? \nz.mem [0] : 
                            (N165)? \nz.mem [80] : 
                            (N167)? \nz.mem [160] : 
                            (N169)? \nz.mem [240] : 
                            (N171)? \nz.mem [320] : 
                            (N173)? \nz.mem [400] : 
                            (N175)? \nz.mem [480] : 
                            (N177)? \nz.mem [560] : 
                            (N179)? \nz.mem [640] : 
                            (N181)? \nz.mem [720] : 
                            (N183)? \nz.mem [800] : 
                            (N185)? \nz.mem [880] : 
                            (N187)? \nz.mem [960] : 
                            (N189)? \nz.mem [1040] : 
                            (N191)? \nz.mem [1120] : 
                            (N193)? \nz.mem [1200] : 
                            (N195)? \nz.mem [1280] : 
                            (N197)? \nz.mem [1360] : 
                            (N199)? \nz.mem [1440] : 
                            (N201)? \nz.mem [1520] : 
                            (N203)? \nz.mem [1600] : 
                            (N205)? \nz.mem [1680] : 
                            (N207)? \nz.mem [1760] : 
                            (N209)? \nz.mem [1840] : 
                            (N211)? \nz.mem [1920] : 
                            (N213)? \nz.mem [2000] : 
                            (N215)? \nz.mem [2080] : 
                            (N217)? \nz.mem [2160] : 
                            (N219)? \nz.mem [2240] : 
                            (N221)? \nz.mem [2320] : 
                            (N223)? \nz.mem [2400] : 
                            (N225)? \nz.mem [2480] : 
                            (N164)? \nz.mem [2560] : 
                            (N166)? \nz.mem [2640] : 
                            (N168)? \nz.mem [2720] : 
                            (N170)? \nz.mem [2800] : 
                            (N172)? \nz.mem [2880] : 
                            (N174)? \nz.mem [2960] : 
                            (N176)? \nz.mem [3040] : 
                            (N178)? \nz.mem [3120] : 
                            (N180)? \nz.mem [3200] : 
                            (N182)? \nz.mem [3280] : 
                            (N184)? \nz.mem [3360] : 
                            (N186)? \nz.mem [3440] : 
                            (N188)? \nz.mem [3520] : 
                            (N190)? \nz.mem [3600] : 
                            (N192)? \nz.mem [3680] : 
                            (N194)? \nz.mem [3760] : 
                            (N196)? \nz.mem [3840] : 
                            (N198)? \nz.mem [3920] : 
                            (N200)? \nz.mem [4000] : 
                            (N202)? \nz.mem [4080] : 
                            (N204)? \nz.mem [4160] : 
                            (N206)? \nz.mem [4240] : 
                            (N208)? \nz.mem [4320] : 
                            (N210)? \nz.mem [4400] : 
                            (N212)? \nz.mem [4480] : 
                            (N214)? \nz.mem [4560] : 
                            (N216)? \nz.mem [4640] : 
                            (N218)? \nz.mem [4720] : 
                            (N220)? \nz.mem [4800] : 
                            (N222)? \nz.mem [4880] : 
                            (N224)? \nz.mem [4960] : 
                            (N226)? \nz.mem [5040] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p80
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N11497 = ~addr_i[5];
  assign N11498 = N11497 & N11539;
  assign N11499 = N11497 & N11540;
  assign N11500 = N11497 & N11541;
  assign N11501 = N11497 & N11542;
  assign N11502 = ~addr_i[2];
  assign N11503 = N11502 & N11551;
  assign N11504 = N11502 & N11552;
  assign N11505 = N11502 & N11553;
  assign N11506 = N11502 & N11554;
  assign N537 = N11507 & N11503;
  assign N536 = N11507 & N11504;
  assign N535 = N11507 & N11505;
  assign N534 = N11507 & N11506;
  assign N533 = N11508 & N11503;
  assign N532 = N11508 & N11504;
  assign N531 = N11508 & N11505;
  assign N530 = N11508 & N11506;
  assign N529 = N11509 & N11503;
  assign N528 = N11509 & N11504;
  assign N527 = N11509 & N11505;
  assign N526 = N11509 & N11506;
  assign N525 = N11546 & N11503;
  assign N524 = N11546 & N11504;
  assign N523 = N11546 & N11505;
  assign N522 = N11546 & N11506;
  assign N521 = N11498 & N11510;
  assign N520 = N11498 & N11511;
  assign N519 = N11498 & N11512;
  assign N518 = N11498 & N11558;
  assign N517 = N11498 & N11503;
  assign N516 = N11498 & N11504;
  assign N515 = N11498 & N11505;
  assign N514 = N11498 & N11506;
  assign N513 = N11499 & N11510;
  assign N512 = N11499 & N11511;
  assign N511 = N11499 & N11512;
  assign N510 = N11499 & N11558;
  assign N509 = N11499 & N11503;
  assign N508 = N11499 & N11504;
  assign N507 = N11499 & N11505;
  assign N506 = N11499 & N11506;
  assign N505 = N11500 & N11510;
  assign N504 = N11500 & N11511;
  assign N503 = N11500 & N11512;
  assign N502 = N11500 & N11558;
  assign N501 = N11500 & N11503;
  assign N500 = N11500 & N11504;
  assign N499 = N11500 & N11505;
  assign N498 = N11500 & N11506;
  assign N497 = N11501 & N11510;
  assign N496 = N11501 & N11511;
  assign N495 = N11501 & N11512;
  assign N494 = N11501 & N11558;
  assign N493 = N11501 & N11503;
  assign N492 = N11501 & N11504;
  assign N491 = N11501 & N11505;
  assign N490 = N11501 & N11506;
  assign N11507 = addr_i[5] & N11539;
  assign N11508 = addr_i[5] & N11540;
  assign N11509 = addr_i[5] & N11541;
  assign N11510 = addr_i[2] & N11551;
  assign N11511 = addr_i[2] & N11552;
  assign N11512 = addr_i[2] & N11553;
  assign N641 = N11507 & N11510;
  assign N640 = N11507 & N11511;
  assign N639 = N11507 & N11512;
  assign N638 = N11507 & N11558;
  assign N637 = N11507 & N11559;
  assign N636 = N11507 & N11560;
  assign N635 = N11507 & N11561;
  assign N634 = N11507 & N11562;
  assign N633 = N11508 & N11510;
  assign N632 = N11508 & N11511;
  assign N631 = N11508 & N11512;
  assign N630 = N11508 & N11558;
  assign N629 = N11508 & N11559;
  assign N628 = N11508 & N11560;
  assign N627 = N11508 & N11561;
  assign N626 = N11508 & N11562;
  assign N625 = N11509 & N11510;
  assign N624 = N11509 & N11511;
  assign N623 = N11509 & N11512;
  assign N622 = N11509 & N11558;
  assign N621 = N11509 & N11559;
  assign N620 = N11509 & N11560;
  assign N619 = N11509 & N11561;
  assign N618 = N11509 & N11562;
  assign N617 = N11546 & N11510;
  assign N616 = N11546 & N11511;
  assign N615 = N11546 & N11512;
  assign N614 = N11547 & N11510;
  assign N613 = N11547 & N11511;
  assign N612 = N11547 & N11512;
  assign N611 = N11548 & N11510;
  assign N610 = N11548 & N11511;
  assign N609 = N11548 & N11512;
  assign N608 = N11549 & N11510;
  assign N607 = N11549 & N11511;
  assign N606 = N11549 & N11512;
  assign N605 = N11550 & N11510;
  assign N604 = N11550 & N11511;
  assign N603 = N11550 & N11512;
  assign N972 = N11513 & N11558;
  assign N971 = N11514 & N11558;
  assign N970 = N11515 & N11558;
  assign N969 = N11546 & N11516;
  assign N968 = N11546 & N11517;
  assign N967 = N11546 & N11518;
  assign N1329 = N11513 & N11559;
  assign N1328 = N11513 & N11560;
  assign N1327 = N11513 & N11561;
  assign N1326 = N11513 & N11562;
  assign N1325 = N11514 & N11559;
  assign N1324 = N11514 & N11560;
  assign N1323 = N11514 & N11561;
  assign N1322 = N11514 & N11562;
  assign N1321 = N11515 & N11559;
  assign N1320 = N11515 & N11560;
  assign N1319 = N11515 & N11561;
  assign N1318 = N11515 & N11562;
  assign N1317 = N11529 & N11559;
  assign N1316 = N11529 & N11560;
  assign N1315 = N11529 & N11561;
  assign N1314 = N11529 & N11562;
  assign N1313 = N11547 & N11516;
  assign N1312 = N11547 & N11517;
  assign N1311 = N11547 & N11518;
  assign N1310 = N11547 & N11534;
  assign N1309 = N11548 & N11516;
  assign N1308 = N11548 & N11517;
  assign N1307 = N11548 & N11518;
  assign N1306 = N11548 & N11534;
  assign N1305 = N11549 & N11516;
  assign N1304 = N11549 & N11517;
  assign N1303 = N11549 & N11518;
  assign N1302 = N11549 & N11534;
  assign N1301 = N11550 & N11516;
  assign N1300 = N11550 & N11517;
  assign N1299 = N11550 & N11518;
  assign N1298 = N11550 & N11534;
  assign N11513 = addr_i[5] & N11539;
  assign N11514 = addr_i[5] & N11540;
  assign N11515 = addr_i[5] & N11541;
  assign N11516 = addr_i[2] & N11551;
  assign N11517 = addr_i[2] & N11552;
  assign N11518 = addr_i[2] & N11553;
  assign N1498 = N11513 & N11516;
  assign N1497 = N11513 & N11517;
  assign N1496 = N11513 & N11518;
  assign N1495 = N11513 & N11534;
  assign N1494 = N11513 & N11535;
  assign N1493 = N11513 & N11536;
  assign N1492 = N11513 & N11537;
  assign N1491 = N11513 & N11538;
  assign N1490 = N11514 & N11516;
  assign N1489 = N11514 & N11517;
  assign N1488 = N11514 & N11518;
  assign N1487 = N11514 & N11534;
  assign N1486 = N11514 & N11535;
  assign N1485 = N11514 & N11536;
  assign N1484 = N11514 & N11537;
  assign N1483 = N11514 & N11538;
  assign N1482 = N11515 & N11516;
  assign N1481 = N11515 & N11517;
  assign N1480 = N11515 & N11518;
  assign N1479 = N11515 & N11534;
  assign N1478 = N11515 & N11535;
  assign N1477 = N11515 & N11536;
  assign N1476 = N11515 & N11537;
  assign N1475 = N11515 & N11538;
  assign N1474 = N11529 & N11516;
  assign N1473 = N11529 & N11517;
  assign N1472 = N11529 & N11518;
  assign N1471 = N11530 & N11516;
  assign N1470 = N11530 & N11517;
  assign N1469 = N11530 & N11518;
  assign N1468 = N11531 & N11516;
  assign N1467 = N11531 & N11517;
  assign N1466 = N11531 & N11518;
  assign N1465 = N11532 & N11516;
  assign N1464 = N11532 & N11517;
  assign N1463 = N11532 & N11518;
  assign N1462 = N11533 & N11516;
  assign N1461 = N11533 & N11517;
  assign N1460 = N11533 & N11518;
  assign N2091 = N11519 & N11535;
  assign N2090 = N11519 & N11536;
  assign N2089 = N11519 & N11537;
  assign N2088 = N11519 & N11538;
  assign N2087 = N11530 & N11524;
  assign N2086 = N11531 & N11524;
  assign N2085 = N11532 & N11524;
  assign N2084 = N11533 & N11524;
  assign N11519 = addr_i[5] & N11542;
  assign N11520 = N11497 & N11539;
  assign N11521 = N11497 & N11540;
  assign N11522 = N11497 & N11541;
  assign N11523 = N11497 & N11542;
  assign N11524 = addr_i[2] & N11554;
  assign N11525 = N11502 & N11551;
  assign N11526 = N11502 & N11552;
  assign N11527 = N11502 & N11553;
  assign N11528 = N11502 & N11554;
  assign N2211 = N11543 & N11524;
  assign N2210 = N11543 & N11525;
  assign N2209 = N11543 & N11526;
  assign N2208 = N11543 & N11527;
  assign N2207 = N11543 & N11528;
  assign N2206 = N11544 & N11524;
  assign N2205 = N11544 & N11525;
  assign N2204 = N11544 & N11526;
  assign N2203 = N11544 & N11527;
  assign N2202 = N11544 & N11528;
  assign N2201 = N11545 & N11524;
  assign N2200 = N11545 & N11525;
  assign N2199 = N11545 & N11526;
  assign N2198 = N11545 & N11527;
  assign N2197 = N11545 & N11528;
  assign N2196 = N11519 & N11555;
  assign N2195 = N11519 & N11556;
  assign N2194 = N11519 & N11557;
  assign N2193 = N11519 & N11524;
  assign N2192 = N11519 & N11525;
  assign N2191 = N11519 & N11526;
  assign N2190 = N11519 & N11527;
  assign N2189 = N11519 & N11528;
  assign N2188 = N11520 & N11555;
  assign N2187 = N11520 & N11556;
  assign N2186 = N11520 & N11557;
  assign N2185 = N11520 & N11524;
  assign N2184 = N11520 & N11525;
  assign N2183 = N11520 & N11526;
  assign N2182 = N11520 & N11527;
  assign N2181 = N11520 & N11528;
  assign N2180 = N11521 & N11555;
  assign N2179 = N11521 & N11556;
  assign N2178 = N11521 & N11557;
  assign N2177 = N11521 & N11524;
  assign N2176 = N11521 & N11525;
  assign N2175 = N11521 & N11526;
  assign N2174 = N11521 & N11527;
  assign N2173 = N11521 & N11528;
  assign N2172 = N11522 & N11555;
  assign N2171 = N11522 & N11556;
  assign N2170 = N11522 & N11557;
  assign N2169 = N11522 & N11524;
  assign N2168 = N11522 & N11525;
  assign N2167 = N11522 & N11526;
  assign N2166 = N11522 & N11527;
  assign N2165 = N11522 & N11528;
  assign N2164 = N11523 & N11555;
  assign N2163 = N11523 & N11556;
  assign N2162 = N11523 & N11557;
  assign N2161 = N11523 & N11524;
  assign N2160 = N11523 & N11525;
  assign N2159 = N11523 & N11526;
  assign N2158 = N11523 & N11527;
  assign N2157 = N11523 & N11528;
  assign N11529 = addr_i[5] & N11542;
  assign N11530 = N11497 & N11539;
  assign N11531 = N11497 & N11540;
  assign N11532 = N11497 & N11541;
  assign N11533 = N11497 & N11542;
  assign N11534 = addr_i[2] & N11554;
  assign N11535 = N11502 & N11551;
  assign N11536 = N11502 & N11552;
  assign N11537 = N11502 & N11553;
  assign N11538 = N11502 & N11554;
  assign N2331 = N11543 & N11534;
  assign N2330 = N11543 & N11535;
  assign N2329 = N11543 & N11536;
  assign N2328 = N11543 & N11537;
  assign N2327 = N11543 & N11538;
  assign N2326 = N11544 & N11534;
  assign N2325 = N11544 & N11535;
  assign N2324 = N11544 & N11536;
  assign N2323 = N11544 & N11537;
  assign N2322 = N11544 & N11538;
  assign N2321 = N11545 & N11534;
  assign N2320 = N11545 & N11535;
  assign N2319 = N11545 & N11536;
  assign N2318 = N11545 & N11537;
  assign N2317 = N11545 & N11538;
  assign N2316 = N11529 & N11555;
  assign N2315 = N11529 & N11556;
  assign N2314 = N11529 & N11557;
  assign N2313 = N11529 & N11534;
  assign N2312 = N11529 & N11535;
  assign N2311 = N11529 & N11536;
  assign N2310 = N11529 & N11537;
  assign N2309 = N11529 & N11538;
  assign N2308 = N11530 & N11555;
  assign N2307 = N11530 & N11556;
  assign N2306 = N11530 & N11557;
  assign N2305 = N11530 & N11534;
  assign N2304 = N11530 & N11535;
  assign N2303 = N11530 & N11536;
  assign N2302 = N11530 & N11537;
  assign N2301 = N11530 & N11538;
  assign N2300 = N11531 & N11555;
  assign N2299 = N11531 & N11556;
  assign N2298 = N11531 & N11557;
  assign N2297 = N11531 & N11534;
  assign N2296 = N11531 & N11535;
  assign N2295 = N11531 & N11536;
  assign N2294 = N11531 & N11537;
  assign N2293 = N11531 & N11538;
  assign N2292 = N11532 & N11555;
  assign N2291 = N11532 & N11556;
  assign N2290 = N11532 & N11557;
  assign N2289 = N11532 & N11534;
  assign N2288 = N11532 & N11535;
  assign N2287 = N11532 & N11536;
  assign N2286 = N11532 & N11537;
  assign N2285 = N11532 & N11538;
  assign N2284 = N11533 & N11555;
  assign N2283 = N11533 & N11556;
  assign N2282 = N11533 & N11557;
  assign N2281 = N11533 & N11534;
  assign N2280 = N11533 & N11535;
  assign N2279 = N11533 & N11536;
  assign N2278 = N11533 & N11537;
  assign N2277 = N11533 & N11538;
  assign N11539 = addr_i[3] & addr_i[4];
  assign N11540 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N11541 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N11542 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N11543 = addr_i[5] & N11539;
  assign N11544 = addr_i[5] & N11540;
  assign N11545 = addr_i[5] & N11541;
  assign N11546 = addr_i[5] & N11542;
  assign N11547 = N11497 & N11539;
  assign N11548 = N11497 & N11540;
  assign N11549 = N11497 & N11541;
  assign N11550 = N11497 & N11542;
  assign N11551 = addr_i[0] & addr_i[1];
  assign N11552 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N11553 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N11554 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N11555 = addr_i[2] & N11551;
  assign N11556 = addr_i[2] & N11552;
  assign N11557 = addr_i[2] & N11553;
  assign N11558 = addr_i[2] & N11554;
  assign N11559 = N11502 & N11551;
  assign N11560 = N11502 & N11552;
  assign N11561 = N11502 & N11553;
  assign N11562 = N11502 & N11554;
  assign N2460 = N11543 & N11555;
  assign N2459 = N11543 & N11556;
  assign N2458 = N11543 & N11557;
  assign N2457 = N11543 & N11558;
  assign N2456 = N11543 & N11559;
  assign N2455 = N11543 & N11560;
  assign N2454 = N11543 & N11561;
  assign N2453 = N11543 & N11562;
  assign N2452 = N11544 & N11555;
  assign N2451 = N11544 & N11556;
  assign N2450 = N11544 & N11557;
  assign N2449 = N11544 & N11558;
  assign N2448 = N11544 & N11559;
  assign N2447 = N11544 & N11560;
  assign N2446 = N11544 & N11561;
  assign N2445 = N11544 & N11562;
  assign N2444 = N11545 & N11555;
  assign N2443 = N11545 & N11556;
  assign N2442 = N11545 & N11557;
  assign N2441 = N11545 & N11558;
  assign N2440 = N11545 & N11559;
  assign N2439 = N11545 & N11560;
  assign N2438 = N11545 & N11561;
  assign N2437 = N11545 & N11562;
  assign N2436 = N11546 & N11555;
  assign N2435 = N11546 & N11556;
  assign N2434 = N11546 & N11557;
  assign N2433 = N11546 & N11558;
  assign N2432 = N11546 & N11559;
  assign N2431 = N11546 & N11560;
  assign N2430 = N11546 & N11561;
  assign N2429 = N11546 & N11562;
  assign N2428 = N11547 & N11555;
  assign N2427 = N11547 & N11556;
  assign N2426 = N11547 & N11557;
  assign N2425 = N11547 & N11558;
  assign N2424 = N11547 & N11559;
  assign N2423 = N11547 & N11560;
  assign N2422 = N11547 & N11561;
  assign N2421 = N11547 & N11562;
  assign N2420 = N11548 & N11555;
  assign N2419 = N11548 & N11556;
  assign N2418 = N11548 & N11557;
  assign N2417 = N11548 & N11558;
  assign N2416 = N11548 & N11559;
  assign N2415 = N11548 & N11560;
  assign N2414 = N11548 & N11561;
  assign N2413 = N11548 & N11562;
  assign N2412 = N11549 & N11555;
  assign N2411 = N11549 & N11556;
  assign N2410 = N11549 & N11557;
  assign N2409 = N11549 & N11558;
  assign N2408 = N11549 & N11559;
  assign N2407 = N11549 & N11560;
  assign N2406 = N11549 & N11561;
  assign N2405 = N11549 & N11562;
  assign N2404 = N11550 & N11555;
  assign N2403 = N11550 & N11556;
  assign N2402 = N11550 & N11557;
  assign N2401 = N11550 & N11558;
  assign N2400 = N11550 & N11559;
  assign N2399 = N11550 & N11560;
  assign N2398 = N11550 & N11561;
  assign N2397 = N11550 & N11562;
  assign N11563 = addr_i[5] & N11635;
  assign N11564 = addr_i[5] & N11636;
  assign N11565 = addr_i[5] & N11637;
  assign N11566 = addr_i[2] & N11647;
  assign N11567 = addr_i[2] & N11648;
  assign N11568 = addr_i[2] & N11649;
  assign N2629 = N11563 & N11566;
  assign N2628 = N11563 & N11567;
  assign N2627 = N11563 & N11568;
  assign N2626 = N11563 & N11654;
  assign N2625 = N11563 & N11595;
  assign N2624 = N11563 & N11596;
  assign N2623 = N11563 & N11597;
  assign N2622 = N11563 & N11598;
  assign N2621 = N11564 & N11566;
  assign N2620 = N11564 & N11567;
  assign N2619 = N11564 & N11568;
  assign N2618 = N11564 & N11654;
  assign N2617 = N11564 & N11595;
  assign N2616 = N11564 & N11596;
  assign N2615 = N11564 & N11597;
  assign N2614 = N11564 & N11598;
  assign N2613 = N11565 & N11566;
  assign N2612 = N11565 & N11567;
  assign N2611 = N11565 & N11568;
  assign N2610 = N11565 & N11654;
  assign N2609 = N11565 & N11595;
  assign N2608 = N11565 & N11596;
  assign N2607 = N11565 & N11597;
  assign N2606 = N11565 & N11598;
  assign N2605 = N11642 & N11566;
  assign N2604 = N11642 & N11567;
  assign N2603 = N11642 & N11568;
  assign N2602 = N11591 & N11566;
  assign N2601 = N11591 & N11567;
  assign N2600 = N11591 & N11568;
  assign N2599 = N11592 & N11566;
  assign N2598 = N11592 & N11567;
  assign N2597 = N11592 & N11568;
  assign N2596 = N11593 & N11566;
  assign N2595 = N11593 & N11567;
  assign N2594 = N11593 & N11568;
  assign N2593 = N11594 & N11566;
  assign N2592 = N11594 & N11567;
  assign N2591 = N11594 & N11568;
  assign N3252 = N11569 & N11654;
  assign N3251 = N11569 & N11595;
  assign N3250 = N11569 & N11596;
  assign N3249 = N11569 & N11597;
  assign N3248 = N11569 & N11598;
  assign N3247 = N11570 & N11654;
  assign N3246 = N11570 & N11595;
  assign N3245 = N11570 & N11596;
  assign N3244 = N11570 & N11597;
  assign N3243 = N11570 & N11598;
  assign N3242 = N11571 & N11654;
  assign N3241 = N11571 & N11595;
  assign N3240 = N11571 & N11596;
  assign N3239 = N11571 & N11597;
  assign N3238 = N11571 & N11598;
  assign N3237 = N11642 & N11572;
  assign N3236 = N11642 & N11573;
  assign N3235 = N11642 & N11574;
  assign N3234 = N11642 & N11595;
  assign N3233 = N11642 & N11596;
  assign N3232 = N11642 & N11597;
  assign N3231 = N11642 & N11598;
  assign N3230 = N11591 & N11572;
  assign N3229 = N11591 & N11573;
  assign N3228 = N11591 & N11574;
  assign N3227 = N11591 & N11654;
  assign N3226 = N11592 & N11572;
  assign N3225 = N11592 & N11573;
  assign N3224 = N11592 & N11574;
  assign N3223 = N11592 & N11654;
  assign N3222 = N11593 & N11572;
  assign N3221 = N11593 & N11573;
  assign N3220 = N11593 & N11574;
  assign N3219 = N11593 & N11654;
  assign N3218 = N11594 & N11572;
  assign N3217 = N11594 & N11573;
  assign N3216 = N11594 & N11574;
  assign N3215 = N11594 & N11654;
  assign N11569 = addr_i[5] & N11635;
  assign N11570 = addr_i[5] & N11636;
  assign N11571 = addr_i[5] & N11637;
  assign N11572 = addr_i[2] & N11647;
  assign N11573 = addr_i[2] & N11648;
  assign N11574 = addr_i[2] & N11649;
  assign N3486 = N11569 & N11572;
  assign N3485 = N11569 & N11573;
  assign N3484 = N11569 & N11574;
  assign N3483 = N11569 & N11630;
  assign N3482 = N11569 & N11587;
  assign N3481 = N11569 & N11588;
  assign N3480 = N11569 & N11589;
  assign N3479 = N11569 & N11590;
  assign N3478 = N11570 & N11572;
  assign N3477 = N11570 & N11573;
  assign N3476 = N11570 & N11574;
  assign N3475 = N11570 & N11630;
  assign N3474 = N11570 & N11587;
  assign N3473 = N11570 & N11588;
  assign N3472 = N11570 & N11589;
  assign N3471 = N11570 & N11590;
  assign N3470 = N11571 & N11572;
  assign N3469 = N11571 & N11573;
  assign N3468 = N11571 & N11574;
  assign N3467 = N11571 & N11630;
  assign N3466 = N11571 & N11587;
  assign N3465 = N11571 & N11588;
  assign N3464 = N11571 & N11589;
  assign N3463 = N11571 & N11590;
  assign N3462 = N11625 & N11572;
  assign N3461 = N11625 & N11573;
  assign N3460 = N11625 & N11574;
  assign N3459 = N11583 & N11572;
  assign N3458 = N11583 & N11573;
  assign N3457 = N11583 & N11574;
  assign N3456 = N11584 & N11572;
  assign N3455 = N11584 & N11573;
  assign N3454 = N11584 & N11574;
  assign N3453 = N11585 & N11572;
  assign N3452 = N11585 & N11573;
  assign N3451 = N11585 & N11574;
  assign N3450 = N11586 & N11572;
  assign N3449 = N11586 & N11573;
  assign N3448 = N11586 & N11574;
  assign N4020 = N11599 & N11630;
  assign N4019 = N11600 & N11630;
  assign N4018 = N11601 & N11630;
  assign N4017 = N11625 & N11602;
  assign N4016 = N11625 & N11603;
  assign N4015 = N11625 & N11604;
  assign N4014 = N11625 & N11587;
  assign N4013 = N11625 & N11588;
  assign N4012 = N11625 & N11589;
  assign N4011 = N11625 & N11590;
  assign N4010 = N11583 & N11630;
  assign N4009 = N11584 & N11630;
  assign N4008 = N11585 & N11630;
  assign N4007 = N11586 & N11630;
  assign N11575 = N11497 & N11635;
  assign N11576 = N11497 & N11636;
  assign N11577 = N11497 & N11637;
  assign N11578 = N11497 & N11638;
  assign N11579 = N11502 & N11647;
  assign N11580 = N11502 & N11648;
  assign N11581 = N11502 & N11649;
  assign N11582 = N11502 & N11650;
  assign N4133 = N11599 & N11579;
  assign N4132 = N11599 & N11580;
  assign N4131 = N11599 & N11581;
  assign N4130 = N11599 & N11582;
  assign N4129 = N11600 & N11579;
  assign N4128 = N11600 & N11580;
  assign N4127 = N11600 & N11581;
  assign N4126 = N11600 & N11582;
  assign N4125 = N11601 & N11579;
  assign N4124 = N11601 & N11580;
  assign N4123 = N11601 & N11581;
  assign N4122 = N11601 & N11582;
  assign N4121 = N11615 & N11579;
  assign N4120 = N11615 & N11580;
  assign N4119 = N11615 & N11581;
  assign N4118 = N11615 & N11582;
  assign N4117 = N11575 & N11602;
  assign N4116 = N11575 & N11603;
  assign N4115 = N11575 & N11604;
  assign N4114 = N11575 & N11620;
  assign N4113 = N11575 & N11579;
  assign N4112 = N11575 & N11580;
  assign N4111 = N11575 & N11581;
  assign N4110 = N11575 & N11582;
  assign N4109 = N11576 & N11602;
  assign N4108 = N11576 & N11603;
  assign N4107 = N11576 & N11604;
  assign N4106 = N11576 & N11620;
  assign N4105 = N11576 & N11579;
  assign N4104 = N11576 & N11580;
  assign N4103 = N11576 & N11581;
  assign N4102 = N11576 & N11582;
  assign N4101 = N11577 & N11602;
  assign N4100 = N11577 & N11603;
  assign N4099 = N11577 & N11604;
  assign N4098 = N11577 & N11620;
  assign N4097 = N11577 & N11579;
  assign N4096 = N11577 & N11580;
  assign N4095 = N11577 & N11581;
  assign N4094 = N11577 & N11582;
  assign N4093 = N11578 & N11602;
  assign N4092 = N11578 & N11603;
  assign N4091 = N11578 & N11604;
  assign N4090 = N11578 & N11620;
  assign N4089 = N11578 & N11579;
  assign N4088 = N11578 & N11580;
  assign N4087 = N11578 & N11581;
  assign N4086 = N11578 & N11582;
  assign N11583 = N11497 & N11635;
  assign N11584 = N11497 & N11636;
  assign N11585 = N11497 & N11637;
  assign N11586 = N11497 & N11638;
  assign N11587 = N11502 & N11647;
  assign N11588 = N11502 & N11648;
  assign N11589 = N11502 & N11649;
  assign N11590 = N11502 & N11650;
  assign N4246 = N11599 & N11587;
  assign N4245 = N11599 & N11588;
  assign N4244 = N11599 & N11589;
  assign N4243 = N11599 & N11590;
  assign N4242 = N11600 & N11587;
  assign N4241 = N11600 & N11588;
  assign N4240 = N11600 & N11589;
  assign N4239 = N11600 & N11590;
  assign N4238 = N11601 & N11587;
  assign N4237 = N11601 & N11588;
  assign N4236 = N11601 & N11589;
  assign N4235 = N11601 & N11590;
  assign N4234 = N11615 & N11587;
  assign N4233 = N11615 & N11588;
  assign N4232 = N11615 & N11589;
  assign N4231 = N11615 & N11590;
  assign N4230 = N11583 & N11602;
  assign N4229 = N11583 & N11603;
  assign N4228 = N11583 & N11604;
  assign N4227 = N11583 & N11620;
  assign N4226 = N11583 & N11587;
  assign N4225 = N11583 & N11588;
  assign N4224 = N11583 & N11589;
  assign N4223 = N11583 & N11590;
  assign N4222 = N11584 & N11602;
  assign N4221 = N11584 & N11603;
  assign N4220 = N11584 & N11604;
  assign N4219 = N11584 & N11620;
  assign N4218 = N11584 & N11587;
  assign N4217 = N11584 & N11588;
  assign N4216 = N11584 & N11589;
  assign N4215 = N11584 & N11590;
  assign N4214 = N11585 & N11602;
  assign N4213 = N11585 & N11603;
  assign N4212 = N11585 & N11604;
  assign N4211 = N11585 & N11620;
  assign N4210 = N11585 & N11587;
  assign N4209 = N11585 & N11588;
  assign N4208 = N11585 & N11589;
  assign N4207 = N11585 & N11590;
  assign N4206 = N11586 & N11602;
  assign N4205 = N11586 & N11603;
  assign N4204 = N11586 & N11604;
  assign N4203 = N11586 & N11620;
  assign N4202 = N11586 & N11587;
  assign N4201 = N11586 & N11588;
  assign N4200 = N11586 & N11589;
  assign N4199 = N11586 & N11590;
  assign N11591 = N11497 & N11635;
  assign N11592 = N11497 & N11636;
  assign N11593 = N11497 & N11637;
  assign N11594 = N11497 & N11638;
  assign N11595 = N11502 & N11647;
  assign N11596 = N11502 & N11648;
  assign N11597 = N11502 & N11649;
  assign N11598 = N11502 & N11650;
  assign N4359 = N11599 & N11595;
  assign N4358 = N11599 & N11596;
  assign N4357 = N11599 & N11597;
  assign N4356 = N11599 & N11598;
  assign N4355 = N11600 & N11595;
  assign N4354 = N11600 & N11596;
  assign N4353 = N11600 & N11597;
  assign N4352 = N11600 & N11598;
  assign N4351 = N11601 & N11595;
  assign N4350 = N11601 & N11596;
  assign N4349 = N11601 & N11597;
  assign N4348 = N11601 & N11598;
  assign N4347 = N11615 & N11595;
  assign N4346 = N11615 & N11596;
  assign N4345 = N11615 & N11597;
  assign N4344 = N11615 & N11598;
  assign N4343 = N11591 & N11602;
  assign N4342 = N11591 & N11603;
  assign N4341 = N11591 & N11604;
  assign N4340 = N11591 & N11620;
  assign N4339 = N11591 & N11595;
  assign N4338 = N11591 & N11596;
  assign N4337 = N11591 & N11597;
  assign N4336 = N11591 & N11598;
  assign N4335 = N11592 & N11602;
  assign N4334 = N11592 & N11603;
  assign N4333 = N11592 & N11604;
  assign N4332 = N11592 & N11620;
  assign N4331 = N11592 & N11595;
  assign N4330 = N11592 & N11596;
  assign N4329 = N11592 & N11597;
  assign N4328 = N11592 & N11598;
  assign N4327 = N11593 & N11602;
  assign N4326 = N11593 & N11603;
  assign N4325 = N11593 & N11604;
  assign N4324 = N11593 & N11620;
  assign N4323 = N11593 & N11595;
  assign N4322 = N11593 & N11596;
  assign N4321 = N11593 & N11597;
  assign N4320 = N11593 & N11598;
  assign N4319 = N11594 & N11602;
  assign N4318 = N11594 & N11603;
  assign N4317 = N11594 & N11604;
  assign N4316 = N11594 & N11620;
  assign N4315 = N11594 & N11595;
  assign N4314 = N11594 & N11596;
  assign N4313 = N11594 & N11597;
  assign N4312 = N11594 & N11598;
  assign N11599 = addr_i[5] & N11635;
  assign N11600 = addr_i[5] & N11636;
  assign N11601 = addr_i[5] & N11637;
  assign N11602 = addr_i[2] & N11647;
  assign N11603 = addr_i[2] & N11648;
  assign N11604 = addr_i[2] & N11649;
  assign N4463 = N11599 & N11602;
  assign N4462 = N11599 & N11603;
  assign N4461 = N11599 & N11604;
  assign N4460 = N11599 & N11620;
  assign N4459 = N11599 & N11655;
  assign N4458 = N11599 & N11656;
  assign N4457 = N11599 & N11657;
  assign N4456 = N11599 & N11658;
  assign N4455 = N11600 & N11602;
  assign N4454 = N11600 & N11603;
  assign N4453 = N11600 & N11604;
  assign N4452 = N11600 & N11620;
  assign N4451 = N11600 & N11655;
  assign N4450 = N11600 & N11656;
  assign N4449 = N11600 & N11657;
  assign N4448 = N11600 & N11658;
  assign N4447 = N11601 & N11602;
  assign N4446 = N11601 & N11603;
  assign N4445 = N11601 & N11604;
  assign N4444 = N11601 & N11620;
  assign N4443 = N11601 & N11655;
  assign N4442 = N11601 & N11656;
  assign N4441 = N11601 & N11657;
  assign N4440 = N11601 & N11658;
  assign N4439 = N11615 & N11602;
  assign N4438 = N11615 & N11603;
  assign N4437 = N11615 & N11604;
  assign N4436 = N11643 & N11602;
  assign N4435 = N11643 & N11603;
  assign N4434 = N11643 & N11604;
  assign N4433 = N11644 & N11602;
  assign N4432 = N11644 & N11603;
  assign N4431 = N11644 & N11604;
  assign N4430 = N11645 & N11602;
  assign N4429 = N11645 & N11603;
  assign N4428 = N11645 & N11604;
  assign N4427 = N11646 & N11602;
  assign N4426 = N11646 & N11603;
  assign N4425 = N11646 & N11604;
  assign N4932 = N11605 & N11620;
  assign N4931 = N11606 & N11620;
  assign N4930 = N11607 & N11620;
  assign N4929 = N11615 & N11608;
  assign N4928 = N11615 & N11609;
  assign N4927 = N11615 & N11610;
  assign N4926 = N11615 & N11655;
  assign N4925 = N11615 & N11656;
  assign N4924 = N11615 & N11657;
  assign N4923 = N11615 & N11658;
  assign N4922 = N11643 & N11620;
  assign N4921 = N11644 & N11620;
  assign N4920 = N11645 & N11620;
  assign N4919 = N11646 & N11620;
  assign N5159 = N11605 & N11655;
  assign N5158 = N11605 & N11656;
  assign N5157 = N11605 & N11657;
  assign N5156 = N11605 & N11658;
  assign N5155 = N11606 & N11655;
  assign N5154 = N11606 & N11656;
  assign N5153 = N11606 & N11657;
  assign N5152 = N11606 & N11658;
  assign N5151 = N11607 & N11655;
  assign N5150 = N11607 & N11656;
  assign N5149 = N11607 & N11657;
  assign N5148 = N11607 & N11658;
  assign N5147 = N11613 & N11655;
  assign N5146 = N11613 & N11656;
  assign N5145 = N11613 & N11657;
  assign N5144 = N11613 & N11658;
  assign N5143 = N11643 & N11608;
  assign N5142 = N11643 & N11609;
  assign N5141 = N11643 & N11610;
  assign N5140 = N11643 & N11614;
  assign N5139 = N11644 & N11608;
  assign N5138 = N11644 & N11609;
  assign N5137 = N11644 & N11610;
  assign N5136 = N11644 & N11614;
  assign N5135 = N11645 & N11608;
  assign N5134 = N11645 & N11609;
  assign N5133 = N11645 & N11610;
  assign N5132 = N11645 & N11614;
  assign N5131 = N11646 & N11608;
  assign N5130 = N11646 & N11609;
  assign N5129 = N11646 & N11610;
  assign N5128 = N11646 & N11614;
  assign N11605 = addr_i[5] & N11635;
  assign N11606 = addr_i[5] & N11636;
  assign N11607 = addr_i[5] & N11637;
  assign N11608 = addr_i[2] & N11647;
  assign N11609 = addr_i[2] & N11648;
  assign N11610 = addr_i[2] & N11649;
  assign N5328 = N11605 & N11608;
  assign N5327 = N11605 & N11609;
  assign N5326 = N11605 & N11610;
  assign N5325 = N11605 & N11614;
  assign N5324 = N11605 & N11631;
  assign N5323 = N11605 & N11632;
  assign N5322 = N11605 & N11633;
  assign N5321 = N11605 & N11634;
  assign N5320 = N11606 & N11608;
  assign N5319 = N11606 & N11609;
  assign N5318 = N11606 & N11610;
  assign N5317 = N11606 & N11614;
  assign N5316 = N11606 & N11631;
  assign N5315 = N11606 & N11632;
  assign N5314 = N11606 & N11633;
  assign N5313 = N11606 & N11634;
  assign N5312 = N11607 & N11608;
  assign N5311 = N11607 & N11609;
  assign N5310 = N11607 & N11610;
  assign N5309 = N11607 & N11614;
  assign N5308 = N11607 & N11631;
  assign N5307 = N11607 & N11632;
  assign N5306 = N11607 & N11633;
  assign N5305 = N11607 & N11634;
  assign N5304 = N11613 & N11608;
  assign N5303 = N11613 & N11609;
  assign N5302 = N11613 & N11610;
  assign N5301 = N11626 & N11608;
  assign N5300 = N11626 & N11609;
  assign N5299 = N11626 & N11610;
  assign N5298 = N11627 & N11608;
  assign N5297 = N11627 & N11609;
  assign N5296 = N11627 & N11610;
  assign N5295 = N11628 & N11608;
  assign N5294 = N11628 & N11609;
  assign N5293 = N11628 & N11610;
  assign N5292 = N11629 & N11608;
  assign N5291 = N11629 & N11609;
  assign N5290 = N11629 & N11610;
  assign N11611 = addr_i[5] & N11638;
  assign N11612 = addr_i[2] & N11650;
  assign N5863 = N11639 & N11612;
  assign N5862 = N11640 & N11612;
  assign N5861 = N11641 & N11612;
  assign N5860 = N11611 & N11651;
  assign N5859 = N11611 & N11652;
  assign N5858 = N11611 & N11653;
  assign N5857 = N11611 & N11612;
  assign N5856 = N11611 & N11631;
  assign N5855 = N11611 & N11632;
  assign N5854 = N11611 & N11633;
  assign N5853 = N11611 & N11634;
  assign N5852 = N11626 & N11612;
  assign N5851 = N11627 & N11612;
  assign N5850 = N11628 & N11612;
  assign N5849 = N11629 & N11612;
  assign N11613 = addr_i[5] & N11638;
  assign N11614 = addr_i[2] & N11650;
  assign N5943 = N11639 & N11614;
  assign N5942 = N11640 & N11614;
  assign N5941 = N11641 & N11614;
  assign N5940 = N11613 & N11651;
  assign N5939 = N11613 & N11652;
  assign N5938 = N11613 & N11653;
  assign N5937 = N11613 & N11614;
  assign N5936 = N11613 & N11631;
  assign N5935 = N11613 & N11632;
  assign N5934 = N11613 & N11633;
  assign N5933 = N11613 & N11634;
  assign N5932 = N11626 & N11614;
  assign N5931 = N11627 & N11614;
  assign N5930 = N11628 & N11614;
  assign N5929 = N11629 & N11614;
  assign N11615 = addr_i[5] & N11638;
  assign N11616 = N11497 & N11635;
  assign N11617 = N11497 & N11636;
  assign N11618 = N11497 & N11637;
  assign N11619 = N11497 & N11638;
  assign N11620 = addr_i[2] & N11650;
  assign N11621 = N11502 & N11647;
  assign N11622 = N11502 & N11648;
  assign N11623 = N11502 & N11649;
  assign N11624 = N11502 & N11650;
  assign N6063 = N11639 & N11620;
  assign N6062 = N11639 & N11621;
  assign N6061 = N11639 & N11622;
  assign N6060 = N11639 & N11623;
  assign N6059 = N11639 & N11624;
  assign N6058 = N11640 & N11620;
  assign N6057 = N11640 & N11621;
  assign N6056 = N11640 & N11622;
  assign N6055 = N11640 & N11623;
  assign N6054 = N11640 & N11624;
  assign N6053 = N11641 & N11620;
  assign N6052 = N11641 & N11621;
  assign N6051 = N11641 & N11622;
  assign N6050 = N11641 & N11623;
  assign N6049 = N11641 & N11624;
  assign N6048 = N11615 & N11651;
  assign N6047 = N11615 & N11652;
  assign N6046 = N11615 & N11653;
  assign N6045 = N11615 & N11620;
  assign N6044 = N11615 & N11621;
  assign N6043 = N11615 & N11622;
  assign N6042 = N11615 & N11623;
  assign N6041 = N11615 & N11624;
  assign N6040 = N11616 & N11651;
  assign N6039 = N11616 & N11652;
  assign N6038 = N11616 & N11653;
  assign N6037 = N11616 & N11620;
  assign N6036 = N11616 & N11621;
  assign N6035 = N11616 & N11622;
  assign N6034 = N11616 & N11623;
  assign N6033 = N11616 & N11624;
  assign N6032 = N11617 & N11651;
  assign N6031 = N11617 & N11652;
  assign N6030 = N11617 & N11653;
  assign N6029 = N11617 & N11620;
  assign N6028 = N11617 & N11621;
  assign N6027 = N11617 & N11622;
  assign N6026 = N11617 & N11623;
  assign N6025 = N11617 & N11624;
  assign N6024 = N11618 & N11651;
  assign N6023 = N11618 & N11652;
  assign N6022 = N11618 & N11653;
  assign N6021 = N11618 & N11620;
  assign N6020 = N11618 & N11621;
  assign N6019 = N11618 & N11622;
  assign N6018 = N11618 & N11623;
  assign N6017 = N11618 & N11624;
  assign N6016 = N11619 & N11651;
  assign N6015 = N11619 & N11652;
  assign N6014 = N11619 & N11653;
  assign N6013 = N11619 & N11620;
  assign N6012 = N11619 & N11621;
  assign N6011 = N11619 & N11622;
  assign N6010 = N11619 & N11623;
  assign N6009 = N11619 & N11624;
  assign N11625 = addr_i[5] & N11638;
  assign N11626 = N11497 & N11635;
  assign N11627 = N11497 & N11636;
  assign N11628 = N11497 & N11637;
  assign N11629 = N11497 & N11638;
  assign N11630 = addr_i[2] & N11650;
  assign N11631 = N11502 & N11647;
  assign N11632 = N11502 & N11648;
  assign N11633 = N11502 & N11649;
  assign N11634 = N11502 & N11650;
  assign N6183 = N11639 & N11630;
  assign N6182 = N11639 & N11631;
  assign N6181 = N11639 & N11632;
  assign N6180 = N11639 & N11633;
  assign N6179 = N11639 & N11634;
  assign N6178 = N11640 & N11630;
  assign N6177 = N11640 & N11631;
  assign N6176 = N11640 & N11632;
  assign N6175 = N11640 & N11633;
  assign N6174 = N11640 & N11634;
  assign N6173 = N11641 & N11630;
  assign N6172 = N11641 & N11631;
  assign N6171 = N11641 & N11632;
  assign N6170 = N11641 & N11633;
  assign N6169 = N11641 & N11634;
  assign N6168 = N11625 & N11651;
  assign N6167 = N11625 & N11652;
  assign N6166 = N11625 & N11653;
  assign N6165 = N11625 & N11630;
  assign N6164 = N11625 & N11631;
  assign N6163 = N11625 & N11632;
  assign N6162 = N11625 & N11633;
  assign N6161 = N11625 & N11634;
  assign N6160 = N11626 & N11651;
  assign N6159 = N11626 & N11652;
  assign N6158 = N11626 & N11653;
  assign N6157 = N11626 & N11630;
  assign N6156 = N11626 & N11631;
  assign N6155 = N11626 & N11632;
  assign N6154 = N11626 & N11633;
  assign N6153 = N11626 & N11634;
  assign N6152 = N11627 & N11651;
  assign N6151 = N11627 & N11652;
  assign N6150 = N11627 & N11653;
  assign N6149 = N11627 & N11630;
  assign N6148 = N11627 & N11631;
  assign N6147 = N11627 & N11632;
  assign N6146 = N11627 & N11633;
  assign N6145 = N11627 & N11634;
  assign N6144 = N11628 & N11651;
  assign N6143 = N11628 & N11652;
  assign N6142 = N11628 & N11653;
  assign N6141 = N11628 & N11630;
  assign N6140 = N11628 & N11631;
  assign N6139 = N11628 & N11632;
  assign N6138 = N11628 & N11633;
  assign N6137 = N11628 & N11634;
  assign N6136 = N11629 & N11651;
  assign N6135 = N11629 & N11652;
  assign N6134 = N11629 & N11653;
  assign N6133 = N11629 & N11630;
  assign N6132 = N11629 & N11631;
  assign N6131 = N11629 & N11632;
  assign N6130 = N11629 & N11633;
  assign N6129 = N11629 & N11634;
  assign N11635 = addr_i[3] & addr_i[4];
  assign N11636 = N8 & addr_i[4];
  assign N8 = ~addr_i[3];
  assign N11637 = addr_i[3] & N9;
  assign N9 = ~addr_i[4];
  assign N11638 = N10 & N11;
  assign N10 = ~addr_i[3];
  assign N11 = ~addr_i[4];
  assign N11639 = addr_i[5] & N11635;
  assign N11640 = addr_i[5] & N11636;
  assign N11641 = addr_i[5] & N11637;
  assign N11642 = addr_i[5] & N11638;
  assign N11643 = N11497 & N11635;
  assign N11644 = N11497 & N11636;
  assign N11645 = N11497 & N11637;
  assign N11646 = N11497 & N11638;
  assign N11647 = addr_i[0] & addr_i[1];
  assign N11648 = N12 & addr_i[1];
  assign N12 = ~addr_i[0];
  assign N11649 = addr_i[0] & N13;
  assign N13 = ~addr_i[1];
  assign N11650 = N14 & N15;
  assign N14 = ~addr_i[0];
  assign N15 = ~addr_i[1];
  assign N11651 = addr_i[2] & N11647;
  assign N11652 = addr_i[2] & N11648;
  assign N11653 = addr_i[2] & N11649;
  assign N11654 = addr_i[2] & N11650;
  assign N11655 = N11502 & N11647;
  assign N11656 = N11502 & N11648;
  assign N11657 = N11502 & N11649;
  assign N11658 = N11502 & N11650;
  assign N6312 = N11639 & N11651;
  assign N6311 = N11639 & N11652;
  assign N6310 = N11639 & N11653;
  assign N6309 = N11639 & N11654;
  assign N6308 = N11639 & N11655;
  assign N6307 = N11639 & N11656;
  assign N6306 = N11639 & N11657;
  assign N6305 = N11639 & N11658;
  assign N6304 = N11640 & N11651;
  assign N6303 = N11640 & N11652;
  assign N6302 = N11640 & N11653;
  assign N6301 = N11640 & N11654;
  assign N6300 = N11640 & N11655;
  assign N6299 = N11640 & N11656;
  assign N6298 = N11640 & N11657;
  assign N6297 = N11640 & N11658;
  assign N6296 = N11641 & N11651;
  assign N6295 = N11641 & N11652;
  assign N6294 = N11641 & N11653;
  assign N6293 = N11641 & N11654;
  assign N6292 = N11641 & N11655;
  assign N6291 = N11641 & N11656;
  assign N6290 = N11641 & N11657;
  assign N6289 = N11641 & N11658;
  assign N6288 = N11642 & N11651;
  assign N6287 = N11642 & N11652;
  assign N6286 = N11642 & N11653;
  assign N6285 = N11642 & N11654;
  assign N6284 = N11642 & N11655;
  assign N6283 = N11642 & N11656;
  assign N6282 = N11642 & N11657;
  assign N6281 = N11642 & N11658;
  assign N6280 = N11643 & N11651;
  assign N6279 = N11643 & N11652;
  assign N6278 = N11643 & N11653;
  assign N6277 = N11643 & N11654;
  assign N6276 = N11643 & N11655;
  assign N6275 = N11643 & N11656;
  assign N6274 = N11643 & N11657;
  assign N6273 = N11643 & N11658;
  assign N6272 = N11644 & N11651;
  assign N6271 = N11644 & N11652;
  assign N6270 = N11644 & N11653;
  assign N6269 = N11644 & N11654;
  assign N6268 = N11644 & N11655;
  assign N6267 = N11644 & N11656;
  assign N6266 = N11644 & N11657;
  assign N6265 = N11644 & N11658;
  assign N6264 = N11645 & N11651;
  assign N6263 = N11645 & N11652;
  assign N6262 = N11645 & N11653;
  assign N6261 = N11645 & N11654;
  assign N6260 = N11645 & N11655;
  assign N6259 = N11645 & N11656;
  assign N6258 = N11645 & N11657;
  assign N6257 = N11645 & N11658;
  assign N6256 = N11646 & N11651;
  assign N6255 = N11646 & N11652;
  assign N6254 = N11646 & N11653;
  assign N6253 = N11646 & N11654;
  assign N6252 = N11646 & N11655;
  assign N6251 = N11646 & N11656;
  assign N6250 = N11646 & N11657;
  assign N6249 = N11646 & N11658;
  assign { N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230 } = (N16)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N229)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[0];
  assign { N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295 } = (N17)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N294)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[1];
  assign { N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360 } = (N18)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N359)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[2];
  assign { N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425 } = (N19)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N424)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[3];
  assign { N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538 } = (N20)? { N641, N640, N639, N638, N537, N536, N535, N534, N633, N632, N631, N630, N533, N532, N531, N530, N625, N624, N623, N622, N529, N528, N527, N526, N617, N616, N615, N2433, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N489)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[4];
  assign { N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642 } = (N21)? { N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N2433, N2432, N2431, N2430, N2429, N614, N613, N612, N2425, N2424, N2423, N2422, N2421, N611, N610, N609, N2417, N2416, N2415, N2414, N2413, N608, N607, N606, N2409, N2408, N2407, N2406, N2405, N605, N604, N603, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N602)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[5];
  assign { N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707 } = (N22)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N706)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[6];
  assign { N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772 } = (N23)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N771)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = w_mask_i[7];
  assign { N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837 } = (N24)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N836)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N24 = w_mask_i[8];
  assign { N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902 } = (N25)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N901)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = w_mask_i[9];
  assign { N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973 } = (N26)? { N1498, N1497, N1496, N972, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N971, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N970, N1321, N1320, N1319, N1318, N969, N968, N967, N2433, N2432, N2431, N2430, N2429, N1313, N1312, N1311, N2425, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N2417, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N2409, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N966)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = w_mask_i[10];
  assign { N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038 } = (N27)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1037)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = w_mask_i[11];
  assign { N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103 } = (N28)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1102)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N28 = w_mask_i[12];
  assign { N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168 } = (N29)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1167)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = w_mask_i[13];
  assign { N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233 } = (N30)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1232)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = w_mask_i[14];
  assign { N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330 } = (N31)? { N1498, N1497, N1496, N1495, N1329, N1328, N1327, N1326, N1490, N1489, N1488, N1487, N1325, N1324, N1323, N1322, N1482, N1481, N1480, N1479, N1321, N1320, N1319, N1318, N1474, N1473, N1472, N2313, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N2424, N2423, N2422, N2421, N1309, N1308, N1307, N1306, N2416, N2415, N2414, N2413, N1305, N1304, N1303, N1302, N2408, N2407, N2406, N2405, N1301, N1300, N1299, N1298, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1297)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = w_mask_i[15];
  assign { N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395 } = (N32)? { N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N2313, N2312, N2311, N2310, N2309, N1471, N1470, N1469, N2305, N2304, N2303, N2302, N2301, N1468, N1467, N1466, N2297, N2296, N2295, N2294, N2293, N1465, N1464, N1463, N2289, N2288, N2287, N2286, N2285, N1462, N1461, N1460, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1394)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = w_mask_i[16];
  assign { N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499 } = (N33)? { N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N2313, N2312, N2311, N2310, N2309, N1471, N1470, N1469, N2305, N2304, N2303, N2302, N2301, N1468, N1467, N1466, N2297, N2296, N2295, N2294, N2293, N1465, N1464, N1463, N2289, N2288, N2287, N2286, N2285, N1462, N1461, N1460, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = w_mask_i[17];
  assign { N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564 } = (N34)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1563)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = w_mask_i[18];
  assign { N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629 } = (N35)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1628)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = w_mask_i[19];
  assign { N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694 } = (N36)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1693)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = w_mask_i[20];
  assign { N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759 } = (N37)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1758)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N37 = w_mask_i[21];
  assign { N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824 } = (N38)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1823)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N38 = w_mask_i[22];
  assign { N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889 } = (N39)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1888)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N39 = w_mask_i[23];
  assign { N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954 } = (N40)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1953)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = w_mask_i[24];
  assign { N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019 } = (N41)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2018)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = w_mask_i[25];
  assign { N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092 } = (N42)? { N2460, N2459, N2458, N2211, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2206, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2201, N2320, N2319, N2318, N2317, N2196, N2195, N2194, N2193, N2091, N2090, N2089, N2088, N2308, N2307, N2306, N2087, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2086, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2085, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2084, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2083)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = w_mask_i[26];
  assign { N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212 } = (N43)? { N2460, N2459, N2458, N2211, N2210, N2209, N2208, N2207, N2452, N2451, N2450, N2206, N2205, N2204, N2203, N2202, N2444, N2443, N2442, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2156)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N43 = w_mask_i[27];
  assign { N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332 } = (N44)? { N2460, N2459, N2458, N2331, N2330, N2329, N2328, N2327, N2452, N2451, N2450, N2326, N2325, N2324, N2323, N2322, N2444, N2443, N2442, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2276)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = w_mask_i[28];
  assign { N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461 } = (N45)? { N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2396)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = w_mask_i[29];
  assign { N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526 } = (N46)? { N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N6285, N3234, N3233, N3232, N3231, N2602, N2601, N2600, N3227, N4339, N4338, N4337, N4336, N2599, N2598, N2597, N3223, N4331, N4330, N4329, N4328, N2596, N2595, N2594, N3219, N4323, N4322, N4321, N4320, N2593, N2592, N2591, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2525)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N46 = w_mask_i[30];
  assign { N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630 } = (N47)? { N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N6285, N3234, N3233, N3232, N3231, N2602, N2601, N2600, N3227, N4339, N4338, N4337, N4336, N2599, N2598, N2597, N3223, N4331, N4330, N4329, N4328, N2596, N2595, N2594, N3219, N4323, N4322, N4321, N4320, N2593, N2592, N2591, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2590)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N47 = w_mask_i[31];
  assign { N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695 } = (N48)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2694)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = w_mask_i[32];
  assign { N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760 } = (N49)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2759)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N49 = w_mask_i[33];
  assign { N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825 } = (N50)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2824)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = w_mask_i[34];
  assign { N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890 } = (N51)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2889)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N51 = w_mask_i[35];
  assign { N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955 } = (N52)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2954)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = w_mask_i[36];
  assign { N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020 } = (N53)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3019)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N53 = w_mask_i[37];
  assign { N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085 } = (N54)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3084)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N54 = w_mask_i[38];
  assign { N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150 } = (N55)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3149)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N55 = w_mask_i[39];
  assign { N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253 } = (N56)? { N3486, N3485, N3484, N3252, N3251, N3250, N3249, N3248, N3478, N3477, N3476, N3247, N3246, N3245, N3244, N3243, N3470, N3469, N3468, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N6285, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N4339, N4338, N4337, N4336, N3226, N3225, N3224, N3223, N4331, N4330, N4329, N4328, N3222, N3221, N3220, N3219, N4323, N4322, N4321, N4320, N3218, N3217, N3216, N3215, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3214)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = w_mask_i[40];
  assign { N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318 } = (N57)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N6165, N4014, N4013, N4012, N4011, N3459, N3458, N3457, N4010, N4226, N4225, N4224, N4223, N3456, N3455, N3454, N4009, N4218, N4217, N4216, N4215, N3453, N3452, N3451, N4008, N4210, N4209, N4208, N4207, N3450, N3449, N3448, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3317)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N57 = w_mask_i[41];
  assign { N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383 } = (N58)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N6165, N4014, N4013, N4012, N4011, N3459, N3458, N3457, N4010, N4226, N4225, N4224, N4223, N3456, N3455, N3454, N4009, N4218, N4217, N4216, N4215, N3453, N3452, N3451, N4008, N4210, N4209, N4208, N4207, N3450, N3449, N3448, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3382)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N58 = w_mask_i[42];
  assign { N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487 } = (N59)? { N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N6165, N4014, N4013, N4012, N4011, N3459, N3458, N3457, N4010, N4226, N4225, N4224, N4223, N3456, N3455, N3454, N4009, N4218, N4217, N4216, N4215, N3453, N3452, N3451, N4008, N4210, N4209, N4208, N4207, N3450, N3449, N3448, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3447)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N59 = w_mask_i[43];
  assign { N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552 } = (N60)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3551)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = w_mask_i[44];
  assign { N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617 } = (N61)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3616)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N61 = w_mask_i[45];
  assign { N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682 } = (N62)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3681)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N62 = w_mask_i[46];
  assign { N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747 } = (N63)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3746)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N63 = w_mask_i[47];
  assign { N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812 } = (N64)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3811)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N64 = w_mask_i[48];
  assign { N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877 } = (N65)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3876)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N65 = w_mask_i[49];
  assign { N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942 } = (N66)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3941)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N66 = w_mask_i[50];
  assign { N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, N4072, N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021 } = (N67)? { N4463, N4462, N4461, N4020, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4019, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4018, N4238, N4237, N4236, N4235, N4017, N4016, N4015, N6165, N4014, N4013, N4012, N4011, N4230, N4229, N4228, N4010, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4009, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4008, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4007, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4006)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N67 = w_mask_i[51];
  assign { N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134 } = (N68)? { N4463, N4462, N4461, N4460, N4133, N4132, N4131, N4130, N4455, N4454, N4453, N4452, N4129, N4128, N4127, N4126, N4447, N4446, N4445, N4444, N4125, N4124, N4123, N4122, N4439, N4438, N4437, N6045, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4085)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N68 = w_mask_i[52];
  assign { N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247 } = (N69)? { N4463, N4462, N4461, N4460, N4246, N4245, N4244, N4243, N4455, N4454, N4453, N4452, N4242, N4241, N4240, N4239, N4447, N4446, N4445, N4444, N4238, N4237, N4236, N4235, N4439, N4438, N4437, N6045, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4198)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N69 = w_mask_i[53];
  assign { N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360 } = (N70)? { N4463, N4462, N4461, N4460, N4359, N4358, N4357, N4356, N4455, N4454, N4453, N4452, N4355, N4354, N4353, N4352, N4447, N4446, N4445, N4444, N4351, N4350, N4349, N4348, N4439, N4438, N4437, N6045, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4311)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = w_mask_i[54];
  assign { N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464 } = (N71)? { N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N6045, N4926, N4925, N4924, N4923, N4436, N4435, N4434, N4922, N6276, N6275, N6274, N6273, N4433, N4432, N4431, N4921, N6268, N6267, N6266, N6265, N4430, N4429, N4428, N4920, N6260, N6259, N6258, N6257, N4427, N4426, N4425, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4424)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N71 = w_mask_i[55];
  assign { N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529 } = (N72)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4528)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N72 = w_mask_i[56];
  assign { N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594 } = (N73)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4593)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N73 = w_mask_i[57];
  assign { N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659 } = (N74)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4658)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N74 = w_mask_i[58];
  assign { N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724 } = (N75)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4723)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N75 = w_mask_i[59];
  assign { N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789 } = (N76)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4788)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N76 = w_mask_i[60];
  assign { N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854 } = (N77)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4853)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N77 = w_mask_i[61];
  assign { N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933 } = (N78)? { N5328, N5327, N5326, N4932, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N4931, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N4930, N5151, N5150, N5149, N5148, N4929, N4928, N4927, N6045, N4926, N4925, N4924, N4923, N5143, N5142, N5141, N4922, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N4921, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N4920, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N4919, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4918)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N78 = w_mask_i[62];
  assign { N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998 } = (N79)? { N5328, N5327, N5326, N5325, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N5317, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N5309, N5151, N5150, N5149, N5148, N5304, N5303, N5302, N5937, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N5136, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N5132, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N5128, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4997)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N79 = w_mask_i[63];
  assign { N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063 } = (N80)? { N5328, N5327, N5326, N5325, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N5317, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N5309, N5151, N5150, N5149, N5148, N5304, N5303, N5302, N5937, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N5136, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N5132, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N5128, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5062)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N80 = w_mask_i[64];
  assign { N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160 } = (N81)? { N5328, N5327, N5326, N5325, N5159, N5158, N5157, N5156, N5320, N5319, N5318, N5317, N5155, N5154, N5153, N5152, N5312, N5311, N5310, N5309, N5151, N5150, N5149, N5148, N5304, N5303, N5302, N5937, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N6276, N6275, N6274, N6273, N5139, N5138, N5137, N5136, N6268, N6267, N6266, N6265, N5135, N5134, N5133, N5132, N6260, N6259, N6258, N6257, N5131, N5130, N5129, N5128, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5127)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N81 = w_mask_i[65];
  assign { N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225 } = (N82)? { N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5937, N5936, N5935, N5934, N5933, N5301, N5300, N5299, N5932, N6156, N6155, N6154, N6153, N5298, N5297, N5296, N5931, N6148, N6147, N6146, N6145, N5295, N5294, N5293, N5930, N6140, N6139, N6138, N6137, N5292, N5291, N5290, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5224)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N82 = w_mask_i[66];
  assign { N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329 } = (N83)? { N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5937, N5936, N5935, N5934, N5933, N5301, N5300, N5299, N5932, N6156, N6155, N6154, N6153, N5298, N5297, N5296, N5931, N6148, N6147, N6146, N6145, N5295, N5294, N5293, N5930, N6140, N6139, N6138, N6137, N5292, N5291, N5290, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5289)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N83 = w_mask_i[67];
  assign { N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394 } = (N84)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5393)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N84 = w_mask_i[68];
  assign { N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459 } = (N85)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5458)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N85 = w_mask_i[69];
  assign { N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562, N5561, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524 } = (N86)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5523)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N86 = w_mask_i[70];
  assign { N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, N5626, N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589 } = (N87)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5588)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N87 = w_mask_i[71];
  assign { N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654 } = (N88)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5653)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N88 = w_mask_i[72];
  assign { N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719 } = (N89)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5718)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N89 = w_mask_i[73];
  assign { N5847, N5846, N5845, N5844, N5843, N5842, N5841, N5840, N5839, N5838, N5837, N5836, N5835, N5834, N5833, N5832, N5831, N5830, N5829, N5828, N5827, N5826, N5825, N5824, N5823, N5822, N5821, N5820, N5819, N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784 } = (N90)? { N6312, N6311, N6310, N5863, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5862, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5861, N6172, N6171, N6170, N6169, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N6160, N6159, N6158, N5852, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5851, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5850, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5849, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5783)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N90 = w_mask_i[74];
  assign { N5927, N5926, N5925, N5924, N5923, N5922, N5921, N5920, N5919, N5918, N5917, N5916, N5915, N5914, N5913, N5912, N5911, N5910, N5909, N5908, N5907, N5906, N5905, N5904, N5903, N5902, N5901, N5900, N5899, N5898, N5897, N5896, N5895, N5894, N5893, N5892, N5891, N5890, N5889, N5888, N5887, N5886, N5885, N5884, N5883, N5882, N5881, N5880, N5879, N5878, N5877, N5876, N5875, N5874, N5873, N5872, N5871, N5870, N5869, N5868, N5867, N5866, N5865, N5864 } = (N91)? { N6312, N6311, N6310, N5863, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5862, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5861, N6172, N6171, N6170, N6169, N5860, N5859, N5858, N5857, N5856, N5855, N5854, N5853, N6160, N6159, N6158, N5852, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5851, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5850, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5849, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5848)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N91 = w_mask_i[75];
  assign { N6007, N6006, N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998, N5997, N5996, N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, N5986, N5985, N5984, N5983, N5982, N5981, N5980, N5979, N5978, N5977, N5976, N5975, N5974, N5973, N5972, N5971, N5970, N5969, N5968, N5967, N5966, N5965, N5964, N5963, N5962, N5961, N5960, N5959, N5958, N5957, N5956, N5955, N5954, N5953, N5952, N5951, N5950, N5949, N5948, N5947, N5946, N5945, N5944 } = (N92)? { N6312, N6311, N6310, N5943, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N5942, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N5941, N6172, N6171, N6170, N6169, N5940, N5939, N5938, N5937, N5936, N5935, N5934, N5933, N6160, N6159, N6158, N5932, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N5931, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N5930, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N5929, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N5928)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N92 = w_mask_i[76];
  assign { N6127, N6126, N6125, N6124, N6123, N6122, N6121, N6120, N6119, N6118, N6117, N6116, N6115, N6114, N6113, N6112, N6111, N6110, N6109, N6108, N6107, N6106, N6105, N6104, N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, N6093, N6092, N6091, N6090, N6089, N6088, N6087, N6086, N6085, N6084, N6083, N6082, N6081, N6080, N6079, N6078, N6077, N6076, N6075, N6074, N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064 } = (N93)? { N6312, N6311, N6310, N6063, N6062, N6061, N6060, N6059, N6304, N6303, N6302, N6058, N6057, N6056, N6055, N6054, N6296, N6295, N6294, N6053, N6052, N6051, N6050, N6049, N6048, N6047, N6046, N6045, N6044, N6043, N6042, N6041, N6040, N6039, N6038, N6037, N6036, N6035, N6034, N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025, N6024, N6023, N6022, N6021, N6020, N6019, N6018, N6017, N6016, N6015, N6014, N6013, N6012, N6011, N6010, N6009 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6008)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N93 = w_mask_i[77];
  assign { N6247, N6246, N6245, N6244, N6243, N6242, N6241, N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, N6231, N6230, N6229, N6228, N6227, N6226, N6225, N6224, N6223, N6222, N6221, N6220, N6219, N6218, N6217, N6216, N6215, N6214, N6213, N6212, N6211, N6210, N6209, N6208, N6207, N6206, N6205, N6204, N6203, N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184 } = (N94)? { N6312, N6311, N6310, N6183, N6182, N6181, N6180, N6179, N6304, N6303, N6302, N6178, N6177, N6176, N6175, N6174, N6296, N6295, N6294, N6173, N6172, N6171, N6170, N6169, N6168, N6167, N6166, N6165, N6164, N6163, N6162, N6161, N6160, N6159, N6158, N6157, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N6149, N6148, N6147, N6146, N6145, N6144, N6143, N6142, N6141, N6140, N6139, N6138, N6137, N6136, N6135, N6134, N6133, N6132, N6131, N6130, N6129 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6128)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N94 = w_mask_i[78];
  assign { N6376, N6375, N6374, N6373, N6372, N6371, N6370, N6369, N6368, N6367, N6366, N6365, N6364, N6363, N6362, N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, N6351, N6350, N6349, N6348, N6347, N6346, N6345, N6344, N6343, N6342, N6341, N6340, N6339, N6338, N6337, N6336, N6335, N6334, N6333, N6332, N6331, N6330, N6329, N6328, N6327, N6326, N6325, N6324, N6323, N6322, N6321, N6320, N6319, N6318, N6317, N6316, N6315, N6314, N6313 } = (N95)? { N6312, N6311, N6310, N6309, N6308, N6307, N6306, N6305, N6304, N6303, N6302, N6301, N6300, N6299, N6298, N6297, N6296, N6295, N6294, N6293, N6292, N6291, N6290, N6289, N6288, N6287, N6286, N6285, N6284, N6283, N6282, N6281, N6280, N6279, N6278, N6277, N6276, N6275, N6274, N6273, N6272, N6271, N6270, N6269, N6268, N6267, N6266, N6265, N6264, N6263, N6262, N6261, N6260, N6259, N6258, N6257, N6256, N6255, N6254, N6253, N6252, N6251, N6250, N6249 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N6248)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N95 = w_mask_i[79];
  assign { N11496, N11495, N11494, N11493, N11492, N11491, N11490, N11489, N11488, N11487, N11486, N11485, N11484, N11483, N11482, N11481, N11480, N11479, N11478, N11477, N11476, N11475, N11474, N11473, N11472, N11471, N11470, N11469, N11468, N11467, N11466, N11465, N11464, N11463, N11462, N11461, N11460, N11459, N11458, N11457, N11456, N11455, N11454, N11453, N11452, N11451, N11450, N11449, N11448, N11447, N11446, N11445, N11444, N11443, N11442, N11441, N11440, N11439, N11438, N11437, N11436, N11435, N11434, N11433, N11432, N11431, N11430, N11429, N11428, N11427, N11426, N11425, N11424, N11423, N11422, N11421, N11420, N11419, N11418, N11417, N11416, N11415, N11414, N11413, N11412, N11411, N11410, N11409, N11408, N11407, N11406, N11405, N11404, N11403, N11402, N11401, N11400, N11399, N11398, N11397, N11396, N11395, N11394, N11393, N11392, N11391, N11390, N11389, N11388, N11387, N11386, N11385, N11384, N11383, N11382, N11381, N11380, N11379, N11378, N11377, N11376, N11375, N11374, N11373, N11372, N11371, N11370, N11369, N11368, N11367, N11366, N11365, N11364, N11363, N11362, N11361, N11360, N11359, N11358, N11357, N11356, N11355, N11354, N11353, N11352, N11351, N11350, N11349, N11348, N11347, N11346, N11345, N11344, N11343, N11342, N11341, N11340, N11339, N11338, N11337, N11336, N11335, N11334, N11333, N11332, N11331, N11330, N11329, N11328, N11327, N11326, N11325, N11324, N11323, N11322, N11321, N11320, N11319, N11318, N11317, N11316, N11315, N11314, N11313, N11312, N11311, N11310, N11309, N11308, N11307, N11306, N11305, N11304, N11303, N11302, N11301, N11300, N11299, N11298, N11297, N11296, N11295, N11294, N11293, N11292, N11291, N11290, N11289, N11288, N11287, N11286, N11285, N11284, N11283, N11282, N11281, N11280, N11279, N11278, N11277, N11276, N11275, N11274, N11273, N11272, N11271, N11270, N11269, N11268, N11267, N11266, N11265, N11264, N11263, N11262, N11261, N11260, N11259, N11258, N11257, N11256, N11255, N11254, N11253, N11252, N11251, N11250, N11249, N11248, N11247, N11246, N11245, N11244, N11243, N11242, N11241, N11240, N11239, N11238, N11237, N11236, N11235, N11234, N11233, N11232, N11231, N11230, N11229, N11228, N11227, N11226, N11225, N11224, N11223, N11222, N11221, N11220, N11219, N11218, N11217, N11216, N11215, N11214, N11213, N11212, N11211, N11210, N11209, N11208, N11207, N11206, N11205, N11204, N11203, N11202, N11201, N11200, N11199, N11198, N11197, N11196, N11195, N11194, N11193, N11192, N11191, N11190, N11189, N11188, N11187, N11186, N11185, N11184, N11183, N11182, N11181, N11180, N11179, N11178, N11177, N11176, N11175, N11174, N11173, N11172, N11171, N11170, N11169, N11168, N11167, N11166, N11165, N11164, N11163, N11162, N11161, N11160, N11159, N11158, N11157, N11156, N11155, N11154, N11153, N11152, N11151, N11150, N11149, N11148, N11147, N11146, N11145, N11144, N11143, N11142, N11141, N11140, N11139, N11138, N11137, N11136, N11135, N11134, N11133, N11132, N11131, N11130, N11129, N11128, N11127, N11126, N11125, N11124, N11123, N11122, N11121, N11120, N11119, N11118, N11117, N11116, N11115, N11114, N11113, N11112, N11111, N11110, N11109, N11108, N11107, N11106, N11105, N11104, N11103, N11102, N11101, N11100, N11099, N11098, N11097, N11096, N11095, N11094, N11093, N11092, N11091, N11090, N11089, N11088, N11087, N11086, N11085, N11084, N11083, N11082, N11081, N11080, N11079, N11078, N11077, N11076, N11075, N11074, N11073, N11072, N11071, N11070, N11069, N11068, N11067, N11066, N11065, N11064, N11063, N11062, N11061, N11060, N11059, N11058, N11057, N11056, N11055, N11054, N11053, N11052, N11051, N11050, N11049, N11048, N11047, N11046, N11045, N11044, N11043, N11042, N11041, N11040, N11039, N11038, N11037, N11036, N11035, N11034, N11033, N11032, N11031, N11030, N11029, N11028, N11027, N11026, N11025, N11024, N11023, N11022, N11021, N11020, N11019, N11018, N11017, N11016, N11015, N11014, N11013, N11012, N11011, N11010, N11009, N11008, N11007, N11006, N11005, N11004, N11003, N11002, N11001, N11000, N10999, N10998, N10997, N10996, N10995, N10994, N10993, N10992, N10991, N10990, N10989, N10988, N10987, N10986, N10985, N10984, N10983, N10982, N10981, N10980, N10979, N10978, N10977, N10976, N10975, N10974, N10973, N10972, N10971, N10970, N10969, N10968, N10967, N10966, N10965, N10964, N10963, N10962, N10961, N10960, N10959, N10958, N10957, N10956, N10955, N10954, N10953, N10952, N10951, N10950, N10949, N10948, N10947, N10946, N10945, N10944, N10943, N10942, N10941, N10940, N10939, N10938, N10937, N10936, N10935, N10934, N10933, N10932, N10931, N10930, N10929, N10928, N10927, N10926, N10925, N10924, N10923, N10922, N10921, N10920, N10919, N10918, N10917, N10916, N10915, N10914, N10913, N10912, N10911, N10910, N10909, N10908, N10907, N10906, N10905, N10904, N10903, N10902, N10901, N10900, N10899, N10898, N10897, N10896, N10895, N10894, N10893, N10892, N10891, N10890, N10889, N10888, N10887, N10886, N10885, N10884, N10883, N10882, N10881, N10880, N10879, N10878, N10877, N10876, N10875, N10874, N10873, N10872, N10871, N10870, N10869, N10868, N10867, N10866, N10865, N10864, N10863, N10862, N10861, N10860, N10859, N10858, N10857, N10856, N10855, N10854, N10853, N10852, N10851, N10850, N10849, N10848, N10847, N10846, N10845, N10844, N10843, N10842, N10841, N10840, N10839, N10838, N10837, N10836, N10835, N10834, N10833, N10832, N10831, N10830, N10829, N10828, N10827, N10826, N10825, N10824, N10823, N10822, N10821, N10820, N10819, N10818, N10817, N10816, N10815, N10814, N10813, N10812, N10811, N10810, N10809, N10808, N10807, N10806, N10805, N10804, N10803, N10802, N10801, N10800, N10799, N10798, N10797, N10796, N10795, N10794, N10793, N10792, N10791, N10790, N10789, N10788, N10787, N10786, N10785, N10784, N10783, N10782, N10781, N10780, N10779, N10778, N10777, N10776, N10775, N10774, N10773, N10772, N10771, N10770, N10769, N10768, N10767, N10766, N10765, N10764, N10763, N10762, N10761, N10760, N10759, N10758, N10757, N10756, N10755, N10754, N10753, N10752, N10751, N10750, N10749, N10748, N10747, N10746, N10745, N10744, N10743, N10742, N10741, N10740, N10739, N10738, N10737, N10736, N10735, N10734, N10733, N10732, N10731, N10730, N10729, N10728, N10727, N10726, N10725, N10724, N10723, N10722, N10721, N10720, N10719, N10718, N10717, N10716, N10715, N10714, N10713, N10712, N10711, N10710, N10709, N10708, N10707, N10706, N10705, N10704, N10703, N10702, N10701, N10700, N10699, N10698, N10697, N10696, N10695, N10694, N10693, N10692, N10691, N10690, N10689, N10688, N10687, N10686, N10685, N10684, N10683, N10682, N10681, N10680, N10679, N10678, N10677, N10676, N10675, N10674, N10673, N10672, N10671, N10670, N10669, N10668, N10667, N10666, N10665, N10664, N10663, N10662, N10661, N10660, N10659, N10658, N10657, N10656, N10655, N10654, N10653, N10652, N10651, N10650, N10649, N10648, N10647, N10646, N10645, N10644, N10643, N10642, N10641, N10640, N10639, N10638, N10637, N10636, N10635, N10634, N10633, N10632, N10631, N10630, N10629, N10628, N10627, N10626, N10625, N10624, N10623, N10622, N10621, N10620, N10619, N10618, N10617, N10616, N10615, N10614, N10613, N10612, N10611, N10610, N10609, N10608, N10607, N10606, N10605, N10604, N10603, N10602, N10601, N10600, N10599, N10598, N10597, N10596, N10595, N10594, N10593, N10592, N10591, N10590, N10589, N10588, N10587, N10586, N10585, N10584, N10583, N10582, N10581, N10580, N10579, N10578, N10577, N10576, N10575, N10574, N10573, N10572, N10571, N10570, N10569, N10568, N10567, N10566, N10565, N10564, N10563, N10562, N10561, N10560, N10559, N10558, N10557, N10556, N10555, N10554, N10553, N10552, N10551, N10550, N10549, N10548, N10547, N10546, N10545, N10544, N10543, N10542, N10541, N10540, N10539, N10538, N10537, N10536, N10535, N10534, N10533, N10532, N10531, N10530, N10529, N10528, N10527, N10526, N10525, N10524, N10523, N10522, N10521, N10520, N10519, N10518, N10517, N10516, N10515, N10514, N10513, N10512, N10511, N10510, N10509, N10508, N10507, N10506, N10505, N10504, N10503, N10502, N10501, N10500, N10499, N10498, N10497, N10496, N10495, N10494, N10493, N10492, N10491, N10490, N10489, N10488, N10487, N10486, N10485, N10484, N10483, N10482, N10481, N10480, N10479, N10478, N10477, N10476, N10475, N10474, N10473, N10472, N10471, N10470, N10469, N10468, N10467, N10466, N10465, N10464, N10463, N10462, N10461, N10460, N10459, N10458, N10457, N10456, N10455, N10454, N10453, N10452, N10451, N10450, N10449, N10448, N10447, N10446, N10445, N10444, N10443, N10442, N10441, N10440, N10439, N10438, N10437, N10436, N10435, N10434, N10433, N10432, N10431, N10430, N10429, N10428, N10427, N10426, N10425, N10424, N10423, N10422, N10421, N10420, N10419, N10418, N10417, N10416, N10415, N10414, N10413, N10412, N10411, N10410, N10409, N10408, N10407, N10406, N10405, N10404, N10403, N10402, N10401, N10400, N10399, N10398, N10397, N10396, N10395, N10394, N10393, N10392, N10391, N10390, N10389, N10388, N10387, N10386, N10385, N10384, N10383, N10382, N10381, N10380, N10379, N10378, N10377, N10376, N10375, N10374, N10373, N10372, N10371, N10370, N10369, N10368, N10367, N10366, N10365, N10364, N10363, N10362, N10361, N10360, N10359, N10358, N10357, N10356, N10355, N10354, N10353, N10352, N10351, N10350, N10349, N10348, N10347, N10346, N10345, N10344, N10343, N10342, N10341, N10340, N10339, N10338, N10337, N10336, N10335, N10334, N10333, N10332, N10331, N10330, N10329, N10328, N10327, N10326, N10325, N10324, N10323, N10322, N10321, N10320, N10319, N10318, N10317, N10316, N10315, N10314, N10313, N10312, N10311, N10310, N10309, N10308, N10307, N10306, N10305, N10304, N10303, N10302, N10301, N10300, N10299, N10298, N10297, N10296, N10295, N10294, N10293, N10292, N10291, N10290, N10289, N10288, N10287, N10286, N10285, N10284, N10283, N10282, N10281, N10280, N10279, N10278, N10277, N10276, N10275, N10274, N10273, N10272, N10271, N10270, N10269, N10268, N10267, N10266, N10265, N10264, N10263, N10262, N10261, N10260, N10259, N10258, N10257, N10256, N10255, N10254, N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742, N9741, N9740, N9739, N9738, N9737, N9736, N9735, N9734, N9733, N9732, N9731, N9730, N9729, N9728, N9727, N9726, N9725, N9724, N9723, N9722, N9721, N9720, N9719, N9718, N9717, N9716, N9715, N9714, N9713, N9712, N9711, N9710, N9709, N9708, N9707, N9706, N9705, N9704, N9703, N9702, N9701, N9700, N9699, N9698, N9697, N9696, N9695, N9694, N9693, N9692, N9691, N9690, N9689, N9688, N9687, N9686, N9685, N9684, N9683, N9682, N9681, N9680, N9679, N9678, N9677, N9676, N9675, N9674, N9673, N9672, N9671, N9670, N9669, N9668, N9667, N9666, N9665, N9664, N9663, N9662, N9661, N9660, N9659, N9658, N9657, N9656, N9655, N9654, N9653, N9652, N9651, N9650, N9649, N9648, N9647, N9646, N9645, N9644, N9643, N9642, N9641, N9640, N9639, N9638, N9637, N9636, N9635, N9634, N9633, N9632, N9631, N9630, N9629, N9628, N9627, N9626, N9625, N9624, N9623, N9622, N9621, N9620, N9619, N9618, N9617, N9616, N9615, N9614, N9613, N9612, N9611, N9610, N9609, N9608, N9607, N9606, N9605, N9604, N9603, N9602, N9601, N9600, N9599, N9598, N9597, N9596, N9595, N9594, N9593, N9592, N9591, N9590, N9589, N9588, N9587, N9586, N9585, N9584, N9583, N9582, N9581, N9580, N9579, N9578, N9577, N9576, N9575, N9574, N9573, N9572, N9571, N9570, N9569, N9568, N9567, N9566, N9565, N9564, N9563, N9562, N9561, N9560, N9559, N9558, N9557, N9556, N9555, N9554, N9553, N9552, N9551, N9550, N9549, N9548, N9547, N9546, N9545, N9544, N9543, N9542, N9541, N9540, N9539, N9538, N9537, N9536, N9535, N9534, N9533, N9532, N9531, N9530, N9529, N9528, N9527, N9526, N9525, N9524, N9523, N9522, N9521, N9520, N9519, N9518, N9517, N9516, N9515, N9514, N9513, N9512, N9511, N9510, N9509, N9508, N9507, N9506, N9505, N9504, N9503, N9502, N9501, N9500, N9499, N9498, N9497, N9496, N9495, N9494, N9493, N9492, N9491, N9490, N9489, N9488, N9487, N9486, N9485, N9484, N9483, N9482, N9481, N9480, N9479, N9478, N9477, N9476, N9475, N9474, N9473, N9472, N9471, N9470, N9469, N9468, N9467, N9466, N9465, N9464, N9463, N9462, N9461, N9460, N9459, N9458, N9457, N9456, N9455, N9454, N9453, N9452, N9451, N9450, N9449, N9448, N9447, N9446, N9445, N9444, N9443, N9442, N9441, N9440, N9439, N9438, N9437, N9436, N9435, N9434, N9433, N9432, N9431, N9430, N9429, N9428, N9427, N9426, N9425, N9424, N9423, N9422, N9421, N9420, N9419, N9418, N9417, N9416, N9415, N9414, N9413, N9412, N9411, N9410, N9409, N9408, N9407, N9406, N9405, N9404, N9403, N9402, N9401, N9400, N9399, N9398, N9397, N9396, N9395, N9394, N9393, N9392, N9391, N9390, N9389, N9388, N9387, N9386, N9385, N9384, N9383, N9382, N9381, N9380, N9379, N9378, N9377, N9376, N9375, N9374, N9373, N9372, N9371, N9370, N9369, N9368, N9367, N9366, N9365, N9364, N9363, N9362, N9361, N9360, N9359, N9358, N9357, N9356, N9355, N9354, N9353, N9352, N9351, N9350, N9349, N9348, N9347, N9346, N9345, N9344, N9343, N9342, N9341, N9340, N9339, N9338, N9337, N9336, N9335, N9334, N9333, N9332, N9331, N9330, N9329, N9328, N9327, N9326, N9325, N9324, N9323, N9322, N9321, N9320, N9319, N9318, N9317, N9316, N9315, N9314, N9313, N9312, N9311, N9310, N9309, N9308, N9307, N9306, N9305, N9304, N9303, N9302, N9301, N9300, N9299, N9298, N9297, N9296, N9295, N9294, N9293, N9292, N9291, N9290, N9289, N9288, N9287, N9286, N9285, N9284, N9283, N9282, N9281, N9280, N9279, N9278, N9277, N9276, N9275, N9274, N9273, N9272, N9271, N9270, N9269, N9268, N9267, N9266, N9265, N9264, N9263, N9262, N9261, N9260, N9259, N9258, N9257, N9256, N9255, N9254, N9253, N9252, N9251, N9250, N9249, N9248, N9247, N9246, N9245, N9244, N9243, N9242, N9241, N9240, N9239, N9238, N9237, N9236, N9235, N9234, N9233, N9232, N9231, N9230, N9229, N9228, N9227, N9226, N9225, N9224, N9223, N9222, N9221, N9220, N9219, N9218, N9217, N9216, N9215, N9214, N9213, N9212, N9211, N9210, N9209, N9208, N9207, N9206, N9205, N9204, N9203, N9202, N9201, N9200, N9199, N9198, N9197, N9196, N9195, N9194, N9193, N9192, N9191, N9190, N9189, N9188, N9187, N9186, N9185, N9184, N9183, N9182, N9181, N9180, N9179, N9178, N9177, N9176, N9175, N9174, N9173, N9172, N9171, N9170, N9169, N9168, N9167, N9166, N9165, N9164, N9163, N9162, N9161, N9160, N9159, N9158, N9157, N9156, N9155, N9154, N9153, N9152, N9151, N9150, N9149, N9148, N9147, N9146, N9145, N9144, N9143, N9142, N9141, N9140, N9139, N9138, N9137, N9136, N9135, N9134, N9133, N9132, N9131, N9130, N9129, N9128, N9127, N9126, N9125, N9124, N9123, N9122, N9121, N9120, N9119, N9118, N9117, N9116, N9115, N9114, N9113, N9112, N9111, N9110, N9109, N9108, N9107, N9106, N9105, N9104, N9103, N9102, N9101, N9100, N9099, N9098, N9097, N9096, N9095, N9094, N9093, N9092, N9091, N9090, N9089, N9088, N9087, N9086, N9085, N9084, N9083, N9082, N9081, N9080, N9079, N9078, N9077, N9076, N9075, N9074, N9073, N9072, N9071, N9070, N9069, N9068, N9067, N9066, N9065, N9064, N9063, N9062, N9061, N9060, N9059, N9058, N9057, N9056, N9055, N9054, N9053, N9052, N9051, N9050, N9049, N9048, N9047, N9046, N9045, N9044, N9043, N9042, N9041, N9040, N9039, N9038, N9037, N9036, N9035, N9034, N9033, N9032, N9031, N9030, N9029, N9028, N9027, N9026, N9025, N9024, N9023, N9022, N9021, N9020, N9019, N9018, N9017, N9016, N9015, N9014, N9013, N9012, N9011, N9010, N9009, N9008, N9007, N9006, N9005, N9004, N9003, N9002, N9001, N9000, N8999, N8998, N8997, N8996, N8995, N8994, N8993, N8992, N8991, N8990, N8989, N8988, N8987, N8986, N8985, N8984, N8983, N8982, N8981, N8980, N8979, N8978, N8977, N8976, N8975, N8974, N8973, N8972, N8971, N8970, N8969, N8968, N8967, N8966, N8965, N8964, N8963, N8962, N8961, N8960, N8959, N8958, N8957, N8956, N8955, N8954, N8953, N8952, N8951, N8950, N8949, N8948, N8947, N8946, N8945, N8944, N8943, N8942, N8941, N8940, N8939, N8938, N8937, N8936, N8935, N8934, N8933, N8932, N8931, N8930, N8929, N8928, N8927, N8926, N8925, N8924, N8923, N8922, N8921, N8920, N8919, N8918, N8917, N8916, N8915, N8914, N8913, N8912, N8911, N8910, N8909, N8908, N8907, N8906, N8905, N8904, N8903, N8902, N8901, N8900, N8899, N8898, N8897, N8896, N8895, N8894, N8893, N8892, N8891, N8890, N8889, N8888, N8887, N8886, N8885, N8884, N8883, N8882, N8881, N8880, N8879, N8878, N8877, N8876, N8875, N8874, N8873, N8872, N8871, N8870, N8869, N8868, N8867, N8866, N8865, N8864, N8863, N8862, N8861, N8860, N8859, N8858, N8857, N8856, N8855, N8854, N8853, N8852, N8851, N8850, N8849, N8848, N8847, N8846, N8845, N8844, N8843, N8842, N8841, N8840, N8839, N8838, N8837, N8836, N8835, N8834, N8833, N8832, N8831, N8830, N8829, N8828, N8827, N8826, N8825, N8824, N8823, N8822, N8821, N8820, N8819, N8818, N8817, N8816, N8815, N8814, N8813, N8812, N8811, N8810, N8809, N8808, N8807, N8806, N8805, N8804, N8803, N8802, N8801, N8800, N8799, N8798, N8797, N8796, N8795, N8794, N8793, N8792, N8791, N8790, N8789, N8788, N8787, N8786, N8785, N8784, N8783, N8782, N8781, N8780, N8779, N8778, N8777, N8776, N8775, N8774, N8773, N8772, N8771, N8770, N8769, N8768, N8767, N8766, N8765, N8764, N8763, N8762, N8761, N8760, N8759, N8758, N8757, N8756, N8755, N8754, N8753, N8752, N8751, N8750, N8749, N8748, N8747, N8746, N8745, N8744, N8743, N8742, N8741, N8740, N8739, N8738, N8737, N8736, N8735, N8734, N8733, N8732, N8731, N8730, N8729, N8728, N8727, N8726, N8725, N8724, N8723, N8722, N8721, N8720, N8719, N8718, N8717, N8716, N8715, N8714, N8713, N8712, N8711, N8710, N8709, N8708, N8707, N8706, N8705, N8704, N8703, N8702, N8701, N8700, N8699, N8698, N8697, N8696, N8695, N8694, N8693, N8692, N8691, N8690, N8689, N8688, N8687, N8686, N8685, N8684, N8683, N8682, N8681, N8680, N8679, N8678, N8677, N8676, N8675, N8674, N8673, N8672, N8671, N8670, N8669, N8668, N8667, N8666, N8665, N8664, N8663, N8662, N8661, N8660, N8659, N8658, N8657, N8656, N8655, N8654, N8653, N8652, N8651, N8650, N8649, N8648, N8647, N8646, N8645, N8644, N8643, N8642, N8641, N8640, N8639, N8638, N8637, N8636, N8635, N8634, N8633, N8632, N8631, N8630, N8629, N8628, N8627, N8626, N8625, N8624, N8623, N8622, N8621, N8620, N8619, N8618, N8617, N8616, N8615, N8614, N8613, N8612, N8611, N8610, N8609, N8608, N8607, N8606, N8605, N8604, N8603, N8602, N8601, N8600, N8599, N8598, N8597, N8596, N8595, N8594, N8593, N8592, N8591, N8590, N8589, N8588, N8587, N8586, N8585, N8584, N8583, N8582, N8581, N8580, N8579, N8578, N8577, N8576, N8575, N8574, N8573, N8572, N8571, N8570, N8569, N8568, N8567, N8566, N8565, N8564, N8563, N8562, N8561, N8560, N8559, N8558, N8557, N8556, N8555, N8554, N8553, N8552, N8551, N8550, N8549, N8548, N8547, N8546, N8545, N8544, N8543, N8542, N8541, N8540, N8539, N8538, N8537, N8536, N8535, N8534, N8533, N8532, N8531, N8530, N8529, N8528, N8527, N8526, N8525, N8524, N8523, N8522, N8521, N8520, N8519, N8518, N8517, N8516, N8515, N8514, N8513, N8512, N8511, N8510, N8509, N8508, N8507, N8506, N8505, N8504, N8503, N8502, N8501, N8500, N8499, N8498, N8497, N8496, N8495, N8494, N8493, N8492, N8491, N8490, N8489, N8488, N8487, N8486, N8485, N8484, N8483, N8482, N8481, N8480, N8479, N8478, N8477, N8476, N8475, N8474, N8473, N8472, N8471, N8470, N8469, N8468, N8467, N8466, N8465, N8464, N8463, N8462, N8461, N8460, N8459, N8458, N8457, N8456, N8455, N8454, N8453, N8452, N8451, N8450, N8449, N8448, N8447, N8446, N8445, N8444, N8443, N8442, N8441, N8440, N8439, N8438, N8437, N8436, N8435, N8434, N8433, N8432, N8431, N8430, N8429, N8428, N8427, N8426, N8425, N8424, N8423, N8422, N8421, N8420, N8419, N8418, N8417, N8416, N8415, N8414, N8413, N8412, N8411, N8410, N8409, N8408, N8407, N8406, N8405, N8404, N8403, N8402, N8401, N8400, N8399, N8398, N8397, N8396, N8395, N8394, N8393, N8392, N8391, N8390, N8389, N8388, N8387, N8386, N8385, N8384, N8383, N8382, N8381, N8380, N8379, N8378, N8377, N8376, N8375, N8374, N8373, N8372, N8371, N8370, N8369, N8368, N8367, N8366, N8365, N8364, N8363, N8362, N8361, N8360, N8359, N8358, N8357, N8356, N8355, N8354, N8353, N8352, N8351, N8350, N8349, N8348, N8347, N8346, N8345, N8344, N8343, N8342, N8341, N8340, N8339, N8338, N8337, N8336, N8335, N8334, N8333, N8332, N8331, N8330, N8329, N8328, N8327, N8326, N8325, N8324, N8323, N8322, N8321, N8320, N8319, N8318, N8317, N8316, N8315, N8314, N8313, N8312, N8311, N8310, N8309, N8308, N8307, N8306, N8305, N8304, N8303, N8302, N8301, N8300, N8299, N8298, N8297, N8296, N8295, N8294, N8293, N8292, N8291, N8290, N8289, N8288, N8287, N8286, N8285, N8284, N8283, N8282, N8281, N8280, N8279, N8278, N8277, N8276, N8275, N8274, N8273, N8272, N8271, N8270, N8269, N8268, N8267, N8266, N8265, N8264, N8263, N8262, N8261, N8260, N8259, N8258, N8257, N8256, N8255, N8254, N8253, N8252, N8251, N8250, N8249, N8248, N8247, N8246, N8245, N8244, N8243, N8242, N8241, N8240, N8239, N8238, N8237, N8236, N8235, N8234, N8233, N8232, N8231, N8230, N8229, N8228, N8227, N8226, N8225, N8224, N8223, N8222, N8221, N8220, N8219, N8218, N8217, N8216, N8215, N8214, N8213, N8212, N8211, N8210, N8209, N8208, N8207, N8206, N8205, N8204, N8203, N8202, N8201, N8200, N8199, N8198, N8197, N8196, N8195, N8194, N8193, N8192, N8191, N8190, N8189, N8188, N8187, N8186, N8185, N8184, N8183, N8182, N8181, N8180, N8179, N8178, N8177, N8176, N8175, N8174, N8173, N8172, N8171, N8170, N8169, N8168, N8167, N8166, N8165, N8164, N8163, N8162, N8161, N8160, N8159, N8158, N8157, N8156, N8155, N8154, N8153, N8152, N8151, N8150, N8149, N8148, N8147, N8146, N8145, N8144, N8143, N8142, N8141, N8140, N8139, N8138, N8137, N8136, N8135, N8134, N8133, N8132, N8131, N8130, N8129, N8128, N8127, N8126, N8125, N8124, N8123, N8122, N8121, N8120, N8119, N8118, N8117, N8116, N8115, N8114, N8113, N8112, N8111, N8110, N8109, N8108, N8107, N8106, N8105, N8104, N8103, N8102, N8101, N8100, N8099, N8098, N8097, N8096, N8095, N8094, N8093, N8092, N8091, N8090, N8089, N8088, N8087, N8086, N8085, N8084, N8083, N8082, N8081, N8080, N8079, N8078, N8077, N8076, N8075, N8074, N8073, N8072, N8071, N8070, N8069, N8068, N8067, N8066, N8065, N8064, N8063, N8062, N8061, N8060, N8059, N8058, N8057, N8056, N8055, N8054, N8053, N8052, N8051, N8050, N8049, N8048, N8047, N8046, N8045, N8044, N8043, N8042, N8041, N8040, N8039, N8038, N8037, N8036, N8035, N8034, N8033, N8032, N8031, N8030, N8029, N8028, N8027, N8026, N8025, N8024, N8023, N8022, N8021, N8020, N8019, N8018, N8017, N8016, N8015, N8014, N8013, N8012, N8011, N8010, N8009, N8008, N8007, N8006, N8005, N8004, N8003, N8002, N8001, N8000, N7999, N7998, N7997, N7996, N7995, N7994, N7993, N7992, N7991, N7990, N7989, N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, N7979, N7978, N7977, N7976, N7975, N7974, N7973, N7972, N7971, N7970, N7969, N7968, N7967, N7966, N7965, N7964, N7963, N7962, N7961, N7960, N7959, N7958, N7957, N7956, N7955, N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946, N7945, N7944, N7943, N7942, N7941, N7940, N7939, N7938, N7937, N7936, N7935, N7934, N7933, N7932, N7931, N7930, N7929, N7928, N7927, N7926, N7925, N7924, N7923, N7922, N7921, N7920, N7919, N7918, N7917, N7916, N7915, N7914, N7913, N7912, N7911, N7910, N7909, N7908, N7907, N7906, N7905, N7904, N7903, N7902, N7901, N7900, N7899, N7898, N7897, N7896, N7895, N7894, N7893, N7892, N7891, N7890, N7889, N7888, N7887, N7886, N7885, N7884, N7883, N7882, N7881, N7880, N7879, N7878, N7877, N7876, N7875, N7874, N7873, N7872, N7871, N7870, N7869, N7868, N7867, N7866, N7865, N7864, N7863, N7862, N7861, N7860, N7859, N7858, N7857, N7856, N7855, N7854, N7853, N7852, N7851, N7850, N7849, N7848, N7847, N7846, N7845, N7844, N7843, N7842, N7841, N7840, N7839, N7838, N7837, N7836, N7835, N7834, N7833, N7832, N7831, N7830, N7829, N7828, N7827, N7826, N7825, N7824, N7823, N7822, N7821, N7820, N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, N7809, N7808, N7807, N7806, N7805, N7804, N7803, N7802, N7801, N7800, N7799, N7798, N7797, N7796, N7795, N7794, N7793, N7792, N7791, N7790, N7789, N7788, N7787, N7786, N7785, N7784, N7783, N7782, N7781, N7780, N7779, N7778, N7777, N7776, N7775, N7774, N7773, N7772, N7771, N7770, N7769, N7768, N7767, N7766, N7765, N7764, N7763, N7762, N7761, N7760, N7759, N7758, N7757, N7756, N7755, N7754, N7753, N7752, N7751, N7750, N7749, N7748, N7747, N7746, N7745, N7744, N7743, N7742, N7741, N7740, N7739, N7738, N7737, N7736, N7735, N7734, N7733, N7732, N7731, N7730, N7729, N7728, N7727, N7726, N7725, N7724, N7723, N7722, N7721, N7720, N7719, N7718, N7717, N7716, N7715, N7714, N7713, N7712, N7711, N7710, N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696, N7695, N7694, N7693, N7692, N7691, N7690, N7689, N7688, N7687, N7686, N7685, N7684, N7683, N7682, N7681, N7680, N7679, N7678, N7677, N7676, N7675, N7674, N7673, N7672, N7671, N7670, N7669, N7668, N7667, N7666, N7665, N7664, N7663, N7662, N7661, N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, N7641, N7640, N7639, N7638, N7637, N7636, N7635, N7634, N7633, N7632, N7631, N7630, N7629, N7628, N7627, N7626, N7625, N7624, N7623, N7622, N7621, N7620, N7619, N7618, N7617, N7616, N7615, N7614, N7613, N7612, N7611, N7610, N7609, N7608, N7607, N7606, N7605, N7604, N7603, N7602, N7601, N7600, N7599, N7598, N7597, N7596, N7595, N7594, N7593, N7592, N7591, N7590, N7589, N7588, N7587, N7586, N7585, N7584, N7583, N7582, N7581, N7580, N7579, N7578, N7577, N7576, N7575, N7574, N7573, N7572, N7571, N7570, N7569, N7568, N7567, N7566, N7565, N7564, N7563, N7562, N7561, N7560, N7559, N7558, N7557, N7556, N7555, N7554, N7553, N7552, N7551, N7550, N7549, N7548, N7547, N7546, N7545, N7544, N7543, N7542, N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7533, N7532, N7531, N7530, N7529, N7528, N7527, N7526, N7525, N7524, N7523, N7522, N7521, N7520, N7519, N7518, N7517, N7516, N7515, N7514, N7513, N7512, N7511, N7510, N7509, N7508, N7507, N7506, N7505, N7504, N7503, N7502, N7501, N7500, N7499, N7498, N7497, N7496, N7495, N7494, N7493, N7492, N7491, N7490, N7489, N7488, N7487, N7486, N7485, N7484, N7483, N7482, N7481, N7480, N7479, N7478, N7477, N7476, N7475, N7474, N7473, N7472, N7471, N7470, N7469, N7468, N7467, N7466, N7465, N7464, N7463, N7462, N7461, N7460, N7459, N7458, N7457, N7456, N7455, N7454, N7453, N7452, N7451, N7450, N7449, N7448, N7447, N7446, N7445, N7444, N7443, N7442, N7441, N7440, N7439, N7438, N7437, N7436, N7435, N7434, N7433, N7432, N7431, N7430, N7429, N7428, N7427, N7426, N7425, N7424, N7423, N7422, N7421, N7420, N7419, N7418, N7417, N7416, N7415, N7414, N7413, N7412, N7411, N7410, N7409, N7408, N7407, N7406, N7405, N7404, N7403, N7402, N7401, N7400, N7399, N7398, N7397, N7396, N7395, N7394, N7393, N7392, N7391, N7390, N7389, N7388, N7387, N7386, N7385, N7384, N7383, N7382, N7381, N7380, N7379, N7378, N7377, N7376, N7375, N7374, N7373, N7372, N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360, N7359, N7358, N7357, N7356, N7355, N7354, N7353, N7352, N7351, N7350, N7349, N7348, N7347, N7346, N7345, N7344, N7343, N7342, N7341, N7340, N7339, N7338, N7337, N7336, N7335, N7334, N7333, N7332, N7331, N7330, N7329, N7328, N7327, N7326, N7325, N7324, N7323, N7322, N7321, N7320, N7319, N7318, N7317, N7316, N7315, N7314, N7313, N7312, N7311, N7310, N7309, N7308, N7307, N7306, N7305, N7304, N7303, N7302, N7301, N7300, N7299, N7298, N7297, N7296, N7295, N7294, N7293, N7292, N7291, N7290, N7289, N7288, N7287, N7286, N7285, N7284, N7283, N7282, N7281, N7280, N7279, N7278, N7277, N7276, N7275, N7274, N7273, N7272, N7271, N7270, N7269, N7268, N7267, N7266, N7265, N7264, N7263, N7262, N7261, N7260, N7259, N7258, N7257, N7256, N7255, N7254, N7253, N7252, N7251, N7250, N7249, N7248, N7247, N7246, N7245, N7244, N7243, N7242, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, N7223, N7222, N7221, N7220, N7219, N7218, N7217, N7216, N7215, N7214, N7213, N7212, N7211, N7210, N7209, N7208, N7207, N7206, N7205, N7204, N7203, N7202, N7201, N7200, N7199, N7198, N7197, N7196, N7195, N7194, N7193, N7192, N7191, N7190, N7189, N7188, N7187, N7186, N7185, N7184, N7183, N7182, N7181, N7180, N7179, N7178, N7177, N7176, N7175, N7174, N7173, N7172, N7171, N7170, N7169, N7168, N7167, N7166, N7165, N7164, N7163, N7162, N7161, N7160, N7159, N7158, N7157, N7156, N7155, N7154, N7153, N7152, N7151, N7150, N7149, N7148, N7147, N7146, N7145, N7144, N7143, N7142, N7141, N7140, N7139, N7138, N7137, N7136, N7135, N7134, N7133, N7132, N7131, N7130, N7129, N7128, N7127, N7126, N7125, N7124, N7123, N7122, N7121, N7120, N7119, N7118, N7117, N7116, N7115, N7114, N7113, N7112, N7111, N7110, N7109, N7108, N7107, N7106, N7105, N7104, N7103, N7102, N7101, N7100, N7099, N7098, N7097, N7096, N7095, N7094, N7093, N7092, N7091, N7090, N7089, N7088, N7087, N7086, N7085, N7084, N7083, N7082, N7081, N7080, N7079, N7078, N7077, N7076, N7075, N7074, N7073, N7072, N7071, N7070, N7069, N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, N7049, N7048, N7047, N7046, N7045, N7044, N7043, N7042, N7041, N7040, N7039, N7038, N7037, N7036, N7035, N7034, N7033, N7032, N7031, N7030, N7029, N7028, N7027, N7026, N7025, N7024, N7023, N7022, N7021, N7020, N7019, N7018, N7017, N7016, N7015, N7014, N7013, N7012, N7011, N7010, N7009, N7008, N7007, N7006, N7005, N7004, N7003, N7002, N7001, N7000, N6999, N6998, N6997, N6996, N6995, N6994, N6993, N6992, N6991, N6990, N6989, N6988, N6987, N6986, N6985, N6984, N6983, N6982, N6981, N6980, N6979, N6978, N6977, N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, N6957, N6956, N6955, N6954, N6953, N6952, N6951, N6950, N6949, N6948, N6947, N6946, N6945, N6944, N6943, N6942, N6941, N6940, N6939, N6938, N6937, N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923, N6922, N6921, N6920, N6919, N6918, N6917, N6916, N6915, N6914, N6913, N6912, N6911, N6910, N6909, N6908, N6907, N6906, N6905, N6904, N6903, N6902, N6901, N6900, N6899, N6898, N6897, N6896, N6895, N6894, N6893, N6892, N6891, N6890, N6889, N6888, N6887, N6886, N6885, N6884, N6883, N6882, N6881, N6880, N6879, N6878, N6877, N6876, N6875, N6874, N6873, N6872, N6871, N6870, N6869, N6868, N6867, N6866, N6865, N6864, N6863, N6862, N6861, N6860, N6859, N6858, N6857, N6856, N6855, N6854, N6853, N6852, N6851, N6850, N6849, N6848, N6847, N6846, N6845, N6844, N6843, N6842, N6841, N6840, N6839, N6838, N6837, N6836, N6835, N6834, N6833, N6832, N6831, N6830, N6829, N6828, N6827, N6826, N6825, N6824, N6823, N6822, N6821, N6820, N6819, N6818, N6817, N6816, N6815, N6814, N6813, N6812, N6811, N6810, N6809, N6808, N6807, N6806, N6805, N6804, N6803, N6802, N6801, N6800, N6799, N6798, N6797, N6796, N6795, N6794, N6793, N6792, N6791, N6790, N6789, N6788, N6787, N6786, N6785, N6784, N6783, N6782, N6781, N6780, N6779, N6778, N6777, N6776, N6775, N6774, N6773, N6772, N6771, N6770, N6769, N6768, N6767, N6766, N6765, N6764, N6763, N6762, N6761, N6760, N6759, N6758, N6757, N6756, N6755, N6754, N6753, N6752, N6751, N6750, N6749, N6748, N6747, N6746, N6745, N6744, N6743, N6742, N6741, N6740, N6739, N6738, N6737, N6736, N6735, N6734, N6733, N6732, N6731, N6730, N6729, N6728, N6727, N6726, N6725, N6724, N6723, N6722, N6721, N6720, N6719, N6718, N6717, N6716, N6715, N6714, N6713, N6712, N6711, N6710, N6709, N6708, N6707, N6706, N6705, N6704, N6703, N6702, N6701, N6700, N6699, N6698, N6697, N6696, N6695, N6694, N6693, N6692, N6691, N6690, N6689, N6688, N6687, N6686, N6685, N6684, N6683, N6682, N6681, N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667, N6666, N6665, N6664, N6663, N6662, N6661, N6660, N6659, N6658, N6657, N6656, N6655, N6654, N6653, N6652, N6651, N6650, N6649, N6648, N6647, N6646, N6645, N6644, N6643, N6642, N6641, N6640, N6639, N6638, N6637, N6636, N6635, N6634, N6633, N6632, N6631, N6630, N6629, N6628, N6627, N6626, N6625, N6624, N6623, N6622, N6621, N6620, N6619, N6618, N6617, N6616, N6615, N6614, N6613, N6612, N6611, N6610, N6609, N6608, N6607, N6606, N6605, N6604, N6603, N6602, N6601, N6600, N6599, N6598, N6597, N6596, N6595, N6594, N6593, N6592, N6591, N6590, N6589, N6588, N6587, N6586, N6585, N6584, N6583, N6582, N6581, N6580, N6579, N6578, N6577, N6576, N6575, N6574, N6573, N6572, N6571, N6570, N6569, N6568, N6567, N6566, N6565, N6564, N6563, N6562, N6561, N6560, N6559, N6558, N6557, N6556, N6555, N6554, N6553, N6552, N6551, N6550, N6549, N6548, N6547, N6546, N6545, N6544, N6543, N6542, N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514, N6513, N6512, N6511, N6510, N6509, N6508, N6507, N6506, N6505, N6504, N6503, N6502, N6501, N6500, N6499, N6498, N6497, N6496, N6495, N6494, N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485, N6484, N6483, N6482, N6481, N6480, N6479, N6478, N6477, N6476, N6475, N6474, N6473, N6472, N6471, N6470, N6469, N6468, N6467, N6466, N6465, N6464, N6463, N6462, N6461, N6460, N6459, N6458, N6457, N6456, N6455, N6454, N6453, N6452, N6451, N6450, N6449, N6448, N6447, N6446, N6445, N6444, N6443, N6442, N6441, N6440, N6439, N6438, N6437, N6436, N6435, N6434, N6433, N6432, N6431, N6430, N6429, N6428, N6427, N6426, N6425, N6424, N6423, N6422, N6421, N6420, N6419, N6418, N6417, N6416, N6415, N6414, N6413, N6412, N6411, N6410, N6409, N6408, N6407, N6406, N6405, N6404, N6403, N6402, N6401, N6400, N6399, N6398, N6397, N6396, N6395, N6394, N6393, N6392, N6391, N6390, N6389, N6388, N6387, N6386, N6385, N6384, N6383, N6382, N6381, N6380, N6379, N6378, N6377 } = (N96)? { N6376, N6247, N6127, N6007, N5927, N5847, N5782, N5717, N5652, N5587, N5522, N5457, N5392, N5288, N5223, N5126, N5061, N4996, N4917, N4852, N4787, N4722, N4657, N4592, N4527, N4423, N4310, N4197, N4084, N4005, N3940, N3875, N3810, N3745, N3680, N3615, N3550, N3446, N3381, N3316, N3213, N3148, N3083, N3018, N2953, N2888, N2823, N2758, N2693, N2589, N2524, N2395, N2275, N2155, N2082, N2017, N1952, N1887, N1822, N1757, N1692, N1627, N1562, N1458, N1393, N1296, N1231, N1166, N1101, N1036, N965, N900, N835, N770, N705, N601, N488, N423, N358, N293, N6375, N6246, N6126, N6006, N5926, N5846, N5781, N5716, N5651, N5586, N5521, N5456, N5391, N5287, N5222, N5125, N5060, N4995, N4916, N4851, N4786, N4721, N4656, N4591, N4526, N4422, N4309, N4196, N4083, N4004, N3939, N3874, N3809, N3744, N3679, N3614, N3549, N3445, N3380, N3315, N3212, N3147, N3082, N3017, N2952, N2887, N2822, N2757, N2692, N2588, N2523, N2394, N2274, N2154, N2081, N2016, N1951, N1886, N1821, N1756, N1691, N1626, N1561, N1457, N1392, N1295, N1230, N1165, N1100, N1035, N964, N899, N834, N769, N704, N600, N487, N422, N357, N292, N6374, N6245, N6125, N6005, N5925, N5845, N5780, N5715, N5650, N5585, N5520, N5455, N5390, N5286, N5221, N5124, N5059, N4994, N4915, N4850, N4785, N4720, N4655, N4590, N4525, N4421, N4308, N4195, N4082, N4003, N3938, N3873, N3808, N3743, N3678, N3613, N3548, N3444, N3379, N3314, N3211, N3146, N3081, N3016, N2951, N2886, N2821, N2756, N2691, N2587, N2522, N2393, N2273, N2153, N2080, N2015, N1950, N1885, N1820, N1755, N1690, N1625, N1560, N1456, N1391, N1294, N1229, N1164, N1099, N1034, N963, N898, N833, N768, N703, N599, N486, N421, N356, N291, N6373, N6244, N6124, N6004, N5924, N5844, N5779, N5714, N5649, N5584, N5519, N5454, N5389, N5285, N5220, N5123, N5058, N4993, N4914, N4849, N4784, N4719, N4654, N4589, N4524, N4420, N4307, N4194, N4081, N4002, N3937, N3872, N3807, N3742, N3677, N3612, N3547, N3443, N3378, N3313, N3210, N3145, N3080, N3015, N2950, N2885, N2820, N2755, N2690, N2586, N2521, N2392, N2272, N2152, N2079, N2014, N1949, N1884, N1819, N1754, N1689, N1624, N1559, N1455, N1390, N1293, N1228, N1163, N1098, N1033, N962, N897, N832, N767, N702, N598, N485, N420, N355, N290, N6372, N6243, N6123, N6003, N5923, N5843, N5778, N5713, N5648, N5583, N5518, N5453, N5388, N5284, N5219, N5122, N5057, N4992, N4913, N4848, N4783, N4718, N4653, N4588, N4523, N4419, N4306, N4193, N4080, N4001, N3936, N3871, N3806, N3741, N3676, N3611, N3546, N3442, N3377, N3312, N3209, N3144, N3079, N3014, N2949, N2884, N2819, N2754, N2689, N2585, N2520, N2391, N2271, N2151, N2078, N2013, N1948, N1883, N1818, N1753, N1688, N1623, N1558, N1454, N1389, N1292, N1227, N1162, N1097, N1032, N961, N896, N831, N766, N701, N597, N484, N419, N354, N289, N6371, N6242, N6122, N6002, N5922, N5842, N5777, N5712, N5647, N5582, N5517, N5452, N5387, N5283, N5218, N5121, N5056, N4991, N4912, N4847, N4782, N4717, N4652, N4587, N4522, N4418, N4305, N4192, N4079, N4000, N3935, N3870, N3805, N3740, N3675, N3610, N3545, N3441, N3376, N3311, N3208, N3143, N3078, N3013, N2948, N2883, N2818, N2753, N2688, N2584, N2519, N2390, N2270, N2150, N2077, N2012, N1947, N1882, N1817, N1752, N1687, N1622, N1557, N1453, N1388, N1291, N1226, N1161, N1096, N1031, N960, N895, N830, N765, N700, N596, N483, N418, N353, N288, N6370, N6241, N6121, N6001, N5921, N5841, N5776, N5711, N5646, N5581, N5516, N5451, N5386, N5282, N5217, N5120, N5055, N4990, N4911, N4846, N4781, N4716, N4651, N4586, N4521, N4417, N4304, N4191, N4078, N3999, N3934, N3869, N3804, N3739, N3674, N3609, N3544, N3440, N3375, N3310, N3207, N3142, N3077, N3012, N2947, N2882, N2817, N2752, N2687, N2583, N2518, N2389, N2269, N2149, N2076, N2011, N1946, N1881, N1816, N1751, N1686, N1621, N1556, N1452, N1387, N1290, N1225, N1160, N1095, N1030, N959, N894, N829, N764, N699, N595, N482, N417, N352, N287, N6369, N6240, N6120, N6000, N5920, N5840, N5775, N5710, N5645, N5580, N5515, N5450, N5385, N5281, N5216, N5119, N5054, N4989, N4910, N4845, N4780, N4715, N4650, N4585, N4520, N4416, N4303, N4190, N4077, N3998, N3933, N3868, N3803, N3738, N3673, N3608, N3543, N3439, N3374, N3309, N3206, N3141, N3076, N3011, N2946, N2881, N2816, N2751, N2686, N2582, N2517, N2388, N2268, N2148, N2075, N2010, N1945, N1880, N1815, N1750, N1685, N1620, N1555, N1451, N1386, N1289, N1224, N1159, N1094, N1029, N958, N893, N828, N763, N698, N594, N481, N416, N351, N286, N6368, N6239, N6119, N5999, N5919, N5839, N5774, N5709, N5644, N5579, N5514, N5449, N5384, N5280, N5215, N5118, N5053, N4988, N4909, N4844, N4779, N4714, N4649, N4584, N4519, N4415, N4302, N4189, N4076, N3997, N3932, N3867, N3802, N3737, N3672, N3607, N3542, N3438, N3373, N3308, N3205, N3140, N3075, N3010, N2945, N2880, N2815, N2750, N2685, N2581, N2516, N2387, N2267, N2147, N2074, N2009, N1944, N1879, N1814, N1749, N1684, N1619, N1554, N1450, N1385, N1288, N1223, N1158, N1093, N1028, N957, N892, N827, N762, N697, N593, N480, N415, N350, N285, N6367, N6238, N6118, N5998, N5918, N5838, N5773, N5708, N5643, N5578, N5513, N5448, N5383, N5279, N5214, N5117, N5052, N4987, N4908, N4843, N4778, N4713, N4648, N4583, N4518, N4414, N4301, N4188, N4075, N3996, N3931, N3866, N3801, N3736, N3671, N3606, N3541, N3437, N3372, N3307, N3204, N3139, N3074, N3009, N2944, N2879, N2814, N2749, N2684, N2580, N2515, N2386, N2266, N2146, N2073, N2008, N1943, N1878, N1813, N1748, N1683, N1618, N1553, N1449, N1384, N1287, N1222, N1157, N1092, N1027, N956, N891, N826, N761, N696, N592, N479, N414, N349, N284, N6366, N6237, N6117, N5997, N5917, N5837, N5772, N5707, N5642, N5577, N5512, N5447, N5382, N5278, N5213, N5116, N5051, N4986, N4907, N4842, N4777, N4712, N4647, N4582, N4517, N4413, N4300, N4187, N4074, N3995, N3930, N3865, N3800, N3735, N3670, N3605, N3540, N3436, N3371, N3306, N3203, N3138, N3073, N3008, N2943, N2878, N2813, N2748, N2683, N2579, N2514, N2385, N2265, N2145, N2072, N2007, N1942, N1877, N1812, N1747, N1682, N1617, N1552, N1448, N1383, N1286, N1221, N1156, N1091, N1026, N955, N890, N825, N760, N695, N591, N478, N413, N348, N283, N6365, N6236, N6116, N5996, N5916, N5836, N5771, N5706, N5641, N5576, N5511, N5446, N5381, N5277, N5212, N5115, N5050, N4985, N4906, N4841, N4776, N4711, N4646, N4581, N4516, N4412, N4299, N4186, N4073, N3994, N3929, N3864, N3799, N3734, N3669, N3604, N3539, N3435, N3370, N3305, N3202, N3137, N3072, N3007, N2942, N2877, N2812, N2747, N2682, N2578, N2513, N2384, N2264, N2144, N2071, N2006, N1941, N1876, N1811, N1746, N1681, N1616, N1551, N1447, N1382, N1285, N1220, N1155, N1090, N1025, N954, N889, N824, N759, N694, N590, N477, N412, N347, N282, N6364, N6235, N6115, N5995, N5915, N5835, N5770, N5705, N5640, N5575, N5510, N5445, N5380, N5276, N5211, N5114, N5049, N4984, N4905, N4840, N4775, N4710, N4645, N4580, N4515, N4411, N4298, N4185, N4072, N3993, N3928, N3863, N3798, N3733, N3668, N3603, N3538, N3434, N3369, N3304, N3201, N3136, N3071, N3006, N2941, N2876, N2811, N2746, N2681, N2577, N2512, N2383, N2263, N2143, N2070, N2005, N1940, N1875, N1810, N1745, N1680, N1615, N1550, N1446, N1381, N1284, N1219, N1154, N1089, N1024, N953, N888, N823, N758, N693, N589, N476, N411, N346, N281, N6363, N6234, N6114, N5994, N5914, N5834, N5769, N5704, N5639, N5574, N5509, N5444, N5379, N5275, N5210, N5113, N5048, N4983, N4904, N4839, N4774, N4709, N4644, N4579, N4514, N4410, N4297, N4184, N4071, N3992, N3927, N3862, N3797, N3732, N3667, N3602, N3537, N3433, N3368, N3303, N3200, N3135, N3070, N3005, N2940, N2875, N2810, N2745, N2680, N2576, N2511, N2382, N2262, N2142, N2069, N2004, N1939, N1874, N1809, N1744, N1679, N1614, N1549, N1445, N1380, N1283, N1218, N1153, N1088, N1023, N952, N887, N822, N757, N692, N588, N475, N410, N345, N280, N6362, N6233, N6113, N5993, N5913, N5833, N5768, N5703, N5638, N5573, N5508, N5443, N5378, N5274, N5209, N5112, N5047, N4982, N4903, N4838, N4773, N4708, N4643, N4578, N4513, N4409, N4296, N4183, N4070, N3991, N3926, N3861, N3796, N3731, N3666, N3601, N3536, N3432, N3367, N3302, N3199, N3134, N3069, N3004, N2939, N2874, N2809, N2744, N2679, N2575, N2510, N2381, N2261, N2141, N2068, N2003, N1938, N1873, N1808, N1743, N1678, N1613, N1548, N1444, N1379, N1282, N1217, N1152, N1087, N1022, N951, N886, N821, N756, N691, N587, N474, N409, N344, N279, N6361, N6232, N6112, N5992, N5912, N5832, N5767, N5702, N5637, N5572, N5507, N5442, N5377, N5273, N5208, N5111, N5046, N4981, N4902, N4837, N4772, N4707, N4642, N4577, N4512, N4408, N4295, N4182, N4069, N3990, N3925, N3860, N3795, N3730, N3665, N3600, N3535, N3431, N3366, N3301, N3198, N3133, N3068, N3003, N2938, N2873, N2808, N2743, N2678, N2574, N2509, N2380, N2260, N2140, N2067, N2002, N1937, N1872, N1807, N1742, N1677, N1612, N1547, N1443, N1378, N1281, N1216, N1151, N1086, N1021, N950, N885, N820, N755, N690, N586, N473, N408, N343, N278, N6360, N6231, N6111, N5991, N5911, N5831, N5766, N5701, N5636, N5571, N5506, N5441, N5376, N5272, N5207, N5110, N5045, N4980, N4901, N4836, N4771, N4706, N4641, N4576, N4511, N4407, N4294, N4181, N4068, N3989, N3924, N3859, N3794, N3729, N3664, N3599, N3534, N3430, N3365, N3300, N3197, N3132, N3067, N3002, N2937, N2872, N2807, N2742, N2677, N2573, N2508, N2379, N2259, N2139, N2066, N2001, N1936, N1871, N1806, N1741, N1676, N1611, N1546, N1442, N1377, N1280, N1215, N1150, N1085, N1020, N949, N884, N819, N754, N689, N585, N472, N407, N342, N277, N6359, N6230, N6110, N5990, N5910, N5830, N5765, N5700, N5635, N5570, N5505, N5440, N5375, N5271, N5206, N5109, N5044, N4979, N4900, N4835, N4770, N4705, N4640, N4575, N4510, N4406, N4293, N4180, N4067, N3988, N3923, N3858, N3793, N3728, N3663, N3598, N3533, N3429, N3364, N3299, N3196, N3131, N3066, N3001, N2936, N2871, N2806, N2741, N2676, N2572, N2507, N2378, N2258, N2138, N2065, N2000, N1935, N1870, N1805, N1740, N1675, N1610, N1545, N1441, N1376, N1279, N1214, N1149, N1084, N1019, N948, N883, N818, N753, N688, N584, N471, N406, N341, N276, N6358, N6229, N6109, N5989, N5909, N5829, N5764, N5699, N5634, N5569, N5504, N5439, N5374, N5270, N5205, N5108, N5043, N4978, N4899, N4834, N4769, N4704, N4639, N4574, N4509, N4405, N4292, N4179, N4066, N3987, N3922, N3857, N3792, N3727, N3662, N3597, N3532, N3428, N3363, N3298, N3195, N3130, N3065, N3000, N2935, N2870, N2805, N2740, N2675, N2571, N2506, N2377, N2257, N2137, N2064, N1999, N1934, N1869, N1804, N1739, N1674, N1609, N1544, N1440, N1375, N1278, N1213, N1148, N1083, N1018, N947, N882, N817, N752, N687, N583, N470, N405, N340, N275, N6357, N6228, N6108, N5988, N5908, N5828, N5763, N5698, N5633, N5568, N5503, N5438, N5373, N5269, N5204, N5107, N5042, N4977, N4898, N4833, N4768, N4703, N4638, N4573, N4508, N4404, N4291, N4178, N4065, N3986, N3921, N3856, N3791, N3726, N3661, N3596, N3531, N3427, N3362, N3297, N3194, N3129, N3064, N2999, N2934, N2869, N2804, N2739, N2674, N2570, N2505, N2376, N2256, N2136, N2063, N1998, N1933, N1868, N1803, N1738, N1673, N1608, N1543, N1439, N1374, N1277, N1212, N1147, N1082, N1017, N946, N881, N816, N751, N686, N582, N469, N404, N339, N274, N6356, N6227, N6107, N5987, N5907, N5827, N5762, N5697, N5632, N5567, N5502, N5437, N5372, N5268, N5203, N5106, N5041, N4976, N4897, N4832, N4767, N4702, N4637, N4572, N4507, N4403, N4290, N4177, N4064, N3985, N3920, N3855, N3790, N3725, N3660, N3595, N3530, N3426, N3361, N3296, N3193, N3128, N3063, N2998, N2933, N2868, N2803, N2738, N2673, N2569, N2504, N2375, N2255, N2135, N2062, N1997, N1932, N1867, N1802, N1737, N1672, N1607, N1542, N1438, N1373, N1276, N1211, N1146, N1081, N1016, N945, N880, N815, N750, N685, N581, N468, N403, N338, N273, N6355, N6226, N6106, N5986, N5906, N5826, N5761, N5696, N5631, N5566, N5501, N5436, N5371, N5267, N5202, N5105, N5040, N4975, N4896, N4831, N4766, N4701, N4636, N4571, N4506, N4402, N4289, N4176, N4063, N3984, N3919, N3854, N3789, N3724, N3659, N3594, N3529, N3425, N3360, N3295, N3192, N3127, N3062, N2997, N2932, N2867, N2802, N2737, N2672, N2568, N2503, N2374, N2254, N2134, N2061, N1996, N1931, N1866, N1801, N1736, N1671, N1606, N1541, N1437, N1372, N1275, N1210, N1145, N1080, N1015, N944, N879, N814, N749, N684, N580, N467, N402, N337, N272, N6354, N6225, N6105, N5985, N5905, N5825, N5760, N5695, N5630, N5565, N5500, N5435, N5370, N5266, N5201, N5104, N5039, N4974, N4895, N4830, N4765, N4700, N4635, N4570, N4505, N4401, N4288, N4175, N4062, N3983, N3918, N3853, N3788, N3723, N3658, N3593, N3528, N3424, N3359, N3294, N3191, N3126, N3061, N2996, N2931, N2866, N2801, N2736, N2671, N2567, N2502, N2373, N2253, N2133, N2060, N1995, N1930, N1865, N1800, N1735, N1670, N1605, N1540, N1436, N1371, N1274, N1209, N1144, N1079, N1014, N943, N878, N813, N748, N683, N579, N466, N401, N336, N271, N6353, N6224, N6104, N5984, N5904, N5824, N5759, N5694, N5629, N5564, N5499, N5434, N5369, N5265, N5200, N5103, N5038, N4973, N4894, N4829, N4764, N4699, N4634, N4569, N4504, N4400, N4287, N4174, N4061, N3982, N3917, N3852, N3787, N3722, N3657, N3592, N3527, N3423, N3358, N3293, N3190, N3125, N3060, N2995, N2930, N2865, N2800, N2735, N2670, N2566, N2501, N2372, N2252, N2132, N2059, N1994, N1929, N1864, N1799, N1734, N1669, N1604, N1539, N1435, N1370, N1273, N1208, N1143, N1078, N1013, N942, N877, N812, N747, N682, N578, N465, N400, N335, N270, N6352, N6223, N6103, N5983, N5903, N5823, N5758, N5693, N5628, N5563, N5498, N5433, N5368, N5264, N5199, N5102, N5037, N4972, N4893, N4828, N4763, N4698, N4633, N4568, N4503, N4399, N4286, N4173, N4060, N3981, N3916, N3851, N3786, N3721, N3656, N3591, N3526, N3422, N3357, N3292, N3189, N3124, N3059, N2994, N2929, N2864, N2799, N2734, N2669, N2565, N2500, N2371, N2251, N2131, N2058, N1993, N1928, N1863, N1798, N1733, N1668, N1603, N1538, N1434, N1369, N1272, N1207, N1142, N1077, N1012, N941, N876, N811, N746, N681, N577, N464, N399, N334, N269, N6351, N6222, N6102, N5982, N5902, N5822, N5757, N5692, N5627, N5562, N5497, N5432, N5367, N5263, N5198, N5101, N5036, N4971, N4892, N4827, N4762, N4697, N4632, N4567, N4502, N4398, N4285, N4172, N4059, N3980, N3915, N3850, N3785, N3720, N3655, N3590, N3525, N3421, N3356, N3291, N3188, N3123, N3058, N2993, N2928, N2863, N2798, N2733, N2668, N2564, N2499, N2370, N2250, N2130, N2057, N1992, N1927, N1862, N1797, N1732, N1667, N1602, N1537, N1433, N1368, N1271, N1206, N1141, N1076, N1011, N940, N875, N810, N745, N680, N576, N463, N398, N333, N268, N6350, N6221, N6101, N5981, N5901, N5821, N5756, N5691, N5626, N5561, N5496, N5431, N5366, N5262, N5197, N5100, N5035, N4970, N4891, N4826, N4761, N4696, N4631, N4566, N4501, N4397, N4284, N4171, N4058, N3979, N3914, N3849, N3784, N3719, N3654, N3589, N3524, N3420, N3355, N3290, N3187, N3122, N3057, N2992, N2927, N2862, N2797, N2732, N2667, N2563, N2498, N2369, N2249, N2129, N2056, N1991, N1926, N1861, N1796, N1731, N1666, N1601, N1536, N1432, N1367, N1270, N1205, N1140, N1075, N1010, N939, N874, N809, N744, N679, N575, N462, N397, N332, N267, N6349, N6220, N6100, N5980, N5900, N5820, N5755, N5690, N5625, N5560, N5495, N5430, N5365, N5261, N5196, N5099, N5034, N4969, N4890, N4825, N4760, N4695, N4630, N4565, N4500, N4396, N4283, N4170, N4057, N3978, N3913, N3848, N3783, N3718, N3653, N3588, N3523, N3419, N3354, N3289, N3186, N3121, N3056, N2991, N2926, N2861, N2796, N2731, N2666, N2562, N2497, N2368, N2248, N2128, N2055, N1990, N1925, N1860, N1795, N1730, N1665, N1600, N1535, N1431, N1366, N1269, N1204, N1139, N1074, N1009, N938, N873, N808, N743, N678, N574, N461, N396, N331, N266, N6348, N6219, N6099, N5979, N5899, N5819, N5754, N5689, N5624, N5559, N5494, N5429, N5364, N5260, N5195, N5098, N5033, N4968, N4889, N4824, N4759, N4694, N4629, N4564, N4499, N4395, N4282, N4169, N4056, N3977, N3912, N3847, N3782, N3717, N3652, N3587, N3522, N3418, N3353, N3288, N3185, N3120, N3055, N2990, N2925, N2860, N2795, N2730, N2665, N2561, N2496, N2367, N2247, N2127, N2054, N1989, N1924, N1859, N1794, N1729, N1664, N1599, N1534, N1430, N1365, N1268, N1203, N1138, N1073, N1008, N937, N872, N807, N742, N677, N573, N460, N395, N330, N265, N6347, N6218, N6098, N5978, N5898, N5818, N5753, N5688, N5623, N5558, N5493, N5428, N5363, N5259, N5194, N5097, N5032, N4967, N4888, N4823, N4758, N4693, N4628, N4563, N4498, N4394, N4281, N4168, N4055, N3976, N3911, N3846, N3781, N3716, N3651, N3586, N3521, N3417, N3352, N3287, N3184, N3119, N3054, N2989, N2924, N2859, N2794, N2729, N2664, N2560, N2495, N2366, N2246, N2126, N2053, N1988, N1923, N1858, N1793, N1728, N1663, N1598, N1533, N1429, N1364, N1267, N1202, N1137, N1072, N1007, N936, N871, N806, N741, N676, N572, N459, N394, N329, N264, N6346, N6217, N6097, N5977, N5897, N5817, N5752, N5687, N5622, N5557, N5492, N5427, N5362, N5258, N5193, N5096, N5031, N4966, N4887, N4822, N4757, N4692, N4627, N4562, N4497, N4393, N4280, N4167, N4054, N3975, N3910, N3845, N3780, N3715, N3650, N3585, N3520, N3416, N3351, N3286, N3183, N3118, N3053, N2988, N2923, N2858, N2793, N2728, N2663, N2559, N2494, N2365, N2245, N2125, N2052, N1987, N1922, N1857, N1792, N1727, N1662, N1597, N1532, N1428, N1363, N1266, N1201, N1136, N1071, N1006, N935, N870, N805, N740, N675, N571, N458, N393, N328, N263, N6345, N6216, N6096, N5976, N5896, N5816, N5751, N5686, N5621, N5556, N5491, N5426, N5361, N5257, N5192, N5095, N5030, N4965, N4886, N4821, N4756, N4691, N4626, N4561, N4496, N4392, N4279, N4166, N4053, N3974, N3909, N3844, N3779, N3714, N3649, N3584, N3519, N3415, N3350, N3285, N3182, N3117, N3052, N2987, N2922, N2857, N2792, N2727, N2662, N2558, N2493, N2364, N2244, N2124, N2051, N1986, N1921, N1856, N1791, N1726, N1661, N1596, N1531, N1427, N1362, N1265, N1200, N1135, N1070, N1005, N934, N869, N804, N739, N674, N570, N457, N392, N327, N262, N6344, N6215, N6095, N5975, N5895, N5815, N5750, N5685, N5620, N5555, N5490, N5425, N5360, N5256, N5191, N5094, N5029, N4964, N4885, N4820, N4755, N4690, N4625, N4560, N4495, N4391, N4278, N4165, N4052, N3973, N3908, N3843, N3778, N3713, N3648, N3583, N3518, N3414, N3349, N3284, N3181, N3116, N3051, N2986, N2921, N2856, N2791, N2726, N2661, N2557, N2492, N2363, N2243, N2123, N2050, N1985, N1920, N1855, N1790, N1725, N1660, N1595, N1530, N1426, N1361, N1264, N1199, N1134, N1069, N1004, N933, N868, N803, N738, N673, N569, N456, N391, N326, N261, N6343, N6214, N6094, N5974, N5894, N5814, N5749, N5684, N5619, N5554, N5489, N5424, N5359, N5255, N5190, N5093, N5028, N4963, N4884, N4819, N4754, N4689, N4624, N4559, N4494, N4390, N4277, N4164, N4051, N3972, N3907, N3842, N3777, N3712, N3647, N3582, N3517, N3413, N3348, N3283, N3180, N3115, N3050, N2985, N2920, N2855, N2790, N2725, N2660, N2556, N2491, N2362, N2242, N2122, N2049, N1984, N1919, N1854, N1789, N1724, N1659, N1594, N1529, N1425, N1360, N1263, N1198, N1133, N1068, N1003, N932, N867, N802, N737, N672, N568, N455, N390, N325, N260, N6342, N6213, N6093, N5973, N5893, N5813, N5748, N5683, N5618, N5553, N5488, N5423, N5358, N5254, N5189, N5092, N5027, N4962, N4883, N4818, N4753, N4688, N4623, N4558, N4493, N4389, N4276, N4163, N4050, N3971, N3906, N3841, N3776, N3711, N3646, N3581, N3516, N3412, N3347, N3282, N3179, N3114, N3049, N2984, N2919, N2854, N2789, N2724, N2659, N2555, N2490, N2361, N2241, N2121, N2048, N1983, N1918, N1853, N1788, N1723, N1658, N1593, N1528, N1424, N1359, N1262, N1197, N1132, N1067, N1002, N931, N866, N801, N736, N671, N567, N454, N389, N324, N259, N6341, N6212, N6092, N5972, N5892, N5812, N5747, N5682, N5617, N5552, N5487, N5422, N5357, N5253, N5188, N5091, N5026, N4961, N4882, N4817, N4752, N4687, N4622, N4557, N4492, N4388, N4275, N4162, N4049, N3970, N3905, N3840, N3775, N3710, N3645, N3580, N3515, N3411, N3346, N3281, N3178, N3113, N3048, N2983, N2918, N2853, N2788, N2723, N2658, N2554, N2489, N2360, N2240, N2120, N2047, N1982, N1917, N1852, N1787, N1722, N1657, N1592, N1527, N1423, N1358, N1261, N1196, N1131, N1066, N1001, N930, N865, N800, N735, N670, N566, N453, N388, N323, N258, N6340, N6211, N6091, N5971, N5891, N5811, N5746, N5681, N5616, N5551, N5486, N5421, N5356, N5252, N5187, N5090, N5025, N4960, N4881, N4816, N4751, N4686, N4621, N4556, N4491, N4387, N4274, N4161, N4048, N3969, N3904, N3839, N3774, N3709, N3644, N3579, N3514, N3410, N3345, N3280, N3177, N3112, N3047, N2982, N2917, N2852, N2787, N2722, N2657, N2553, N2488, N2359, N2239, N2119, N2046, N1981, N1916, N1851, N1786, N1721, N1656, N1591, N1526, N1422, N1357, N1260, N1195, N1130, N1065, N1000, N929, N864, N799, N734, N669, N565, N452, N387, N322, N257, N6339, N6210, N6090, N5970, N5890, N5810, N5745, N5680, N5615, N5550, N5485, N5420, N5355, N5251, N5186, N5089, N5024, N4959, N4880, N4815, N4750, N4685, N4620, N4555, N4490, N4386, N4273, N4160, N4047, N3968, N3903, N3838, N3773, N3708, N3643, N3578, N3513, N3409, N3344, N3279, N3176, N3111, N3046, N2981, N2916, N2851, N2786, N2721, N2656, N2552, N2487, N2358, N2238, N2118, N2045, N1980, N1915, N1850, N1785, N1720, N1655, N1590, N1525, N1421, N1356, N1259, N1194, N1129, N1064, N999, N928, N863, N798, N733, N668, N564, N451, N386, N321, N256, N6338, N6209, N6089, N5969, N5889, N5809, N5744, N5679, N5614, N5549, N5484, N5419, N5354, N5250, N5185, N5088, N5023, N4958, N4879, N4814, N4749, N4684, N4619, N4554, N4489, N4385, N4272, N4159, N4046, N3967, N3902, N3837, N3772, N3707, N3642, N3577, N3512, N3408, N3343, N3278, N3175, N3110, N3045, N2980, N2915, N2850, N2785, N2720, N2655, N2551, N2486, N2357, N2237, N2117, N2044, N1979, N1914, N1849, N1784, N1719, N1654, N1589, N1524, N1420, N1355, N1258, N1193, N1128, N1063, N998, N927, N862, N797, N732, N667, N563, N450, N385, N320, N255, N6337, N6208, N6088, N5968, N5888, N5808, N5743, N5678, N5613, N5548, N5483, N5418, N5353, N5249, N5184, N5087, N5022, N4957, N4878, N4813, N4748, N4683, N4618, N4553, N4488, N4384, N4271, N4158, N4045, N3966, N3901, N3836, N3771, N3706, N3641, N3576, N3511, N3407, N3342, N3277, N3174, N3109, N3044, N2979, N2914, N2849, N2784, N2719, N2654, N2550, N2485, N2356, N2236, N2116, N2043, N1978, N1913, N1848, N1783, N1718, N1653, N1588, N1523, N1419, N1354, N1257, N1192, N1127, N1062, N997, N926, N861, N796, N731, N666, N562, N449, N384, N319, N254, N6336, N6207, N6087, N5967, N5887, N5807, N5742, N5677, N5612, N5547, N5482, N5417, N5352, N5248, N5183, N5086, N5021, N4956, N4877, N4812, N4747, N4682, N4617, N4552, N4487, N4383, N4270, N4157, N4044, N3965, N3900, N3835, N3770, N3705, N3640, N3575, N3510, N3406, N3341, N3276, N3173, N3108, N3043, N2978, N2913, N2848, N2783, N2718, N2653, N2549, N2484, N2355, N2235, N2115, N2042, N1977, N1912, N1847, N1782, N1717, N1652, N1587, N1522, N1418, N1353, N1256, N1191, N1126, N1061, N996, N925, N860, N795, N730, N665, N561, N448, N383, N318, N253, N6335, N6206, N6086, N5966, N5886, N5806, N5741, N5676, N5611, N5546, N5481, N5416, N5351, N5247, N5182, N5085, N5020, N4955, N4876, N4811, N4746, N4681, N4616, N4551, N4486, N4382, N4269, N4156, N4043, N3964, N3899, N3834, N3769, N3704, N3639, N3574, N3509, N3405, N3340, N3275, N3172, N3107, N3042, N2977, N2912, N2847, N2782, N2717, N2652, N2548, N2483, N2354, N2234, N2114, N2041, N1976, N1911, N1846, N1781, N1716, N1651, N1586, N1521, N1417, N1352, N1255, N1190, N1125, N1060, N995, N924, N859, N794, N729, N664, N560, N447, N382, N317, N252, N6334, N6205, N6085, N5965, N5885, N5805, N5740, N5675, N5610, N5545, N5480, N5415, N5350, N5246, N5181, N5084, N5019, N4954, N4875, N4810, N4745, N4680, N4615, N4550, N4485, N4381, N4268, N4155, N4042, N3963, N3898, N3833, N3768, N3703, N3638, N3573, N3508, N3404, N3339, N3274, N3171, N3106, N3041, N2976, N2911, N2846, N2781, N2716, N2651, N2547, N2482, N2353, N2233, N2113, N2040, N1975, N1910, N1845, N1780, N1715, N1650, N1585, N1520, N1416, N1351, N1254, N1189, N1124, N1059, N994, N923, N858, N793, N728, N663, N559, N446, N381, N316, N251, N6333, N6204, N6084, N5964, N5884, N5804, N5739, N5674, N5609, N5544, N5479, N5414, N5349, N5245, N5180, N5083, N5018, N4953, N4874, N4809, N4744, N4679, N4614, N4549, N4484, N4380, N4267, N4154, N4041, N3962, N3897, N3832, N3767, N3702, N3637, N3572, N3507, N3403, N3338, N3273, N3170, N3105, N3040, N2975, N2910, N2845, N2780, N2715, N2650, N2546, N2481, N2352, N2232, N2112, N2039, N1974, N1909, N1844, N1779, N1714, N1649, N1584, N1519, N1415, N1350, N1253, N1188, N1123, N1058, N993, N922, N857, N792, N727, N662, N558, N445, N380, N315, N250, N6332, N6203, N6083, N5963, N5883, N5803, N5738, N5673, N5608, N5543, N5478, N5413, N5348, N5244, N5179, N5082, N5017, N4952, N4873, N4808, N4743, N4678, N4613, N4548, N4483, N4379, N4266, N4153, N4040, N3961, N3896, N3831, N3766, N3701, N3636, N3571, N3506, N3402, N3337, N3272, N3169, N3104, N3039, N2974, N2909, N2844, N2779, N2714, N2649, N2545, N2480, N2351, N2231, N2111, N2038, N1973, N1908, N1843, N1778, N1713, N1648, N1583, N1518, N1414, N1349, N1252, N1187, N1122, N1057, N992, N921, N856, N791, N726, N661, N557, N444, N379, N314, N249, N6331, N6202, N6082, N5962, N5882, N5802, N5737, N5672, N5607, N5542, N5477, N5412, N5347, N5243, N5178, N5081, N5016, N4951, N4872, N4807, N4742, N4677, N4612, N4547, N4482, N4378, N4265, N4152, N4039, N3960, N3895, N3830, N3765, N3700, N3635, N3570, N3505, N3401, N3336, N3271, N3168, N3103, N3038, N2973, N2908, N2843, N2778, N2713, N2648, N2544, N2479, N2350, N2230, N2110, N2037, N1972, N1907, N1842, N1777, N1712, N1647, N1582, N1517, N1413, N1348, N1251, N1186, N1121, N1056, N991, N920, N855, N790, N725, N660, N556, N443, N378, N313, N248, N6330, N6201, N6081, N5961, N5881, N5801, N5736, N5671, N5606, N5541, N5476, N5411, N5346, N5242, N5177, N5080, N5015, N4950, N4871, N4806, N4741, N4676, N4611, N4546, N4481, N4377, N4264, N4151, N4038, N3959, N3894, N3829, N3764, N3699, N3634, N3569, N3504, N3400, N3335, N3270, N3167, N3102, N3037, N2972, N2907, N2842, N2777, N2712, N2647, N2543, N2478, N2349, N2229, N2109, N2036, N1971, N1906, N1841, N1776, N1711, N1646, N1581, N1516, N1412, N1347, N1250, N1185, N1120, N1055, N990, N919, N854, N789, N724, N659, N555, N442, N377, N312, N247, N6329, N6200, N6080, N5960, N5880, N5800, N5735, N5670, N5605, N5540, N5475, N5410, N5345, N5241, N5176, N5079, N5014, N4949, N4870, N4805, N4740, N4675, N4610, N4545, N4480, N4376, N4263, N4150, N4037, N3958, N3893, N3828, N3763, N3698, N3633, N3568, N3503, N3399, N3334, N3269, N3166, N3101, N3036, N2971, N2906, N2841, N2776, N2711, N2646, N2542, N2477, N2348, N2228, N2108, N2035, N1970, N1905, N1840, N1775, N1710, N1645, N1580, N1515, N1411, N1346, N1249, N1184, N1119, N1054, N989, N918, N853, N788, N723, N658, N554, N441, N376, N311, N246, N6328, N6199, N6079, N5959, N5879, N5799, N5734, N5669, N5604, N5539, N5474, N5409, N5344, N5240, N5175, N5078, N5013, N4948, N4869, N4804, N4739, N4674, N4609, N4544, N4479, N4375, N4262, N4149, N4036, N3957, N3892, N3827, N3762, N3697, N3632, N3567, N3502, N3398, N3333, N3268, N3165, N3100, N3035, N2970, N2905, N2840, N2775, N2710, N2645, N2541, N2476, N2347, N2227, N2107, N2034, N1969, N1904, N1839, N1774, N1709, N1644, N1579, N1514, N1410, N1345, N1248, N1183, N1118, N1053, N988, N917, N852, N787, N722, N657, N553, N440, N375, N310, N245, N6327, N6198, N6078, N5958, N5878, N5798, N5733, N5668, N5603, N5538, N5473, N5408, N5343, N5239, N5174, N5077, N5012, N4947, N4868, N4803, N4738, N4673, N4608, N4543, N4478, N4374, N4261, N4148, N4035, N3956, N3891, N3826, N3761, N3696, N3631, N3566, N3501, N3397, N3332, N3267, N3164, N3099, N3034, N2969, N2904, N2839, N2774, N2709, N2644, N2540, N2475, N2346, N2226, N2106, N2033, N1968, N1903, N1838, N1773, N1708, N1643, N1578, N1513, N1409, N1344, N1247, N1182, N1117, N1052, N987, N916, N851, N786, N721, N656, N552, N439, N374, N309, N244, N6326, N6197, N6077, N5957, N5877, N5797, N5732, N5667, N5602, N5537, N5472, N5407, N5342, N5238, N5173, N5076, N5011, N4946, N4867, N4802, N4737, N4672, N4607, N4542, N4477, N4373, N4260, N4147, N4034, N3955, N3890, N3825, N3760, N3695, N3630, N3565, N3500, N3396, N3331, N3266, N3163, N3098, N3033, N2968, N2903, N2838, N2773, N2708, N2643, N2539, N2474, N2345, N2225, N2105, N2032, N1967, N1902, N1837, N1772, N1707, N1642, N1577, N1512, N1408, N1343, N1246, N1181, N1116, N1051, N986, N915, N850, N785, N720, N655, N551, N438, N373, N308, N243, N6325, N6196, N6076, N5956, N5876, N5796, N5731, N5666, N5601, N5536, N5471, N5406, N5341, N5237, N5172, N5075, N5010, N4945, N4866, N4801, N4736, N4671, N4606, N4541, N4476, N4372, N4259, N4146, N4033, N3954, N3889, N3824, N3759, N3694, N3629, N3564, N3499, N3395, N3330, N3265, N3162, N3097, N3032, N2967, N2902, N2837, N2772, N2707, N2642, N2538, N2473, N2344, N2224, N2104, N2031, N1966, N1901, N1836, N1771, N1706, N1641, N1576, N1511, N1407, N1342, N1245, N1180, N1115, N1050, N985, N914, N849, N784, N719, N654, N550, N437, N372, N307, N242, N6324, N6195, N6075, N5955, N5875, N5795, N5730, N5665, N5600, N5535, N5470, N5405, N5340, N5236, N5171, N5074, N5009, N4944, N4865, N4800, N4735, N4670, N4605, N4540, N4475, N4371, N4258, N4145, N4032, N3953, N3888, N3823, N3758, N3693, N3628, N3563, N3498, N3394, N3329, N3264, N3161, N3096, N3031, N2966, N2901, N2836, N2771, N2706, N2641, N2537, N2472, N2343, N2223, N2103, N2030, N1965, N1900, N1835, N1770, N1705, N1640, N1575, N1510, N1406, N1341, N1244, N1179, N1114, N1049, N984, N913, N848, N783, N718, N653, N549, N436, N371, N306, N241, N6323, N6194, N6074, N5954, N5874, N5794, N5729, N5664, N5599, N5534, N5469, N5404, N5339, N5235, N5170, N5073, N5008, N4943, N4864, N4799, N4734, N4669, N4604, N4539, N4474, N4370, N4257, N4144, N4031, N3952, N3887, N3822, N3757, N3692, N3627, N3562, N3497, N3393, N3328, N3263, N3160, N3095, N3030, N2965, N2900, N2835, N2770, N2705, N2640, N2536, N2471, N2342, N2222, N2102, N2029, N1964, N1899, N1834, N1769, N1704, N1639, N1574, N1509, N1405, N1340, N1243, N1178, N1113, N1048, N983, N912, N847, N782, N717, N652, N548, N435, N370, N305, N240, N6322, N6193, N6073, N5953, N5873, N5793, N5728, N5663, N5598, N5533, N5468, N5403, N5338, N5234, N5169, N5072, N5007, N4942, N4863, N4798, N4733, N4668, N4603, N4538, N4473, N4369, N4256, N4143, N4030, N3951, N3886, N3821, N3756, N3691, N3626, N3561, N3496, N3392, N3327, N3262, N3159, N3094, N3029, N2964, N2899, N2834, N2769, N2704, N2639, N2535, N2470, N2341, N2221, N2101, N2028, N1963, N1898, N1833, N1768, N1703, N1638, N1573, N1508, N1404, N1339, N1242, N1177, N1112, N1047, N982, N911, N846, N781, N716, N651, N547, N434, N369, N304, N239, N6321, N6192, N6072, N5952, N5872, N5792, N5727, N5662, N5597, N5532, N5467, N5402, N5337, N5233, N5168, N5071, N5006, N4941, N4862, N4797, N4732, N4667, N4602, N4537, N4472, N4368, N4255, N4142, N4029, N3950, N3885, N3820, N3755, N3690, N3625, N3560, N3495, N3391, N3326, N3261, N3158, N3093, N3028, N2963, N2898, N2833, N2768, N2703, N2638, N2534, N2469, N2340, N2220, N2100, N2027, N1962, N1897, N1832, N1767, N1702, N1637, N1572, N1507, N1403, N1338, N1241, N1176, N1111, N1046, N981, N910, N845, N780, N715, N650, N546, N433, N368, N303, N238, N6320, N6191, N6071, N5951, N5871, N5791, N5726, N5661, N5596, N5531, N5466, N5401, N5336, N5232, N5167, N5070, N5005, N4940, N4861, N4796, N4731, N4666, N4601, N4536, N4471, N4367, N4254, N4141, N4028, N3949, N3884, N3819, N3754, N3689, N3624, N3559, N3494, N3390, N3325, N3260, N3157, N3092, N3027, N2962, N2897, N2832, N2767, N2702, N2637, N2533, N2468, N2339, N2219, N2099, N2026, N1961, N1896, N1831, N1766, N1701, N1636, N1571, N1506, N1402, N1337, N1240, N1175, N1110, N1045, N980, N909, N844, N779, N714, N649, N545, N432, N367, N302, N237, N6319, N6190, N6070, N5950, N5870, N5790, N5725, N5660, N5595, N5530, N5465, N5400, N5335, N5231, N5166, N5069, N5004, N4939, N4860, N4795, N4730, N4665, N4600, N4535, N4470, N4366, N4253, N4140, N4027, N3948, N3883, N3818, N3753, N3688, N3623, N3558, N3493, N3389, N3324, N3259, N3156, N3091, N3026, N2961, N2896, N2831, N2766, N2701, N2636, N2532, N2467, N2338, N2218, N2098, N2025, N1960, N1895, N1830, N1765, N1700, N1635, N1570, N1505, N1401, N1336, N1239, N1174, N1109, N1044, N979, N908, N843, N778, N713, N648, N544, N431, N366, N301, N236, N6318, N6189, N6069, N5949, N5869, N5789, N5724, N5659, N5594, N5529, N5464, N5399, N5334, N5230, N5165, N5068, N5003, N4938, N4859, N4794, N4729, N4664, N4599, N4534, N4469, N4365, N4252, N4139, N4026, N3947, N3882, N3817, N3752, N3687, N3622, N3557, N3492, N3388, N3323, N3258, N3155, N3090, N3025, N2960, N2895, N2830, N2765, N2700, N2635, N2531, N2466, N2337, N2217, N2097, N2024, N1959, N1894, N1829, N1764, N1699, N1634, N1569, N1504, N1400, N1335, N1238, N1173, N1108, N1043, N978, N907, N842, N777, N712, N647, N543, N430, N365, N300, N235, N6317, N6188, N6068, N5948, N5868, N5788, N5723, N5658, N5593, N5528, N5463, N5398, N5333, N5229, N5164, N5067, N5002, N4937, N4858, N4793, N4728, N4663, N4598, N4533, N4468, N4364, N4251, N4138, N4025, N3946, N3881, N3816, N3751, N3686, N3621, N3556, N3491, N3387, N3322, N3257, N3154, N3089, N3024, N2959, N2894, N2829, N2764, N2699, N2634, N2530, N2465, N2336, N2216, N2096, N2023, N1958, N1893, N1828, N1763, N1698, N1633, N1568, N1503, N1399, N1334, N1237, N1172, N1107, N1042, N977, N906, N841, N776, N711, N646, N542, N429, N364, N299, N234, N6316, N6187, N6067, N5947, N5867, N5787, N5722, N5657, N5592, N5527, N5462, N5397, N5332, N5228, N5163, N5066, N5001, N4936, N4857, N4792, N4727, N4662, N4597, N4532, N4467, N4363, N4250, N4137, N4024, N3945, N3880, N3815, N3750, N3685, N3620, N3555, N3490, N3386, N3321, N3256, N3153, N3088, N3023, N2958, N2893, N2828, N2763, N2698, N2633, N2529, N2464, N2335, N2215, N2095, N2022, N1957, N1892, N1827, N1762, N1697, N1632, N1567, N1502, N1398, N1333, N1236, N1171, N1106, N1041, N976, N905, N840, N775, N710, N645, N541, N428, N363, N298, N233, N6315, N6186, N6066, N5946, N5866, N5786, N5721, N5656, N5591, N5526, N5461, N5396, N5331, N5227, N5162, N5065, N5000, N4935, N4856, N4791, N4726, N4661, N4596, N4531, N4466, N4362, N4249, N4136, N4023, N3944, N3879, N3814, N3749, N3684, N3619, N3554, N3489, N3385, N3320, N3255, N3152, N3087, N3022, N2957, N2892, N2827, N2762, N2697, N2632, N2528, N2463, N2334, N2214, N2094, N2021, N1956, N1891, N1826, N1761, N1696, N1631, N1566, N1501, N1397, N1332, N1235, N1170, N1105, N1040, N975, N904, N839, N774, N709, N644, N540, N427, N362, N297, N232, N6314, N6185, N6065, N5945, N5865, N5785, N5720, N5655, N5590, N5525, N5460, N5395, N5330, N5226, N5161, N5064, N4999, N4934, N4855, N4790, N4725, N4660, N4595, N4530, N4465, N4361, N4248, N4135, N4022, N3943, N3878, N3813, N3748, N3683, N3618, N3553, N3488, N3384, N3319, N3254, N3151, N3086, N3021, N2956, N2891, N2826, N2761, N2696, N2631, N2527, N2462, N2333, N2213, N2093, N2020, N1955, N1890, N1825, N1760, N1695, N1630, N1565, N1500, N1396, N1331, N1234, N1169, N1104, N1039, N974, N903, N838, N773, N708, N643, N539, N426, N361, N296, N231, N6313, N6184, N6064, N5944, N5864, N5784, N5719, N5654, N5589, N5524, N5459, N5394, N5329, N5225, N5160, N5063, N4998, N4933, N4854, N4789, N4724, N4659, N4594, N4529, N4464, N4360, N4247, N4134, N4021, N3942, N3877, N3812, N3747, N3682, N3617, N3552, N3487, N3383, N3318, N3253, N3150, N3085, N3020, N2955, N2890, N2825, N2760, N2695, N2630, N2526, N2461, N2332, N2212, N2092, N2019, N1954, N1889, N1824, N1759, N1694, N1629, N1564, N1499, N1395, N1330, N1233, N1168, N1103, N1038, N973, N902, N837, N772, N707, N642, N538, N425, N360, N295, N230 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N228)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N96 = N227;
  assign \nz.read_en  = v_i & N11659;
  assign N11659 = ~w_i;
  assign N97 = ~\nz.addr_r [0];
  assign N98 = ~\nz.addr_r [1];
  assign N99 = N97 & N98;
  assign N100 = N97 & \nz.addr_r [1];
  assign N101 = \nz.addr_r [0] & N98;
  assign N102 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N103 = ~\nz.addr_r [2];
  assign N104 = N99 & N103;
  assign N105 = N99 & \nz.addr_r [2];
  assign N106 = N101 & N103;
  assign N107 = N101 & \nz.addr_r [2];
  assign N108 = N100 & N103;
  assign N109 = N100 & \nz.addr_r [2];
  assign N110 = N102 & N103;
  assign N111 = N102 & \nz.addr_r [2];
  assign N112 = ~\nz.addr_r [3];
  assign N113 = N104 & N112;
  assign N114 = N104 & \nz.addr_r [3];
  assign N115 = N106 & N112;
  assign N116 = N106 & \nz.addr_r [3];
  assign N117 = N108 & N112;
  assign N118 = N108 & \nz.addr_r [3];
  assign N119 = N110 & N112;
  assign N120 = N110 & \nz.addr_r [3];
  assign N121 = N105 & N112;
  assign N122 = N105 & \nz.addr_r [3];
  assign N123 = N107 & N112;
  assign N124 = N107 & \nz.addr_r [3];
  assign N125 = N109 & N112;
  assign N126 = N109 & \nz.addr_r [3];
  assign N127 = N111 & N112;
  assign N128 = N111 & \nz.addr_r [3];
  assign N129 = ~\nz.addr_r [4];
  assign N130 = N113 & N129;
  assign N131 = N113 & \nz.addr_r [4];
  assign N132 = N115 & N129;
  assign N133 = N115 & \nz.addr_r [4];
  assign N134 = N117 & N129;
  assign N135 = N117 & \nz.addr_r [4];
  assign N136 = N119 & N129;
  assign N137 = N119 & \nz.addr_r [4];
  assign N138 = N121 & N129;
  assign N139 = N121 & \nz.addr_r [4];
  assign N140 = N123 & N129;
  assign N141 = N123 & \nz.addr_r [4];
  assign N142 = N125 & N129;
  assign N143 = N125 & \nz.addr_r [4];
  assign N144 = N127 & N129;
  assign N145 = N127 & \nz.addr_r [4];
  assign N146 = N114 & N129;
  assign N147 = N114 & \nz.addr_r [4];
  assign N148 = N116 & N129;
  assign N149 = N116 & \nz.addr_r [4];
  assign N150 = N118 & N129;
  assign N151 = N118 & \nz.addr_r [4];
  assign N152 = N120 & N129;
  assign N153 = N120 & \nz.addr_r [4];
  assign N154 = N122 & N129;
  assign N155 = N122 & \nz.addr_r [4];
  assign N156 = N124 & N129;
  assign N157 = N124 & \nz.addr_r [4];
  assign N158 = N126 & N129;
  assign N159 = N126 & \nz.addr_r [4];
  assign N160 = N128 & N129;
  assign N161 = N128 & \nz.addr_r [4];
  assign N162 = ~\nz.addr_r [5];
  assign N163 = N130 & N162;
  assign N164 = N130 & \nz.addr_r [5];
  assign N165 = N132 & N162;
  assign N166 = N132 & \nz.addr_r [5];
  assign N167 = N134 & N162;
  assign N168 = N134 & \nz.addr_r [5];
  assign N169 = N136 & N162;
  assign N170 = N136 & \nz.addr_r [5];
  assign N171 = N138 & N162;
  assign N172 = N138 & \nz.addr_r [5];
  assign N173 = N140 & N162;
  assign N174 = N140 & \nz.addr_r [5];
  assign N175 = N142 & N162;
  assign N176 = N142 & \nz.addr_r [5];
  assign N177 = N144 & N162;
  assign N178 = N144 & \nz.addr_r [5];
  assign N179 = N146 & N162;
  assign N180 = N146 & \nz.addr_r [5];
  assign N181 = N148 & N162;
  assign N182 = N148 & \nz.addr_r [5];
  assign N183 = N150 & N162;
  assign N184 = N150 & \nz.addr_r [5];
  assign N185 = N152 & N162;
  assign N186 = N152 & \nz.addr_r [5];
  assign N187 = N154 & N162;
  assign N188 = N154 & \nz.addr_r [5];
  assign N189 = N156 & N162;
  assign N190 = N156 & \nz.addr_r [5];
  assign N191 = N158 & N162;
  assign N192 = N158 & \nz.addr_r [5];
  assign N193 = N160 & N162;
  assign N194 = N160 & \nz.addr_r [5];
  assign N195 = N131 & N162;
  assign N196 = N131 & \nz.addr_r [5];
  assign N197 = N133 & N162;
  assign N198 = N133 & \nz.addr_r [5];
  assign N199 = N135 & N162;
  assign N200 = N135 & \nz.addr_r [5];
  assign N201 = N137 & N162;
  assign N202 = N137 & \nz.addr_r [5];
  assign N203 = N139 & N162;
  assign N204 = N139 & \nz.addr_r [5];
  assign N205 = N141 & N162;
  assign N206 = N141 & \nz.addr_r [5];
  assign N207 = N143 & N162;
  assign N208 = N143 & \nz.addr_r [5];
  assign N209 = N145 & N162;
  assign N210 = N145 & \nz.addr_r [5];
  assign N211 = N147 & N162;
  assign N212 = N147 & \nz.addr_r [5];
  assign N213 = N149 & N162;
  assign N214 = N149 & \nz.addr_r [5];
  assign N215 = N151 & N162;
  assign N216 = N151 & \nz.addr_r [5];
  assign N217 = N153 & N162;
  assign N218 = N153 & \nz.addr_r [5];
  assign N219 = N155 & N162;
  assign N220 = N155 & \nz.addr_r [5];
  assign N221 = N157 & N162;
  assign N222 = N157 & \nz.addr_r [5];
  assign N223 = N159 & N162;
  assign N224 = N159 & \nz.addr_r [5];
  assign N225 = N161 & N162;
  assign N226 = N161 & \nz.addr_r [5];
  assign N227 = v_i & w_i;
  assign N228 = ~N227;
  assign N229 = ~w_mask_i[0];
  assign N294 = ~w_mask_i[1];
  assign N359 = ~w_mask_i[2];
  assign N424 = ~w_mask_i[3];
  assign N489 = ~w_mask_i[4];
  assign N602 = ~w_mask_i[5];
  assign N706 = ~w_mask_i[6];
  assign N771 = ~w_mask_i[7];
  assign N836 = ~w_mask_i[8];
  assign N901 = ~w_mask_i[9];
  assign N966 = ~w_mask_i[10];
  assign N1037 = ~w_mask_i[11];
  assign N1102 = ~w_mask_i[12];
  assign N1167 = ~w_mask_i[13];
  assign N1232 = ~w_mask_i[14];
  assign N1297 = ~w_mask_i[15];
  assign N1394 = ~w_mask_i[16];
  assign N1459 = ~w_mask_i[17];
  assign N1563 = ~w_mask_i[18];
  assign N1628 = ~w_mask_i[19];
  assign N1693 = ~w_mask_i[20];
  assign N1758 = ~w_mask_i[21];
  assign N1823 = ~w_mask_i[22];
  assign N1888 = ~w_mask_i[23];
  assign N1953 = ~w_mask_i[24];
  assign N2018 = ~w_mask_i[25];
  assign N2083 = ~w_mask_i[26];
  assign N2156 = ~w_mask_i[27];
  assign N2276 = ~w_mask_i[28];
  assign N2396 = ~w_mask_i[29];
  assign N2525 = ~w_mask_i[30];
  assign N2590 = ~w_mask_i[31];
  assign N2694 = ~w_mask_i[32];
  assign N2759 = ~w_mask_i[33];
  assign N2824 = ~w_mask_i[34];
  assign N2889 = ~w_mask_i[35];
  assign N2954 = ~w_mask_i[36];
  assign N3019 = ~w_mask_i[37];
  assign N3084 = ~w_mask_i[38];
  assign N3149 = ~w_mask_i[39];
  assign N3214 = ~w_mask_i[40];
  assign N3317 = ~w_mask_i[41];
  assign N3382 = ~w_mask_i[42];
  assign N3447 = ~w_mask_i[43];
  assign N3551 = ~w_mask_i[44];
  assign N3616 = ~w_mask_i[45];
  assign N3681 = ~w_mask_i[46];
  assign N3746 = ~w_mask_i[47];
  assign N3811 = ~w_mask_i[48];
  assign N3876 = ~w_mask_i[49];
  assign N3941 = ~w_mask_i[50];
  assign N4006 = ~w_mask_i[51];
  assign N4085 = ~w_mask_i[52];
  assign N4198 = ~w_mask_i[53];
  assign N4311 = ~w_mask_i[54];
  assign N4424 = ~w_mask_i[55];
  assign N4528 = ~w_mask_i[56];
  assign N4593 = ~w_mask_i[57];
  assign N4658 = ~w_mask_i[58];
  assign N4723 = ~w_mask_i[59];
  assign N4788 = ~w_mask_i[60];
  assign N4853 = ~w_mask_i[61];
  assign N4918 = ~w_mask_i[62];
  assign N4997 = ~w_mask_i[63];
  assign N5062 = ~w_mask_i[64];
  assign N5127 = ~w_mask_i[65];
  assign N5224 = ~w_mask_i[66];
  assign N5289 = ~w_mask_i[67];
  assign N5393 = ~w_mask_i[68];
  assign N5458 = ~w_mask_i[69];
  assign N5523 = ~w_mask_i[70];
  assign N5588 = ~w_mask_i[71];
  assign N5653 = ~w_mask_i[72];
  assign N5718 = ~w_mask_i[73];
  assign N5783 = ~w_mask_i[74];
  assign N5848 = ~w_mask_i[75];
  assign N5928 = ~w_mask_i[76];
  assign N6008 = ~w_mask_i[77];
  assign N6128 = ~w_mask_i[78];
  assign N6248 = ~w_mask_i[79];

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N11496) begin
      \nz.mem_5119_sv2v_reg  <= data_i[79];
    end 
    if(N11495) begin
      \nz.mem_5118_sv2v_reg  <= data_i[78];
    end 
    if(N11494) begin
      \nz.mem_5117_sv2v_reg  <= data_i[77];
    end 
    if(N11493) begin
      \nz.mem_5116_sv2v_reg  <= data_i[76];
    end 
    if(N11492) begin
      \nz.mem_5115_sv2v_reg  <= data_i[75];
    end 
    if(N11491) begin
      \nz.mem_5114_sv2v_reg  <= data_i[74];
    end 
    if(N11490) begin
      \nz.mem_5113_sv2v_reg  <= data_i[73];
    end 
    if(N11489) begin
      \nz.mem_5112_sv2v_reg  <= data_i[72];
    end 
    if(N11488) begin
      \nz.mem_5111_sv2v_reg  <= data_i[71];
    end 
    if(N11487) begin
      \nz.mem_5110_sv2v_reg  <= data_i[70];
    end 
    if(N11486) begin
      \nz.mem_5109_sv2v_reg  <= data_i[69];
    end 
    if(N11485) begin
      \nz.mem_5108_sv2v_reg  <= data_i[68];
    end 
    if(N11484) begin
      \nz.mem_5107_sv2v_reg  <= data_i[67];
    end 
    if(N11483) begin
      \nz.mem_5106_sv2v_reg  <= data_i[66];
    end 
    if(N11482) begin
      \nz.mem_5105_sv2v_reg  <= data_i[65];
    end 
    if(N11481) begin
      \nz.mem_5104_sv2v_reg  <= data_i[64];
    end 
    if(N11480) begin
      \nz.mem_5103_sv2v_reg  <= data_i[63];
    end 
    if(N11479) begin
      \nz.mem_5102_sv2v_reg  <= data_i[62];
    end 
    if(N11478) begin
      \nz.mem_5101_sv2v_reg  <= data_i[61];
    end 
    if(N11477) begin
      \nz.mem_5100_sv2v_reg  <= data_i[60];
    end 
    if(N11476) begin
      \nz.mem_5099_sv2v_reg  <= data_i[59];
    end 
    if(N11475) begin
      \nz.mem_5098_sv2v_reg  <= data_i[58];
    end 
    if(N11474) begin
      \nz.mem_5097_sv2v_reg  <= data_i[57];
    end 
    if(N11473) begin
      \nz.mem_5096_sv2v_reg  <= data_i[56];
    end 
    if(N11472) begin
      \nz.mem_5095_sv2v_reg  <= data_i[55];
    end 
    if(N11471) begin
      \nz.mem_5094_sv2v_reg  <= data_i[54];
    end 
    if(N11470) begin
      \nz.mem_5093_sv2v_reg  <= data_i[53];
    end 
    if(N11469) begin
      \nz.mem_5092_sv2v_reg  <= data_i[52];
    end 
    if(N11468) begin
      \nz.mem_5091_sv2v_reg  <= data_i[51];
    end 
    if(N11467) begin
      \nz.mem_5090_sv2v_reg  <= data_i[50];
    end 
    if(N11466) begin
      \nz.mem_5089_sv2v_reg  <= data_i[49];
    end 
    if(N11465) begin
      \nz.mem_5088_sv2v_reg  <= data_i[48];
    end 
    if(N11464) begin
      \nz.mem_5087_sv2v_reg  <= data_i[47];
    end 
    if(N11463) begin
      \nz.mem_5086_sv2v_reg  <= data_i[46];
    end 
    if(N11462) begin
      \nz.mem_5085_sv2v_reg  <= data_i[45];
    end 
    if(N11461) begin
      \nz.mem_5084_sv2v_reg  <= data_i[44];
    end 
    if(N11460) begin
      \nz.mem_5083_sv2v_reg  <= data_i[43];
    end 
    if(N11459) begin
      \nz.mem_5082_sv2v_reg  <= data_i[42];
    end 
    if(N11458) begin
      \nz.mem_5081_sv2v_reg  <= data_i[41];
    end 
    if(N11457) begin
      \nz.mem_5080_sv2v_reg  <= data_i[40];
    end 
    if(N11456) begin
      \nz.mem_5079_sv2v_reg  <= data_i[39];
    end 
    if(N11455) begin
      \nz.mem_5078_sv2v_reg  <= data_i[38];
    end 
    if(N11454) begin
      \nz.mem_5077_sv2v_reg  <= data_i[37];
    end 
    if(N11453) begin
      \nz.mem_5076_sv2v_reg  <= data_i[36];
    end 
    if(N11452) begin
      \nz.mem_5075_sv2v_reg  <= data_i[35];
    end 
    if(N11451) begin
      \nz.mem_5074_sv2v_reg  <= data_i[34];
    end 
    if(N11450) begin
      \nz.mem_5073_sv2v_reg  <= data_i[33];
    end 
    if(N11449) begin
      \nz.mem_5072_sv2v_reg  <= data_i[32];
    end 
    if(N11448) begin
      \nz.mem_5071_sv2v_reg  <= data_i[31];
    end 
    if(N11447) begin
      \nz.mem_5070_sv2v_reg  <= data_i[30];
    end 
    if(N11446) begin
      \nz.mem_5069_sv2v_reg  <= data_i[29];
    end 
    if(N11445) begin
      \nz.mem_5068_sv2v_reg  <= data_i[28];
    end 
    if(N11444) begin
      \nz.mem_5067_sv2v_reg  <= data_i[27];
    end 
    if(N11443) begin
      \nz.mem_5066_sv2v_reg  <= data_i[26];
    end 
    if(N11442) begin
      \nz.mem_5065_sv2v_reg  <= data_i[25];
    end 
    if(N11441) begin
      \nz.mem_5064_sv2v_reg  <= data_i[24];
    end 
    if(N11440) begin
      \nz.mem_5063_sv2v_reg  <= data_i[23];
    end 
    if(N11439) begin
      \nz.mem_5062_sv2v_reg  <= data_i[22];
    end 
    if(N11438) begin
      \nz.mem_5061_sv2v_reg  <= data_i[21];
    end 
    if(N11437) begin
      \nz.mem_5060_sv2v_reg  <= data_i[20];
    end 
    if(N11436) begin
      \nz.mem_5059_sv2v_reg  <= data_i[19];
    end 
    if(N11435) begin
      \nz.mem_5058_sv2v_reg  <= data_i[18];
    end 
    if(N11434) begin
      \nz.mem_5057_sv2v_reg  <= data_i[17];
    end 
    if(N11433) begin
      \nz.mem_5056_sv2v_reg  <= data_i[16];
    end 
    if(N11432) begin
      \nz.mem_5055_sv2v_reg  <= data_i[15];
    end 
    if(N11431) begin
      \nz.mem_5054_sv2v_reg  <= data_i[14];
    end 
    if(N11430) begin
      \nz.mem_5053_sv2v_reg  <= data_i[13];
    end 
    if(N11429) begin
      \nz.mem_5052_sv2v_reg  <= data_i[12];
    end 
    if(N11428) begin
      \nz.mem_5051_sv2v_reg  <= data_i[11];
    end 
    if(N11427) begin
      \nz.mem_5050_sv2v_reg  <= data_i[10];
    end 
    if(N11426) begin
      \nz.mem_5049_sv2v_reg  <= data_i[9];
    end 
    if(N11425) begin
      \nz.mem_5048_sv2v_reg  <= data_i[8];
    end 
    if(N11424) begin
      \nz.mem_5047_sv2v_reg  <= data_i[7];
    end 
    if(N11423) begin
      \nz.mem_5046_sv2v_reg  <= data_i[6];
    end 
    if(N11422) begin
      \nz.mem_5045_sv2v_reg  <= data_i[5];
    end 
    if(N11421) begin
      \nz.mem_5044_sv2v_reg  <= data_i[4];
    end 
    if(N11420) begin
      \nz.mem_5043_sv2v_reg  <= data_i[3];
    end 
    if(N11419) begin
      \nz.mem_5042_sv2v_reg  <= data_i[2];
    end 
    if(N11418) begin
      \nz.mem_5041_sv2v_reg  <= data_i[1];
    end 
    if(N11417) begin
      \nz.mem_5040_sv2v_reg  <= data_i[0];
    end 
    if(N11416) begin
      \nz.mem_5039_sv2v_reg  <= data_i[79];
    end 
    if(N11415) begin
      \nz.mem_5038_sv2v_reg  <= data_i[78];
    end 
    if(N11414) begin
      \nz.mem_5037_sv2v_reg  <= data_i[77];
    end 
    if(N11413) begin
      \nz.mem_5036_sv2v_reg  <= data_i[76];
    end 
    if(N11412) begin
      \nz.mem_5035_sv2v_reg  <= data_i[75];
    end 
    if(N11411) begin
      \nz.mem_5034_sv2v_reg  <= data_i[74];
    end 
    if(N11410) begin
      \nz.mem_5033_sv2v_reg  <= data_i[73];
    end 
    if(N11409) begin
      \nz.mem_5032_sv2v_reg  <= data_i[72];
    end 
    if(N11408) begin
      \nz.mem_5031_sv2v_reg  <= data_i[71];
    end 
    if(N11407) begin
      \nz.mem_5030_sv2v_reg  <= data_i[70];
    end 
    if(N11406) begin
      \nz.mem_5029_sv2v_reg  <= data_i[69];
    end 
    if(N11405) begin
      \nz.mem_5028_sv2v_reg  <= data_i[68];
    end 
    if(N11404) begin
      \nz.mem_5027_sv2v_reg  <= data_i[67];
    end 
    if(N11403) begin
      \nz.mem_5026_sv2v_reg  <= data_i[66];
    end 
    if(N11402) begin
      \nz.mem_5025_sv2v_reg  <= data_i[65];
    end 
    if(N11401) begin
      \nz.mem_5024_sv2v_reg  <= data_i[64];
    end 
    if(N11400) begin
      \nz.mem_5023_sv2v_reg  <= data_i[63];
    end 
    if(N11399) begin
      \nz.mem_5022_sv2v_reg  <= data_i[62];
    end 
    if(N11398) begin
      \nz.mem_5021_sv2v_reg  <= data_i[61];
    end 
    if(N11397) begin
      \nz.mem_5020_sv2v_reg  <= data_i[60];
    end 
    if(N11396) begin
      \nz.mem_5019_sv2v_reg  <= data_i[59];
    end 
    if(N11395) begin
      \nz.mem_5018_sv2v_reg  <= data_i[58];
    end 
    if(N11394) begin
      \nz.mem_5017_sv2v_reg  <= data_i[57];
    end 
    if(N11393) begin
      \nz.mem_5016_sv2v_reg  <= data_i[56];
    end 
    if(N11392) begin
      \nz.mem_5015_sv2v_reg  <= data_i[55];
    end 
    if(N11391) begin
      \nz.mem_5014_sv2v_reg  <= data_i[54];
    end 
    if(N11390) begin
      \nz.mem_5013_sv2v_reg  <= data_i[53];
    end 
    if(N11389) begin
      \nz.mem_5012_sv2v_reg  <= data_i[52];
    end 
    if(N11388) begin
      \nz.mem_5011_sv2v_reg  <= data_i[51];
    end 
    if(N11387) begin
      \nz.mem_5010_sv2v_reg  <= data_i[50];
    end 
    if(N11386) begin
      \nz.mem_5009_sv2v_reg  <= data_i[49];
    end 
    if(N11385) begin
      \nz.mem_5008_sv2v_reg  <= data_i[48];
    end 
    if(N11384) begin
      \nz.mem_5007_sv2v_reg  <= data_i[47];
    end 
    if(N11383) begin
      \nz.mem_5006_sv2v_reg  <= data_i[46];
    end 
    if(N11382) begin
      \nz.mem_5005_sv2v_reg  <= data_i[45];
    end 
    if(N11381) begin
      \nz.mem_5004_sv2v_reg  <= data_i[44];
    end 
    if(N11380) begin
      \nz.mem_5003_sv2v_reg  <= data_i[43];
    end 
    if(N11379) begin
      \nz.mem_5002_sv2v_reg  <= data_i[42];
    end 
    if(N11378) begin
      \nz.mem_5001_sv2v_reg  <= data_i[41];
    end 
    if(N11377) begin
      \nz.mem_5000_sv2v_reg  <= data_i[40];
    end 
    if(N11376) begin
      \nz.mem_4999_sv2v_reg  <= data_i[39];
    end 
    if(N11375) begin
      \nz.mem_4998_sv2v_reg  <= data_i[38];
    end 
    if(N11374) begin
      \nz.mem_4997_sv2v_reg  <= data_i[37];
    end 
    if(N11373) begin
      \nz.mem_4996_sv2v_reg  <= data_i[36];
    end 
    if(N11372) begin
      \nz.mem_4995_sv2v_reg  <= data_i[35];
    end 
    if(N11371) begin
      \nz.mem_4994_sv2v_reg  <= data_i[34];
    end 
    if(N11370) begin
      \nz.mem_4993_sv2v_reg  <= data_i[33];
    end 
    if(N11369) begin
      \nz.mem_4992_sv2v_reg  <= data_i[32];
    end 
    if(N11368) begin
      \nz.mem_4991_sv2v_reg  <= data_i[31];
    end 
    if(N11367) begin
      \nz.mem_4990_sv2v_reg  <= data_i[30];
    end 
    if(N11366) begin
      \nz.mem_4989_sv2v_reg  <= data_i[29];
    end 
    if(N11365) begin
      \nz.mem_4988_sv2v_reg  <= data_i[28];
    end 
    if(N11364) begin
      \nz.mem_4987_sv2v_reg  <= data_i[27];
    end 
    if(N11363) begin
      \nz.mem_4986_sv2v_reg  <= data_i[26];
    end 
    if(N11362) begin
      \nz.mem_4985_sv2v_reg  <= data_i[25];
    end 
    if(N11361) begin
      \nz.mem_4984_sv2v_reg  <= data_i[24];
    end 
    if(N11360) begin
      \nz.mem_4983_sv2v_reg  <= data_i[23];
    end 
    if(N11359) begin
      \nz.mem_4982_sv2v_reg  <= data_i[22];
    end 
    if(N11358) begin
      \nz.mem_4981_sv2v_reg  <= data_i[21];
    end 
    if(N11357) begin
      \nz.mem_4980_sv2v_reg  <= data_i[20];
    end 
    if(N11356) begin
      \nz.mem_4979_sv2v_reg  <= data_i[19];
    end 
    if(N11355) begin
      \nz.mem_4978_sv2v_reg  <= data_i[18];
    end 
    if(N11354) begin
      \nz.mem_4977_sv2v_reg  <= data_i[17];
    end 
    if(N11353) begin
      \nz.mem_4976_sv2v_reg  <= data_i[16];
    end 
    if(N11352) begin
      \nz.mem_4975_sv2v_reg  <= data_i[15];
    end 
    if(N11351) begin
      \nz.mem_4974_sv2v_reg  <= data_i[14];
    end 
    if(N11350) begin
      \nz.mem_4973_sv2v_reg  <= data_i[13];
    end 
    if(N11349) begin
      \nz.mem_4972_sv2v_reg  <= data_i[12];
    end 
    if(N11348) begin
      \nz.mem_4971_sv2v_reg  <= data_i[11];
    end 
    if(N11347) begin
      \nz.mem_4970_sv2v_reg  <= data_i[10];
    end 
    if(N11346) begin
      \nz.mem_4969_sv2v_reg  <= data_i[9];
    end 
    if(N11345) begin
      \nz.mem_4968_sv2v_reg  <= data_i[8];
    end 
    if(N11344) begin
      \nz.mem_4967_sv2v_reg  <= data_i[7];
    end 
    if(N11343) begin
      \nz.mem_4966_sv2v_reg  <= data_i[6];
    end 
    if(N11342) begin
      \nz.mem_4965_sv2v_reg  <= data_i[5];
    end 
    if(N11341) begin
      \nz.mem_4964_sv2v_reg  <= data_i[4];
    end 
    if(N11340) begin
      \nz.mem_4963_sv2v_reg  <= data_i[3];
    end 
    if(N11339) begin
      \nz.mem_4962_sv2v_reg  <= data_i[2];
    end 
    if(N11338) begin
      \nz.mem_4961_sv2v_reg  <= data_i[1];
    end 
    if(N11337) begin
      \nz.mem_4960_sv2v_reg  <= data_i[0];
    end 
    if(N11336) begin
      \nz.mem_4959_sv2v_reg  <= data_i[79];
    end 
    if(N11335) begin
      \nz.mem_4958_sv2v_reg  <= data_i[78];
    end 
    if(N11334) begin
      \nz.mem_4957_sv2v_reg  <= data_i[77];
    end 
    if(N11333) begin
      \nz.mem_4956_sv2v_reg  <= data_i[76];
    end 
    if(N11332) begin
      \nz.mem_4955_sv2v_reg  <= data_i[75];
    end 
    if(N11331) begin
      \nz.mem_4954_sv2v_reg  <= data_i[74];
    end 
    if(N11330) begin
      \nz.mem_4953_sv2v_reg  <= data_i[73];
    end 
    if(N11329) begin
      \nz.mem_4952_sv2v_reg  <= data_i[72];
    end 
    if(N11328) begin
      \nz.mem_4951_sv2v_reg  <= data_i[71];
    end 
    if(N11327) begin
      \nz.mem_4950_sv2v_reg  <= data_i[70];
    end 
    if(N11326) begin
      \nz.mem_4949_sv2v_reg  <= data_i[69];
    end 
    if(N11325) begin
      \nz.mem_4948_sv2v_reg  <= data_i[68];
    end 
    if(N11324) begin
      \nz.mem_4947_sv2v_reg  <= data_i[67];
    end 
    if(N11323) begin
      \nz.mem_4946_sv2v_reg  <= data_i[66];
    end 
    if(N11322) begin
      \nz.mem_4945_sv2v_reg  <= data_i[65];
    end 
    if(N11321) begin
      \nz.mem_4944_sv2v_reg  <= data_i[64];
    end 
    if(N11320) begin
      \nz.mem_4943_sv2v_reg  <= data_i[63];
    end 
    if(N11319) begin
      \nz.mem_4942_sv2v_reg  <= data_i[62];
    end 
    if(N11318) begin
      \nz.mem_4941_sv2v_reg  <= data_i[61];
    end 
    if(N11317) begin
      \nz.mem_4940_sv2v_reg  <= data_i[60];
    end 
    if(N11316) begin
      \nz.mem_4939_sv2v_reg  <= data_i[59];
    end 
    if(N11315) begin
      \nz.mem_4938_sv2v_reg  <= data_i[58];
    end 
    if(N11314) begin
      \nz.mem_4937_sv2v_reg  <= data_i[57];
    end 
    if(N11313) begin
      \nz.mem_4936_sv2v_reg  <= data_i[56];
    end 
    if(N11312) begin
      \nz.mem_4935_sv2v_reg  <= data_i[55];
    end 
    if(N11311) begin
      \nz.mem_4934_sv2v_reg  <= data_i[54];
    end 
    if(N11310) begin
      \nz.mem_4933_sv2v_reg  <= data_i[53];
    end 
    if(N11309) begin
      \nz.mem_4932_sv2v_reg  <= data_i[52];
    end 
    if(N11308) begin
      \nz.mem_4931_sv2v_reg  <= data_i[51];
    end 
    if(N11307) begin
      \nz.mem_4930_sv2v_reg  <= data_i[50];
    end 
    if(N11306) begin
      \nz.mem_4929_sv2v_reg  <= data_i[49];
    end 
    if(N11305) begin
      \nz.mem_4928_sv2v_reg  <= data_i[48];
    end 
    if(N11304) begin
      \nz.mem_4927_sv2v_reg  <= data_i[47];
    end 
    if(N11303) begin
      \nz.mem_4926_sv2v_reg  <= data_i[46];
    end 
    if(N11302) begin
      \nz.mem_4925_sv2v_reg  <= data_i[45];
    end 
    if(N11301) begin
      \nz.mem_4924_sv2v_reg  <= data_i[44];
    end 
    if(N11300) begin
      \nz.mem_4923_sv2v_reg  <= data_i[43];
    end 
    if(N11299) begin
      \nz.mem_4922_sv2v_reg  <= data_i[42];
    end 
    if(N11298) begin
      \nz.mem_4921_sv2v_reg  <= data_i[41];
    end 
    if(N11297) begin
      \nz.mem_4920_sv2v_reg  <= data_i[40];
    end 
    if(N11296) begin
      \nz.mem_4919_sv2v_reg  <= data_i[39];
    end 
    if(N11295) begin
      \nz.mem_4918_sv2v_reg  <= data_i[38];
    end 
    if(N11294) begin
      \nz.mem_4917_sv2v_reg  <= data_i[37];
    end 
    if(N11293) begin
      \nz.mem_4916_sv2v_reg  <= data_i[36];
    end 
    if(N11292) begin
      \nz.mem_4915_sv2v_reg  <= data_i[35];
    end 
    if(N11291) begin
      \nz.mem_4914_sv2v_reg  <= data_i[34];
    end 
    if(N11290) begin
      \nz.mem_4913_sv2v_reg  <= data_i[33];
    end 
    if(N11289) begin
      \nz.mem_4912_sv2v_reg  <= data_i[32];
    end 
    if(N11288) begin
      \nz.mem_4911_sv2v_reg  <= data_i[31];
    end 
    if(N11287) begin
      \nz.mem_4910_sv2v_reg  <= data_i[30];
    end 
    if(N11286) begin
      \nz.mem_4909_sv2v_reg  <= data_i[29];
    end 
    if(N11285) begin
      \nz.mem_4908_sv2v_reg  <= data_i[28];
    end 
    if(N11284) begin
      \nz.mem_4907_sv2v_reg  <= data_i[27];
    end 
    if(N11283) begin
      \nz.mem_4906_sv2v_reg  <= data_i[26];
    end 
    if(N11282) begin
      \nz.mem_4905_sv2v_reg  <= data_i[25];
    end 
    if(N11281) begin
      \nz.mem_4904_sv2v_reg  <= data_i[24];
    end 
    if(N11280) begin
      \nz.mem_4903_sv2v_reg  <= data_i[23];
    end 
    if(N11279) begin
      \nz.mem_4902_sv2v_reg  <= data_i[22];
    end 
    if(N11278) begin
      \nz.mem_4901_sv2v_reg  <= data_i[21];
    end 
    if(N11277) begin
      \nz.mem_4900_sv2v_reg  <= data_i[20];
    end 
    if(N11276) begin
      \nz.mem_4899_sv2v_reg  <= data_i[19];
    end 
    if(N11275) begin
      \nz.mem_4898_sv2v_reg  <= data_i[18];
    end 
    if(N11274) begin
      \nz.mem_4897_sv2v_reg  <= data_i[17];
    end 
    if(N11273) begin
      \nz.mem_4896_sv2v_reg  <= data_i[16];
    end 
    if(N11272) begin
      \nz.mem_4895_sv2v_reg  <= data_i[15];
    end 
    if(N11271) begin
      \nz.mem_4894_sv2v_reg  <= data_i[14];
    end 
    if(N11270) begin
      \nz.mem_4893_sv2v_reg  <= data_i[13];
    end 
    if(N11269) begin
      \nz.mem_4892_sv2v_reg  <= data_i[12];
    end 
    if(N11268) begin
      \nz.mem_4891_sv2v_reg  <= data_i[11];
    end 
    if(N11267) begin
      \nz.mem_4890_sv2v_reg  <= data_i[10];
    end 
    if(N11266) begin
      \nz.mem_4889_sv2v_reg  <= data_i[9];
    end 
    if(N11265) begin
      \nz.mem_4888_sv2v_reg  <= data_i[8];
    end 
    if(N11264) begin
      \nz.mem_4887_sv2v_reg  <= data_i[7];
    end 
    if(N11263) begin
      \nz.mem_4886_sv2v_reg  <= data_i[6];
    end 
    if(N11262) begin
      \nz.mem_4885_sv2v_reg  <= data_i[5];
    end 
    if(N11261) begin
      \nz.mem_4884_sv2v_reg  <= data_i[4];
    end 
    if(N11260) begin
      \nz.mem_4883_sv2v_reg  <= data_i[3];
    end 
    if(N11259) begin
      \nz.mem_4882_sv2v_reg  <= data_i[2];
    end 
    if(N11258) begin
      \nz.mem_4881_sv2v_reg  <= data_i[1];
    end 
    if(N11257) begin
      \nz.mem_4880_sv2v_reg  <= data_i[0];
    end 
    if(N11256) begin
      \nz.mem_4879_sv2v_reg  <= data_i[79];
    end 
    if(N11255) begin
      \nz.mem_4878_sv2v_reg  <= data_i[78];
    end 
    if(N11254) begin
      \nz.mem_4877_sv2v_reg  <= data_i[77];
    end 
    if(N11253) begin
      \nz.mem_4876_sv2v_reg  <= data_i[76];
    end 
    if(N11252) begin
      \nz.mem_4875_sv2v_reg  <= data_i[75];
    end 
    if(N11251) begin
      \nz.mem_4874_sv2v_reg  <= data_i[74];
    end 
    if(N11250) begin
      \nz.mem_4873_sv2v_reg  <= data_i[73];
    end 
    if(N11249) begin
      \nz.mem_4872_sv2v_reg  <= data_i[72];
    end 
    if(N11248) begin
      \nz.mem_4871_sv2v_reg  <= data_i[71];
    end 
    if(N11247) begin
      \nz.mem_4870_sv2v_reg  <= data_i[70];
    end 
    if(N11246) begin
      \nz.mem_4869_sv2v_reg  <= data_i[69];
    end 
    if(N11245) begin
      \nz.mem_4868_sv2v_reg  <= data_i[68];
    end 
    if(N11244) begin
      \nz.mem_4867_sv2v_reg  <= data_i[67];
    end 
    if(N11243) begin
      \nz.mem_4866_sv2v_reg  <= data_i[66];
    end 
    if(N11242) begin
      \nz.mem_4865_sv2v_reg  <= data_i[65];
    end 
    if(N11241) begin
      \nz.mem_4864_sv2v_reg  <= data_i[64];
    end 
    if(N11240) begin
      \nz.mem_4863_sv2v_reg  <= data_i[63];
    end 
    if(N11239) begin
      \nz.mem_4862_sv2v_reg  <= data_i[62];
    end 
    if(N11238) begin
      \nz.mem_4861_sv2v_reg  <= data_i[61];
    end 
    if(N11237) begin
      \nz.mem_4860_sv2v_reg  <= data_i[60];
    end 
    if(N11236) begin
      \nz.mem_4859_sv2v_reg  <= data_i[59];
    end 
    if(N11235) begin
      \nz.mem_4858_sv2v_reg  <= data_i[58];
    end 
    if(N11234) begin
      \nz.mem_4857_sv2v_reg  <= data_i[57];
    end 
    if(N11233) begin
      \nz.mem_4856_sv2v_reg  <= data_i[56];
    end 
    if(N11232) begin
      \nz.mem_4855_sv2v_reg  <= data_i[55];
    end 
    if(N11231) begin
      \nz.mem_4854_sv2v_reg  <= data_i[54];
    end 
    if(N11230) begin
      \nz.mem_4853_sv2v_reg  <= data_i[53];
    end 
    if(N11229) begin
      \nz.mem_4852_sv2v_reg  <= data_i[52];
    end 
    if(N11228) begin
      \nz.mem_4851_sv2v_reg  <= data_i[51];
    end 
    if(N11227) begin
      \nz.mem_4850_sv2v_reg  <= data_i[50];
    end 
    if(N11226) begin
      \nz.mem_4849_sv2v_reg  <= data_i[49];
    end 
    if(N11225) begin
      \nz.mem_4848_sv2v_reg  <= data_i[48];
    end 
    if(N11224) begin
      \nz.mem_4847_sv2v_reg  <= data_i[47];
    end 
    if(N11223) begin
      \nz.mem_4846_sv2v_reg  <= data_i[46];
    end 
    if(N11222) begin
      \nz.mem_4845_sv2v_reg  <= data_i[45];
    end 
    if(N11221) begin
      \nz.mem_4844_sv2v_reg  <= data_i[44];
    end 
    if(N11220) begin
      \nz.mem_4843_sv2v_reg  <= data_i[43];
    end 
    if(N11219) begin
      \nz.mem_4842_sv2v_reg  <= data_i[42];
    end 
    if(N11218) begin
      \nz.mem_4841_sv2v_reg  <= data_i[41];
    end 
    if(N11217) begin
      \nz.mem_4840_sv2v_reg  <= data_i[40];
    end 
    if(N11216) begin
      \nz.mem_4839_sv2v_reg  <= data_i[39];
    end 
    if(N11215) begin
      \nz.mem_4838_sv2v_reg  <= data_i[38];
    end 
    if(N11214) begin
      \nz.mem_4837_sv2v_reg  <= data_i[37];
    end 
    if(N11213) begin
      \nz.mem_4836_sv2v_reg  <= data_i[36];
    end 
    if(N11212) begin
      \nz.mem_4835_sv2v_reg  <= data_i[35];
    end 
    if(N11211) begin
      \nz.mem_4834_sv2v_reg  <= data_i[34];
    end 
    if(N11210) begin
      \nz.mem_4833_sv2v_reg  <= data_i[33];
    end 
    if(N11209) begin
      \nz.mem_4832_sv2v_reg  <= data_i[32];
    end 
    if(N11208) begin
      \nz.mem_4831_sv2v_reg  <= data_i[31];
    end 
    if(N11207) begin
      \nz.mem_4830_sv2v_reg  <= data_i[30];
    end 
    if(N11206) begin
      \nz.mem_4829_sv2v_reg  <= data_i[29];
    end 
    if(N11205) begin
      \nz.mem_4828_sv2v_reg  <= data_i[28];
    end 
    if(N11204) begin
      \nz.mem_4827_sv2v_reg  <= data_i[27];
    end 
    if(N11203) begin
      \nz.mem_4826_sv2v_reg  <= data_i[26];
    end 
    if(N11202) begin
      \nz.mem_4825_sv2v_reg  <= data_i[25];
    end 
    if(N11201) begin
      \nz.mem_4824_sv2v_reg  <= data_i[24];
    end 
    if(N11200) begin
      \nz.mem_4823_sv2v_reg  <= data_i[23];
    end 
    if(N11199) begin
      \nz.mem_4822_sv2v_reg  <= data_i[22];
    end 
    if(N11198) begin
      \nz.mem_4821_sv2v_reg  <= data_i[21];
    end 
    if(N11197) begin
      \nz.mem_4820_sv2v_reg  <= data_i[20];
    end 
    if(N11196) begin
      \nz.mem_4819_sv2v_reg  <= data_i[19];
    end 
    if(N11195) begin
      \nz.mem_4818_sv2v_reg  <= data_i[18];
    end 
    if(N11194) begin
      \nz.mem_4817_sv2v_reg  <= data_i[17];
    end 
    if(N11193) begin
      \nz.mem_4816_sv2v_reg  <= data_i[16];
    end 
    if(N11192) begin
      \nz.mem_4815_sv2v_reg  <= data_i[15];
    end 
    if(N11191) begin
      \nz.mem_4814_sv2v_reg  <= data_i[14];
    end 
    if(N11190) begin
      \nz.mem_4813_sv2v_reg  <= data_i[13];
    end 
    if(N11189) begin
      \nz.mem_4812_sv2v_reg  <= data_i[12];
    end 
    if(N11188) begin
      \nz.mem_4811_sv2v_reg  <= data_i[11];
    end 
    if(N11187) begin
      \nz.mem_4810_sv2v_reg  <= data_i[10];
    end 
    if(N11186) begin
      \nz.mem_4809_sv2v_reg  <= data_i[9];
    end 
    if(N11185) begin
      \nz.mem_4808_sv2v_reg  <= data_i[8];
    end 
    if(N11184) begin
      \nz.mem_4807_sv2v_reg  <= data_i[7];
    end 
    if(N11183) begin
      \nz.mem_4806_sv2v_reg  <= data_i[6];
    end 
    if(N11182) begin
      \nz.mem_4805_sv2v_reg  <= data_i[5];
    end 
    if(N11181) begin
      \nz.mem_4804_sv2v_reg  <= data_i[4];
    end 
    if(N11180) begin
      \nz.mem_4803_sv2v_reg  <= data_i[3];
    end 
    if(N11179) begin
      \nz.mem_4802_sv2v_reg  <= data_i[2];
    end 
    if(N11178) begin
      \nz.mem_4801_sv2v_reg  <= data_i[1];
    end 
    if(N11177) begin
      \nz.mem_4800_sv2v_reg  <= data_i[0];
    end 
    if(N11176) begin
      \nz.mem_4799_sv2v_reg  <= data_i[79];
    end 
    if(N11175) begin
      \nz.mem_4798_sv2v_reg  <= data_i[78];
    end 
    if(N11174) begin
      \nz.mem_4797_sv2v_reg  <= data_i[77];
    end 
    if(N11173) begin
      \nz.mem_4796_sv2v_reg  <= data_i[76];
    end 
    if(N11172) begin
      \nz.mem_4795_sv2v_reg  <= data_i[75];
    end 
    if(N11171) begin
      \nz.mem_4794_sv2v_reg  <= data_i[74];
    end 
    if(N11170) begin
      \nz.mem_4793_sv2v_reg  <= data_i[73];
    end 
    if(N11169) begin
      \nz.mem_4792_sv2v_reg  <= data_i[72];
    end 
    if(N11168) begin
      \nz.mem_4791_sv2v_reg  <= data_i[71];
    end 
    if(N11167) begin
      \nz.mem_4790_sv2v_reg  <= data_i[70];
    end 
    if(N11166) begin
      \nz.mem_4789_sv2v_reg  <= data_i[69];
    end 
    if(N11165) begin
      \nz.mem_4788_sv2v_reg  <= data_i[68];
    end 
    if(N11164) begin
      \nz.mem_4787_sv2v_reg  <= data_i[67];
    end 
    if(N11163) begin
      \nz.mem_4786_sv2v_reg  <= data_i[66];
    end 
    if(N11162) begin
      \nz.mem_4785_sv2v_reg  <= data_i[65];
    end 
    if(N11161) begin
      \nz.mem_4784_sv2v_reg  <= data_i[64];
    end 
    if(N11160) begin
      \nz.mem_4783_sv2v_reg  <= data_i[63];
    end 
    if(N11159) begin
      \nz.mem_4782_sv2v_reg  <= data_i[62];
    end 
    if(N11158) begin
      \nz.mem_4781_sv2v_reg  <= data_i[61];
    end 
    if(N11157) begin
      \nz.mem_4780_sv2v_reg  <= data_i[60];
    end 
    if(N11156) begin
      \nz.mem_4779_sv2v_reg  <= data_i[59];
    end 
    if(N11155) begin
      \nz.mem_4778_sv2v_reg  <= data_i[58];
    end 
    if(N11154) begin
      \nz.mem_4777_sv2v_reg  <= data_i[57];
    end 
    if(N11153) begin
      \nz.mem_4776_sv2v_reg  <= data_i[56];
    end 
    if(N11152) begin
      \nz.mem_4775_sv2v_reg  <= data_i[55];
    end 
    if(N11151) begin
      \nz.mem_4774_sv2v_reg  <= data_i[54];
    end 
    if(N11150) begin
      \nz.mem_4773_sv2v_reg  <= data_i[53];
    end 
    if(N11149) begin
      \nz.mem_4772_sv2v_reg  <= data_i[52];
    end 
    if(N11148) begin
      \nz.mem_4771_sv2v_reg  <= data_i[51];
    end 
    if(N11147) begin
      \nz.mem_4770_sv2v_reg  <= data_i[50];
    end 
    if(N11146) begin
      \nz.mem_4769_sv2v_reg  <= data_i[49];
    end 
    if(N11145) begin
      \nz.mem_4768_sv2v_reg  <= data_i[48];
    end 
    if(N11144) begin
      \nz.mem_4767_sv2v_reg  <= data_i[47];
    end 
    if(N11143) begin
      \nz.mem_4766_sv2v_reg  <= data_i[46];
    end 
    if(N11142) begin
      \nz.mem_4765_sv2v_reg  <= data_i[45];
    end 
    if(N11141) begin
      \nz.mem_4764_sv2v_reg  <= data_i[44];
    end 
    if(N11140) begin
      \nz.mem_4763_sv2v_reg  <= data_i[43];
    end 
    if(N11139) begin
      \nz.mem_4762_sv2v_reg  <= data_i[42];
    end 
    if(N11138) begin
      \nz.mem_4761_sv2v_reg  <= data_i[41];
    end 
    if(N11137) begin
      \nz.mem_4760_sv2v_reg  <= data_i[40];
    end 
    if(N11136) begin
      \nz.mem_4759_sv2v_reg  <= data_i[39];
    end 
    if(N11135) begin
      \nz.mem_4758_sv2v_reg  <= data_i[38];
    end 
    if(N11134) begin
      \nz.mem_4757_sv2v_reg  <= data_i[37];
    end 
    if(N11133) begin
      \nz.mem_4756_sv2v_reg  <= data_i[36];
    end 
    if(N11132) begin
      \nz.mem_4755_sv2v_reg  <= data_i[35];
    end 
    if(N11131) begin
      \nz.mem_4754_sv2v_reg  <= data_i[34];
    end 
    if(N11130) begin
      \nz.mem_4753_sv2v_reg  <= data_i[33];
    end 
    if(N11129) begin
      \nz.mem_4752_sv2v_reg  <= data_i[32];
    end 
    if(N11128) begin
      \nz.mem_4751_sv2v_reg  <= data_i[31];
    end 
    if(N11127) begin
      \nz.mem_4750_sv2v_reg  <= data_i[30];
    end 
    if(N11126) begin
      \nz.mem_4749_sv2v_reg  <= data_i[29];
    end 
    if(N11125) begin
      \nz.mem_4748_sv2v_reg  <= data_i[28];
    end 
    if(N11124) begin
      \nz.mem_4747_sv2v_reg  <= data_i[27];
    end 
    if(N11123) begin
      \nz.mem_4746_sv2v_reg  <= data_i[26];
    end 
    if(N11122) begin
      \nz.mem_4745_sv2v_reg  <= data_i[25];
    end 
    if(N11121) begin
      \nz.mem_4744_sv2v_reg  <= data_i[24];
    end 
    if(N11120) begin
      \nz.mem_4743_sv2v_reg  <= data_i[23];
    end 
    if(N11119) begin
      \nz.mem_4742_sv2v_reg  <= data_i[22];
    end 
    if(N11118) begin
      \nz.mem_4741_sv2v_reg  <= data_i[21];
    end 
    if(N11117) begin
      \nz.mem_4740_sv2v_reg  <= data_i[20];
    end 
    if(N11116) begin
      \nz.mem_4739_sv2v_reg  <= data_i[19];
    end 
    if(N11115) begin
      \nz.mem_4738_sv2v_reg  <= data_i[18];
    end 
    if(N11114) begin
      \nz.mem_4737_sv2v_reg  <= data_i[17];
    end 
    if(N11113) begin
      \nz.mem_4736_sv2v_reg  <= data_i[16];
    end 
    if(N11112) begin
      \nz.mem_4735_sv2v_reg  <= data_i[15];
    end 
    if(N11111) begin
      \nz.mem_4734_sv2v_reg  <= data_i[14];
    end 
    if(N11110) begin
      \nz.mem_4733_sv2v_reg  <= data_i[13];
    end 
    if(N11109) begin
      \nz.mem_4732_sv2v_reg  <= data_i[12];
    end 
    if(N11108) begin
      \nz.mem_4731_sv2v_reg  <= data_i[11];
    end 
    if(N11107) begin
      \nz.mem_4730_sv2v_reg  <= data_i[10];
    end 
    if(N11106) begin
      \nz.mem_4729_sv2v_reg  <= data_i[9];
    end 
    if(N11105) begin
      \nz.mem_4728_sv2v_reg  <= data_i[8];
    end 
    if(N11104) begin
      \nz.mem_4727_sv2v_reg  <= data_i[7];
    end 
    if(N11103) begin
      \nz.mem_4726_sv2v_reg  <= data_i[6];
    end 
    if(N11102) begin
      \nz.mem_4725_sv2v_reg  <= data_i[5];
    end 
    if(N11101) begin
      \nz.mem_4724_sv2v_reg  <= data_i[4];
    end 
    if(N11100) begin
      \nz.mem_4723_sv2v_reg  <= data_i[3];
    end 
    if(N11099) begin
      \nz.mem_4722_sv2v_reg  <= data_i[2];
    end 
    if(N11098) begin
      \nz.mem_4721_sv2v_reg  <= data_i[1];
    end 
    if(N11097) begin
      \nz.mem_4720_sv2v_reg  <= data_i[0];
    end 
    if(N11096) begin
      \nz.mem_4719_sv2v_reg  <= data_i[79];
    end 
    if(N11095) begin
      \nz.mem_4718_sv2v_reg  <= data_i[78];
    end 
    if(N11094) begin
      \nz.mem_4717_sv2v_reg  <= data_i[77];
    end 
    if(N11093) begin
      \nz.mem_4716_sv2v_reg  <= data_i[76];
    end 
    if(N11092) begin
      \nz.mem_4715_sv2v_reg  <= data_i[75];
    end 
    if(N11091) begin
      \nz.mem_4714_sv2v_reg  <= data_i[74];
    end 
    if(N11090) begin
      \nz.mem_4713_sv2v_reg  <= data_i[73];
    end 
    if(N11089) begin
      \nz.mem_4712_sv2v_reg  <= data_i[72];
    end 
    if(N11088) begin
      \nz.mem_4711_sv2v_reg  <= data_i[71];
    end 
    if(N11087) begin
      \nz.mem_4710_sv2v_reg  <= data_i[70];
    end 
    if(N11086) begin
      \nz.mem_4709_sv2v_reg  <= data_i[69];
    end 
    if(N11085) begin
      \nz.mem_4708_sv2v_reg  <= data_i[68];
    end 
    if(N11084) begin
      \nz.mem_4707_sv2v_reg  <= data_i[67];
    end 
    if(N11083) begin
      \nz.mem_4706_sv2v_reg  <= data_i[66];
    end 
    if(N11082) begin
      \nz.mem_4705_sv2v_reg  <= data_i[65];
    end 
    if(N11081) begin
      \nz.mem_4704_sv2v_reg  <= data_i[64];
    end 
    if(N11080) begin
      \nz.mem_4703_sv2v_reg  <= data_i[63];
    end 
    if(N11079) begin
      \nz.mem_4702_sv2v_reg  <= data_i[62];
    end 
    if(N11078) begin
      \nz.mem_4701_sv2v_reg  <= data_i[61];
    end 
    if(N11077) begin
      \nz.mem_4700_sv2v_reg  <= data_i[60];
    end 
    if(N11076) begin
      \nz.mem_4699_sv2v_reg  <= data_i[59];
    end 
    if(N11075) begin
      \nz.mem_4698_sv2v_reg  <= data_i[58];
    end 
    if(N11074) begin
      \nz.mem_4697_sv2v_reg  <= data_i[57];
    end 
    if(N11073) begin
      \nz.mem_4696_sv2v_reg  <= data_i[56];
    end 
    if(N11072) begin
      \nz.mem_4695_sv2v_reg  <= data_i[55];
    end 
    if(N11071) begin
      \nz.mem_4694_sv2v_reg  <= data_i[54];
    end 
    if(N11070) begin
      \nz.mem_4693_sv2v_reg  <= data_i[53];
    end 
    if(N11069) begin
      \nz.mem_4692_sv2v_reg  <= data_i[52];
    end 
    if(N11068) begin
      \nz.mem_4691_sv2v_reg  <= data_i[51];
    end 
    if(N11067) begin
      \nz.mem_4690_sv2v_reg  <= data_i[50];
    end 
    if(N11066) begin
      \nz.mem_4689_sv2v_reg  <= data_i[49];
    end 
    if(N11065) begin
      \nz.mem_4688_sv2v_reg  <= data_i[48];
    end 
    if(N11064) begin
      \nz.mem_4687_sv2v_reg  <= data_i[47];
    end 
    if(N11063) begin
      \nz.mem_4686_sv2v_reg  <= data_i[46];
    end 
    if(N11062) begin
      \nz.mem_4685_sv2v_reg  <= data_i[45];
    end 
    if(N11061) begin
      \nz.mem_4684_sv2v_reg  <= data_i[44];
    end 
    if(N11060) begin
      \nz.mem_4683_sv2v_reg  <= data_i[43];
    end 
    if(N11059) begin
      \nz.mem_4682_sv2v_reg  <= data_i[42];
    end 
    if(N11058) begin
      \nz.mem_4681_sv2v_reg  <= data_i[41];
    end 
    if(N11057) begin
      \nz.mem_4680_sv2v_reg  <= data_i[40];
    end 
    if(N11056) begin
      \nz.mem_4679_sv2v_reg  <= data_i[39];
    end 
    if(N11055) begin
      \nz.mem_4678_sv2v_reg  <= data_i[38];
    end 
    if(N11054) begin
      \nz.mem_4677_sv2v_reg  <= data_i[37];
    end 
    if(N11053) begin
      \nz.mem_4676_sv2v_reg  <= data_i[36];
    end 
    if(N11052) begin
      \nz.mem_4675_sv2v_reg  <= data_i[35];
    end 
    if(N11051) begin
      \nz.mem_4674_sv2v_reg  <= data_i[34];
    end 
    if(N11050) begin
      \nz.mem_4673_sv2v_reg  <= data_i[33];
    end 
    if(N11049) begin
      \nz.mem_4672_sv2v_reg  <= data_i[32];
    end 
    if(N11048) begin
      \nz.mem_4671_sv2v_reg  <= data_i[31];
    end 
    if(N11047) begin
      \nz.mem_4670_sv2v_reg  <= data_i[30];
    end 
    if(N11046) begin
      \nz.mem_4669_sv2v_reg  <= data_i[29];
    end 
    if(N11045) begin
      \nz.mem_4668_sv2v_reg  <= data_i[28];
    end 
    if(N11044) begin
      \nz.mem_4667_sv2v_reg  <= data_i[27];
    end 
    if(N11043) begin
      \nz.mem_4666_sv2v_reg  <= data_i[26];
    end 
    if(N11042) begin
      \nz.mem_4665_sv2v_reg  <= data_i[25];
    end 
    if(N11041) begin
      \nz.mem_4664_sv2v_reg  <= data_i[24];
    end 
    if(N11040) begin
      \nz.mem_4663_sv2v_reg  <= data_i[23];
    end 
    if(N11039) begin
      \nz.mem_4662_sv2v_reg  <= data_i[22];
    end 
    if(N11038) begin
      \nz.mem_4661_sv2v_reg  <= data_i[21];
    end 
    if(N11037) begin
      \nz.mem_4660_sv2v_reg  <= data_i[20];
    end 
    if(N11036) begin
      \nz.mem_4659_sv2v_reg  <= data_i[19];
    end 
    if(N11035) begin
      \nz.mem_4658_sv2v_reg  <= data_i[18];
    end 
    if(N11034) begin
      \nz.mem_4657_sv2v_reg  <= data_i[17];
    end 
    if(N11033) begin
      \nz.mem_4656_sv2v_reg  <= data_i[16];
    end 
    if(N11032) begin
      \nz.mem_4655_sv2v_reg  <= data_i[15];
    end 
    if(N11031) begin
      \nz.mem_4654_sv2v_reg  <= data_i[14];
    end 
    if(N11030) begin
      \nz.mem_4653_sv2v_reg  <= data_i[13];
    end 
    if(N11029) begin
      \nz.mem_4652_sv2v_reg  <= data_i[12];
    end 
    if(N11028) begin
      \nz.mem_4651_sv2v_reg  <= data_i[11];
    end 
    if(N11027) begin
      \nz.mem_4650_sv2v_reg  <= data_i[10];
    end 
    if(N11026) begin
      \nz.mem_4649_sv2v_reg  <= data_i[9];
    end 
    if(N11025) begin
      \nz.mem_4648_sv2v_reg  <= data_i[8];
    end 
    if(N11024) begin
      \nz.mem_4647_sv2v_reg  <= data_i[7];
    end 
    if(N11023) begin
      \nz.mem_4646_sv2v_reg  <= data_i[6];
    end 
    if(N11022) begin
      \nz.mem_4645_sv2v_reg  <= data_i[5];
    end 
    if(N11021) begin
      \nz.mem_4644_sv2v_reg  <= data_i[4];
    end 
    if(N11020) begin
      \nz.mem_4643_sv2v_reg  <= data_i[3];
    end 
    if(N11019) begin
      \nz.mem_4642_sv2v_reg  <= data_i[2];
    end 
    if(N11018) begin
      \nz.mem_4641_sv2v_reg  <= data_i[1];
    end 
    if(N11017) begin
      \nz.mem_4640_sv2v_reg  <= data_i[0];
    end 
    if(N11016) begin
      \nz.mem_4639_sv2v_reg  <= data_i[79];
    end 
    if(N11015) begin
      \nz.mem_4638_sv2v_reg  <= data_i[78];
    end 
    if(N11014) begin
      \nz.mem_4637_sv2v_reg  <= data_i[77];
    end 
    if(N11013) begin
      \nz.mem_4636_sv2v_reg  <= data_i[76];
    end 
    if(N11012) begin
      \nz.mem_4635_sv2v_reg  <= data_i[75];
    end 
    if(N11011) begin
      \nz.mem_4634_sv2v_reg  <= data_i[74];
    end 
    if(N11010) begin
      \nz.mem_4633_sv2v_reg  <= data_i[73];
    end 
    if(N11009) begin
      \nz.mem_4632_sv2v_reg  <= data_i[72];
    end 
    if(N11008) begin
      \nz.mem_4631_sv2v_reg  <= data_i[71];
    end 
    if(N11007) begin
      \nz.mem_4630_sv2v_reg  <= data_i[70];
    end 
    if(N11006) begin
      \nz.mem_4629_sv2v_reg  <= data_i[69];
    end 
    if(N11005) begin
      \nz.mem_4628_sv2v_reg  <= data_i[68];
    end 
    if(N11004) begin
      \nz.mem_4627_sv2v_reg  <= data_i[67];
    end 
    if(N11003) begin
      \nz.mem_4626_sv2v_reg  <= data_i[66];
    end 
    if(N11002) begin
      \nz.mem_4625_sv2v_reg  <= data_i[65];
    end 
    if(N11001) begin
      \nz.mem_4624_sv2v_reg  <= data_i[64];
    end 
    if(N11000) begin
      \nz.mem_4623_sv2v_reg  <= data_i[63];
    end 
    if(N10999) begin
      \nz.mem_4622_sv2v_reg  <= data_i[62];
    end 
    if(N10998) begin
      \nz.mem_4621_sv2v_reg  <= data_i[61];
    end 
    if(N10997) begin
      \nz.mem_4620_sv2v_reg  <= data_i[60];
    end 
    if(N10996) begin
      \nz.mem_4619_sv2v_reg  <= data_i[59];
    end 
    if(N10995) begin
      \nz.mem_4618_sv2v_reg  <= data_i[58];
    end 
    if(N10994) begin
      \nz.mem_4617_sv2v_reg  <= data_i[57];
    end 
    if(N10993) begin
      \nz.mem_4616_sv2v_reg  <= data_i[56];
    end 
    if(N10992) begin
      \nz.mem_4615_sv2v_reg  <= data_i[55];
    end 
    if(N10991) begin
      \nz.mem_4614_sv2v_reg  <= data_i[54];
    end 
    if(N10990) begin
      \nz.mem_4613_sv2v_reg  <= data_i[53];
    end 
    if(N10989) begin
      \nz.mem_4612_sv2v_reg  <= data_i[52];
    end 
    if(N10988) begin
      \nz.mem_4611_sv2v_reg  <= data_i[51];
    end 
    if(N10987) begin
      \nz.mem_4610_sv2v_reg  <= data_i[50];
    end 
    if(N10986) begin
      \nz.mem_4609_sv2v_reg  <= data_i[49];
    end 
    if(N10985) begin
      \nz.mem_4608_sv2v_reg  <= data_i[48];
    end 
    if(N10984) begin
      \nz.mem_4607_sv2v_reg  <= data_i[47];
    end 
    if(N10983) begin
      \nz.mem_4606_sv2v_reg  <= data_i[46];
    end 
    if(N10982) begin
      \nz.mem_4605_sv2v_reg  <= data_i[45];
    end 
    if(N10981) begin
      \nz.mem_4604_sv2v_reg  <= data_i[44];
    end 
    if(N10980) begin
      \nz.mem_4603_sv2v_reg  <= data_i[43];
    end 
    if(N10979) begin
      \nz.mem_4602_sv2v_reg  <= data_i[42];
    end 
    if(N10978) begin
      \nz.mem_4601_sv2v_reg  <= data_i[41];
    end 
    if(N10977) begin
      \nz.mem_4600_sv2v_reg  <= data_i[40];
    end 
    if(N10976) begin
      \nz.mem_4599_sv2v_reg  <= data_i[39];
    end 
    if(N10975) begin
      \nz.mem_4598_sv2v_reg  <= data_i[38];
    end 
    if(N10974) begin
      \nz.mem_4597_sv2v_reg  <= data_i[37];
    end 
    if(N10973) begin
      \nz.mem_4596_sv2v_reg  <= data_i[36];
    end 
    if(N10972) begin
      \nz.mem_4595_sv2v_reg  <= data_i[35];
    end 
    if(N10971) begin
      \nz.mem_4594_sv2v_reg  <= data_i[34];
    end 
    if(N10970) begin
      \nz.mem_4593_sv2v_reg  <= data_i[33];
    end 
    if(N10969) begin
      \nz.mem_4592_sv2v_reg  <= data_i[32];
    end 
    if(N10968) begin
      \nz.mem_4591_sv2v_reg  <= data_i[31];
    end 
    if(N10967) begin
      \nz.mem_4590_sv2v_reg  <= data_i[30];
    end 
    if(N10966) begin
      \nz.mem_4589_sv2v_reg  <= data_i[29];
    end 
    if(N10965) begin
      \nz.mem_4588_sv2v_reg  <= data_i[28];
    end 
    if(N10964) begin
      \nz.mem_4587_sv2v_reg  <= data_i[27];
    end 
    if(N10963) begin
      \nz.mem_4586_sv2v_reg  <= data_i[26];
    end 
    if(N10962) begin
      \nz.mem_4585_sv2v_reg  <= data_i[25];
    end 
    if(N10961) begin
      \nz.mem_4584_sv2v_reg  <= data_i[24];
    end 
    if(N10960) begin
      \nz.mem_4583_sv2v_reg  <= data_i[23];
    end 
    if(N10959) begin
      \nz.mem_4582_sv2v_reg  <= data_i[22];
    end 
    if(N10958) begin
      \nz.mem_4581_sv2v_reg  <= data_i[21];
    end 
    if(N10957) begin
      \nz.mem_4580_sv2v_reg  <= data_i[20];
    end 
    if(N10956) begin
      \nz.mem_4579_sv2v_reg  <= data_i[19];
    end 
    if(N10955) begin
      \nz.mem_4578_sv2v_reg  <= data_i[18];
    end 
    if(N10954) begin
      \nz.mem_4577_sv2v_reg  <= data_i[17];
    end 
    if(N10953) begin
      \nz.mem_4576_sv2v_reg  <= data_i[16];
    end 
    if(N10952) begin
      \nz.mem_4575_sv2v_reg  <= data_i[15];
    end 
    if(N10951) begin
      \nz.mem_4574_sv2v_reg  <= data_i[14];
    end 
    if(N10950) begin
      \nz.mem_4573_sv2v_reg  <= data_i[13];
    end 
    if(N10949) begin
      \nz.mem_4572_sv2v_reg  <= data_i[12];
    end 
    if(N10948) begin
      \nz.mem_4571_sv2v_reg  <= data_i[11];
    end 
    if(N10947) begin
      \nz.mem_4570_sv2v_reg  <= data_i[10];
    end 
    if(N10946) begin
      \nz.mem_4569_sv2v_reg  <= data_i[9];
    end 
    if(N10945) begin
      \nz.mem_4568_sv2v_reg  <= data_i[8];
    end 
    if(N10944) begin
      \nz.mem_4567_sv2v_reg  <= data_i[7];
    end 
    if(N10943) begin
      \nz.mem_4566_sv2v_reg  <= data_i[6];
    end 
    if(N10942) begin
      \nz.mem_4565_sv2v_reg  <= data_i[5];
    end 
    if(N10941) begin
      \nz.mem_4564_sv2v_reg  <= data_i[4];
    end 
    if(N10940) begin
      \nz.mem_4563_sv2v_reg  <= data_i[3];
    end 
    if(N10939) begin
      \nz.mem_4562_sv2v_reg  <= data_i[2];
    end 
    if(N10938) begin
      \nz.mem_4561_sv2v_reg  <= data_i[1];
    end 
    if(N10937) begin
      \nz.mem_4560_sv2v_reg  <= data_i[0];
    end 
    if(N10936) begin
      \nz.mem_4559_sv2v_reg  <= data_i[79];
    end 
    if(N10935) begin
      \nz.mem_4558_sv2v_reg  <= data_i[78];
    end 
    if(N10934) begin
      \nz.mem_4557_sv2v_reg  <= data_i[77];
    end 
    if(N10933) begin
      \nz.mem_4556_sv2v_reg  <= data_i[76];
    end 
    if(N10932) begin
      \nz.mem_4555_sv2v_reg  <= data_i[75];
    end 
    if(N10931) begin
      \nz.mem_4554_sv2v_reg  <= data_i[74];
    end 
    if(N10930) begin
      \nz.mem_4553_sv2v_reg  <= data_i[73];
    end 
    if(N10929) begin
      \nz.mem_4552_sv2v_reg  <= data_i[72];
    end 
    if(N10928) begin
      \nz.mem_4551_sv2v_reg  <= data_i[71];
    end 
    if(N10927) begin
      \nz.mem_4550_sv2v_reg  <= data_i[70];
    end 
    if(N10926) begin
      \nz.mem_4549_sv2v_reg  <= data_i[69];
    end 
    if(N10925) begin
      \nz.mem_4548_sv2v_reg  <= data_i[68];
    end 
    if(N10924) begin
      \nz.mem_4547_sv2v_reg  <= data_i[67];
    end 
    if(N10923) begin
      \nz.mem_4546_sv2v_reg  <= data_i[66];
    end 
    if(N10922) begin
      \nz.mem_4545_sv2v_reg  <= data_i[65];
    end 
    if(N10921) begin
      \nz.mem_4544_sv2v_reg  <= data_i[64];
    end 
    if(N10920) begin
      \nz.mem_4543_sv2v_reg  <= data_i[63];
    end 
    if(N10919) begin
      \nz.mem_4542_sv2v_reg  <= data_i[62];
    end 
    if(N10918) begin
      \nz.mem_4541_sv2v_reg  <= data_i[61];
    end 
    if(N10917) begin
      \nz.mem_4540_sv2v_reg  <= data_i[60];
    end 
    if(N10916) begin
      \nz.mem_4539_sv2v_reg  <= data_i[59];
    end 
    if(N10915) begin
      \nz.mem_4538_sv2v_reg  <= data_i[58];
    end 
    if(N10914) begin
      \nz.mem_4537_sv2v_reg  <= data_i[57];
    end 
    if(N10913) begin
      \nz.mem_4536_sv2v_reg  <= data_i[56];
    end 
    if(N10912) begin
      \nz.mem_4535_sv2v_reg  <= data_i[55];
    end 
    if(N10911) begin
      \nz.mem_4534_sv2v_reg  <= data_i[54];
    end 
    if(N10910) begin
      \nz.mem_4533_sv2v_reg  <= data_i[53];
    end 
    if(N10909) begin
      \nz.mem_4532_sv2v_reg  <= data_i[52];
    end 
    if(N10908) begin
      \nz.mem_4531_sv2v_reg  <= data_i[51];
    end 
    if(N10907) begin
      \nz.mem_4530_sv2v_reg  <= data_i[50];
    end 
    if(N10906) begin
      \nz.mem_4529_sv2v_reg  <= data_i[49];
    end 
    if(N10905) begin
      \nz.mem_4528_sv2v_reg  <= data_i[48];
    end 
    if(N10904) begin
      \nz.mem_4527_sv2v_reg  <= data_i[47];
    end 
    if(N10903) begin
      \nz.mem_4526_sv2v_reg  <= data_i[46];
    end 
    if(N10902) begin
      \nz.mem_4525_sv2v_reg  <= data_i[45];
    end 
    if(N10901) begin
      \nz.mem_4524_sv2v_reg  <= data_i[44];
    end 
    if(N10900) begin
      \nz.mem_4523_sv2v_reg  <= data_i[43];
    end 
    if(N10899) begin
      \nz.mem_4522_sv2v_reg  <= data_i[42];
    end 
    if(N10898) begin
      \nz.mem_4521_sv2v_reg  <= data_i[41];
    end 
    if(N10897) begin
      \nz.mem_4520_sv2v_reg  <= data_i[40];
    end 
    if(N10896) begin
      \nz.mem_4519_sv2v_reg  <= data_i[39];
    end 
    if(N10895) begin
      \nz.mem_4518_sv2v_reg  <= data_i[38];
    end 
    if(N10894) begin
      \nz.mem_4517_sv2v_reg  <= data_i[37];
    end 
    if(N10893) begin
      \nz.mem_4516_sv2v_reg  <= data_i[36];
    end 
    if(N10892) begin
      \nz.mem_4515_sv2v_reg  <= data_i[35];
    end 
    if(N10891) begin
      \nz.mem_4514_sv2v_reg  <= data_i[34];
    end 
    if(N10890) begin
      \nz.mem_4513_sv2v_reg  <= data_i[33];
    end 
    if(N10889) begin
      \nz.mem_4512_sv2v_reg  <= data_i[32];
    end 
    if(N10888) begin
      \nz.mem_4511_sv2v_reg  <= data_i[31];
    end 
    if(N10887) begin
      \nz.mem_4510_sv2v_reg  <= data_i[30];
    end 
    if(N10886) begin
      \nz.mem_4509_sv2v_reg  <= data_i[29];
    end 
    if(N10885) begin
      \nz.mem_4508_sv2v_reg  <= data_i[28];
    end 
    if(N10884) begin
      \nz.mem_4507_sv2v_reg  <= data_i[27];
    end 
    if(N10883) begin
      \nz.mem_4506_sv2v_reg  <= data_i[26];
    end 
    if(N10882) begin
      \nz.mem_4505_sv2v_reg  <= data_i[25];
    end 
    if(N10881) begin
      \nz.mem_4504_sv2v_reg  <= data_i[24];
    end 
    if(N10880) begin
      \nz.mem_4503_sv2v_reg  <= data_i[23];
    end 
    if(N10879) begin
      \nz.mem_4502_sv2v_reg  <= data_i[22];
    end 
    if(N10878) begin
      \nz.mem_4501_sv2v_reg  <= data_i[21];
    end 
    if(N10877) begin
      \nz.mem_4500_sv2v_reg  <= data_i[20];
    end 
    if(N10876) begin
      \nz.mem_4499_sv2v_reg  <= data_i[19];
    end 
    if(N10875) begin
      \nz.mem_4498_sv2v_reg  <= data_i[18];
    end 
    if(N10874) begin
      \nz.mem_4497_sv2v_reg  <= data_i[17];
    end 
    if(N10873) begin
      \nz.mem_4496_sv2v_reg  <= data_i[16];
    end 
    if(N10872) begin
      \nz.mem_4495_sv2v_reg  <= data_i[15];
    end 
    if(N10871) begin
      \nz.mem_4494_sv2v_reg  <= data_i[14];
    end 
    if(N10870) begin
      \nz.mem_4493_sv2v_reg  <= data_i[13];
    end 
    if(N10869) begin
      \nz.mem_4492_sv2v_reg  <= data_i[12];
    end 
    if(N10868) begin
      \nz.mem_4491_sv2v_reg  <= data_i[11];
    end 
    if(N10867) begin
      \nz.mem_4490_sv2v_reg  <= data_i[10];
    end 
    if(N10866) begin
      \nz.mem_4489_sv2v_reg  <= data_i[9];
    end 
    if(N10865) begin
      \nz.mem_4488_sv2v_reg  <= data_i[8];
    end 
    if(N10864) begin
      \nz.mem_4487_sv2v_reg  <= data_i[7];
    end 
    if(N10863) begin
      \nz.mem_4486_sv2v_reg  <= data_i[6];
    end 
    if(N10862) begin
      \nz.mem_4485_sv2v_reg  <= data_i[5];
    end 
    if(N10861) begin
      \nz.mem_4484_sv2v_reg  <= data_i[4];
    end 
    if(N10860) begin
      \nz.mem_4483_sv2v_reg  <= data_i[3];
    end 
    if(N10859) begin
      \nz.mem_4482_sv2v_reg  <= data_i[2];
    end 
    if(N10858) begin
      \nz.mem_4481_sv2v_reg  <= data_i[1];
    end 
    if(N10857) begin
      \nz.mem_4480_sv2v_reg  <= data_i[0];
    end 
    if(N10856) begin
      \nz.mem_4479_sv2v_reg  <= data_i[79];
    end 
    if(N10855) begin
      \nz.mem_4478_sv2v_reg  <= data_i[78];
    end 
    if(N10854) begin
      \nz.mem_4477_sv2v_reg  <= data_i[77];
    end 
    if(N10853) begin
      \nz.mem_4476_sv2v_reg  <= data_i[76];
    end 
    if(N10852) begin
      \nz.mem_4475_sv2v_reg  <= data_i[75];
    end 
    if(N10851) begin
      \nz.mem_4474_sv2v_reg  <= data_i[74];
    end 
    if(N10850) begin
      \nz.mem_4473_sv2v_reg  <= data_i[73];
    end 
    if(N10849) begin
      \nz.mem_4472_sv2v_reg  <= data_i[72];
    end 
    if(N10848) begin
      \nz.mem_4471_sv2v_reg  <= data_i[71];
    end 
    if(N10847) begin
      \nz.mem_4470_sv2v_reg  <= data_i[70];
    end 
    if(N10846) begin
      \nz.mem_4469_sv2v_reg  <= data_i[69];
    end 
    if(N10845) begin
      \nz.mem_4468_sv2v_reg  <= data_i[68];
    end 
    if(N10844) begin
      \nz.mem_4467_sv2v_reg  <= data_i[67];
    end 
    if(N10843) begin
      \nz.mem_4466_sv2v_reg  <= data_i[66];
    end 
    if(N10842) begin
      \nz.mem_4465_sv2v_reg  <= data_i[65];
    end 
    if(N10841) begin
      \nz.mem_4464_sv2v_reg  <= data_i[64];
    end 
    if(N10840) begin
      \nz.mem_4463_sv2v_reg  <= data_i[63];
    end 
    if(N10839) begin
      \nz.mem_4462_sv2v_reg  <= data_i[62];
    end 
    if(N10838) begin
      \nz.mem_4461_sv2v_reg  <= data_i[61];
    end 
    if(N10837) begin
      \nz.mem_4460_sv2v_reg  <= data_i[60];
    end 
    if(N10836) begin
      \nz.mem_4459_sv2v_reg  <= data_i[59];
    end 
    if(N10835) begin
      \nz.mem_4458_sv2v_reg  <= data_i[58];
    end 
    if(N10834) begin
      \nz.mem_4457_sv2v_reg  <= data_i[57];
    end 
    if(N10833) begin
      \nz.mem_4456_sv2v_reg  <= data_i[56];
    end 
    if(N10832) begin
      \nz.mem_4455_sv2v_reg  <= data_i[55];
    end 
    if(N10831) begin
      \nz.mem_4454_sv2v_reg  <= data_i[54];
    end 
    if(N10830) begin
      \nz.mem_4453_sv2v_reg  <= data_i[53];
    end 
    if(N10829) begin
      \nz.mem_4452_sv2v_reg  <= data_i[52];
    end 
    if(N10828) begin
      \nz.mem_4451_sv2v_reg  <= data_i[51];
    end 
    if(N10827) begin
      \nz.mem_4450_sv2v_reg  <= data_i[50];
    end 
    if(N10826) begin
      \nz.mem_4449_sv2v_reg  <= data_i[49];
    end 
    if(N10825) begin
      \nz.mem_4448_sv2v_reg  <= data_i[48];
    end 
    if(N10824) begin
      \nz.mem_4447_sv2v_reg  <= data_i[47];
    end 
    if(N10823) begin
      \nz.mem_4446_sv2v_reg  <= data_i[46];
    end 
    if(N10822) begin
      \nz.mem_4445_sv2v_reg  <= data_i[45];
    end 
    if(N10821) begin
      \nz.mem_4444_sv2v_reg  <= data_i[44];
    end 
    if(N10820) begin
      \nz.mem_4443_sv2v_reg  <= data_i[43];
    end 
    if(N10819) begin
      \nz.mem_4442_sv2v_reg  <= data_i[42];
    end 
    if(N10818) begin
      \nz.mem_4441_sv2v_reg  <= data_i[41];
    end 
    if(N10817) begin
      \nz.mem_4440_sv2v_reg  <= data_i[40];
    end 
    if(N10816) begin
      \nz.mem_4439_sv2v_reg  <= data_i[39];
    end 
    if(N10815) begin
      \nz.mem_4438_sv2v_reg  <= data_i[38];
    end 
    if(N10814) begin
      \nz.mem_4437_sv2v_reg  <= data_i[37];
    end 
    if(N10813) begin
      \nz.mem_4436_sv2v_reg  <= data_i[36];
    end 
    if(N10812) begin
      \nz.mem_4435_sv2v_reg  <= data_i[35];
    end 
    if(N10811) begin
      \nz.mem_4434_sv2v_reg  <= data_i[34];
    end 
    if(N10810) begin
      \nz.mem_4433_sv2v_reg  <= data_i[33];
    end 
    if(N10809) begin
      \nz.mem_4432_sv2v_reg  <= data_i[32];
    end 
    if(N10808) begin
      \nz.mem_4431_sv2v_reg  <= data_i[31];
    end 
    if(N10807) begin
      \nz.mem_4430_sv2v_reg  <= data_i[30];
    end 
    if(N10806) begin
      \nz.mem_4429_sv2v_reg  <= data_i[29];
    end 
    if(N10805) begin
      \nz.mem_4428_sv2v_reg  <= data_i[28];
    end 
    if(N10804) begin
      \nz.mem_4427_sv2v_reg  <= data_i[27];
    end 
    if(N10803) begin
      \nz.mem_4426_sv2v_reg  <= data_i[26];
    end 
    if(N10802) begin
      \nz.mem_4425_sv2v_reg  <= data_i[25];
    end 
    if(N10801) begin
      \nz.mem_4424_sv2v_reg  <= data_i[24];
    end 
    if(N10800) begin
      \nz.mem_4423_sv2v_reg  <= data_i[23];
    end 
    if(N10799) begin
      \nz.mem_4422_sv2v_reg  <= data_i[22];
    end 
    if(N10798) begin
      \nz.mem_4421_sv2v_reg  <= data_i[21];
    end 
    if(N10797) begin
      \nz.mem_4420_sv2v_reg  <= data_i[20];
    end 
    if(N10796) begin
      \nz.mem_4419_sv2v_reg  <= data_i[19];
    end 
    if(N10795) begin
      \nz.mem_4418_sv2v_reg  <= data_i[18];
    end 
    if(N10794) begin
      \nz.mem_4417_sv2v_reg  <= data_i[17];
    end 
    if(N10793) begin
      \nz.mem_4416_sv2v_reg  <= data_i[16];
    end 
    if(N10792) begin
      \nz.mem_4415_sv2v_reg  <= data_i[15];
    end 
    if(N10791) begin
      \nz.mem_4414_sv2v_reg  <= data_i[14];
    end 
    if(N10790) begin
      \nz.mem_4413_sv2v_reg  <= data_i[13];
    end 
    if(N10789) begin
      \nz.mem_4412_sv2v_reg  <= data_i[12];
    end 
    if(N10788) begin
      \nz.mem_4411_sv2v_reg  <= data_i[11];
    end 
    if(N10787) begin
      \nz.mem_4410_sv2v_reg  <= data_i[10];
    end 
    if(N10786) begin
      \nz.mem_4409_sv2v_reg  <= data_i[9];
    end 
    if(N10785) begin
      \nz.mem_4408_sv2v_reg  <= data_i[8];
    end 
    if(N10784) begin
      \nz.mem_4407_sv2v_reg  <= data_i[7];
    end 
    if(N10783) begin
      \nz.mem_4406_sv2v_reg  <= data_i[6];
    end 
    if(N10782) begin
      \nz.mem_4405_sv2v_reg  <= data_i[5];
    end 
    if(N10781) begin
      \nz.mem_4404_sv2v_reg  <= data_i[4];
    end 
    if(N10780) begin
      \nz.mem_4403_sv2v_reg  <= data_i[3];
    end 
    if(N10779) begin
      \nz.mem_4402_sv2v_reg  <= data_i[2];
    end 
    if(N10778) begin
      \nz.mem_4401_sv2v_reg  <= data_i[1];
    end 
    if(N10777) begin
      \nz.mem_4400_sv2v_reg  <= data_i[0];
    end 
    if(N10776) begin
      \nz.mem_4399_sv2v_reg  <= data_i[79];
    end 
    if(N10775) begin
      \nz.mem_4398_sv2v_reg  <= data_i[78];
    end 
    if(N10774) begin
      \nz.mem_4397_sv2v_reg  <= data_i[77];
    end 
    if(N10773) begin
      \nz.mem_4396_sv2v_reg  <= data_i[76];
    end 
    if(N10772) begin
      \nz.mem_4395_sv2v_reg  <= data_i[75];
    end 
    if(N10771) begin
      \nz.mem_4394_sv2v_reg  <= data_i[74];
    end 
    if(N10770) begin
      \nz.mem_4393_sv2v_reg  <= data_i[73];
    end 
    if(N10769) begin
      \nz.mem_4392_sv2v_reg  <= data_i[72];
    end 
    if(N10768) begin
      \nz.mem_4391_sv2v_reg  <= data_i[71];
    end 
    if(N10767) begin
      \nz.mem_4390_sv2v_reg  <= data_i[70];
    end 
    if(N10766) begin
      \nz.mem_4389_sv2v_reg  <= data_i[69];
    end 
    if(N10765) begin
      \nz.mem_4388_sv2v_reg  <= data_i[68];
    end 
    if(N10764) begin
      \nz.mem_4387_sv2v_reg  <= data_i[67];
    end 
    if(N10763) begin
      \nz.mem_4386_sv2v_reg  <= data_i[66];
    end 
    if(N10762) begin
      \nz.mem_4385_sv2v_reg  <= data_i[65];
    end 
    if(N10761) begin
      \nz.mem_4384_sv2v_reg  <= data_i[64];
    end 
    if(N10760) begin
      \nz.mem_4383_sv2v_reg  <= data_i[63];
    end 
    if(N10759) begin
      \nz.mem_4382_sv2v_reg  <= data_i[62];
    end 
    if(N10758) begin
      \nz.mem_4381_sv2v_reg  <= data_i[61];
    end 
    if(N10757) begin
      \nz.mem_4380_sv2v_reg  <= data_i[60];
    end 
    if(N10756) begin
      \nz.mem_4379_sv2v_reg  <= data_i[59];
    end 
    if(N10755) begin
      \nz.mem_4378_sv2v_reg  <= data_i[58];
    end 
    if(N10754) begin
      \nz.mem_4377_sv2v_reg  <= data_i[57];
    end 
    if(N10753) begin
      \nz.mem_4376_sv2v_reg  <= data_i[56];
    end 
    if(N10752) begin
      \nz.mem_4375_sv2v_reg  <= data_i[55];
    end 
    if(N10751) begin
      \nz.mem_4374_sv2v_reg  <= data_i[54];
    end 
    if(N10750) begin
      \nz.mem_4373_sv2v_reg  <= data_i[53];
    end 
    if(N10749) begin
      \nz.mem_4372_sv2v_reg  <= data_i[52];
    end 
    if(N10748) begin
      \nz.mem_4371_sv2v_reg  <= data_i[51];
    end 
    if(N10747) begin
      \nz.mem_4370_sv2v_reg  <= data_i[50];
    end 
    if(N10746) begin
      \nz.mem_4369_sv2v_reg  <= data_i[49];
    end 
    if(N10745) begin
      \nz.mem_4368_sv2v_reg  <= data_i[48];
    end 
    if(N10744) begin
      \nz.mem_4367_sv2v_reg  <= data_i[47];
    end 
    if(N10743) begin
      \nz.mem_4366_sv2v_reg  <= data_i[46];
    end 
    if(N10742) begin
      \nz.mem_4365_sv2v_reg  <= data_i[45];
    end 
    if(N10741) begin
      \nz.mem_4364_sv2v_reg  <= data_i[44];
    end 
    if(N10740) begin
      \nz.mem_4363_sv2v_reg  <= data_i[43];
    end 
    if(N10739) begin
      \nz.mem_4362_sv2v_reg  <= data_i[42];
    end 
    if(N10738) begin
      \nz.mem_4361_sv2v_reg  <= data_i[41];
    end 
    if(N10737) begin
      \nz.mem_4360_sv2v_reg  <= data_i[40];
    end 
    if(N10736) begin
      \nz.mem_4359_sv2v_reg  <= data_i[39];
    end 
    if(N10735) begin
      \nz.mem_4358_sv2v_reg  <= data_i[38];
    end 
    if(N10734) begin
      \nz.mem_4357_sv2v_reg  <= data_i[37];
    end 
    if(N10733) begin
      \nz.mem_4356_sv2v_reg  <= data_i[36];
    end 
    if(N10732) begin
      \nz.mem_4355_sv2v_reg  <= data_i[35];
    end 
    if(N10731) begin
      \nz.mem_4354_sv2v_reg  <= data_i[34];
    end 
    if(N10730) begin
      \nz.mem_4353_sv2v_reg  <= data_i[33];
    end 
    if(N10729) begin
      \nz.mem_4352_sv2v_reg  <= data_i[32];
    end 
    if(N10728) begin
      \nz.mem_4351_sv2v_reg  <= data_i[31];
    end 
    if(N10727) begin
      \nz.mem_4350_sv2v_reg  <= data_i[30];
    end 
    if(N10726) begin
      \nz.mem_4349_sv2v_reg  <= data_i[29];
    end 
    if(N10725) begin
      \nz.mem_4348_sv2v_reg  <= data_i[28];
    end 
    if(N10724) begin
      \nz.mem_4347_sv2v_reg  <= data_i[27];
    end 
    if(N10723) begin
      \nz.mem_4346_sv2v_reg  <= data_i[26];
    end 
    if(N10722) begin
      \nz.mem_4345_sv2v_reg  <= data_i[25];
    end 
    if(N10721) begin
      \nz.mem_4344_sv2v_reg  <= data_i[24];
    end 
    if(N10720) begin
      \nz.mem_4343_sv2v_reg  <= data_i[23];
    end 
    if(N10719) begin
      \nz.mem_4342_sv2v_reg  <= data_i[22];
    end 
    if(N10718) begin
      \nz.mem_4341_sv2v_reg  <= data_i[21];
    end 
    if(N10717) begin
      \nz.mem_4340_sv2v_reg  <= data_i[20];
    end 
    if(N10716) begin
      \nz.mem_4339_sv2v_reg  <= data_i[19];
    end 
    if(N10715) begin
      \nz.mem_4338_sv2v_reg  <= data_i[18];
    end 
    if(N10714) begin
      \nz.mem_4337_sv2v_reg  <= data_i[17];
    end 
    if(N10713) begin
      \nz.mem_4336_sv2v_reg  <= data_i[16];
    end 
    if(N10712) begin
      \nz.mem_4335_sv2v_reg  <= data_i[15];
    end 
    if(N10711) begin
      \nz.mem_4334_sv2v_reg  <= data_i[14];
    end 
    if(N10710) begin
      \nz.mem_4333_sv2v_reg  <= data_i[13];
    end 
    if(N10709) begin
      \nz.mem_4332_sv2v_reg  <= data_i[12];
    end 
    if(N10708) begin
      \nz.mem_4331_sv2v_reg  <= data_i[11];
    end 
    if(N10707) begin
      \nz.mem_4330_sv2v_reg  <= data_i[10];
    end 
    if(N10706) begin
      \nz.mem_4329_sv2v_reg  <= data_i[9];
    end 
    if(N10705) begin
      \nz.mem_4328_sv2v_reg  <= data_i[8];
    end 
    if(N10704) begin
      \nz.mem_4327_sv2v_reg  <= data_i[7];
    end 
    if(N10703) begin
      \nz.mem_4326_sv2v_reg  <= data_i[6];
    end 
    if(N10702) begin
      \nz.mem_4325_sv2v_reg  <= data_i[5];
    end 
    if(N10701) begin
      \nz.mem_4324_sv2v_reg  <= data_i[4];
    end 
    if(N10700) begin
      \nz.mem_4323_sv2v_reg  <= data_i[3];
    end 
    if(N10699) begin
      \nz.mem_4322_sv2v_reg  <= data_i[2];
    end 
    if(N10698) begin
      \nz.mem_4321_sv2v_reg  <= data_i[1];
    end 
    if(N10697) begin
      \nz.mem_4320_sv2v_reg  <= data_i[0];
    end 
    if(N10696) begin
      \nz.mem_4319_sv2v_reg  <= data_i[79];
    end 
    if(N10695) begin
      \nz.mem_4318_sv2v_reg  <= data_i[78];
    end 
    if(N10694) begin
      \nz.mem_4317_sv2v_reg  <= data_i[77];
    end 
    if(N10693) begin
      \nz.mem_4316_sv2v_reg  <= data_i[76];
    end 
    if(N10692) begin
      \nz.mem_4315_sv2v_reg  <= data_i[75];
    end 
    if(N10691) begin
      \nz.mem_4314_sv2v_reg  <= data_i[74];
    end 
    if(N10690) begin
      \nz.mem_4313_sv2v_reg  <= data_i[73];
    end 
    if(N10689) begin
      \nz.mem_4312_sv2v_reg  <= data_i[72];
    end 
    if(N10688) begin
      \nz.mem_4311_sv2v_reg  <= data_i[71];
    end 
    if(N10687) begin
      \nz.mem_4310_sv2v_reg  <= data_i[70];
    end 
    if(N10686) begin
      \nz.mem_4309_sv2v_reg  <= data_i[69];
    end 
    if(N10685) begin
      \nz.mem_4308_sv2v_reg  <= data_i[68];
    end 
    if(N10684) begin
      \nz.mem_4307_sv2v_reg  <= data_i[67];
    end 
    if(N10683) begin
      \nz.mem_4306_sv2v_reg  <= data_i[66];
    end 
    if(N10682) begin
      \nz.mem_4305_sv2v_reg  <= data_i[65];
    end 
    if(N10681) begin
      \nz.mem_4304_sv2v_reg  <= data_i[64];
    end 
    if(N10680) begin
      \nz.mem_4303_sv2v_reg  <= data_i[63];
    end 
    if(N10679) begin
      \nz.mem_4302_sv2v_reg  <= data_i[62];
    end 
    if(N10678) begin
      \nz.mem_4301_sv2v_reg  <= data_i[61];
    end 
    if(N10677) begin
      \nz.mem_4300_sv2v_reg  <= data_i[60];
    end 
    if(N10676) begin
      \nz.mem_4299_sv2v_reg  <= data_i[59];
    end 
    if(N10675) begin
      \nz.mem_4298_sv2v_reg  <= data_i[58];
    end 
    if(N10674) begin
      \nz.mem_4297_sv2v_reg  <= data_i[57];
    end 
    if(N10673) begin
      \nz.mem_4296_sv2v_reg  <= data_i[56];
    end 
    if(N10672) begin
      \nz.mem_4295_sv2v_reg  <= data_i[55];
    end 
    if(N10671) begin
      \nz.mem_4294_sv2v_reg  <= data_i[54];
    end 
    if(N10670) begin
      \nz.mem_4293_sv2v_reg  <= data_i[53];
    end 
    if(N10669) begin
      \nz.mem_4292_sv2v_reg  <= data_i[52];
    end 
    if(N10668) begin
      \nz.mem_4291_sv2v_reg  <= data_i[51];
    end 
    if(N10667) begin
      \nz.mem_4290_sv2v_reg  <= data_i[50];
    end 
    if(N10666) begin
      \nz.mem_4289_sv2v_reg  <= data_i[49];
    end 
    if(N10665) begin
      \nz.mem_4288_sv2v_reg  <= data_i[48];
    end 
    if(N10664) begin
      \nz.mem_4287_sv2v_reg  <= data_i[47];
    end 
    if(N10663) begin
      \nz.mem_4286_sv2v_reg  <= data_i[46];
    end 
    if(N10662) begin
      \nz.mem_4285_sv2v_reg  <= data_i[45];
    end 
    if(N10661) begin
      \nz.mem_4284_sv2v_reg  <= data_i[44];
    end 
    if(N10660) begin
      \nz.mem_4283_sv2v_reg  <= data_i[43];
    end 
    if(N10659) begin
      \nz.mem_4282_sv2v_reg  <= data_i[42];
    end 
    if(N10658) begin
      \nz.mem_4281_sv2v_reg  <= data_i[41];
    end 
    if(N10657) begin
      \nz.mem_4280_sv2v_reg  <= data_i[40];
    end 
    if(N10656) begin
      \nz.mem_4279_sv2v_reg  <= data_i[39];
    end 
    if(N10655) begin
      \nz.mem_4278_sv2v_reg  <= data_i[38];
    end 
    if(N10654) begin
      \nz.mem_4277_sv2v_reg  <= data_i[37];
    end 
    if(N10653) begin
      \nz.mem_4276_sv2v_reg  <= data_i[36];
    end 
    if(N10652) begin
      \nz.mem_4275_sv2v_reg  <= data_i[35];
    end 
    if(N10651) begin
      \nz.mem_4274_sv2v_reg  <= data_i[34];
    end 
    if(N10650) begin
      \nz.mem_4273_sv2v_reg  <= data_i[33];
    end 
    if(N10649) begin
      \nz.mem_4272_sv2v_reg  <= data_i[32];
    end 
    if(N10648) begin
      \nz.mem_4271_sv2v_reg  <= data_i[31];
    end 
    if(N10647) begin
      \nz.mem_4270_sv2v_reg  <= data_i[30];
    end 
    if(N10646) begin
      \nz.mem_4269_sv2v_reg  <= data_i[29];
    end 
    if(N10645) begin
      \nz.mem_4268_sv2v_reg  <= data_i[28];
    end 
    if(N10644) begin
      \nz.mem_4267_sv2v_reg  <= data_i[27];
    end 
    if(N10643) begin
      \nz.mem_4266_sv2v_reg  <= data_i[26];
    end 
    if(N10642) begin
      \nz.mem_4265_sv2v_reg  <= data_i[25];
    end 
    if(N10641) begin
      \nz.mem_4264_sv2v_reg  <= data_i[24];
    end 
    if(N10640) begin
      \nz.mem_4263_sv2v_reg  <= data_i[23];
    end 
    if(N10639) begin
      \nz.mem_4262_sv2v_reg  <= data_i[22];
    end 
    if(N10638) begin
      \nz.mem_4261_sv2v_reg  <= data_i[21];
    end 
    if(N10637) begin
      \nz.mem_4260_sv2v_reg  <= data_i[20];
    end 
    if(N10636) begin
      \nz.mem_4259_sv2v_reg  <= data_i[19];
    end 
    if(N10635) begin
      \nz.mem_4258_sv2v_reg  <= data_i[18];
    end 
    if(N10634) begin
      \nz.mem_4257_sv2v_reg  <= data_i[17];
    end 
    if(N10633) begin
      \nz.mem_4256_sv2v_reg  <= data_i[16];
    end 
    if(N10632) begin
      \nz.mem_4255_sv2v_reg  <= data_i[15];
    end 
    if(N10631) begin
      \nz.mem_4254_sv2v_reg  <= data_i[14];
    end 
    if(N10630) begin
      \nz.mem_4253_sv2v_reg  <= data_i[13];
    end 
    if(N10629) begin
      \nz.mem_4252_sv2v_reg  <= data_i[12];
    end 
    if(N10628) begin
      \nz.mem_4251_sv2v_reg  <= data_i[11];
    end 
    if(N10627) begin
      \nz.mem_4250_sv2v_reg  <= data_i[10];
    end 
    if(N10626) begin
      \nz.mem_4249_sv2v_reg  <= data_i[9];
    end 
    if(N10625) begin
      \nz.mem_4248_sv2v_reg  <= data_i[8];
    end 
    if(N10624) begin
      \nz.mem_4247_sv2v_reg  <= data_i[7];
    end 
    if(N10623) begin
      \nz.mem_4246_sv2v_reg  <= data_i[6];
    end 
    if(N10622) begin
      \nz.mem_4245_sv2v_reg  <= data_i[5];
    end 
    if(N10621) begin
      \nz.mem_4244_sv2v_reg  <= data_i[4];
    end 
    if(N10620) begin
      \nz.mem_4243_sv2v_reg  <= data_i[3];
    end 
    if(N10619) begin
      \nz.mem_4242_sv2v_reg  <= data_i[2];
    end 
    if(N10618) begin
      \nz.mem_4241_sv2v_reg  <= data_i[1];
    end 
    if(N10617) begin
      \nz.mem_4240_sv2v_reg  <= data_i[0];
    end 
    if(N10616) begin
      \nz.mem_4239_sv2v_reg  <= data_i[79];
    end 
    if(N10615) begin
      \nz.mem_4238_sv2v_reg  <= data_i[78];
    end 
    if(N10614) begin
      \nz.mem_4237_sv2v_reg  <= data_i[77];
    end 
    if(N10613) begin
      \nz.mem_4236_sv2v_reg  <= data_i[76];
    end 
    if(N10612) begin
      \nz.mem_4235_sv2v_reg  <= data_i[75];
    end 
    if(N10611) begin
      \nz.mem_4234_sv2v_reg  <= data_i[74];
    end 
    if(N10610) begin
      \nz.mem_4233_sv2v_reg  <= data_i[73];
    end 
    if(N10609) begin
      \nz.mem_4232_sv2v_reg  <= data_i[72];
    end 
    if(N10608) begin
      \nz.mem_4231_sv2v_reg  <= data_i[71];
    end 
    if(N10607) begin
      \nz.mem_4230_sv2v_reg  <= data_i[70];
    end 
    if(N10606) begin
      \nz.mem_4229_sv2v_reg  <= data_i[69];
    end 
    if(N10605) begin
      \nz.mem_4228_sv2v_reg  <= data_i[68];
    end 
    if(N10604) begin
      \nz.mem_4227_sv2v_reg  <= data_i[67];
    end 
    if(N10603) begin
      \nz.mem_4226_sv2v_reg  <= data_i[66];
    end 
    if(N10602) begin
      \nz.mem_4225_sv2v_reg  <= data_i[65];
    end 
    if(N10601) begin
      \nz.mem_4224_sv2v_reg  <= data_i[64];
    end 
    if(N10600) begin
      \nz.mem_4223_sv2v_reg  <= data_i[63];
    end 
    if(N10599) begin
      \nz.mem_4222_sv2v_reg  <= data_i[62];
    end 
    if(N10598) begin
      \nz.mem_4221_sv2v_reg  <= data_i[61];
    end 
    if(N10597) begin
      \nz.mem_4220_sv2v_reg  <= data_i[60];
    end 
    if(N10596) begin
      \nz.mem_4219_sv2v_reg  <= data_i[59];
    end 
    if(N10595) begin
      \nz.mem_4218_sv2v_reg  <= data_i[58];
    end 
    if(N10594) begin
      \nz.mem_4217_sv2v_reg  <= data_i[57];
    end 
    if(N10593) begin
      \nz.mem_4216_sv2v_reg  <= data_i[56];
    end 
    if(N10592) begin
      \nz.mem_4215_sv2v_reg  <= data_i[55];
    end 
    if(N10591) begin
      \nz.mem_4214_sv2v_reg  <= data_i[54];
    end 
    if(N10590) begin
      \nz.mem_4213_sv2v_reg  <= data_i[53];
    end 
    if(N10589) begin
      \nz.mem_4212_sv2v_reg  <= data_i[52];
    end 
    if(N10588) begin
      \nz.mem_4211_sv2v_reg  <= data_i[51];
    end 
    if(N10587) begin
      \nz.mem_4210_sv2v_reg  <= data_i[50];
    end 
    if(N10586) begin
      \nz.mem_4209_sv2v_reg  <= data_i[49];
    end 
    if(N10585) begin
      \nz.mem_4208_sv2v_reg  <= data_i[48];
    end 
    if(N10584) begin
      \nz.mem_4207_sv2v_reg  <= data_i[47];
    end 
    if(N10583) begin
      \nz.mem_4206_sv2v_reg  <= data_i[46];
    end 
    if(N10582) begin
      \nz.mem_4205_sv2v_reg  <= data_i[45];
    end 
    if(N10581) begin
      \nz.mem_4204_sv2v_reg  <= data_i[44];
    end 
    if(N10580) begin
      \nz.mem_4203_sv2v_reg  <= data_i[43];
    end 
    if(N10579) begin
      \nz.mem_4202_sv2v_reg  <= data_i[42];
    end 
    if(N10578) begin
      \nz.mem_4201_sv2v_reg  <= data_i[41];
    end 
    if(N10577) begin
      \nz.mem_4200_sv2v_reg  <= data_i[40];
    end 
    if(N10576) begin
      \nz.mem_4199_sv2v_reg  <= data_i[39];
    end 
    if(N10575) begin
      \nz.mem_4198_sv2v_reg  <= data_i[38];
    end 
    if(N10574) begin
      \nz.mem_4197_sv2v_reg  <= data_i[37];
    end 
    if(N10573) begin
      \nz.mem_4196_sv2v_reg  <= data_i[36];
    end 
    if(N10572) begin
      \nz.mem_4195_sv2v_reg  <= data_i[35];
    end 
    if(N10571) begin
      \nz.mem_4194_sv2v_reg  <= data_i[34];
    end 
    if(N10570) begin
      \nz.mem_4193_sv2v_reg  <= data_i[33];
    end 
    if(N10569) begin
      \nz.mem_4192_sv2v_reg  <= data_i[32];
    end 
    if(N10568) begin
      \nz.mem_4191_sv2v_reg  <= data_i[31];
    end 
    if(N10567) begin
      \nz.mem_4190_sv2v_reg  <= data_i[30];
    end 
    if(N10566) begin
      \nz.mem_4189_sv2v_reg  <= data_i[29];
    end 
    if(N10565) begin
      \nz.mem_4188_sv2v_reg  <= data_i[28];
    end 
    if(N10564) begin
      \nz.mem_4187_sv2v_reg  <= data_i[27];
    end 
    if(N10563) begin
      \nz.mem_4186_sv2v_reg  <= data_i[26];
    end 
    if(N10562) begin
      \nz.mem_4185_sv2v_reg  <= data_i[25];
    end 
    if(N10561) begin
      \nz.mem_4184_sv2v_reg  <= data_i[24];
    end 
    if(N10560) begin
      \nz.mem_4183_sv2v_reg  <= data_i[23];
    end 
    if(N10559) begin
      \nz.mem_4182_sv2v_reg  <= data_i[22];
    end 
    if(N10558) begin
      \nz.mem_4181_sv2v_reg  <= data_i[21];
    end 
    if(N10557) begin
      \nz.mem_4180_sv2v_reg  <= data_i[20];
    end 
    if(N10556) begin
      \nz.mem_4179_sv2v_reg  <= data_i[19];
    end 
    if(N10555) begin
      \nz.mem_4178_sv2v_reg  <= data_i[18];
    end 
    if(N10554) begin
      \nz.mem_4177_sv2v_reg  <= data_i[17];
    end 
    if(N10553) begin
      \nz.mem_4176_sv2v_reg  <= data_i[16];
    end 
    if(N10552) begin
      \nz.mem_4175_sv2v_reg  <= data_i[15];
    end 
    if(N10551) begin
      \nz.mem_4174_sv2v_reg  <= data_i[14];
    end 
    if(N10550) begin
      \nz.mem_4173_sv2v_reg  <= data_i[13];
    end 
    if(N10549) begin
      \nz.mem_4172_sv2v_reg  <= data_i[12];
    end 
    if(N10548) begin
      \nz.mem_4171_sv2v_reg  <= data_i[11];
    end 
    if(N10547) begin
      \nz.mem_4170_sv2v_reg  <= data_i[10];
    end 
    if(N10546) begin
      \nz.mem_4169_sv2v_reg  <= data_i[9];
    end 
    if(N10545) begin
      \nz.mem_4168_sv2v_reg  <= data_i[8];
    end 
    if(N10544) begin
      \nz.mem_4167_sv2v_reg  <= data_i[7];
    end 
    if(N10543) begin
      \nz.mem_4166_sv2v_reg  <= data_i[6];
    end 
    if(N10542) begin
      \nz.mem_4165_sv2v_reg  <= data_i[5];
    end 
    if(N10541) begin
      \nz.mem_4164_sv2v_reg  <= data_i[4];
    end 
    if(N10540) begin
      \nz.mem_4163_sv2v_reg  <= data_i[3];
    end 
    if(N10539) begin
      \nz.mem_4162_sv2v_reg  <= data_i[2];
    end 
    if(N10538) begin
      \nz.mem_4161_sv2v_reg  <= data_i[1];
    end 
    if(N10537) begin
      \nz.mem_4160_sv2v_reg  <= data_i[0];
    end 
    if(N10536) begin
      \nz.mem_4159_sv2v_reg  <= data_i[79];
    end 
    if(N10535) begin
      \nz.mem_4158_sv2v_reg  <= data_i[78];
    end 
    if(N10534) begin
      \nz.mem_4157_sv2v_reg  <= data_i[77];
    end 
    if(N10533) begin
      \nz.mem_4156_sv2v_reg  <= data_i[76];
    end 
    if(N10532) begin
      \nz.mem_4155_sv2v_reg  <= data_i[75];
    end 
    if(N10531) begin
      \nz.mem_4154_sv2v_reg  <= data_i[74];
    end 
    if(N10530) begin
      \nz.mem_4153_sv2v_reg  <= data_i[73];
    end 
    if(N10529) begin
      \nz.mem_4152_sv2v_reg  <= data_i[72];
    end 
    if(N10528) begin
      \nz.mem_4151_sv2v_reg  <= data_i[71];
    end 
    if(N10527) begin
      \nz.mem_4150_sv2v_reg  <= data_i[70];
    end 
    if(N10526) begin
      \nz.mem_4149_sv2v_reg  <= data_i[69];
    end 
    if(N10525) begin
      \nz.mem_4148_sv2v_reg  <= data_i[68];
    end 
    if(N10524) begin
      \nz.mem_4147_sv2v_reg  <= data_i[67];
    end 
    if(N10523) begin
      \nz.mem_4146_sv2v_reg  <= data_i[66];
    end 
    if(N10522) begin
      \nz.mem_4145_sv2v_reg  <= data_i[65];
    end 
    if(N10521) begin
      \nz.mem_4144_sv2v_reg  <= data_i[64];
    end 
    if(N10520) begin
      \nz.mem_4143_sv2v_reg  <= data_i[63];
    end 
    if(N10519) begin
      \nz.mem_4142_sv2v_reg  <= data_i[62];
    end 
    if(N10518) begin
      \nz.mem_4141_sv2v_reg  <= data_i[61];
    end 
    if(N10517) begin
      \nz.mem_4140_sv2v_reg  <= data_i[60];
    end 
    if(N10516) begin
      \nz.mem_4139_sv2v_reg  <= data_i[59];
    end 
    if(N10515) begin
      \nz.mem_4138_sv2v_reg  <= data_i[58];
    end 
    if(N10514) begin
      \nz.mem_4137_sv2v_reg  <= data_i[57];
    end 
    if(N10513) begin
      \nz.mem_4136_sv2v_reg  <= data_i[56];
    end 
    if(N10512) begin
      \nz.mem_4135_sv2v_reg  <= data_i[55];
    end 
    if(N10511) begin
      \nz.mem_4134_sv2v_reg  <= data_i[54];
    end 
    if(N10510) begin
      \nz.mem_4133_sv2v_reg  <= data_i[53];
    end 
    if(N10509) begin
      \nz.mem_4132_sv2v_reg  <= data_i[52];
    end 
    if(N10508) begin
      \nz.mem_4131_sv2v_reg  <= data_i[51];
    end 
    if(N10507) begin
      \nz.mem_4130_sv2v_reg  <= data_i[50];
    end 
    if(N10506) begin
      \nz.mem_4129_sv2v_reg  <= data_i[49];
    end 
    if(N10505) begin
      \nz.mem_4128_sv2v_reg  <= data_i[48];
    end 
    if(N10504) begin
      \nz.mem_4127_sv2v_reg  <= data_i[47];
    end 
    if(N10503) begin
      \nz.mem_4126_sv2v_reg  <= data_i[46];
    end 
    if(N10502) begin
      \nz.mem_4125_sv2v_reg  <= data_i[45];
    end 
    if(N10501) begin
      \nz.mem_4124_sv2v_reg  <= data_i[44];
    end 
    if(N10500) begin
      \nz.mem_4123_sv2v_reg  <= data_i[43];
    end 
    if(N10499) begin
      \nz.mem_4122_sv2v_reg  <= data_i[42];
    end 
    if(N10498) begin
      \nz.mem_4121_sv2v_reg  <= data_i[41];
    end 
    if(N10497) begin
      \nz.mem_4120_sv2v_reg  <= data_i[40];
    end 
    if(N10496) begin
      \nz.mem_4119_sv2v_reg  <= data_i[39];
    end 
    if(N10495) begin
      \nz.mem_4118_sv2v_reg  <= data_i[38];
    end 
    if(N10494) begin
      \nz.mem_4117_sv2v_reg  <= data_i[37];
    end 
    if(N10493) begin
      \nz.mem_4116_sv2v_reg  <= data_i[36];
    end 
    if(N10492) begin
      \nz.mem_4115_sv2v_reg  <= data_i[35];
    end 
    if(N10491) begin
      \nz.mem_4114_sv2v_reg  <= data_i[34];
    end 
    if(N10490) begin
      \nz.mem_4113_sv2v_reg  <= data_i[33];
    end 
    if(N10489) begin
      \nz.mem_4112_sv2v_reg  <= data_i[32];
    end 
    if(N10488) begin
      \nz.mem_4111_sv2v_reg  <= data_i[31];
    end 
    if(N10487) begin
      \nz.mem_4110_sv2v_reg  <= data_i[30];
    end 
    if(N10486) begin
      \nz.mem_4109_sv2v_reg  <= data_i[29];
    end 
    if(N10485) begin
      \nz.mem_4108_sv2v_reg  <= data_i[28];
    end 
    if(N10484) begin
      \nz.mem_4107_sv2v_reg  <= data_i[27];
    end 
    if(N10483) begin
      \nz.mem_4106_sv2v_reg  <= data_i[26];
    end 
    if(N10482) begin
      \nz.mem_4105_sv2v_reg  <= data_i[25];
    end 
    if(N10481) begin
      \nz.mem_4104_sv2v_reg  <= data_i[24];
    end 
    if(N10480) begin
      \nz.mem_4103_sv2v_reg  <= data_i[23];
    end 
    if(N10479) begin
      \nz.mem_4102_sv2v_reg  <= data_i[22];
    end 
    if(N10478) begin
      \nz.mem_4101_sv2v_reg  <= data_i[21];
    end 
    if(N10477) begin
      \nz.mem_4100_sv2v_reg  <= data_i[20];
    end 
    if(N10476) begin
      \nz.mem_4099_sv2v_reg  <= data_i[19];
    end 
    if(N10475) begin
      \nz.mem_4098_sv2v_reg  <= data_i[18];
    end 
    if(N10474) begin
      \nz.mem_4097_sv2v_reg  <= data_i[17];
    end 
    if(N10473) begin
      \nz.mem_4096_sv2v_reg  <= data_i[16];
    end 
    if(N10472) begin
      \nz.mem_4095_sv2v_reg  <= data_i[15];
    end 
    if(N10471) begin
      \nz.mem_4094_sv2v_reg  <= data_i[14];
    end 
    if(N10470) begin
      \nz.mem_4093_sv2v_reg  <= data_i[13];
    end 
    if(N10469) begin
      \nz.mem_4092_sv2v_reg  <= data_i[12];
    end 
    if(N10468) begin
      \nz.mem_4091_sv2v_reg  <= data_i[11];
    end 
    if(N10467) begin
      \nz.mem_4090_sv2v_reg  <= data_i[10];
    end 
    if(N10466) begin
      \nz.mem_4089_sv2v_reg  <= data_i[9];
    end 
    if(N10465) begin
      \nz.mem_4088_sv2v_reg  <= data_i[8];
    end 
    if(N10464) begin
      \nz.mem_4087_sv2v_reg  <= data_i[7];
    end 
    if(N10463) begin
      \nz.mem_4086_sv2v_reg  <= data_i[6];
    end 
    if(N10462) begin
      \nz.mem_4085_sv2v_reg  <= data_i[5];
    end 
    if(N10461) begin
      \nz.mem_4084_sv2v_reg  <= data_i[4];
    end 
    if(N10460) begin
      \nz.mem_4083_sv2v_reg  <= data_i[3];
    end 
    if(N10459) begin
      \nz.mem_4082_sv2v_reg  <= data_i[2];
    end 
    if(N10458) begin
      \nz.mem_4081_sv2v_reg  <= data_i[1];
    end 
    if(N10457) begin
      \nz.mem_4080_sv2v_reg  <= data_i[0];
    end 
    if(N10456) begin
      \nz.mem_4079_sv2v_reg  <= data_i[79];
    end 
    if(N10455) begin
      \nz.mem_4078_sv2v_reg  <= data_i[78];
    end 
    if(N10454) begin
      \nz.mem_4077_sv2v_reg  <= data_i[77];
    end 
    if(N10453) begin
      \nz.mem_4076_sv2v_reg  <= data_i[76];
    end 
    if(N10452) begin
      \nz.mem_4075_sv2v_reg  <= data_i[75];
    end 
    if(N10451) begin
      \nz.mem_4074_sv2v_reg  <= data_i[74];
    end 
    if(N10450) begin
      \nz.mem_4073_sv2v_reg  <= data_i[73];
    end 
    if(N10449) begin
      \nz.mem_4072_sv2v_reg  <= data_i[72];
    end 
    if(N10448) begin
      \nz.mem_4071_sv2v_reg  <= data_i[71];
    end 
    if(N10447) begin
      \nz.mem_4070_sv2v_reg  <= data_i[70];
    end 
    if(N10446) begin
      \nz.mem_4069_sv2v_reg  <= data_i[69];
    end 
    if(N10445) begin
      \nz.mem_4068_sv2v_reg  <= data_i[68];
    end 
    if(N10444) begin
      \nz.mem_4067_sv2v_reg  <= data_i[67];
    end 
    if(N10443) begin
      \nz.mem_4066_sv2v_reg  <= data_i[66];
    end 
    if(N10442) begin
      \nz.mem_4065_sv2v_reg  <= data_i[65];
    end 
    if(N10441) begin
      \nz.mem_4064_sv2v_reg  <= data_i[64];
    end 
    if(N10440) begin
      \nz.mem_4063_sv2v_reg  <= data_i[63];
    end 
    if(N10439) begin
      \nz.mem_4062_sv2v_reg  <= data_i[62];
    end 
    if(N10438) begin
      \nz.mem_4061_sv2v_reg  <= data_i[61];
    end 
    if(N10437) begin
      \nz.mem_4060_sv2v_reg  <= data_i[60];
    end 
    if(N10436) begin
      \nz.mem_4059_sv2v_reg  <= data_i[59];
    end 
    if(N10435) begin
      \nz.mem_4058_sv2v_reg  <= data_i[58];
    end 
    if(N10434) begin
      \nz.mem_4057_sv2v_reg  <= data_i[57];
    end 
    if(N10433) begin
      \nz.mem_4056_sv2v_reg  <= data_i[56];
    end 
    if(N10432) begin
      \nz.mem_4055_sv2v_reg  <= data_i[55];
    end 
    if(N10431) begin
      \nz.mem_4054_sv2v_reg  <= data_i[54];
    end 
    if(N10430) begin
      \nz.mem_4053_sv2v_reg  <= data_i[53];
    end 
    if(N10429) begin
      \nz.mem_4052_sv2v_reg  <= data_i[52];
    end 
    if(N10428) begin
      \nz.mem_4051_sv2v_reg  <= data_i[51];
    end 
    if(N10427) begin
      \nz.mem_4050_sv2v_reg  <= data_i[50];
    end 
    if(N10426) begin
      \nz.mem_4049_sv2v_reg  <= data_i[49];
    end 
    if(N10425) begin
      \nz.mem_4048_sv2v_reg  <= data_i[48];
    end 
    if(N10424) begin
      \nz.mem_4047_sv2v_reg  <= data_i[47];
    end 
    if(N10423) begin
      \nz.mem_4046_sv2v_reg  <= data_i[46];
    end 
    if(N10422) begin
      \nz.mem_4045_sv2v_reg  <= data_i[45];
    end 
    if(N10421) begin
      \nz.mem_4044_sv2v_reg  <= data_i[44];
    end 
    if(N10420) begin
      \nz.mem_4043_sv2v_reg  <= data_i[43];
    end 
    if(N10419) begin
      \nz.mem_4042_sv2v_reg  <= data_i[42];
    end 
    if(N10418) begin
      \nz.mem_4041_sv2v_reg  <= data_i[41];
    end 
    if(N10417) begin
      \nz.mem_4040_sv2v_reg  <= data_i[40];
    end 
    if(N10416) begin
      \nz.mem_4039_sv2v_reg  <= data_i[39];
    end 
    if(N10415) begin
      \nz.mem_4038_sv2v_reg  <= data_i[38];
    end 
    if(N10414) begin
      \nz.mem_4037_sv2v_reg  <= data_i[37];
    end 
    if(N10413) begin
      \nz.mem_4036_sv2v_reg  <= data_i[36];
    end 
    if(N10412) begin
      \nz.mem_4035_sv2v_reg  <= data_i[35];
    end 
    if(N10411) begin
      \nz.mem_4034_sv2v_reg  <= data_i[34];
    end 
    if(N10410) begin
      \nz.mem_4033_sv2v_reg  <= data_i[33];
    end 
    if(N10409) begin
      \nz.mem_4032_sv2v_reg  <= data_i[32];
    end 
    if(N10408) begin
      \nz.mem_4031_sv2v_reg  <= data_i[31];
    end 
    if(N10407) begin
      \nz.mem_4030_sv2v_reg  <= data_i[30];
    end 
    if(N10406) begin
      \nz.mem_4029_sv2v_reg  <= data_i[29];
    end 
    if(N10405) begin
      \nz.mem_4028_sv2v_reg  <= data_i[28];
    end 
    if(N10404) begin
      \nz.mem_4027_sv2v_reg  <= data_i[27];
    end 
    if(N10403) begin
      \nz.mem_4026_sv2v_reg  <= data_i[26];
    end 
    if(N10402) begin
      \nz.mem_4025_sv2v_reg  <= data_i[25];
    end 
    if(N10401) begin
      \nz.mem_4024_sv2v_reg  <= data_i[24];
    end 
    if(N10400) begin
      \nz.mem_4023_sv2v_reg  <= data_i[23];
    end 
    if(N10399) begin
      \nz.mem_4022_sv2v_reg  <= data_i[22];
    end 
    if(N10398) begin
      \nz.mem_4021_sv2v_reg  <= data_i[21];
    end 
    if(N10397) begin
      \nz.mem_4020_sv2v_reg  <= data_i[20];
    end 
    if(N10396) begin
      \nz.mem_4019_sv2v_reg  <= data_i[19];
    end 
    if(N10395) begin
      \nz.mem_4018_sv2v_reg  <= data_i[18];
    end 
    if(N10394) begin
      \nz.mem_4017_sv2v_reg  <= data_i[17];
    end 
    if(N10393) begin
      \nz.mem_4016_sv2v_reg  <= data_i[16];
    end 
    if(N10392) begin
      \nz.mem_4015_sv2v_reg  <= data_i[15];
    end 
    if(N10391) begin
      \nz.mem_4014_sv2v_reg  <= data_i[14];
    end 
    if(N10390) begin
      \nz.mem_4013_sv2v_reg  <= data_i[13];
    end 
    if(N10389) begin
      \nz.mem_4012_sv2v_reg  <= data_i[12];
    end 
    if(N10388) begin
      \nz.mem_4011_sv2v_reg  <= data_i[11];
    end 
    if(N10387) begin
      \nz.mem_4010_sv2v_reg  <= data_i[10];
    end 
    if(N10386) begin
      \nz.mem_4009_sv2v_reg  <= data_i[9];
    end 
    if(N10385) begin
      \nz.mem_4008_sv2v_reg  <= data_i[8];
    end 
    if(N10384) begin
      \nz.mem_4007_sv2v_reg  <= data_i[7];
    end 
    if(N10383) begin
      \nz.mem_4006_sv2v_reg  <= data_i[6];
    end 
    if(N10382) begin
      \nz.mem_4005_sv2v_reg  <= data_i[5];
    end 
    if(N10381) begin
      \nz.mem_4004_sv2v_reg  <= data_i[4];
    end 
    if(N10380) begin
      \nz.mem_4003_sv2v_reg  <= data_i[3];
    end 
    if(N10379) begin
      \nz.mem_4002_sv2v_reg  <= data_i[2];
    end 
    if(N10378) begin
      \nz.mem_4001_sv2v_reg  <= data_i[1];
    end 
    if(N10377) begin
      \nz.mem_4000_sv2v_reg  <= data_i[0];
    end 
    if(N10376) begin
      \nz.mem_3999_sv2v_reg  <= data_i[79];
    end 
    if(N10375) begin
      \nz.mem_3998_sv2v_reg  <= data_i[78];
    end 
    if(N10374) begin
      \nz.mem_3997_sv2v_reg  <= data_i[77];
    end 
    if(N10373) begin
      \nz.mem_3996_sv2v_reg  <= data_i[76];
    end 
    if(N10372) begin
      \nz.mem_3995_sv2v_reg  <= data_i[75];
    end 
    if(N10371) begin
      \nz.mem_3994_sv2v_reg  <= data_i[74];
    end 
    if(N10370) begin
      \nz.mem_3993_sv2v_reg  <= data_i[73];
    end 
    if(N10369) begin
      \nz.mem_3992_sv2v_reg  <= data_i[72];
    end 
    if(N10368) begin
      \nz.mem_3991_sv2v_reg  <= data_i[71];
    end 
    if(N10367) begin
      \nz.mem_3990_sv2v_reg  <= data_i[70];
    end 
    if(N10366) begin
      \nz.mem_3989_sv2v_reg  <= data_i[69];
    end 
    if(N10365) begin
      \nz.mem_3988_sv2v_reg  <= data_i[68];
    end 
    if(N10364) begin
      \nz.mem_3987_sv2v_reg  <= data_i[67];
    end 
    if(N10363) begin
      \nz.mem_3986_sv2v_reg  <= data_i[66];
    end 
    if(N10362) begin
      \nz.mem_3985_sv2v_reg  <= data_i[65];
    end 
    if(N10361) begin
      \nz.mem_3984_sv2v_reg  <= data_i[64];
    end 
    if(N10360) begin
      \nz.mem_3983_sv2v_reg  <= data_i[63];
    end 
    if(N10359) begin
      \nz.mem_3982_sv2v_reg  <= data_i[62];
    end 
    if(N10358) begin
      \nz.mem_3981_sv2v_reg  <= data_i[61];
    end 
    if(N10357) begin
      \nz.mem_3980_sv2v_reg  <= data_i[60];
    end 
    if(N10356) begin
      \nz.mem_3979_sv2v_reg  <= data_i[59];
    end 
    if(N10355) begin
      \nz.mem_3978_sv2v_reg  <= data_i[58];
    end 
    if(N10354) begin
      \nz.mem_3977_sv2v_reg  <= data_i[57];
    end 
    if(N10353) begin
      \nz.mem_3976_sv2v_reg  <= data_i[56];
    end 
    if(N10352) begin
      \nz.mem_3975_sv2v_reg  <= data_i[55];
    end 
    if(N10351) begin
      \nz.mem_3974_sv2v_reg  <= data_i[54];
    end 
    if(N10350) begin
      \nz.mem_3973_sv2v_reg  <= data_i[53];
    end 
    if(N10349) begin
      \nz.mem_3972_sv2v_reg  <= data_i[52];
    end 
    if(N10348) begin
      \nz.mem_3971_sv2v_reg  <= data_i[51];
    end 
    if(N10347) begin
      \nz.mem_3970_sv2v_reg  <= data_i[50];
    end 
    if(N10346) begin
      \nz.mem_3969_sv2v_reg  <= data_i[49];
    end 
    if(N10345) begin
      \nz.mem_3968_sv2v_reg  <= data_i[48];
    end 
    if(N10344) begin
      \nz.mem_3967_sv2v_reg  <= data_i[47];
    end 
    if(N10343) begin
      \nz.mem_3966_sv2v_reg  <= data_i[46];
    end 
    if(N10342) begin
      \nz.mem_3965_sv2v_reg  <= data_i[45];
    end 
    if(N10341) begin
      \nz.mem_3964_sv2v_reg  <= data_i[44];
    end 
    if(N10340) begin
      \nz.mem_3963_sv2v_reg  <= data_i[43];
    end 
    if(N10339) begin
      \nz.mem_3962_sv2v_reg  <= data_i[42];
    end 
    if(N10338) begin
      \nz.mem_3961_sv2v_reg  <= data_i[41];
    end 
    if(N10337) begin
      \nz.mem_3960_sv2v_reg  <= data_i[40];
    end 
    if(N10336) begin
      \nz.mem_3959_sv2v_reg  <= data_i[39];
    end 
    if(N10335) begin
      \nz.mem_3958_sv2v_reg  <= data_i[38];
    end 
    if(N10334) begin
      \nz.mem_3957_sv2v_reg  <= data_i[37];
    end 
    if(N10333) begin
      \nz.mem_3956_sv2v_reg  <= data_i[36];
    end 
    if(N10332) begin
      \nz.mem_3955_sv2v_reg  <= data_i[35];
    end 
    if(N10331) begin
      \nz.mem_3954_sv2v_reg  <= data_i[34];
    end 
    if(N10330) begin
      \nz.mem_3953_sv2v_reg  <= data_i[33];
    end 
    if(N10329) begin
      \nz.mem_3952_sv2v_reg  <= data_i[32];
    end 
    if(N10328) begin
      \nz.mem_3951_sv2v_reg  <= data_i[31];
    end 
    if(N10327) begin
      \nz.mem_3950_sv2v_reg  <= data_i[30];
    end 
    if(N10326) begin
      \nz.mem_3949_sv2v_reg  <= data_i[29];
    end 
    if(N10325) begin
      \nz.mem_3948_sv2v_reg  <= data_i[28];
    end 
    if(N10324) begin
      \nz.mem_3947_sv2v_reg  <= data_i[27];
    end 
    if(N10323) begin
      \nz.mem_3946_sv2v_reg  <= data_i[26];
    end 
    if(N10322) begin
      \nz.mem_3945_sv2v_reg  <= data_i[25];
    end 
    if(N10321) begin
      \nz.mem_3944_sv2v_reg  <= data_i[24];
    end 
    if(N10320) begin
      \nz.mem_3943_sv2v_reg  <= data_i[23];
    end 
    if(N10319) begin
      \nz.mem_3942_sv2v_reg  <= data_i[22];
    end 
    if(N10318) begin
      \nz.mem_3941_sv2v_reg  <= data_i[21];
    end 
    if(N10317) begin
      \nz.mem_3940_sv2v_reg  <= data_i[20];
    end 
    if(N10316) begin
      \nz.mem_3939_sv2v_reg  <= data_i[19];
    end 
    if(N10315) begin
      \nz.mem_3938_sv2v_reg  <= data_i[18];
    end 
    if(N10314) begin
      \nz.mem_3937_sv2v_reg  <= data_i[17];
    end 
    if(N10313) begin
      \nz.mem_3936_sv2v_reg  <= data_i[16];
    end 
    if(N10312) begin
      \nz.mem_3935_sv2v_reg  <= data_i[15];
    end 
    if(N10311) begin
      \nz.mem_3934_sv2v_reg  <= data_i[14];
    end 
    if(N10310) begin
      \nz.mem_3933_sv2v_reg  <= data_i[13];
    end 
    if(N10309) begin
      \nz.mem_3932_sv2v_reg  <= data_i[12];
    end 
    if(N10308) begin
      \nz.mem_3931_sv2v_reg  <= data_i[11];
    end 
    if(N10307) begin
      \nz.mem_3930_sv2v_reg  <= data_i[10];
    end 
    if(N10306) begin
      \nz.mem_3929_sv2v_reg  <= data_i[9];
    end 
    if(N10305) begin
      \nz.mem_3928_sv2v_reg  <= data_i[8];
    end 
    if(N10304) begin
      \nz.mem_3927_sv2v_reg  <= data_i[7];
    end 
    if(N10303) begin
      \nz.mem_3926_sv2v_reg  <= data_i[6];
    end 
    if(N10302) begin
      \nz.mem_3925_sv2v_reg  <= data_i[5];
    end 
    if(N10301) begin
      \nz.mem_3924_sv2v_reg  <= data_i[4];
    end 
    if(N10300) begin
      \nz.mem_3923_sv2v_reg  <= data_i[3];
    end 
    if(N10299) begin
      \nz.mem_3922_sv2v_reg  <= data_i[2];
    end 
    if(N10298) begin
      \nz.mem_3921_sv2v_reg  <= data_i[1];
    end 
    if(N10297) begin
      \nz.mem_3920_sv2v_reg  <= data_i[0];
    end 
    if(N10296) begin
      \nz.mem_3919_sv2v_reg  <= data_i[79];
    end 
    if(N10295) begin
      \nz.mem_3918_sv2v_reg  <= data_i[78];
    end 
    if(N10294) begin
      \nz.mem_3917_sv2v_reg  <= data_i[77];
    end 
    if(N10293) begin
      \nz.mem_3916_sv2v_reg  <= data_i[76];
    end 
    if(N10292) begin
      \nz.mem_3915_sv2v_reg  <= data_i[75];
    end 
    if(N10291) begin
      \nz.mem_3914_sv2v_reg  <= data_i[74];
    end 
    if(N10290) begin
      \nz.mem_3913_sv2v_reg  <= data_i[73];
    end 
    if(N10289) begin
      \nz.mem_3912_sv2v_reg  <= data_i[72];
    end 
    if(N10288) begin
      \nz.mem_3911_sv2v_reg  <= data_i[71];
    end 
    if(N10287) begin
      \nz.mem_3910_sv2v_reg  <= data_i[70];
    end 
    if(N10286) begin
      \nz.mem_3909_sv2v_reg  <= data_i[69];
    end 
    if(N10285) begin
      \nz.mem_3908_sv2v_reg  <= data_i[68];
    end 
    if(N10284) begin
      \nz.mem_3907_sv2v_reg  <= data_i[67];
    end 
    if(N10283) begin
      \nz.mem_3906_sv2v_reg  <= data_i[66];
    end 
    if(N10282) begin
      \nz.mem_3905_sv2v_reg  <= data_i[65];
    end 
    if(N10281) begin
      \nz.mem_3904_sv2v_reg  <= data_i[64];
    end 
    if(N10280) begin
      \nz.mem_3903_sv2v_reg  <= data_i[63];
    end 
    if(N10279) begin
      \nz.mem_3902_sv2v_reg  <= data_i[62];
    end 
    if(N10278) begin
      \nz.mem_3901_sv2v_reg  <= data_i[61];
    end 
    if(N10277) begin
      \nz.mem_3900_sv2v_reg  <= data_i[60];
    end 
    if(N10276) begin
      \nz.mem_3899_sv2v_reg  <= data_i[59];
    end 
    if(N10275) begin
      \nz.mem_3898_sv2v_reg  <= data_i[58];
    end 
    if(N10274) begin
      \nz.mem_3897_sv2v_reg  <= data_i[57];
    end 
    if(N10273) begin
      \nz.mem_3896_sv2v_reg  <= data_i[56];
    end 
    if(N10272) begin
      \nz.mem_3895_sv2v_reg  <= data_i[55];
    end 
    if(N10271) begin
      \nz.mem_3894_sv2v_reg  <= data_i[54];
    end 
    if(N10270) begin
      \nz.mem_3893_sv2v_reg  <= data_i[53];
    end 
    if(N10269) begin
      \nz.mem_3892_sv2v_reg  <= data_i[52];
    end 
    if(N10268) begin
      \nz.mem_3891_sv2v_reg  <= data_i[51];
    end 
    if(N10267) begin
      \nz.mem_3890_sv2v_reg  <= data_i[50];
    end 
    if(N10266) begin
      \nz.mem_3889_sv2v_reg  <= data_i[49];
    end 
    if(N10265) begin
      \nz.mem_3888_sv2v_reg  <= data_i[48];
    end 
    if(N10264) begin
      \nz.mem_3887_sv2v_reg  <= data_i[47];
    end 
    if(N10263) begin
      \nz.mem_3886_sv2v_reg  <= data_i[46];
    end 
    if(N10262) begin
      \nz.mem_3885_sv2v_reg  <= data_i[45];
    end 
    if(N10261) begin
      \nz.mem_3884_sv2v_reg  <= data_i[44];
    end 
    if(N10260) begin
      \nz.mem_3883_sv2v_reg  <= data_i[43];
    end 
    if(N10259) begin
      \nz.mem_3882_sv2v_reg  <= data_i[42];
    end 
    if(N10258) begin
      \nz.mem_3881_sv2v_reg  <= data_i[41];
    end 
    if(N10257) begin
      \nz.mem_3880_sv2v_reg  <= data_i[40];
    end 
    if(N10256) begin
      \nz.mem_3879_sv2v_reg  <= data_i[39];
    end 
    if(N10255) begin
      \nz.mem_3878_sv2v_reg  <= data_i[38];
    end 
    if(N10254) begin
      \nz.mem_3877_sv2v_reg  <= data_i[37];
    end 
    if(N10253) begin
      \nz.mem_3876_sv2v_reg  <= data_i[36];
    end 
    if(N10252) begin
      \nz.mem_3875_sv2v_reg  <= data_i[35];
    end 
    if(N10251) begin
      \nz.mem_3874_sv2v_reg  <= data_i[34];
    end 
    if(N10250) begin
      \nz.mem_3873_sv2v_reg  <= data_i[33];
    end 
    if(N10249) begin
      \nz.mem_3872_sv2v_reg  <= data_i[32];
    end 
    if(N10248) begin
      \nz.mem_3871_sv2v_reg  <= data_i[31];
    end 
    if(N10247) begin
      \nz.mem_3870_sv2v_reg  <= data_i[30];
    end 
    if(N10246) begin
      \nz.mem_3869_sv2v_reg  <= data_i[29];
    end 
    if(N10245) begin
      \nz.mem_3868_sv2v_reg  <= data_i[28];
    end 
    if(N10244) begin
      \nz.mem_3867_sv2v_reg  <= data_i[27];
    end 
    if(N10243) begin
      \nz.mem_3866_sv2v_reg  <= data_i[26];
    end 
    if(N10242) begin
      \nz.mem_3865_sv2v_reg  <= data_i[25];
    end 
    if(N10241) begin
      \nz.mem_3864_sv2v_reg  <= data_i[24];
    end 
    if(N10240) begin
      \nz.mem_3863_sv2v_reg  <= data_i[23];
    end 
    if(N10239) begin
      \nz.mem_3862_sv2v_reg  <= data_i[22];
    end 
    if(N10238) begin
      \nz.mem_3861_sv2v_reg  <= data_i[21];
    end 
    if(N10237) begin
      \nz.mem_3860_sv2v_reg  <= data_i[20];
    end 
    if(N10236) begin
      \nz.mem_3859_sv2v_reg  <= data_i[19];
    end 
    if(N10235) begin
      \nz.mem_3858_sv2v_reg  <= data_i[18];
    end 
    if(N10234) begin
      \nz.mem_3857_sv2v_reg  <= data_i[17];
    end 
    if(N10233) begin
      \nz.mem_3856_sv2v_reg  <= data_i[16];
    end 
    if(N10232) begin
      \nz.mem_3855_sv2v_reg  <= data_i[15];
    end 
    if(N10231) begin
      \nz.mem_3854_sv2v_reg  <= data_i[14];
    end 
    if(N10230) begin
      \nz.mem_3853_sv2v_reg  <= data_i[13];
    end 
    if(N10229) begin
      \nz.mem_3852_sv2v_reg  <= data_i[12];
    end 
    if(N10228) begin
      \nz.mem_3851_sv2v_reg  <= data_i[11];
    end 
    if(N10227) begin
      \nz.mem_3850_sv2v_reg  <= data_i[10];
    end 
    if(N10226) begin
      \nz.mem_3849_sv2v_reg  <= data_i[9];
    end 
    if(N10225) begin
      \nz.mem_3848_sv2v_reg  <= data_i[8];
    end 
    if(N10224) begin
      \nz.mem_3847_sv2v_reg  <= data_i[7];
    end 
    if(N10223) begin
      \nz.mem_3846_sv2v_reg  <= data_i[6];
    end 
    if(N10222) begin
      \nz.mem_3845_sv2v_reg  <= data_i[5];
    end 
    if(N10221) begin
      \nz.mem_3844_sv2v_reg  <= data_i[4];
    end 
    if(N10220) begin
      \nz.mem_3843_sv2v_reg  <= data_i[3];
    end 
    if(N10219) begin
      \nz.mem_3842_sv2v_reg  <= data_i[2];
    end 
    if(N10218) begin
      \nz.mem_3841_sv2v_reg  <= data_i[1];
    end 
    if(N10217) begin
      \nz.mem_3840_sv2v_reg  <= data_i[0];
    end 
    if(N10216) begin
      \nz.mem_3839_sv2v_reg  <= data_i[79];
    end 
    if(N10215) begin
      \nz.mem_3838_sv2v_reg  <= data_i[78];
    end 
    if(N10214) begin
      \nz.mem_3837_sv2v_reg  <= data_i[77];
    end 
    if(N10213) begin
      \nz.mem_3836_sv2v_reg  <= data_i[76];
    end 
    if(N10212) begin
      \nz.mem_3835_sv2v_reg  <= data_i[75];
    end 
    if(N10211) begin
      \nz.mem_3834_sv2v_reg  <= data_i[74];
    end 
    if(N10210) begin
      \nz.mem_3833_sv2v_reg  <= data_i[73];
    end 
    if(N10209) begin
      \nz.mem_3832_sv2v_reg  <= data_i[72];
    end 
    if(N10208) begin
      \nz.mem_3831_sv2v_reg  <= data_i[71];
    end 
    if(N10207) begin
      \nz.mem_3830_sv2v_reg  <= data_i[70];
    end 
    if(N10206) begin
      \nz.mem_3829_sv2v_reg  <= data_i[69];
    end 
    if(N10205) begin
      \nz.mem_3828_sv2v_reg  <= data_i[68];
    end 
    if(N10204) begin
      \nz.mem_3827_sv2v_reg  <= data_i[67];
    end 
    if(N10203) begin
      \nz.mem_3826_sv2v_reg  <= data_i[66];
    end 
    if(N10202) begin
      \nz.mem_3825_sv2v_reg  <= data_i[65];
    end 
    if(N10201) begin
      \nz.mem_3824_sv2v_reg  <= data_i[64];
    end 
    if(N10200) begin
      \nz.mem_3823_sv2v_reg  <= data_i[63];
    end 
    if(N10199) begin
      \nz.mem_3822_sv2v_reg  <= data_i[62];
    end 
    if(N10198) begin
      \nz.mem_3821_sv2v_reg  <= data_i[61];
    end 
    if(N10197) begin
      \nz.mem_3820_sv2v_reg  <= data_i[60];
    end 
    if(N10196) begin
      \nz.mem_3819_sv2v_reg  <= data_i[59];
    end 
    if(N10195) begin
      \nz.mem_3818_sv2v_reg  <= data_i[58];
    end 
    if(N10194) begin
      \nz.mem_3817_sv2v_reg  <= data_i[57];
    end 
    if(N10193) begin
      \nz.mem_3816_sv2v_reg  <= data_i[56];
    end 
    if(N10192) begin
      \nz.mem_3815_sv2v_reg  <= data_i[55];
    end 
    if(N10191) begin
      \nz.mem_3814_sv2v_reg  <= data_i[54];
    end 
    if(N10190) begin
      \nz.mem_3813_sv2v_reg  <= data_i[53];
    end 
    if(N10189) begin
      \nz.mem_3812_sv2v_reg  <= data_i[52];
    end 
    if(N10188) begin
      \nz.mem_3811_sv2v_reg  <= data_i[51];
    end 
    if(N10187) begin
      \nz.mem_3810_sv2v_reg  <= data_i[50];
    end 
    if(N10186) begin
      \nz.mem_3809_sv2v_reg  <= data_i[49];
    end 
    if(N10185) begin
      \nz.mem_3808_sv2v_reg  <= data_i[48];
    end 
    if(N10184) begin
      \nz.mem_3807_sv2v_reg  <= data_i[47];
    end 
    if(N10183) begin
      \nz.mem_3806_sv2v_reg  <= data_i[46];
    end 
    if(N10182) begin
      \nz.mem_3805_sv2v_reg  <= data_i[45];
    end 
    if(N10181) begin
      \nz.mem_3804_sv2v_reg  <= data_i[44];
    end 
    if(N10180) begin
      \nz.mem_3803_sv2v_reg  <= data_i[43];
    end 
    if(N10179) begin
      \nz.mem_3802_sv2v_reg  <= data_i[42];
    end 
    if(N10178) begin
      \nz.mem_3801_sv2v_reg  <= data_i[41];
    end 
    if(N10177) begin
      \nz.mem_3800_sv2v_reg  <= data_i[40];
    end 
    if(N10176) begin
      \nz.mem_3799_sv2v_reg  <= data_i[39];
    end 
    if(N10175) begin
      \nz.mem_3798_sv2v_reg  <= data_i[38];
    end 
    if(N10174) begin
      \nz.mem_3797_sv2v_reg  <= data_i[37];
    end 
    if(N10173) begin
      \nz.mem_3796_sv2v_reg  <= data_i[36];
    end 
    if(N10172) begin
      \nz.mem_3795_sv2v_reg  <= data_i[35];
    end 
    if(N10171) begin
      \nz.mem_3794_sv2v_reg  <= data_i[34];
    end 
    if(N10170) begin
      \nz.mem_3793_sv2v_reg  <= data_i[33];
    end 
    if(N10169) begin
      \nz.mem_3792_sv2v_reg  <= data_i[32];
    end 
    if(N10168) begin
      \nz.mem_3791_sv2v_reg  <= data_i[31];
    end 
    if(N10167) begin
      \nz.mem_3790_sv2v_reg  <= data_i[30];
    end 
    if(N10166) begin
      \nz.mem_3789_sv2v_reg  <= data_i[29];
    end 
    if(N10165) begin
      \nz.mem_3788_sv2v_reg  <= data_i[28];
    end 
    if(N10164) begin
      \nz.mem_3787_sv2v_reg  <= data_i[27];
    end 
    if(N10163) begin
      \nz.mem_3786_sv2v_reg  <= data_i[26];
    end 
    if(N10162) begin
      \nz.mem_3785_sv2v_reg  <= data_i[25];
    end 
    if(N10161) begin
      \nz.mem_3784_sv2v_reg  <= data_i[24];
    end 
    if(N10160) begin
      \nz.mem_3783_sv2v_reg  <= data_i[23];
    end 
    if(N10159) begin
      \nz.mem_3782_sv2v_reg  <= data_i[22];
    end 
    if(N10158) begin
      \nz.mem_3781_sv2v_reg  <= data_i[21];
    end 
    if(N10157) begin
      \nz.mem_3780_sv2v_reg  <= data_i[20];
    end 
    if(N10156) begin
      \nz.mem_3779_sv2v_reg  <= data_i[19];
    end 
    if(N10155) begin
      \nz.mem_3778_sv2v_reg  <= data_i[18];
    end 
    if(N10154) begin
      \nz.mem_3777_sv2v_reg  <= data_i[17];
    end 
    if(N10153) begin
      \nz.mem_3776_sv2v_reg  <= data_i[16];
    end 
    if(N10152) begin
      \nz.mem_3775_sv2v_reg  <= data_i[15];
    end 
    if(N10151) begin
      \nz.mem_3774_sv2v_reg  <= data_i[14];
    end 
    if(N10150) begin
      \nz.mem_3773_sv2v_reg  <= data_i[13];
    end 
    if(N10149) begin
      \nz.mem_3772_sv2v_reg  <= data_i[12];
    end 
    if(N10148) begin
      \nz.mem_3771_sv2v_reg  <= data_i[11];
    end 
    if(N10147) begin
      \nz.mem_3770_sv2v_reg  <= data_i[10];
    end 
    if(N10146) begin
      \nz.mem_3769_sv2v_reg  <= data_i[9];
    end 
    if(N10145) begin
      \nz.mem_3768_sv2v_reg  <= data_i[8];
    end 
    if(N10144) begin
      \nz.mem_3767_sv2v_reg  <= data_i[7];
    end 
    if(N10143) begin
      \nz.mem_3766_sv2v_reg  <= data_i[6];
    end 
    if(N10142) begin
      \nz.mem_3765_sv2v_reg  <= data_i[5];
    end 
    if(N10141) begin
      \nz.mem_3764_sv2v_reg  <= data_i[4];
    end 
    if(N10140) begin
      \nz.mem_3763_sv2v_reg  <= data_i[3];
    end 
    if(N10139) begin
      \nz.mem_3762_sv2v_reg  <= data_i[2];
    end 
    if(N10138) begin
      \nz.mem_3761_sv2v_reg  <= data_i[1];
    end 
    if(N10137) begin
      \nz.mem_3760_sv2v_reg  <= data_i[0];
    end 
    if(N10136) begin
      \nz.mem_3759_sv2v_reg  <= data_i[79];
    end 
    if(N10135) begin
      \nz.mem_3758_sv2v_reg  <= data_i[78];
    end 
    if(N10134) begin
      \nz.mem_3757_sv2v_reg  <= data_i[77];
    end 
    if(N10133) begin
      \nz.mem_3756_sv2v_reg  <= data_i[76];
    end 
    if(N10132) begin
      \nz.mem_3755_sv2v_reg  <= data_i[75];
    end 
    if(N10131) begin
      \nz.mem_3754_sv2v_reg  <= data_i[74];
    end 
    if(N10130) begin
      \nz.mem_3753_sv2v_reg  <= data_i[73];
    end 
    if(N10129) begin
      \nz.mem_3752_sv2v_reg  <= data_i[72];
    end 
    if(N10128) begin
      \nz.mem_3751_sv2v_reg  <= data_i[71];
    end 
    if(N10127) begin
      \nz.mem_3750_sv2v_reg  <= data_i[70];
    end 
    if(N10126) begin
      \nz.mem_3749_sv2v_reg  <= data_i[69];
    end 
    if(N10125) begin
      \nz.mem_3748_sv2v_reg  <= data_i[68];
    end 
    if(N10124) begin
      \nz.mem_3747_sv2v_reg  <= data_i[67];
    end 
    if(N10123) begin
      \nz.mem_3746_sv2v_reg  <= data_i[66];
    end 
    if(N10122) begin
      \nz.mem_3745_sv2v_reg  <= data_i[65];
    end 
    if(N10121) begin
      \nz.mem_3744_sv2v_reg  <= data_i[64];
    end 
    if(N10120) begin
      \nz.mem_3743_sv2v_reg  <= data_i[63];
    end 
    if(N10119) begin
      \nz.mem_3742_sv2v_reg  <= data_i[62];
    end 
    if(N10118) begin
      \nz.mem_3741_sv2v_reg  <= data_i[61];
    end 
    if(N10117) begin
      \nz.mem_3740_sv2v_reg  <= data_i[60];
    end 
    if(N10116) begin
      \nz.mem_3739_sv2v_reg  <= data_i[59];
    end 
    if(N10115) begin
      \nz.mem_3738_sv2v_reg  <= data_i[58];
    end 
    if(N10114) begin
      \nz.mem_3737_sv2v_reg  <= data_i[57];
    end 
    if(N10113) begin
      \nz.mem_3736_sv2v_reg  <= data_i[56];
    end 
    if(N10112) begin
      \nz.mem_3735_sv2v_reg  <= data_i[55];
    end 
    if(N10111) begin
      \nz.mem_3734_sv2v_reg  <= data_i[54];
    end 
    if(N10110) begin
      \nz.mem_3733_sv2v_reg  <= data_i[53];
    end 
    if(N10109) begin
      \nz.mem_3732_sv2v_reg  <= data_i[52];
    end 
    if(N10108) begin
      \nz.mem_3731_sv2v_reg  <= data_i[51];
    end 
    if(N10107) begin
      \nz.mem_3730_sv2v_reg  <= data_i[50];
    end 
    if(N10106) begin
      \nz.mem_3729_sv2v_reg  <= data_i[49];
    end 
    if(N10105) begin
      \nz.mem_3728_sv2v_reg  <= data_i[48];
    end 
    if(N10104) begin
      \nz.mem_3727_sv2v_reg  <= data_i[47];
    end 
    if(N10103) begin
      \nz.mem_3726_sv2v_reg  <= data_i[46];
    end 
    if(N10102) begin
      \nz.mem_3725_sv2v_reg  <= data_i[45];
    end 
    if(N10101) begin
      \nz.mem_3724_sv2v_reg  <= data_i[44];
    end 
    if(N10100) begin
      \nz.mem_3723_sv2v_reg  <= data_i[43];
    end 
    if(N10099) begin
      \nz.mem_3722_sv2v_reg  <= data_i[42];
    end 
    if(N10098) begin
      \nz.mem_3721_sv2v_reg  <= data_i[41];
    end 
    if(N10097) begin
      \nz.mem_3720_sv2v_reg  <= data_i[40];
    end 
    if(N10096) begin
      \nz.mem_3719_sv2v_reg  <= data_i[39];
    end 
    if(N10095) begin
      \nz.mem_3718_sv2v_reg  <= data_i[38];
    end 
    if(N10094) begin
      \nz.mem_3717_sv2v_reg  <= data_i[37];
    end 
    if(N10093) begin
      \nz.mem_3716_sv2v_reg  <= data_i[36];
    end 
    if(N10092) begin
      \nz.mem_3715_sv2v_reg  <= data_i[35];
    end 
    if(N10091) begin
      \nz.mem_3714_sv2v_reg  <= data_i[34];
    end 
    if(N10090) begin
      \nz.mem_3713_sv2v_reg  <= data_i[33];
    end 
    if(N10089) begin
      \nz.mem_3712_sv2v_reg  <= data_i[32];
    end 
    if(N10088) begin
      \nz.mem_3711_sv2v_reg  <= data_i[31];
    end 
    if(N10087) begin
      \nz.mem_3710_sv2v_reg  <= data_i[30];
    end 
    if(N10086) begin
      \nz.mem_3709_sv2v_reg  <= data_i[29];
    end 
    if(N10085) begin
      \nz.mem_3708_sv2v_reg  <= data_i[28];
    end 
    if(N10084) begin
      \nz.mem_3707_sv2v_reg  <= data_i[27];
    end 
    if(N10083) begin
      \nz.mem_3706_sv2v_reg  <= data_i[26];
    end 
    if(N10082) begin
      \nz.mem_3705_sv2v_reg  <= data_i[25];
    end 
    if(N10081) begin
      \nz.mem_3704_sv2v_reg  <= data_i[24];
    end 
    if(N10080) begin
      \nz.mem_3703_sv2v_reg  <= data_i[23];
    end 
    if(N10079) begin
      \nz.mem_3702_sv2v_reg  <= data_i[22];
    end 
    if(N10078) begin
      \nz.mem_3701_sv2v_reg  <= data_i[21];
    end 
    if(N10077) begin
      \nz.mem_3700_sv2v_reg  <= data_i[20];
    end 
    if(N10076) begin
      \nz.mem_3699_sv2v_reg  <= data_i[19];
    end 
    if(N10075) begin
      \nz.mem_3698_sv2v_reg  <= data_i[18];
    end 
    if(N10074) begin
      \nz.mem_3697_sv2v_reg  <= data_i[17];
    end 
    if(N10073) begin
      \nz.mem_3696_sv2v_reg  <= data_i[16];
    end 
    if(N10072) begin
      \nz.mem_3695_sv2v_reg  <= data_i[15];
    end 
    if(N10071) begin
      \nz.mem_3694_sv2v_reg  <= data_i[14];
    end 
    if(N10070) begin
      \nz.mem_3693_sv2v_reg  <= data_i[13];
    end 
    if(N10069) begin
      \nz.mem_3692_sv2v_reg  <= data_i[12];
    end 
    if(N10068) begin
      \nz.mem_3691_sv2v_reg  <= data_i[11];
    end 
    if(N10067) begin
      \nz.mem_3690_sv2v_reg  <= data_i[10];
    end 
    if(N10066) begin
      \nz.mem_3689_sv2v_reg  <= data_i[9];
    end 
    if(N10065) begin
      \nz.mem_3688_sv2v_reg  <= data_i[8];
    end 
    if(N10064) begin
      \nz.mem_3687_sv2v_reg  <= data_i[7];
    end 
    if(N10063) begin
      \nz.mem_3686_sv2v_reg  <= data_i[6];
    end 
    if(N10062) begin
      \nz.mem_3685_sv2v_reg  <= data_i[5];
    end 
    if(N10061) begin
      \nz.mem_3684_sv2v_reg  <= data_i[4];
    end 
    if(N10060) begin
      \nz.mem_3683_sv2v_reg  <= data_i[3];
    end 
    if(N10059) begin
      \nz.mem_3682_sv2v_reg  <= data_i[2];
    end 
    if(N10058) begin
      \nz.mem_3681_sv2v_reg  <= data_i[1];
    end 
    if(N10057) begin
      \nz.mem_3680_sv2v_reg  <= data_i[0];
    end 
    if(N10056) begin
      \nz.mem_3679_sv2v_reg  <= data_i[79];
    end 
    if(N10055) begin
      \nz.mem_3678_sv2v_reg  <= data_i[78];
    end 
    if(N10054) begin
      \nz.mem_3677_sv2v_reg  <= data_i[77];
    end 
    if(N10053) begin
      \nz.mem_3676_sv2v_reg  <= data_i[76];
    end 
    if(N10052) begin
      \nz.mem_3675_sv2v_reg  <= data_i[75];
    end 
    if(N10051) begin
      \nz.mem_3674_sv2v_reg  <= data_i[74];
    end 
    if(N10050) begin
      \nz.mem_3673_sv2v_reg  <= data_i[73];
    end 
    if(N10049) begin
      \nz.mem_3672_sv2v_reg  <= data_i[72];
    end 
    if(N10048) begin
      \nz.mem_3671_sv2v_reg  <= data_i[71];
    end 
    if(N10047) begin
      \nz.mem_3670_sv2v_reg  <= data_i[70];
    end 
    if(N10046) begin
      \nz.mem_3669_sv2v_reg  <= data_i[69];
    end 
    if(N10045) begin
      \nz.mem_3668_sv2v_reg  <= data_i[68];
    end 
    if(N10044) begin
      \nz.mem_3667_sv2v_reg  <= data_i[67];
    end 
    if(N10043) begin
      \nz.mem_3666_sv2v_reg  <= data_i[66];
    end 
    if(N10042) begin
      \nz.mem_3665_sv2v_reg  <= data_i[65];
    end 
    if(N10041) begin
      \nz.mem_3664_sv2v_reg  <= data_i[64];
    end 
    if(N10040) begin
      \nz.mem_3663_sv2v_reg  <= data_i[63];
    end 
    if(N10039) begin
      \nz.mem_3662_sv2v_reg  <= data_i[62];
    end 
    if(N10038) begin
      \nz.mem_3661_sv2v_reg  <= data_i[61];
    end 
    if(N10037) begin
      \nz.mem_3660_sv2v_reg  <= data_i[60];
    end 
    if(N10036) begin
      \nz.mem_3659_sv2v_reg  <= data_i[59];
    end 
    if(N10035) begin
      \nz.mem_3658_sv2v_reg  <= data_i[58];
    end 
    if(N10034) begin
      \nz.mem_3657_sv2v_reg  <= data_i[57];
    end 
    if(N10033) begin
      \nz.mem_3656_sv2v_reg  <= data_i[56];
    end 
    if(N10032) begin
      \nz.mem_3655_sv2v_reg  <= data_i[55];
    end 
    if(N10031) begin
      \nz.mem_3654_sv2v_reg  <= data_i[54];
    end 
    if(N10030) begin
      \nz.mem_3653_sv2v_reg  <= data_i[53];
    end 
    if(N10029) begin
      \nz.mem_3652_sv2v_reg  <= data_i[52];
    end 
    if(N10028) begin
      \nz.mem_3651_sv2v_reg  <= data_i[51];
    end 
    if(N10027) begin
      \nz.mem_3650_sv2v_reg  <= data_i[50];
    end 
    if(N10026) begin
      \nz.mem_3649_sv2v_reg  <= data_i[49];
    end 
    if(N10025) begin
      \nz.mem_3648_sv2v_reg  <= data_i[48];
    end 
    if(N10024) begin
      \nz.mem_3647_sv2v_reg  <= data_i[47];
    end 
    if(N10023) begin
      \nz.mem_3646_sv2v_reg  <= data_i[46];
    end 
    if(N10022) begin
      \nz.mem_3645_sv2v_reg  <= data_i[45];
    end 
    if(N10021) begin
      \nz.mem_3644_sv2v_reg  <= data_i[44];
    end 
    if(N10020) begin
      \nz.mem_3643_sv2v_reg  <= data_i[43];
    end 
    if(N10019) begin
      \nz.mem_3642_sv2v_reg  <= data_i[42];
    end 
    if(N10018) begin
      \nz.mem_3641_sv2v_reg  <= data_i[41];
    end 
    if(N10017) begin
      \nz.mem_3640_sv2v_reg  <= data_i[40];
    end 
    if(N10016) begin
      \nz.mem_3639_sv2v_reg  <= data_i[39];
    end 
    if(N10015) begin
      \nz.mem_3638_sv2v_reg  <= data_i[38];
    end 
    if(N10014) begin
      \nz.mem_3637_sv2v_reg  <= data_i[37];
    end 
    if(N10013) begin
      \nz.mem_3636_sv2v_reg  <= data_i[36];
    end 
    if(N10012) begin
      \nz.mem_3635_sv2v_reg  <= data_i[35];
    end 
    if(N10011) begin
      \nz.mem_3634_sv2v_reg  <= data_i[34];
    end 
    if(N10010) begin
      \nz.mem_3633_sv2v_reg  <= data_i[33];
    end 
    if(N10009) begin
      \nz.mem_3632_sv2v_reg  <= data_i[32];
    end 
    if(N10008) begin
      \nz.mem_3631_sv2v_reg  <= data_i[31];
    end 
    if(N10007) begin
      \nz.mem_3630_sv2v_reg  <= data_i[30];
    end 
    if(N10006) begin
      \nz.mem_3629_sv2v_reg  <= data_i[29];
    end 
    if(N10005) begin
      \nz.mem_3628_sv2v_reg  <= data_i[28];
    end 
    if(N10004) begin
      \nz.mem_3627_sv2v_reg  <= data_i[27];
    end 
    if(N10003) begin
      \nz.mem_3626_sv2v_reg  <= data_i[26];
    end 
    if(N10002) begin
      \nz.mem_3625_sv2v_reg  <= data_i[25];
    end 
    if(N10001) begin
      \nz.mem_3624_sv2v_reg  <= data_i[24];
    end 
    if(N10000) begin
      \nz.mem_3623_sv2v_reg  <= data_i[23];
    end 
    if(N9999) begin
      \nz.mem_3622_sv2v_reg  <= data_i[22];
    end 
    if(N9998) begin
      \nz.mem_3621_sv2v_reg  <= data_i[21];
    end 
    if(N9997) begin
      \nz.mem_3620_sv2v_reg  <= data_i[20];
    end 
    if(N9996) begin
      \nz.mem_3619_sv2v_reg  <= data_i[19];
    end 
    if(N9995) begin
      \nz.mem_3618_sv2v_reg  <= data_i[18];
    end 
    if(N9994) begin
      \nz.mem_3617_sv2v_reg  <= data_i[17];
    end 
    if(N9993) begin
      \nz.mem_3616_sv2v_reg  <= data_i[16];
    end 
    if(N9992) begin
      \nz.mem_3615_sv2v_reg  <= data_i[15];
    end 
    if(N9991) begin
      \nz.mem_3614_sv2v_reg  <= data_i[14];
    end 
    if(N9990) begin
      \nz.mem_3613_sv2v_reg  <= data_i[13];
    end 
    if(N9989) begin
      \nz.mem_3612_sv2v_reg  <= data_i[12];
    end 
    if(N9988) begin
      \nz.mem_3611_sv2v_reg  <= data_i[11];
    end 
    if(N9987) begin
      \nz.mem_3610_sv2v_reg  <= data_i[10];
    end 
    if(N9986) begin
      \nz.mem_3609_sv2v_reg  <= data_i[9];
    end 
    if(N9985) begin
      \nz.mem_3608_sv2v_reg  <= data_i[8];
    end 
    if(N9984) begin
      \nz.mem_3607_sv2v_reg  <= data_i[7];
    end 
    if(N9983) begin
      \nz.mem_3606_sv2v_reg  <= data_i[6];
    end 
    if(N9982) begin
      \nz.mem_3605_sv2v_reg  <= data_i[5];
    end 
    if(N9981) begin
      \nz.mem_3604_sv2v_reg  <= data_i[4];
    end 
    if(N9980) begin
      \nz.mem_3603_sv2v_reg  <= data_i[3];
    end 
    if(N9979) begin
      \nz.mem_3602_sv2v_reg  <= data_i[2];
    end 
    if(N9978) begin
      \nz.mem_3601_sv2v_reg  <= data_i[1];
    end 
    if(N9977) begin
      \nz.mem_3600_sv2v_reg  <= data_i[0];
    end 
    if(N9976) begin
      \nz.mem_3599_sv2v_reg  <= data_i[79];
    end 
    if(N9975) begin
      \nz.mem_3598_sv2v_reg  <= data_i[78];
    end 
    if(N9974) begin
      \nz.mem_3597_sv2v_reg  <= data_i[77];
    end 
    if(N9973) begin
      \nz.mem_3596_sv2v_reg  <= data_i[76];
    end 
    if(N9972) begin
      \nz.mem_3595_sv2v_reg  <= data_i[75];
    end 
    if(N9971) begin
      \nz.mem_3594_sv2v_reg  <= data_i[74];
    end 
    if(N9970) begin
      \nz.mem_3593_sv2v_reg  <= data_i[73];
    end 
    if(N9969) begin
      \nz.mem_3592_sv2v_reg  <= data_i[72];
    end 
    if(N9968) begin
      \nz.mem_3591_sv2v_reg  <= data_i[71];
    end 
    if(N9967) begin
      \nz.mem_3590_sv2v_reg  <= data_i[70];
    end 
    if(N9966) begin
      \nz.mem_3589_sv2v_reg  <= data_i[69];
    end 
    if(N9965) begin
      \nz.mem_3588_sv2v_reg  <= data_i[68];
    end 
    if(N9964) begin
      \nz.mem_3587_sv2v_reg  <= data_i[67];
    end 
    if(N9963) begin
      \nz.mem_3586_sv2v_reg  <= data_i[66];
    end 
    if(N9962) begin
      \nz.mem_3585_sv2v_reg  <= data_i[65];
    end 
    if(N9961) begin
      \nz.mem_3584_sv2v_reg  <= data_i[64];
    end 
    if(N9960) begin
      \nz.mem_3583_sv2v_reg  <= data_i[63];
    end 
    if(N9959) begin
      \nz.mem_3582_sv2v_reg  <= data_i[62];
    end 
    if(N9958) begin
      \nz.mem_3581_sv2v_reg  <= data_i[61];
    end 
    if(N9957) begin
      \nz.mem_3580_sv2v_reg  <= data_i[60];
    end 
    if(N9956) begin
      \nz.mem_3579_sv2v_reg  <= data_i[59];
    end 
    if(N9955) begin
      \nz.mem_3578_sv2v_reg  <= data_i[58];
    end 
    if(N9954) begin
      \nz.mem_3577_sv2v_reg  <= data_i[57];
    end 
    if(N9953) begin
      \nz.mem_3576_sv2v_reg  <= data_i[56];
    end 
    if(N9952) begin
      \nz.mem_3575_sv2v_reg  <= data_i[55];
    end 
    if(N9951) begin
      \nz.mem_3574_sv2v_reg  <= data_i[54];
    end 
    if(N9950) begin
      \nz.mem_3573_sv2v_reg  <= data_i[53];
    end 
    if(N9949) begin
      \nz.mem_3572_sv2v_reg  <= data_i[52];
    end 
    if(N9948) begin
      \nz.mem_3571_sv2v_reg  <= data_i[51];
    end 
    if(N9947) begin
      \nz.mem_3570_sv2v_reg  <= data_i[50];
    end 
    if(N9946) begin
      \nz.mem_3569_sv2v_reg  <= data_i[49];
    end 
    if(N9945) begin
      \nz.mem_3568_sv2v_reg  <= data_i[48];
    end 
    if(N9944) begin
      \nz.mem_3567_sv2v_reg  <= data_i[47];
    end 
    if(N9943) begin
      \nz.mem_3566_sv2v_reg  <= data_i[46];
    end 
    if(N9942) begin
      \nz.mem_3565_sv2v_reg  <= data_i[45];
    end 
    if(N9941) begin
      \nz.mem_3564_sv2v_reg  <= data_i[44];
    end 
    if(N9940) begin
      \nz.mem_3563_sv2v_reg  <= data_i[43];
    end 
    if(N9939) begin
      \nz.mem_3562_sv2v_reg  <= data_i[42];
    end 
    if(N9938) begin
      \nz.mem_3561_sv2v_reg  <= data_i[41];
    end 
    if(N9937) begin
      \nz.mem_3560_sv2v_reg  <= data_i[40];
    end 
    if(N9936) begin
      \nz.mem_3559_sv2v_reg  <= data_i[39];
    end 
    if(N9935) begin
      \nz.mem_3558_sv2v_reg  <= data_i[38];
    end 
    if(N9934) begin
      \nz.mem_3557_sv2v_reg  <= data_i[37];
    end 
    if(N9933) begin
      \nz.mem_3556_sv2v_reg  <= data_i[36];
    end 
    if(N9932) begin
      \nz.mem_3555_sv2v_reg  <= data_i[35];
    end 
    if(N9931) begin
      \nz.mem_3554_sv2v_reg  <= data_i[34];
    end 
    if(N9930) begin
      \nz.mem_3553_sv2v_reg  <= data_i[33];
    end 
    if(N9929) begin
      \nz.mem_3552_sv2v_reg  <= data_i[32];
    end 
    if(N9928) begin
      \nz.mem_3551_sv2v_reg  <= data_i[31];
    end 
    if(N9927) begin
      \nz.mem_3550_sv2v_reg  <= data_i[30];
    end 
    if(N9926) begin
      \nz.mem_3549_sv2v_reg  <= data_i[29];
    end 
    if(N9925) begin
      \nz.mem_3548_sv2v_reg  <= data_i[28];
    end 
    if(N9924) begin
      \nz.mem_3547_sv2v_reg  <= data_i[27];
    end 
    if(N9923) begin
      \nz.mem_3546_sv2v_reg  <= data_i[26];
    end 
    if(N9922) begin
      \nz.mem_3545_sv2v_reg  <= data_i[25];
    end 
    if(N9921) begin
      \nz.mem_3544_sv2v_reg  <= data_i[24];
    end 
    if(N9920) begin
      \nz.mem_3543_sv2v_reg  <= data_i[23];
    end 
    if(N9919) begin
      \nz.mem_3542_sv2v_reg  <= data_i[22];
    end 
    if(N9918) begin
      \nz.mem_3541_sv2v_reg  <= data_i[21];
    end 
    if(N9917) begin
      \nz.mem_3540_sv2v_reg  <= data_i[20];
    end 
    if(N9916) begin
      \nz.mem_3539_sv2v_reg  <= data_i[19];
    end 
    if(N9915) begin
      \nz.mem_3538_sv2v_reg  <= data_i[18];
    end 
    if(N9914) begin
      \nz.mem_3537_sv2v_reg  <= data_i[17];
    end 
    if(N9913) begin
      \nz.mem_3536_sv2v_reg  <= data_i[16];
    end 
    if(N9912) begin
      \nz.mem_3535_sv2v_reg  <= data_i[15];
    end 
    if(N9911) begin
      \nz.mem_3534_sv2v_reg  <= data_i[14];
    end 
    if(N9910) begin
      \nz.mem_3533_sv2v_reg  <= data_i[13];
    end 
    if(N9909) begin
      \nz.mem_3532_sv2v_reg  <= data_i[12];
    end 
    if(N9908) begin
      \nz.mem_3531_sv2v_reg  <= data_i[11];
    end 
    if(N9907) begin
      \nz.mem_3530_sv2v_reg  <= data_i[10];
    end 
    if(N9906) begin
      \nz.mem_3529_sv2v_reg  <= data_i[9];
    end 
    if(N9905) begin
      \nz.mem_3528_sv2v_reg  <= data_i[8];
    end 
    if(N9904) begin
      \nz.mem_3527_sv2v_reg  <= data_i[7];
    end 
    if(N9903) begin
      \nz.mem_3526_sv2v_reg  <= data_i[6];
    end 
    if(N9902) begin
      \nz.mem_3525_sv2v_reg  <= data_i[5];
    end 
    if(N9901) begin
      \nz.mem_3524_sv2v_reg  <= data_i[4];
    end 
    if(N9900) begin
      \nz.mem_3523_sv2v_reg  <= data_i[3];
    end 
    if(N9899) begin
      \nz.mem_3522_sv2v_reg  <= data_i[2];
    end 
    if(N9898) begin
      \nz.mem_3521_sv2v_reg  <= data_i[1];
    end 
    if(N9897) begin
      \nz.mem_3520_sv2v_reg  <= data_i[0];
    end 
    if(N9896) begin
      \nz.mem_3519_sv2v_reg  <= data_i[79];
    end 
    if(N9895) begin
      \nz.mem_3518_sv2v_reg  <= data_i[78];
    end 
    if(N9894) begin
      \nz.mem_3517_sv2v_reg  <= data_i[77];
    end 
    if(N9893) begin
      \nz.mem_3516_sv2v_reg  <= data_i[76];
    end 
    if(N9892) begin
      \nz.mem_3515_sv2v_reg  <= data_i[75];
    end 
    if(N9891) begin
      \nz.mem_3514_sv2v_reg  <= data_i[74];
    end 
    if(N9890) begin
      \nz.mem_3513_sv2v_reg  <= data_i[73];
    end 
    if(N9889) begin
      \nz.mem_3512_sv2v_reg  <= data_i[72];
    end 
    if(N9888) begin
      \nz.mem_3511_sv2v_reg  <= data_i[71];
    end 
    if(N9887) begin
      \nz.mem_3510_sv2v_reg  <= data_i[70];
    end 
    if(N9886) begin
      \nz.mem_3509_sv2v_reg  <= data_i[69];
    end 
    if(N9885) begin
      \nz.mem_3508_sv2v_reg  <= data_i[68];
    end 
    if(N9884) begin
      \nz.mem_3507_sv2v_reg  <= data_i[67];
    end 
    if(N9883) begin
      \nz.mem_3506_sv2v_reg  <= data_i[66];
    end 
    if(N9882) begin
      \nz.mem_3505_sv2v_reg  <= data_i[65];
    end 
    if(N9881) begin
      \nz.mem_3504_sv2v_reg  <= data_i[64];
    end 
    if(N9880) begin
      \nz.mem_3503_sv2v_reg  <= data_i[63];
    end 
    if(N9879) begin
      \nz.mem_3502_sv2v_reg  <= data_i[62];
    end 
    if(N9878) begin
      \nz.mem_3501_sv2v_reg  <= data_i[61];
    end 
    if(N9877) begin
      \nz.mem_3500_sv2v_reg  <= data_i[60];
    end 
    if(N9876) begin
      \nz.mem_3499_sv2v_reg  <= data_i[59];
    end 
    if(N9875) begin
      \nz.mem_3498_sv2v_reg  <= data_i[58];
    end 
    if(N9874) begin
      \nz.mem_3497_sv2v_reg  <= data_i[57];
    end 
    if(N9873) begin
      \nz.mem_3496_sv2v_reg  <= data_i[56];
    end 
    if(N9872) begin
      \nz.mem_3495_sv2v_reg  <= data_i[55];
    end 
    if(N9871) begin
      \nz.mem_3494_sv2v_reg  <= data_i[54];
    end 
    if(N9870) begin
      \nz.mem_3493_sv2v_reg  <= data_i[53];
    end 
    if(N9869) begin
      \nz.mem_3492_sv2v_reg  <= data_i[52];
    end 
    if(N9868) begin
      \nz.mem_3491_sv2v_reg  <= data_i[51];
    end 
    if(N9867) begin
      \nz.mem_3490_sv2v_reg  <= data_i[50];
    end 
    if(N9866) begin
      \nz.mem_3489_sv2v_reg  <= data_i[49];
    end 
    if(N9865) begin
      \nz.mem_3488_sv2v_reg  <= data_i[48];
    end 
    if(N9864) begin
      \nz.mem_3487_sv2v_reg  <= data_i[47];
    end 
    if(N9863) begin
      \nz.mem_3486_sv2v_reg  <= data_i[46];
    end 
    if(N9862) begin
      \nz.mem_3485_sv2v_reg  <= data_i[45];
    end 
    if(N9861) begin
      \nz.mem_3484_sv2v_reg  <= data_i[44];
    end 
    if(N9860) begin
      \nz.mem_3483_sv2v_reg  <= data_i[43];
    end 
    if(N9859) begin
      \nz.mem_3482_sv2v_reg  <= data_i[42];
    end 
    if(N9858) begin
      \nz.mem_3481_sv2v_reg  <= data_i[41];
    end 
    if(N9857) begin
      \nz.mem_3480_sv2v_reg  <= data_i[40];
    end 
    if(N9856) begin
      \nz.mem_3479_sv2v_reg  <= data_i[39];
    end 
    if(N9855) begin
      \nz.mem_3478_sv2v_reg  <= data_i[38];
    end 
    if(N9854) begin
      \nz.mem_3477_sv2v_reg  <= data_i[37];
    end 
    if(N9853) begin
      \nz.mem_3476_sv2v_reg  <= data_i[36];
    end 
    if(N9852) begin
      \nz.mem_3475_sv2v_reg  <= data_i[35];
    end 
    if(N9851) begin
      \nz.mem_3474_sv2v_reg  <= data_i[34];
    end 
    if(N9850) begin
      \nz.mem_3473_sv2v_reg  <= data_i[33];
    end 
    if(N9849) begin
      \nz.mem_3472_sv2v_reg  <= data_i[32];
    end 
    if(N9848) begin
      \nz.mem_3471_sv2v_reg  <= data_i[31];
    end 
    if(N9847) begin
      \nz.mem_3470_sv2v_reg  <= data_i[30];
    end 
    if(N9846) begin
      \nz.mem_3469_sv2v_reg  <= data_i[29];
    end 
    if(N9845) begin
      \nz.mem_3468_sv2v_reg  <= data_i[28];
    end 
    if(N9844) begin
      \nz.mem_3467_sv2v_reg  <= data_i[27];
    end 
    if(N9843) begin
      \nz.mem_3466_sv2v_reg  <= data_i[26];
    end 
    if(N9842) begin
      \nz.mem_3465_sv2v_reg  <= data_i[25];
    end 
    if(N9841) begin
      \nz.mem_3464_sv2v_reg  <= data_i[24];
    end 
    if(N9840) begin
      \nz.mem_3463_sv2v_reg  <= data_i[23];
    end 
    if(N9839) begin
      \nz.mem_3462_sv2v_reg  <= data_i[22];
    end 
    if(N9838) begin
      \nz.mem_3461_sv2v_reg  <= data_i[21];
    end 
    if(N9837) begin
      \nz.mem_3460_sv2v_reg  <= data_i[20];
    end 
    if(N9836) begin
      \nz.mem_3459_sv2v_reg  <= data_i[19];
    end 
    if(N9835) begin
      \nz.mem_3458_sv2v_reg  <= data_i[18];
    end 
    if(N9834) begin
      \nz.mem_3457_sv2v_reg  <= data_i[17];
    end 
    if(N9833) begin
      \nz.mem_3456_sv2v_reg  <= data_i[16];
    end 
    if(N9832) begin
      \nz.mem_3455_sv2v_reg  <= data_i[15];
    end 
    if(N9831) begin
      \nz.mem_3454_sv2v_reg  <= data_i[14];
    end 
    if(N9830) begin
      \nz.mem_3453_sv2v_reg  <= data_i[13];
    end 
    if(N9829) begin
      \nz.mem_3452_sv2v_reg  <= data_i[12];
    end 
    if(N9828) begin
      \nz.mem_3451_sv2v_reg  <= data_i[11];
    end 
    if(N9827) begin
      \nz.mem_3450_sv2v_reg  <= data_i[10];
    end 
    if(N9826) begin
      \nz.mem_3449_sv2v_reg  <= data_i[9];
    end 
    if(N9825) begin
      \nz.mem_3448_sv2v_reg  <= data_i[8];
    end 
    if(N9824) begin
      \nz.mem_3447_sv2v_reg  <= data_i[7];
    end 
    if(N9823) begin
      \nz.mem_3446_sv2v_reg  <= data_i[6];
    end 
    if(N9822) begin
      \nz.mem_3445_sv2v_reg  <= data_i[5];
    end 
    if(N9821) begin
      \nz.mem_3444_sv2v_reg  <= data_i[4];
    end 
    if(N9820) begin
      \nz.mem_3443_sv2v_reg  <= data_i[3];
    end 
    if(N9819) begin
      \nz.mem_3442_sv2v_reg  <= data_i[2];
    end 
    if(N9818) begin
      \nz.mem_3441_sv2v_reg  <= data_i[1];
    end 
    if(N9817) begin
      \nz.mem_3440_sv2v_reg  <= data_i[0];
    end 
    if(N9816) begin
      \nz.mem_3439_sv2v_reg  <= data_i[79];
    end 
    if(N9815) begin
      \nz.mem_3438_sv2v_reg  <= data_i[78];
    end 
    if(N9814) begin
      \nz.mem_3437_sv2v_reg  <= data_i[77];
    end 
    if(N9813) begin
      \nz.mem_3436_sv2v_reg  <= data_i[76];
    end 
    if(N9812) begin
      \nz.mem_3435_sv2v_reg  <= data_i[75];
    end 
    if(N9811) begin
      \nz.mem_3434_sv2v_reg  <= data_i[74];
    end 
    if(N9810) begin
      \nz.mem_3433_sv2v_reg  <= data_i[73];
    end 
    if(N9809) begin
      \nz.mem_3432_sv2v_reg  <= data_i[72];
    end 
    if(N9808) begin
      \nz.mem_3431_sv2v_reg  <= data_i[71];
    end 
    if(N9807) begin
      \nz.mem_3430_sv2v_reg  <= data_i[70];
    end 
    if(N9806) begin
      \nz.mem_3429_sv2v_reg  <= data_i[69];
    end 
    if(N9805) begin
      \nz.mem_3428_sv2v_reg  <= data_i[68];
    end 
    if(N9804) begin
      \nz.mem_3427_sv2v_reg  <= data_i[67];
    end 
    if(N9803) begin
      \nz.mem_3426_sv2v_reg  <= data_i[66];
    end 
    if(N9802) begin
      \nz.mem_3425_sv2v_reg  <= data_i[65];
    end 
    if(N9801) begin
      \nz.mem_3424_sv2v_reg  <= data_i[64];
    end 
    if(N9800) begin
      \nz.mem_3423_sv2v_reg  <= data_i[63];
    end 
    if(N9799) begin
      \nz.mem_3422_sv2v_reg  <= data_i[62];
    end 
    if(N9798) begin
      \nz.mem_3421_sv2v_reg  <= data_i[61];
    end 
    if(N9797) begin
      \nz.mem_3420_sv2v_reg  <= data_i[60];
    end 
    if(N9796) begin
      \nz.mem_3419_sv2v_reg  <= data_i[59];
    end 
    if(N9795) begin
      \nz.mem_3418_sv2v_reg  <= data_i[58];
    end 
    if(N9794) begin
      \nz.mem_3417_sv2v_reg  <= data_i[57];
    end 
    if(N9793) begin
      \nz.mem_3416_sv2v_reg  <= data_i[56];
    end 
    if(N9792) begin
      \nz.mem_3415_sv2v_reg  <= data_i[55];
    end 
    if(N9791) begin
      \nz.mem_3414_sv2v_reg  <= data_i[54];
    end 
    if(N9790) begin
      \nz.mem_3413_sv2v_reg  <= data_i[53];
    end 
    if(N9789) begin
      \nz.mem_3412_sv2v_reg  <= data_i[52];
    end 
    if(N9788) begin
      \nz.mem_3411_sv2v_reg  <= data_i[51];
    end 
    if(N9787) begin
      \nz.mem_3410_sv2v_reg  <= data_i[50];
    end 
    if(N9786) begin
      \nz.mem_3409_sv2v_reg  <= data_i[49];
    end 
    if(N9785) begin
      \nz.mem_3408_sv2v_reg  <= data_i[48];
    end 
    if(N9784) begin
      \nz.mem_3407_sv2v_reg  <= data_i[47];
    end 
    if(N9783) begin
      \nz.mem_3406_sv2v_reg  <= data_i[46];
    end 
    if(N9782) begin
      \nz.mem_3405_sv2v_reg  <= data_i[45];
    end 
    if(N9781) begin
      \nz.mem_3404_sv2v_reg  <= data_i[44];
    end 
    if(N9780) begin
      \nz.mem_3403_sv2v_reg  <= data_i[43];
    end 
    if(N9779) begin
      \nz.mem_3402_sv2v_reg  <= data_i[42];
    end 
    if(N9778) begin
      \nz.mem_3401_sv2v_reg  <= data_i[41];
    end 
    if(N9777) begin
      \nz.mem_3400_sv2v_reg  <= data_i[40];
    end 
    if(N9776) begin
      \nz.mem_3399_sv2v_reg  <= data_i[39];
    end 
    if(N9775) begin
      \nz.mem_3398_sv2v_reg  <= data_i[38];
    end 
    if(N9774) begin
      \nz.mem_3397_sv2v_reg  <= data_i[37];
    end 
    if(N9773) begin
      \nz.mem_3396_sv2v_reg  <= data_i[36];
    end 
    if(N9772) begin
      \nz.mem_3395_sv2v_reg  <= data_i[35];
    end 
    if(N9771) begin
      \nz.mem_3394_sv2v_reg  <= data_i[34];
    end 
    if(N9770) begin
      \nz.mem_3393_sv2v_reg  <= data_i[33];
    end 
    if(N9769) begin
      \nz.mem_3392_sv2v_reg  <= data_i[32];
    end 
    if(N9768) begin
      \nz.mem_3391_sv2v_reg  <= data_i[31];
    end 
    if(N9767) begin
      \nz.mem_3390_sv2v_reg  <= data_i[30];
    end 
    if(N9766) begin
      \nz.mem_3389_sv2v_reg  <= data_i[29];
    end 
    if(N9765) begin
      \nz.mem_3388_sv2v_reg  <= data_i[28];
    end 
    if(N9764) begin
      \nz.mem_3387_sv2v_reg  <= data_i[27];
    end 
    if(N9763) begin
      \nz.mem_3386_sv2v_reg  <= data_i[26];
    end 
    if(N9762) begin
      \nz.mem_3385_sv2v_reg  <= data_i[25];
    end 
    if(N9761) begin
      \nz.mem_3384_sv2v_reg  <= data_i[24];
    end 
    if(N9760) begin
      \nz.mem_3383_sv2v_reg  <= data_i[23];
    end 
    if(N9759) begin
      \nz.mem_3382_sv2v_reg  <= data_i[22];
    end 
    if(N9758) begin
      \nz.mem_3381_sv2v_reg  <= data_i[21];
    end 
    if(N9757) begin
      \nz.mem_3380_sv2v_reg  <= data_i[20];
    end 
    if(N9756) begin
      \nz.mem_3379_sv2v_reg  <= data_i[19];
    end 
    if(N9755) begin
      \nz.mem_3378_sv2v_reg  <= data_i[18];
    end 
    if(N9754) begin
      \nz.mem_3377_sv2v_reg  <= data_i[17];
    end 
    if(N9753) begin
      \nz.mem_3376_sv2v_reg  <= data_i[16];
    end 
    if(N9752) begin
      \nz.mem_3375_sv2v_reg  <= data_i[15];
    end 
    if(N9751) begin
      \nz.mem_3374_sv2v_reg  <= data_i[14];
    end 
    if(N9750) begin
      \nz.mem_3373_sv2v_reg  <= data_i[13];
    end 
    if(N9749) begin
      \nz.mem_3372_sv2v_reg  <= data_i[12];
    end 
    if(N9748) begin
      \nz.mem_3371_sv2v_reg  <= data_i[11];
    end 
    if(N9747) begin
      \nz.mem_3370_sv2v_reg  <= data_i[10];
    end 
    if(N9746) begin
      \nz.mem_3369_sv2v_reg  <= data_i[9];
    end 
    if(N9745) begin
      \nz.mem_3368_sv2v_reg  <= data_i[8];
    end 
    if(N9744) begin
      \nz.mem_3367_sv2v_reg  <= data_i[7];
    end 
    if(N9743) begin
      \nz.mem_3366_sv2v_reg  <= data_i[6];
    end 
    if(N9742) begin
      \nz.mem_3365_sv2v_reg  <= data_i[5];
    end 
    if(N9741) begin
      \nz.mem_3364_sv2v_reg  <= data_i[4];
    end 
    if(N9740) begin
      \nz.mem_3363_sv2v_reg  <= data_i[3];
    end 
    if(N9739) begin
      \nz.mem_3362_sv2v_reg  <= data_i[2];
    end 
    if(N9738) begin
      \nz.mem_3361_sv2v_reg  <= data_i[1];
    end 
    if(N9737) begin
      \nz.mem_3360_sv2v_reg  <= data_i[0];
    end 
    if(N9736) begin
      \nz.mem_3359_sv2v_reg  <= data_i[79];
    end 
    if(N9735) begin
      \nz.mem_3358_sv2v_reg  <= data_i[78];
    end 
    if(N9734) begin
      \nz.mem_3357_sv2v_reg  <= data_i[77];
    end 
    if(N9733) begin
      \nz.mem_3356_sv2v_reg  <= data_i[76];
    end 
    if(N9732) begin
      \nz.mem_3355_sv2v_reg  <= data_i[75];
    end 
    if(N9731) begin
      \nz.mem_3354_sv2v_reg  <= data_i[74];
    end 
    if(N9730) begin
      \nz.mem_3353_sv2v_reg  <= data_i[73];
    end 
    if(N9729) begin
      \nz.mem_3352_sv2v_reg  <= data_i[72];
    end 
    if(N9728) begin
      \nz.mem_3351_sv2v_reg  <= data_i[71];
    end 
    if(N9727) begin
      \nz.mem_3350_sv2v_reg  <= data_i[70];
    end 
    if(N9726) begin
      \nz.mem_3349_sv2v_reg  <= data_i[69];
    end 
    if(N9725) begin
      \nz.mem_3348_sv2v_reg  <= data_i[68];
    end 
    if(N9724) begin
      \nz.mem_3347_sv2v_reg  <= data_i[67];
    end 
    if(N9723) begin
      \nz.mem_3346_sv2v_reg  <= data_i[66];
    end 
    if(N9722) begin
      \nz.mem_3345_sv2v_reg  <= data_i[65];
    end 
    if(N9721) begin
      \nz.mem_3344_sv2v_reg  <= data_i[64];
    end 
    if(N9720) begin
      \nz.mem_3343_sv2v_reg  <= data_i[63];
    end 
    if(N9719) begin
      \nz.mem_3342_sv2v_reg  <= data_i[62];
    end 
    if(N9718) begin
      \nz.mem_3341_sv2v_reg  <= data_i[61];
    end 
    if(N9717) begin
      \nz.mem_3340_sv2v_reg  <= data_i[60];
    end 
    if(N9716) begin
      \nz.mem_3339_sv2v_reg  <= data_i[59];
    end 
    if(N9715) begin
      \nz.mem_3338_sv2v_reg  <= data_i[58];
    end 
    if(N9714) begin
      \nz.mem_3337_sv2v_reg  <= data_i[57];
    end 
    if(N9713) begin
      \nz.mem_3336_sv2v_reg  <= data_i[56];
    end 
    if(N9712) begin
      \nz.mem_3335_sv2v_reg  <= data_i[55];
    end 
    if(N9711) begin
      \nz.mem_3334_sv2v_reg  <= data_i[54];
    end 
    if(N9710) begin
      \nz.mem_3333_sv2v_reg  <= data_i[53];
    end 
    if(N9709) begin
      \nz.mem_3332_sv2v_reg  <= data_i[52];
    end 
    if(N9708) begin
      \nz.mem_3331_sv2v_reg  <= data_i[51];
    end 
    if(N9707) begin
      \nz.mem_3330_sv2v_reg  <= data_i[50];
    end 
    if(N9706) begin
      \nz.mem_3329_sv2v_reg  <= data_i[49];
    end 
    if(N9705) begin
      \nz.mem_3328_sv2v_reg  <= data_i[48];
    end 
    if(N9704) begin
      \nz.mem_3327_sv2v_reg  <= data_i[47];
    end 
    if(N9703) begin
      \nz.mem_3326_sv2v_reg  <= data_i[46];
    end 
    if(N9702) begin
      \nz.mem_3325_sv2v_reg  <= data_i[45];
    end 
    if(N9701) begin
      \nz.mem_3324_sv2v_reg  <= data_i[44];
    end 
    if(N9700) begin
      \nz.mem_3323_sv2v_reg  <= data_i[43];
    end 
    if(N9699) begin
      \nz.mem_3322_sv2v_reg  <= data_i[42];
    end 
    if(N9698) begin
      \nz.mem_3321_sv2v_reg  <= data_i[41];
    end 
    if(N9697) begin
      \nz.mem_3320_sv2v_reg  <= data_i[40];
    end 
    if(N9696) begin
      \nz.mem_3319_sv2v_reg  <= data_i[39];
    end 
    if(N9695) begin
      \nz.mem_3318_sv2v_reg  <= data_i[38];
    end 
    if(N9694) begin
      \nz.mem_3317_sv2v_reg  <= data_i[37];
    end 
    if(N9693) begin
      \nz.mem_3316_sv2v_reg  <= data_i[36];
    end 
    if(N9692) begin
      \nz.mem_3315_sv2v_reg  <= data_i[35];
    end 
    if(N9691) begin
      \nz.mem_3314_sv2v_reg  <= data_i[34];
    end 
    if(N9690) begin
      \nz.mem_3313_sv2v_reg  <= data_i[33];
    end 
    if(N9689) begin
      \nz.mem_3312_sv2v_reg  <= data_i[32];
    end 
    if(N9688) begin
      \nz.mem_3311_sv2v_reg  <= data_i[31];
    end 
    if(N9687) begin
      \nz.mem_3310_sv2v_reg  <= data_i[30];
    end 
    if(N9686) begin
      \nz.mem_3309_sv2v_reg  <= data_i[29];
    end 
    if(N9685) begin
      \nz.mem_3308_sv2v_reg  <= data_i[28];
    end 
    if(N9684) begin
      \nz.mem_3307_sv2v_reg  <= data_i[27];
    end 
    if(N9683) begin
      \nz.mem_3306_sv2v_reg  <= data_i[26];
    end 
    if(N9682) begin
      \nz.mem_3305_sv2v_reg  <= data_i[25];
    end 
    if(N9681) begin
      \nz.mem_3304_sv2v_reg  <= data_i[24];
    end 
    if(N9680) begin
      \nz.mem_3303_sv2v_reg  <= data_i[23];
    end 
    if(N9679) begin
      \nz.mem_3302_sv2v_reg  <= data_i[22];
    end 
    if(N9678) begin
      \nz.mem_3301_sv2v_reg  <= data_i[21];
    end 
    if(N9677) begin
      \nz.mem_3300_sv2v_reg  <= data_i[20];
    end 
    if(N9676) begin
      \nz.mem_3299_sv2v_reg  <= data_i[19];
    end 
    if(N9675) begin
      \nz.mem_3298_sv2v_reg  <= data_i[18];
    end 
    if(N9674) begin
      \nz.mem_3297_sv2v_reg  <= data_i[17];
    end 
    if(N9673) begin
      \nz.mem_3296_sv2v_reg  <= data_i[16];
    end 
    if(N9672) begin
      \nz.mem_3295_sv2v_reg  <= data_i[15];
    end 
    if(N9671) begin
      \nz.mem_3294_sv2v_reg  <= data_i[14];
    end 
    if(N9670) begin
      \nz.mem_3293_sv2v_reg  <= data_i[13];
    end 
    if(N9669) begin
      \nz.mem_3292_sv2v_reg  <= data_i[12];
    end 
    if(N9668) begin
      \nz.mem_3291_sv2v_reg  <= data_i[11];
    end 
    if(N9667) begin
      \nz.mem_3290_sv2v_reg  <= data_i[10];
    end 
    if(N9666) begin
      \nz.mem_3289_sv2v_reg  <= data_i[9];
    end 
    if(N9665) begin
      \nz.mem_3288_sv2v_reg  <= data_i[8];
    end 
    if(N9664) begin
      \nz.mem_3287_sv2v_reg  <= data_i[7];
    end 
    if(N9663) begin
      \nz.mem_3286_sv2v_reg  <= data_i[6];
    end 
    if(N9662) begin
      \nz.mem_3285_sv2v_reg  <= data_i[5];
    end 
    if(N9661) begin
      \nz.mem_3284_sv2v_reg  <= data_i[4];
    end 
    if(N9660) begin
      \nz.mem_3283_sv2v_reg  <= data_i[3];
    end 
    if(N9659) begin
      \nz.mem_3282_sv2v_reg  <= data_i[2];
    end 
    if(N9658) begin
      \nz.mem_3281_sv2v_reg  <= data_i[1];
    end 
    if(N9657) begin
      \nz.mem_3280_sv2v_reg  <= data_i[0];
    end 
    if(N9656) begin
      \nz.mem_3279_sv2v_reg  <= data_i[79];
    end 
    if(N9655) begin
      \nz.mem_3278_sv2v_reg  <= data_i[78];
    end 
    if(N9654) begin
      \nz.mem_3277_sv2v_reg  <= data_i[77];
    end 
    if(N9653) begin
      \nz.mem_3276_sv2v_reg  <= data_i[76];
    end 
    if(N9652) begin
      \nz.mem_3275_sv2v_reg  <= data_i[75];
    end 
    if(N9651) begin
      \nz.mem_3274_sv2v_reg  <= data_i[74];
    end 
    if(N9650) begin
      \nz.mem_3273_sv2v_reg  <= data_i[73];
    end 
    if(N9649) begin
      \nz.mem_3272_sv2v_reg  <= data_i[72];
    end 
    if(N9648) begin
      \nz.mem_3271_sv2v_reg  <= data_i[71];
    end 
    if(N9647) begin
      \nz.mem_3270_sv2v_reg  <= data_i[70];
    end 
    if(N9646) begin
      \nz.mem_3269_sv2v_reg  <= data_i[69];
    end 
    if(N9645) begin
      \nz.mem_3268_sv2v_reg  <= data_i[68];
    end 
    if(N9644) begin
      \nz.mem_3267_sv2v_reg  <= data_i[67];
    end 
    if(N9643) begin
      \nz.mem_3266_sv2v_reg  <= data_i[66];
    end 
    if(N9642) begin
      \nz.mem_3265_sv2v_reg  <= data_i[65];
    end 
    if(N9641) begin
      \nz.mem_3264_sv2v_reg  <= data_i[64];
    end 
    if(N9640) begin
      \nz.mem_3263_sv2v_reg  <= data_i[63];
    end 
    if(N9639) begin
      \nz.mem_3262_sv2v_reg  <= data_i[62];
    end 
    if(N9638) begin
      \nz.mem_3261_sv2v_reg  <= data_i[61];
    end 
    if(N9637) begin
      \nz.mem_3260_sv2v_reg  <= data_i[60];
    end 
    if(N9636) begin
      \nz.mem_3259_sv2v_reg  <= data_i[59];
    end 
    if(N9635) begin
      \nz.mem_3258_sv2v_reg  <= data_i[58];
    end 
    if(N9634) begin
      \nz.mem_3257_sv2v_reg  <= data_i[57];
    end 
    if(N9633) begin
      \nz.mem_3256_sv2v_reg  <= data_i[56];
    end 
    if(N9632) begin
      \nz.mem_3255_sv2v_reg  <= data_i[55];
    end 
    if(N9631) begin
      \nz.mem_3254_sv2v_reg  <= data_i[54];
    end 
    if(N9630) begin
      \nz.mem_3253_sv2v_reg  <= data_i[53];
    end 
    if(N9629) begin
      \nz.mem_3252_sv2v_reg  <= data_i[52];
    end 
    if(N9628) begin
      \nz.mem_3251_sv2v_reg  <= data_i[51];
    end 
    if(N9627) begin
      \nz.mem_3250_sv2v_reg  <= data_i[50];
    end 
    if(N9626) begin
      \nz.mem_3249_sv2v_reg  <= data_i[49];
    end 
    if(N9625) begin
      \nz.mem_3248_sv2v_reg  <= data_i[48];
    end 
    if(N9624) begin
      \nz.mem_3247_sv2v_reg  <= data_i[47];
    end 
    if(N9623) begin
      \nz.mem_3246_sv2v_reg  <= data_i[46];
    end 
    if(N9622) begin
      \nz.mem_3245_sv2v_reg  <= data_i[45];
    end 
    if(N9621) begin
      \nz.mem_3244_sv2v_reg  <= data_i[44];
    end 
    if(N9620) begin
      \nz.mem_3243_sv2v_reg  <= data_i[43];
    end 
    if(N9619) begin
      \nz.mem_3242_sv2v_reg  <= data_i[42];
    end 
    if(N9618) begin
      \nz.mem_3241_sv2v_reg  <= data_i[41];
    end 
    if(N9617) begin
      \nz.mem_3240_sv2v_reg  <= data_i[40];
    end 
    if(N9616) begin
      \nz.mem_3239_sv2v_reg  <= data_i[39];
    end 
    if(N9615) begin
      \nz.mem_3238_sv2v_reg  <= data_i[38];
    end 
    if(N9614) begin
      \nz.mem_3237_sv2v_reg  <= data_i[37];
    end 
    if(N9613) begin
      \nz.mem_3236_sv2v_reg  <= data_i[36];
    end 
    if(N9612) begin
      \nz.mem_3235_sv2v_reg  <= data_i[35];
    end 
    if(N9611) begin
      \nz.mem_3234_sv2v_reg  <= data_i[34];
    end 
    if(N9610) begin
      \nz.mem_3233_sv2v_reg  <= data_i[33];
    end 
    if(N9609) begin
      \nz.mem_3232_sv2v_reg  <= data_i[32];
    end 
    if(N9608) begin
      \nz.mem_3231_sv2v_reg  <= data_i[31];
    end 
    if(N9607) begin
      \nz.mem_3230_sv2v_reg  <= data_i[30];
    end 
    if(N9606) begin
      \nz.mem_3229_sv2v_reg  <= data_i[29];
    end 
    if(N9605) begin
      \nz.mem_3228_sv2v_reg  <= data_i[28];
    end 
    if(N9604) begin
      \nz.mem_3227_sv2v_reg  <= data_i[27];
    end 
    if(N9603) begin
      \nz.mem_3226_sv2v_reg  <= data_i[26];
    end 
    if(N9602) begin
      \nz.mem_3225_sv2v_reg  <= data_i[25];
    end 
    if(N9601) begin
      \nz.mem_3224_sv2v_reg  <= data_i[24];
    end 
    if(N9600) begin
      \nz.mem_3223_sv2v_reg  <= data_i[23];
    end 
    if(N9599) begin
      \nz.mem_3222_sv2v_reg  <= data_i[22];
    end 
    if(N9598) begin
      \nz.mem_3221_sv2v_reg  <= data_i[21];
    end 
    if(N9597) begin
      \nz.mem_3220_sv2v_reg  <= data_i[20];
    end 
    if(N9596) begin
      \nz.mem_3219_sv2v_reg  <= data_i[19];
    end 
    if(N9595) begin
      \nz.mem_3218_sv2v_reg  <= data_i[18];
    end 
    if(N9594) begin
      \nz.mem_3217_sv2v_reg  <= data_i[17];
    end 
    if(N9593) begin
      \nz.mem_3216_sv2v_reg  <= data_i[16];
    end 
    if(N9592) begin
      \nz.mem_3215_sv2v_reg  <= data_i[15];
    end 
    if(N9591) begin
      \nz.mem_3214_sv2v_reg  <= data_i[14];
    end 
    if(N9590) begin
      \nz.mem_3213_sv2v_reg  <= data_i[13];
    end 
    if(N9589) begin
      \nz.mem_3212_sv2v_reg  <= data_i[12];
    end 
    if(N9588) begin
      \nz.mem_3211_sv2v_reg  <= data_i[11];
    end 
    if(N9587) begin
      \nz.mem_3210_sv2v_reg  <= data_i[10];
    end 
    if(N9586) begin
      \nz.mem_3209_sv2v_reg  <= data_i[9];
    end 
    if(N9585) begin
      \nz.mem_3208_sv2v_reg  <= data_i[8];
    end 
    if(N9584) begin
      \nz.mem_3207_sv2v_reg  <= data_i[7];
    end 
    if(N9583) begin
      \nz.mem_3206_sv2v_reg  <= data_i[6];
    end 
    if(N9582) begin
      \nz.mem_3205_sv2v_reg  <= data_i[5];
    end 
    if(N9581) begin
      \nz.mem_3204_sv2v_reg  <= data_i[4];
    end 
    if(N9580) begin
      \nz.mem_3203_sv2v_reg  <= data_i[3];
    end 
    if(N9579) begin
      \nz.mem_3202_sv2v_reg  <= data_i[2];
    end 
    if(N9578) begin
      \nz.mem_3201_sv2v_reg  <= data_i[1];
    end 
    if(N9577) begin
      \nz.mem_3200_sv2v_reg  <= data_i[0];
    end 
    if(N9576) begin
      \nz.mem_3199_sv2v_reg  <= data_i[79];
    end 
    if(N9575) begin
      \nz.mem_3198_sv2v_reg  <= data_i[78];
    end 
    if(N9574) begin
      \nz.mem_3197_sv2v_reg  <= data_i[77];
    end 
    if(N9573) begin
      \nz.mem_3196_sv2v_reg  <= data_i[76];
    end 
    if(N9572) begin
      \nz.mem_3195_sv2v_reg  <= data_i[75];
    end 
    if(N9571) begin
      \nz.mem_3194_sv2v_reg  <= data_i[74];
    end 
    if(N9570) begin
      \nz.mem_3193_sv2v_reg  <= data_i[73];
    end 
    if(N9569) begin
      \nz.mem_3192_sv2v_reg  <= data_i[72];
    end 
    if(N9568) begin
      \nz.mem_3191_sv2v_reg  <= data_i[71];
    end 
    if(N9567) begin
      \nz.mem_3190_sv2v_reg  <= data_i[70];
    end 
    if(N9566) begin
      \nz.mem_3189_sv2v_reg  <= data_i[69];
    end 
    if(N9565) begin
      \nz.mem_3188_sv2v_reg  <= data_i[68];
    end 
    if(N9564) begin
      \nz.mem_3187_sv2v_reg  <= data_i[67];
    end 
    if(N9563) begin
      \nz.mem_3186_sv2v_reg  <= data_i[66];
    end 
    if(N9562) begin
      \nz.mem_3185_sv2v_reg  <= data_i[65];
    end 
    if(N9561) begin
      \nz.mem_3184_sv2v_reg  <= data_i[64];
    end 
    if(N9560) begin
      \nz.mem_3183_sv2v_reg  <= data_i[63];
    end 
    if(N9559) begin
      \nz.mem_3182_sv2v_reg  <= data_i[62];
    end 
    if(N9558) begin
      \nz.mem_3181_sv2v_reg  <= data_i[61];
    end 
    if(N9557) begin
      \nz.mem_3180_sv2v_reg  <= data_i[60];
    end 
    if(N9556) begin
      \nz.mem_3179_sv2v_reg  <= data_i[59];
    end 
    if(N9555) begin
      \nz.mem_3178_sv2v_reg  <= data_i[58];
    end 
    if(N9554) begin
      \nz.mem_3177_sv2v_reg  <= data_i[57];
    end 
    if(N9553) begin
      \nz.mem_3176_sv2v_reg  <= data_i[56];
    end 
    if(N9552) begin
      \nz.mem_3175_sv2v_reg  <= data_i[55];
    end 
    if(N9551) begin
      \nz.mem_3174_sv2v_reg  <= data_i[54];
    end 
    if(N9550) begin
      \nz.mem_3173_sv2v_reg  <= data_i[53];
    end 
    if(N9549) begin
      \nz.mem_3172_sv2v_reg  <= data_i[52];
    end 
    if(N9548) begin
      \nz.mem_3171_sv2v_reg  <= data_i[51];
    end 
    if(N9547) begin
      \nz.mem_3170_sv2v_reg  <= data_i[50];
    end 
    if(N9546) begin
      \nz.mem_3169_sv2v_reg  <= data_i[49];
    end 
    if(N9545) begin
      \nz.mem_3168_sv2v_reg  <= data_i[48];
    end 
    if(N9544) begin
      \nz.mem_3167_sv2v_reg  <= data_i[47];
    end 
    if(N9543) begin
      \nz.mem_3166_sv2v_reg  <= data_i[46];
    end 
    if(N9542) begin
      \nz.mem_3165_sv2v_reg  <= data_i[45];
    end 
    if(N9541) begin
      \nz.mem_3164_sv2v_reg  <= data_i[44];
    end 
    if(N9540) begin
      \nz.mem_3163_sv2v_reg  <= data_i[43];
    end 
    if(N9539) begin
      \nz.mem_3162_sv2v_reg  <= data_i[42];
    end 
    if(N9538) begin
      \nz.mem_3161_sv2v_reg  <= data_i[41];
    end 
    if(N9537) begin
      \nz.mem_3160_sv2v_reg  <= data_i[40];
    end 
    if(N9536) begin
      \nz.mem_3159_sv2v_reg  <= data_i[39];
    end 
    if(N9535) begin
      \nz.mem_3158_sv2v_reg  <= data_i[38];
    end 
    if(N9534) begin
      \nz.mem_3157_sv2v_reg  <= data_i[37];
    end 
    if(N9533) begin
      \nz.mem_3156_sv2v_reg  <= data_i[36];
    end 
    if(N9532) begin
      \nz.mem_3155_sv2v_reg  <= data_i[35];
    end 
    if(N9531) begin
      \nz.mem_3154_sv2v_reg  <= data_i[34];
    end 
    if(N9530) begin
      \nz.mem_3153_sv2v_reg  <= data_i[33];
    end 
    if(N9529) begin
      \nz.mem_3152_sv2v_reg  <= data_i[32];
    end 
    if(N9528) begin
      \nz.mem_3151_sv2v_reg  <= data_i[31];
    end 
    if(N9527) begin
      \nz.mem_3150_sv2v_reg  <= data_i[30];
    end 
    if(N9526) begin
      \nz.mem_3149_sv2v_reg  <= data_i[29];
    end 
    if(N9525) begin
      \nz.mem_3148_sv2v_reg  <= data_i[28];
    end 
    if(N9524) begin
      \nz.mem_3147_sv2v_reg  <= data_i[27];
    end 
    if(N9523) begin
      \nz.mem_3146_sv2v_reg  <= data_i[26];
    end 
    if(N9522) begin
      \nz.mem_3145_sv2v_reg  <= data_i[25];
    end 
    if(N9521) begin
      \nz.mem_3144_sv2v_reg  <= data_i[24];
    end 
    if(N9520) begin
      \nz.mem_3143_sv2v_reg  <= data_i[23];
    end 
    if(N9519) begin
      \nz.mem_3142_sv2v_reg  <= data_i[22];
    end 
    if(N9518) begin
      \nz.mem_3141_sv2v_reg  <= data_i[21];
    end 
    if(N9517) begin
      \nz.mem_3140_sv2v_reg  <= data_i[20];
    end 
    if(N9516) begin
      \nz.mem_3139_sv2v_reg  <= data_i[19];
    end 
    if(N9515) begin
      \nz.mem_3138_sv2v_reg  <= data_i[18];
    end 
    if(N9514) begin
      \nz.mem_3137_sv2v_reg  <= data_i[17];
    end 
    if(N9513) begin
      \nz.mem_3136_sv2v_reg  <= data_i[16];
    end 
    if(N9512) begin
      \nz.mem_3135_sv2v_reg  <= data_i[15];
    end 
    if(N9511) begin
      \nz.mem_3134_sv2v_reg  <= data_i[14];
    end 
    if(N9510) begin
      \nz.mem_3133_sv2v_reg  <= data_i[13];
    end 
    if(N9509) begin
      \nz.mem_3132_sv2v_reg  <= data_i[12];
    end 
    if(N9508) begin
      \nz.mem_3131_sv2v_reg  <= data_i[11];
    end 
    if(N9507) begin
      \nz.mem_3130_sv2v_reg  <= data_i[10];
    end 
    if(N9506) begin
      \nz.mem_3129_sv2v_reg  <= data_i[9];
    end 
    if(N9505) begin
      \nz.mem_3128_sv2v_reg  <= data_i[8];
    end 
    if(N9504) begin
      \nz.mem_3127_sv2v_reg  <= data_i[7];
    end 
    if(N9503) begin
      \nz.mem_3126_sv2v_reg  <= data_i[6];
    end 
    if(N9502) begin
      \nz.mem_3125_sv2v_reg  <= data_i[5];
    end 
    if(N9501) begin
      \nz.mem_3124_sv2v_reg  <= data_i[4];
    end 
    if(N9500) begin
      \nz.mem_3123_sv2v_reg  <= data_i[3];
    end 
    if(N9499) begin
      \nz.mem_3122_sv2v_reg  <= data_i[2];
    end 
    if(N9498) begin
      \nz.mem_3121_sv2v_reg  <= data_i[1];
    end 
    if(N9497) begin
      \nz.mem_3120_sv2v_reg  <= data_i[0];
    end 
    if(N9496) begin
      \nz.mem_3119_sv2v_reg  <= data_i[79];
    end 
    if(N9495) begin
      \nz.mem_3118_sv2v_reg  <= data_i[78];
    end 
    if(N9494) begin
      \nz.mem_3117_sv2v_reg  <= data_i[77];
    end 
    if(N9493) begin
      \nz.mem_3116_sv2v_reg  <= data_i[76];
    end 
    if(N9492) begin
      \nz.mem_3115_sv2v_reg  <= data_i[75];
    end 
    if(N9491) begin
      \nz.mem_3114_sv2v_reg  <= data_i[74];
    end 
    if(N9490) begin
      \nz.mem_3113_sv2v_reg  <= data_i[73];
    end 
    if(N9489) begin
      \nz.mem_3112_sv2v_reg  <= data_i[72];
    end 
    if(N9488) begin
      \nz.mem_3111_sv2v_reg  <= data_i[71];
    end 
    if(N9487) begin
      \nz.mem_3110_sv2v_reg  <= data_i[70];
    end 
    if(N9486) begin
      \nz.mem_3109_sv2v_reg  <= data_i[69];
    end 
    if(N9485) begin
      \nz.mem_3108_sv2v_reg  <= data_i[68];
    end 
    if(N9484) begin
      \nz.mem_3107_sv2v_reg  <= data_i[67];
    end 
    if(N9483) begin
      \nz.mem_3106_sv2v_reg  <= data_i[66];
    end 
    if(N9482) begin
      \nz.mem_3105_sv2v_reg  <= data_i[65];
    end 
    if(N9481) begin
      \nz.mem_3104_sv2v_reg  <= data_i[64];
    end 
    if(N9480) begin
      \nz.mem_3103_sv2v_reg  <= data_i[63];
    end 
    if(N9479) begin
      \nz.mem_3102_sv2v_reg  <= data_i[62];
    end 
    if(N9478) begin
      \nz.mem_3101_sv2v_reg  <= data_i[61];
    end 
    if(N9477) begin
      \nz.mem_3100_sv2v_reg  <= data_i[60];
    end 
    if(N9476) begin
      \nz.mem_3099_sv2v_reg  <= data_i[59];
    end 
    if(N9475) begin
      \nz.mem_3098_sv2v_reg  <= data_i[58];
    end 
    if(N9474) begin
      \nz.mem_3097_sv2v_reg  <= data_i[57];
    end 
    if(N9473) begin
      \nz.mem_3096_sv2v_reg  <= data_i[56];
    end 
    if(N9472) begin
      \nz.mem_3095_sv2v_reg  <= data_i[55];
    end 
    if(N9471) begin
      \nz.mem_3094_sv2v_reg  <= data_i[54];
    end 
    if(N9470) begin
      \nz.mem_3093_sv2v_reg  <= data_i[53];
    end 
    if(N9469) begin
      \nz.mem_3092_sv2v_reg  <= data_i[52];
    end 
    if(N9468) begin
      \nz.mem_3091_sv2v_reg  <= data_i[51];
    end 
    if(N9467) begin
      \nz.mem_3090_sv2v_reg  <= data_i[50];
    end 
    if(N9466) begin
      \nz.mem_3089_sv2v_reg  <= data_i[49];
    end 
    if(N9465) begin
      \nz.mem_3088_sv2v_reg  <= data_i[48];
    end 
    if(N9464) begin
      \nz.mem_3087_sv2v_reg  <= data_i[47];
    end 
    if(N9463) begin
      \nz.mem_3086_sv2v_reg  <= data_i[46];
    end 
    if(N9462) begin
      \nz.mem_3085_sv2v_reg  <= data_i[45];
    end 
    if(N9461) begin
      \nz.mem_3084_sv2v_reg  <= data_i[44];
    end 
    if(N9460) begin
      \nz.mem_3083_sv2v_reg  <= data_i[43];
    end 
    if(N9459) begin
      \nz.mem_3082_sv2v_reg  <= data_i[42];
    end 
    if(N9458) begin
      \nz.mem_3081_sv2v_reg  <= data_i[41];
    end 
    if(N9457) begin
      \nz.mem_3080_sv2v_reg  <= data_i[40];
    end 
    if(N9456) begin
      \nz.mem_3079_sv2v_reg  <= data_i[39];
    end 
    if(N9455) begin
      \nz.mem_3078_sv2v_reg  <= data_i[38];
    end 
    if(N9454) begin
      \nz.mem_3077_sv2v_reg  <= data_i[37];
    end 
    if(N9453) begin
      \nz.mem_3076_sv2v_reg  <= data_i[36];
    end 
    if(N9452) begin
      \nz.mem_3075_sv2v_reg  <= data_i[35];
    end 
    if(N9451) begin
      \nz.mem_3074_sv2v_reg  <= data_i[34];
    end 
    if(N9450) begin
      \nz.mem_3073_sv2v_reg  <= data_i[33];
    end 
    if(N9449) begin
      \nz.mem_3072_sv2v_reg  <= data_i[32];
    end 
    if(N9448) begin
      \nz.mem_3071_sv2v_reg  <= data_i[31];
    end 
    if(N9447) begin
      \nz.mem_3070_sv2v_reg  <= data_i[30];
    end 
    if(N9446) begin
      \nz.mem_3069_sv2v_reg  <= data_i[29];
    end 
    if(N9445) begin
      \nz.mem_3068_sv2v_reg  <= data_i[28];
    end 
    if(N9444) begin
      \nz.mem_3067_sv2v_reg  <= data_i[27];
    end 
    if(N9443) begin
      \nz.mem_3066_sv2v_reg  <= data_i[26];
    end 
    if(N9442) begin
      \nz.mem_3065_sv2v_reg  <= data_i[25];
    end 
    if(N9441) begin
      \nz.mem_3064_sv2v_reg  <= data_i[24];
    end 
    if(N9440) begin
      \nz.mem_3063_sv2v_reg  <= data_i[23];
    end 
    if(N9439) begin
      \nz.mem_3062_sv2v_reg  <= data_i[22];
    end 
    if(N9438) begin
      \nz.mem_3061_sv2v_reg  <= data_i[21];
    end 
    if(N9437) begin
      \nz.mem_3060_sv2v_reg  <= data_i[20];
    end 
    if(N9436) begin
      \nz.mem_3059_sv2v_reg  <= data_i[19];
    end 
    if(N9435) begin
      \nz.mem_3058_sv2v_reg  <= data_i[18];
    end 
    if(N9434) begin
      \nz.mem_3057_sv2v_reg  <= data_i[17];
    end 
    if(N9433) begin
      \nz.mem_3056_sv2v_reg  <= data_i[16];
    end 
    if(N9432) begin
      \nz.mem_3055_sv2v_reg  <= data_i[15];
    end 
    if(N9431) begin
      \nz.mem_3054_sv2v_reg  <= data_i[14];
    end 
    if(N9430) begin
      \nz.mem_3053_sv2v_reg  <= data_i[13];
    end 
    if(N9429) begin
      \nz.mem_3052_sv2v_reg  <= data_i[12];
    end 
    if(N9428) begin
      \nz.mem_3051_sv2v_reg  <= data_i[11];
    end 
    if(N9427) begin
      \nz.mem_3050_sv2v_reg  <= data_i[10];
    end 
    if(N9426) begin
      \nz.mem_3049_sv2v_reg  <= data_i[9];
    end 
    if(N9425) begin
      \nz.mem_3048_sv2v_reg  <= data_i[8];
    end 
    if(N9424) begin
      \nz.mem_3047_sv2v_reg  <= data_i[7];
    end 
    if(N9423) begin
      \nz.mem_3046_sv2v_reg  <= data_i[6];
    end 
    if(N9422) begin
      \nz.mem_3045_sv2v_reg  <= data_i[5];
    end 
    if(N9421) begin
      \nz.mem_3044_sv2v_reg  <= data_i[4];
    end 
    if(N9420) begin
      \nz.mem_3043_sv2v_reg  <= data_i[3];
    end 
    if(N9419) begin
      \nz.mem_3042_sv2v_reg  <= data_i[2];
    end 
    if(N9418) begin
      \nz.mem_3041_sv2v_reg  <= data_i[1];
    end 
    if(N9417) begin
      \nz.mem_3040_sv2v_reg  <= data_i[0];
    end 
    if(N9416) begin
      \nz.mem_3039_sv2v_reg  <= data_i[79];
    end 
    if(N9415) begin
      \nz.mem_3038_sv2v_reg  <= data_i[78];
    end 
    if(N9414) begin
      \nz.mem_3037_sv2v_reg  <= data_i[77];
    end 
    if(N9413) begin
      \nz.mem_3036_sv2v_reg  <= data_i[76];
    end 
    if(N9412) begin
      \nz.mem_3035_sv2v_reg  <= data_i[75];
    end 
    if(N9411) begin
      \nz.mem_3034_sv2v_reg  <= data_i[74];
    end 
    if(N9410) begin
      \nz.mem_3033_sv2v_reg  <= data_i[73];
    end 
    if(N9409) begin
      \nz.mem_3032_sv2v_reg  <= data_i[72];
    end 
    if(N9408) begin
      \nz.mem_3031_sv2v_reg  <= data_i[71];
    end 
    if(N9407) begin
      \nz.mem_3030_sv2v_reg  <= data_i[70];
    end 
    if(N9406) begin
      \nz.mem_3029_sv2v_reg  <= data_i[69];
    end 
    if(N9405) begin
      \nz.mem_3028_sv2v_reg  <= data_i[68];
    end 
    if(N9404) begin
      \nz.mem_3027_sv2v_reg  <= data_i[67];
    end 
    if(N9403) begin
      \nz.mem_3026_sv2v_reg  <= data_i[66];
    end 
    if(N9402) begin
      \nz.mem_3025_sv2v_reg  <= data_i[65];
    end 
    if(N9401) begin
      \nz.mem_3024_sv2v_reg  <= data_i[64];
    end 
    if(N9400) begin
      \nz.mem_3023_sv2v_reg  <= data_i[63];
    end 
    if(N9399) begin
      \nz.mem_3022_sv2v_reg  <= data_i[62];
    end 
    if(N9398) begin
      \nz.mem_3021_sv2v_reg  <= data_i[61];
    end 
    if(N9397) begin
      \nz.mem_3020_sv2v_reg  <= data_i[60];
    end 
    if(N9396) begin
      \nz.mem_3019_sv2v_reg  <= data_i[59];
    end 
    if(N9395) begin
      \nz.mem_3018_sv2v_reg  <= data_i[58];
    end 
    if(N9394) begin
      \nz.mem_3017_sv2v_reg  <= data_i[57];
    end 
    if(N9393) begin
      \nz.mem_3016_sv2v_reg  <= data_i[56];
    end 
    if(N9392) begin
      \nz.mem_3015_sv2v_reg  <= data_i[55];
    end 
    if(N9391) begin
      \nz.mem_3014_sv2v_reg  <= data_i[54];
    end 
    if(N9390) begin
      \nz.mem_3013_sv2v_reg  <= data_i[53];
    end 
    if(N9389) begin
      \nz.mem_3012_sv2v_reg  <= data_i[52];
    end 
    if(N9388) begin
      \nz.mem_3011_sv2v_reg  <= data_i[51];
    end 
    if(N9387) begin
      \nz.mem_3010_sv2v_reg  <= data_i[50];
    end 
    if(N9386) begin
      \nz.mem_3009_sv2v_reg  <= data_i[49];
    end 
    if(N9385) begin
      \nz.mem_3008_sv2v_reg  <= data_i[48];
    end 
    if(N9384) begin
      \nz.mem_3007_sv2v_reg  <= data_i[47];
    end 
    if(N9383) begin
      \nz.mem_3006_sv2v_reg  <= data_i[46];
    end 
    if(N9382) begin
      \nz.mem_3005_sv2v_reg  <= data_i[45];
    end 
    if(N9381) begin
      \nz.mem_3004_sv2v_reg  <= data_i[44];
    end 
    if(N9380) begin
      \nz.mem_3003_sv2v_reg  <= data_i[43];
    end 
    if(N9379) begin
      \nz.mem_3002_sv2v_reg  <= data_i[42];
    end 
    if(N9378) begin
      \nz.mem_3001_sv2v_reg  <= data_i[41];
    end 
    if(N9377) begin
      \nz.mem_3000_sv2v_reg  <= data_i[40];
    end 
    if(N9376) begin
      \nz.mem_2999_sv2v_reg  <= data_i[39];
    end 
    if(N9375) begin
      \nz.mem_2998_sv2v_reg  <= data_i[38];
    end 
    if(N9374) begin
      \nz.mem_2997_sv2v_reg  <= data_i[37];
    end 
    if(N9373) begin
      \nz.mem_2996_sv2v_reg  <= data_i[36];
    end 
    if(N9372) begin
      \nz.mem_2995_sv2v_reg  <= data_i[35];
    end 
    if(N9371) begin
      \nz.mem_2994_sv2v_reg  <= data_i[34];
    end 
    if(N9370) begin
      \nz.mem_2993_sv2v_reg  <= data_i[33];
    end 
    if(N9369) begin
      \nz.mem_2992_sv2v_reg  <= data_i[32];
    end 
    if(N9368) begin
      \nz.mem_2991_sv2v_reg  <= data_i[31];
    end 
    if(N9367) begin
      \nz.mem_2990_sv2v_reg  <= data_i[30];
    end 
    if(N9366) begin
      \nz.mem_2989_sv2v_reg  <= data_i[29];
    end 
    if(N9365) begin
      \nz.mem_2988_sv2v_reg  <= data_i[28];
    end 
    if(N9364) begin
      \nz.mem_2987_sv2v_reg  <= data_i[27];
    end 
    if(N9363) begin
      \nz.mem_2986_sv2v_reg  <= data_i[26];
    end 
    if(N9362) begin
      \nz.mem_2985_sv2v_reg  <= data_i[25];
    end 
    if(N9361) begin
      \nz.mem_2984_sv2v_reg  <= data_i[24];
    end 
    if(N9360) begin
      \nz.mem_2983_sv2v_reg  <= data_i[23];
    end 
    if(N9359) begin
      \nz.mem_2982_sv2v_reg  <= data_i[22];
    end 
    if(N9358) begin
      \nz.mem_2981_sv2v_reg  <= data_i[21];
    end 
    if(N9357) begin
      \nz.mem_2980_sv2v_reg  <= data_i[20];
    end 
    if(N9356) begin
      \nz.mem_2979_sv2v_reg  <= data_i[19];
    end 
    if(N9355) begin
      \nz.mem_2978_sv2v_reg  <= data_i[18];
    end 
    if(N9354) begin
      \nz.mem_2977_sv2v_reg  <= data_i[17];
    end 
    if(N9353) begin
      \nz.mem_2976_sv2v_reg  <= data_i[16];
    end 
    if(N9352) begin
      \nz.mem_2975_sv2v_reg  <= data_i[15];
    end 
    if(N9351) begin
      \nz.mem_2974_sv2v_reg  <= data_i[14];
    end 
    if(N9350) begin
      \nz.mem_2973_sv2v_reg  <= data_i[13];
    end 
    if(N9349) begin
      \nz.mem_2972_sv2v_reg  <= data_i[12];
    end 
    if(N9348) begin
      \nz.mem_2971_sv2v_reg  <= data_i[11];
    end 
    if(N9347) begin
      \nz.mem_2970_sv2v_reg  <= data_i[10];
    end 
    if(N9346) begin
      \nz.mem_2969_sv2v_reg  <= data_i[9];
    end 
    if(N9345) begin
      \nz.mem_2968_sv2v_reg  <= data_i[8];
    end 
    if(N9344) begin
      \nz.mem_2967_sv2v_reg  <= data_i[7];
    end 
    if(N9343) begin
      \nz.mem_2966_sv2v_reg  <= data_i[6];
    end 
    if(N9342) begin
      \nz.mem_2965_sv2v_reg  <= data_i[5];
    end 
    if(N9341) begin
      \nz.mem_2964_sv2v_reg  <= data_i[4];
    end 
    if(N9340) begin
      \nz.mem_2963_sv2v_reg  <= data_i[3];
    end 
    if(N9339) begin
      \nz.mem_2962_sv2v_reg  <= data_i[2];
    end 
    if(N9338) begin
      \nz.mem_2961_sv2v_reg  <= data_i[1];
    end 
    if(N9337) begin
      \nz.mem_2960_sv2v_reg  <= data_i[0];
    end 
    if(N9336) begin
      \nz.mem_2959_sv2v_reg  <= data_i[79];
    end 
    if(N9335) begin
      \nz.mem_2958_sv2v_reg  <= data_i[78];
    end 
    if(N9334) begin
      \nz.mem_2957_sv2v_reg  <= data_i[77];
    end 
    if(N9333) begin
      \nz.mem_2956_sv2v_reg  <= data_i[76];
    end 
    if(N9332) begin
      \nz.mem_2955_sv2v_reg  <= data_i[75];
    end 
    if(N9331) begin
      \nz.mem_2954_sv2v_reg  <= data_i[74];
    end 
    if(N9330) begin
      \nz.mem_2953_sv2v_reg  <= data_i[73];
    end 
    if(N9329) begin
      \nz.mem_2952_sv2v_reg  <= data_i[72];
    end 
    if(N9328) begin
      \nz.mem_2951_sv2v_reg  <= data_i[71];
    end 
    if(N9327) begin
      \nz.mem_2950_sv2v_reg  <= data_i[70];
    end 
    if(N9326) begin
      \nz.mem_2949_sv2v_reg  <= data_i[69];
    end 
    if(N9325) begin
      \nz.mem_2948_sv2v_reg  <= data_i[68];
    end 
    if(N9324) begin
      \nz.mem_2947_sv2v_reg  <= data_i[67];
    end 
    if(N9323) begin
      \nz.mem_2946_sv2v_reg  <= data_i[66];
    end 
    if(N9322) begin
      \nz.mem_2945_sv2v_reg  <= data_i[65];
    end 
    if(N9321) begin
      \nz.mem_2944_sv2v_reg  <= data_i[64];
    end 
    if(N9320) begin
      \nz.mem_2943_sv2v_reg  <= data_i[63];
    end 
    if(N9319) begin
      \nz.mem_2942_sv2v_reg  <= data_i[62];
    end 
    if(N9318) begin
      \nz.mem_2941_sv2v_reg  <= data_i[61];
    end 
    if(N9317) begin
      \nz.mem_2940_sv2v_reg  <= data_i[60];
    end 
    if(N9316) begin
      \nz.mem_2939_sv2v_reg  <= data_i[59];
    end 
    if(N9315) begin
      \nz.mem_2938_sv2v_reg  <= data_i[58];
    end 
    if(N9314) begin
      \nz.mem_2937_sv2v_reg  <= data_i[57];
    end 
    if(N9313) begin
      \nz.mem_2936_sv2v_reg  <= data_i[56];
    end 
    if(N9312) begin
      \nz.mem_2935_sv2v_reg  <= data_i[55];
    end 
    if(N9311) begin
      \nz.mem_2934_sv2v_reg  <= data_i[54];
    end 
    if(N9310) begin
      \nz.mem_2933_sv2v_reg  <= data_i[53];
    end 
    if(N9309) begin
      \nz.mem_2932_sv2v_reg  <= data_i[52];
    end 
    if(N9308) begin
      \nz.mem_2931_sv2v_reg  <= data_i[51];
    end 
    if(N9307) begin
      \nz.mem_2930_sv2v_reg  <= data_i[50];
    end 
    if(N9306) begin
      \nz.mem_2929_sv2v_reg  <= data_i[49];
    end 
    if(N9305) begin
      \nz.mem_2928_sv2v_reg  <= data_i[48];
    end 
    if(N9304) begin
      \nz.mem_2927_sv2v_reg  <= data_i[47];
    end 
    if(N9303) begin
      \nz.mem_2926_sv2v_reg  <= data_i[46];
    end 
    if(N9302) begin
      \nz.mem_2925_sv2v_reg  <= data_i[45];
    end 
    if(N9301) begin
      \nz.mem_2924_sv2v_reg  <= data_i[44];
    end 
    if(N9300) begin
      \nz.mem_2923_sv2v_reg  <= data_i[43];
    end 
    if(N9299) begin
      \nz.mem_2922_sv2v_reg  <= data_i[42];
    end 
    if(N9298) begin
      \nz.mem_2921_sv2v_reg  <= data_i[41];
    end 
    if(N9297) begin
      \nz.mem_2920_sv2v_reg  <= data_i[40];
    end 
    if(N9296) begin
      \nz.mem_2919_sv2v_reg  <= data_i[39];
    end 
    if(N9295) begin
      \nz.mem_2918_sv2v_reg  <= data_i[38];
    end 
    if(N9294) begin
      \nz.mem_2917_sv2v_reg  <= data_i[37];
    end 
    if(N9293) begin
      \nz.mem_2916_sv2v_reg  <= data_i[36];
    end 
    if(N9292) begin
      \nz.mem_2915_sv2v_reg  <= data_i[35];
    end 
    if(N9291) begin
      \nz.mem_2914_sv2v_reg  <= data_i[34];
    end 
    if(N9290) begin
      \nz.mem_2913_sv2v_reg  <= data_i[33];
    end 
    if(N9289) begin
      \nz.mem_2912_sv2v_reg  <= data_i[32];
    end 
    if(N9288) begin
      \nz.mem_2911_sv2v_reg  <= data_i[31];
    end 
    if(N9287) begin
      \nz.mem_2910_sv2v_reg  <= data_i[30];
    end 
    if(N9286) begin
      \nz.mem_2909_sv2v_reg  <= data_i[29];
    end 
    if(N9285) begin
      \nz.mem_2908_sv2v_reg  <= data_i[28];
    end 
    if(N9284) begin
      \nz.mem_2907_sv2v_reg  <= data_i[27];
    end 
    if(N9283) begin
      \nz.mem_2906_sv2v_reg  <= data_i[26];
    end 
    if(N9282) begin
      \nz.mem_2905_sv2v_reg  <= data_i[25];
    end 
    if(N9281) begin
      \nz.mem_2904_sv2v_reg  <= data_i[24];
    end 
    if(N9280) begin
      \nz.mem_2903_sv2v_reg  <= data_i[23];
    end 
    if(N9279) begin
      \nz.mem_2902_sv2v_reg  <= data_i[22];
    end 
    if(N9278) begin
      \nz.mem_2901_sv2v_reg  <= data_i[21];
    end 
    if(N9277) begin
      \nz.mem_2900_sv2v_reg  <= data_i[20];
    end 
    if(N9276) begin
      \nz.mem_2899_sv2v_reg  <= data_i[19];
    end 
    if(N9275) begin
      \nz.mem_2898_sv2v_reg  <= data_i[18];
    end 
    if(N9274) begin
      \nz.mem_2897_sv2v_reg  <= data_i[17];
    end 
    if(N9273) begin
      \nz.mem_2896_sv2v_reg  <= data_i[16];
    end 
    if(N9272) begin
      \nz.mem_2895_sv2v_reg  <= data_i[15];
    end 
    if(N9271) begin
      \nz.mem_2894_sv2v_reg  <= data_i[14];
    end 
    if(N9270) begin
      \nz.mem_2893_sv2v_reg  <= data_i[13];
    end 
    if(N9269) begin
      \nz.mem_2892_sv2v_reg  <= data_i[12];
    end 
    if(N9268) begin
      \nz.mem_2891_sv2v_reg  <= data_i[11];
    end 
    if(N9267) begin
      \nz.mem_2890_sv2v_reg  <= data_i[10];
    end 
    if(N9266) begin
      \nz.mem_2889_sv2v_reg  <= data_i[9];
    end 
    if(N9265) begin
      \nz.mem_2888_sv2v_reg  <= data_i[8];
    end 
    if(N9264) begin
      \nz.mem_2887_sv2v_reg  <= data_i[7];
    end 
    if(N9263) begin
      \nz.mem_2886_sv2v_reg  <= data_i[6];
    end 
    if(N9262) begin
      \nz.mem_2885_sv2v_reg  <= data_i[5];
    end 
    if(N9261) begin
      \nz.mem_2884_sv2v_reg  <= data_i[4];
    end 
    if(N9260) begin
      \nz.mem_2883_sv2v_reg  <= data_i[3];
    end 
    if(N9259) begin
      \nz.mem_2882_sv2v_reg  <= data_i[2];
    end 
    if(N9258) begin
      \nz.mem_2881_sv2v_reg  <= data_i[1];
    end 
    if(N9257) begin
      \nz.mem_2880_sv2v_reg  <= data_i[0];
    end 
    if(N9256) begin
      \nz.mem_2879_sv2v_reg  <= data_i[79];
    end 
    if(N9255) begin
      \nz.mem_2878_sv2v_reg  <= data_i[78];
    end 
    if(N9254) begin
      \nz.mem_2877_sv2v_reg  <= data_i[77];
    end 
    if(N9253) begin
      \nz.mem_2876_sv2v_reg  <= data_i[76];
    end 
    if(N9252) begin
      \nz.mem_2875_sv2v_reg  <= data_i[75];
    end 
    if(N9251) begin
      \nz.mem_2874_sv2v_reg  <= data_i[74];
    end 
    if(N9250) begin
      \nz.mem_2873_sv2v_reg  <= data_i[73];
    end 
    if(N9249) begin
      \nz.mem_2872_sv2v_reg  <= data_i[72];
    end 
    if(N9248) begin
      \nz.mem_2871_sv2v_reg  <= data_i[71];
    end 
    if(N9247) begin
      \nz.mem_2870_sv2v_reg  <= data_i[70];
    end 
    if(N9246) begin
      \nz.mem_2869_sv2v_reg  <= data_i[69];
    end 
    if(N9245) begin
      \nz.mem_2868_sv2v_reg  <= data_i[68];
    end 
    if(N9244) begin
      \nz.mem_2867_sv2v_reg  <= data_i[67];
    end 
    if(N9243) begin
      \nz.mem_2866_sv2v_reg  <= data_i[66];
    end 
    if(N9242) begin
      \nz.mem_2865_sv2v_reg  <= data_i[65];
    end 
    if(N9241) begin
      \nz.mem_2864_sv2v_reg  <= data_i[64];
    end 
    if(N9240) begin
      \nz.mem_2863_sv2v_reg  <= data_i[63];
    end 
    if(N9239) begin
      \nz.mem_2862_sv2v_reg  <= data_i[62];
    end 
    if(N9238) begin
      \nz.mem_2861_sv2v_reg  <= data_i[61];
    end 
    if(N9237) begin
      \nz.mem_2860_sv2v_reg  <= data_i[60];
    end 
    if(N9236) begin
      \nz.mem_2859_sv2v_reg  <= data_i[59];
    end 
    if(N9235) begin
      \nz.mem_2858_sv2v_reg  <= data_i[58];
    end 
    if(N9234) begin
      \nz.mem_2857_sv2v_reg  <= data_i[57];
    end 
    if(N9233) begin
      \nz.mem_2856_sv2v_reg  <= data_i[56];
    end 
    if(N9232) begin
      \nz.mem_2855_sv2v_reg  <= data_i[55];
    end 
    if(N9231) begin
      \nz.mem_2854_sv2v_reg  <= data_i[54];
    end 
    if(N9230) begin
      \nz.mem_2853_sv2v_reg  <= data_i[53];
    end 
    if(N9229) begin
      \nz.mem_2852_sv2v_reg  <= data_i[52];
    end 
    if(N9228) begin
      \nz.mem_2851_sv2v_reg  <= data_i[51];
    end 
    if(N9227) begin
      \nz.mem_2850_sv2v_reg  <= data_i[50];
    end 
    if(N9226) begin
      \nz.mem_2849_sv2v_reg  <= data_i[49];
    end 
    if(N9225) begin
      \nz.mem_2848_sv2v_reg  <= data_i[48];
    end 
    if(N9224) begin
      \nz.mem_2847_sv2v_reg  <= data_i[47];
    end 
    if(N9223) begin
      \nz.mem_2846_sv2v_reg  <= data_i[46];
    end 
    if(N9222) begin
      \nz.mem_2845_sv2v_reg  <= data_i[45];
    end 
    if(N9221) begin
      \nz.mem_2844_sv2v_reg  <= data_i[44];
    end 
    if(N9220) begin
      \nz.mem_2843_sv2v_reg  <= data_i[43];
    end 
    if(N9219) begin
      \nz.mem_2842_sv2v_reg  <= data_i[42];
    end 
    if(N9218) begin
      \nz.mem_2841_sv2v_reg  <= data_i[41];
    end 
    if(N9217) begin
      \nz.mem_2840_sv2v_reg  <= data_i[40];
    end 
    if(N9216) begin
      \nz.mem_2839_sv2v_reg  <= data_i[39];
    end 
    if(N9215) begin
      \nz.mem_2838_sv2v_reg  <= data_i[38];
    end 
    if(N9214) begin
      \nz.mem_2837_sv2v_reg  <= data_i[37];
    end 
    if(N9213) begin
      \nz.mem_2836_sv2v_reg  <= data_i[36];
    end 
    if(N9212) begin
      \nz.mem_2835_sv2v_reg  <= data_i[35];
    end 
    if(N9211) begin
      \nz.mem_2834_sv2v_reg  <= data_i[34];
    end 
    if(N9210) begin
      \nz.mem_2833_sv2v_reg  <= data_i[33];
    end 
    if(N9209) begin
      \nz.mem_2832_sv2v_reg  <= data_i[32];
    end 
    if(N9208) begin
      \nz.mem_2831_sv2v_reg  <= data_i[31];
    end 
    if(N9207) begin
      \nz.mem_2830_sv2v_reg  <= data_i[30];
    end 
    if(N9206) begin
      \nz.mem_2829_sv2v_reg  <= data_i[29];
    end 
    if(N9205) begin
      \nz.mem_2828_sv2v_reg  <= data_i[28];
    end 
    if(N9204) begin
      \nz.mem_2827_sv2v_reg  <= data_i[27];
    end 
    if(N9203) begin
      \nz.mem_2826_sv2v_reg  <= data_i[26];
    end 
    if(N9202) begin
      \nz.mem_2825_sv2v_reg  <= data_i[25];
    end 
    if(N9201) begin
      \nz.mem_2824_sv2v_reg  <= data_i[24];
    end 
    if(N9200) begin
      \nz.mem_2823_sv2v_reg  <= data_i[23];
    end 
    if(N9199) begin
      \nz.mem_2822_sv2v_reg  <= data_i[22];
    end 
    if(N9198) begin
      \nz.mem_2821_sv2v_reg  <= data_i[21];
    end 
    if(N9197) begin
      \nz.mem_2820_sv2v_reg  <= data_i[20];
    end 
    if(N9196) begin
      \nz.mem_2819_sv2v_reg  <= data_i[19];
    end 
    if(N9195) begin
      \nz.mem_2818_sv2v_reg  <= data_i[18];
    end 
    if(N9194) begin
      \nz.mem_2817_sv2v_reg  <= data_i[17];
    end 
    if(N9193) begin
      \nz.mem_2816_sv2v_reg  <= data_i[16];
    end 
    if(N9192) begin
      \nz.mem_2815_sv2v_reg  <= data_i[15];
    end 
    if(N9191) begin
      \nz.mem_2814_sv2v_reg  <= data_i[14];
    end 
    if(N9190) begin
      \nz.mem_2813_sv2v_reg  <= data_i[13];
    end 
    if(N9189) begin
      \nz.mem_2812_sv2v_reg  <= data_i[12];
    end 
    if(N9188) begin
      \nz.mem_2811_sv2v_reg  <= data_i[11];
    end 
    if(N9187) begin
      \nz.mem_2810_sv2v_reg  <= data_i[10];
    end 
    if(N9186) begin
      \nz.mem_2809_sv2v_reg  <= data_i[9];
    end 
    if(N9185) begin
      \nz.mem_2808_sv2v_reg  <= data_i[8];
    end 
    if(N9184) begin
      \nz.mem_2807_sv2v_reg  <= data_i[7];
    end 
    if(N9183) begin
      \nz.mem_2806_sv2v_reg  <= data_i[6];
    end 
    if(N9182) begin
      \nz.mem_2805_sv2v_reg  <= data_i[5];
    end 
    if(N9181) begin
      \nz.mem_2804_sv2v_reg  <= data_i[4];
    end 
    if(N9180) begin
      \nz.mem_2803_sv2v_reg  <= data_i[3];
    end 
    if(N9179) begin
      \nz.mem_2802_sv2v_reg  <= data_i[2];
    end 
    if(N9178) begin
      \nz.mem_2801_sv2v_reg  <= data_i[1];
    end 
    if(N9177) begin
      \nz.mem_2800_sv2v_reg  <= data_i[0];
    end 
    if(N9176) begin
      \nz.mem_2799_sv2v_reg  <= data_i[79];
    end 
    if(N9175) begin
      \nz.mem_2798_sv2v_reg  <= data_i[78];
    end 
    if(N9174) begin
      \nz.mem_2797_sv2v_reg  <= data_i[77];
    end 
    if(N9173) begin
      \nz.mem_2796_sv2v_reg  <= data_i[76];
    end 
    if(N9172) begin
      \nz.mem_2795_sv2v_reg  <= data_i[75];
    end 
    if(N9171) begin
      \nz.mem_2794_sv2v_reg  <= data_i[74];
    end 
    if(N9170) begin
      \nz.mem_2793_sv2v_reg  <= data_i[73];
    end 
    if(N9169) begin
      \nz.mem_2792_sv2v_reg  <= data_i[72];
    end 
    if(N9168) begin
      \nz.mem_2791_sv2v_reg  <= data_i[71];
    end 
    if(N9167) begin
      \nz.mem_2790_sv2v_reg  <= data_i[70];
    end 
    if(N9166) begin
      \nz.mem_2789_sv2v_reg  <= data_i[69];
    end 
    if(N9165) begin
      \nz.mem_2788_sv2v_reg  <= data_i[68];
    end 
    if(N9164) begin
      \nz.mem_2787_sv2v_reg  <= data_i[67];
    end 
    if(N9163) begin
      \nz.mem_2786_sv2v_reg  <= data_i[66];
    end 
    if(N9162) begin
      \nz.mem_2785_sv2v_reg  <= data_i[65];
    end 
    if(N9161) begin
      \nz.mem_2784_sv2v_reg  <= data_i[64];
    end 
    if(N9160) begin
      \nz.mem_2783_sv2v_reg  <= data_i[63];
    end 
    if(N9159) begin
      \nz.mem_2782_sv2v_reg  <= data_i[62];
    end 
    if(N9158) begin
      \nz.mem_2781_sv2v_reg  <= data_i[61];
    end 
    if(N9157) begin
      \nz.mem_2780_sv2v_reg  <= data_i[60];
    end 
    if(N9156) begin
      \nz.mem_2779_sv2v_reg  <= data_i[59];
    end 
    if(N9155) begin
      \nz.mem_2778_sv2v_reg  <= data_i[58];
    end 
    if(N9154) begin
      \nz.mem_2777_sv2v_reg  <= data_i[57];
    end 
    if(N9153) begin
      \nz.mem_2776_sv2v_reg  <= data_i[56];
    end 
    if(N9152) begin
      \nz.mem_2775_sv2v_reg  <= data_i[55];
    end 
    if(N9151) begin
      \nz.mem_2774_sv2v_reg  <= data_i[54];
    end 
    if(N9150) begin
      \nz.mem_2773_sv2v_reg  <= data_i[53];
    end 
    if(N9149) begin
      \nz.mem_2772_sv2v_reg  <= data_i[52];
    end 
    if(N9148) begin
      \nz.mem_2771_sv2v_reg  <= data_i[51];
    end 
    if(N9147) begin
      \nz.mem_2770_sv2v_reg  <= data_i[50];
    end 
    if(N9146) begin
      \nz.mem_2769_sv2v_reg  <= data_i[49];
    end 
    if(N9145) begin
      \nz.mem_2768_sv2v_reg  <= data_i[48];
    end 
    if(N9144) begin
      \nz.mem_2767_sv2v_reg  <= data_i[47];
    end 
    if(N9143) begin
      \nz.mem_2766_sv2v_reg  <= data_i[46];
    end 
    if(N9142) begin
      \nz.mem_2765_sv2v_reg  <= data_i[45];
    end 
    if(N9141) begin
      \nz.mem_2764_sv2v_reg  <= data_i[44];
    end 
    if(N9140) begin
      \nz.mem_2763_sv2v_reg  <= data_i[43];
    end 
    if(N9139) begin
      \nz.mem_2762_sv2v_reg  <= data_i[42];
    end 
    if(N9138) begin
      \nz.mem_2761_sv2v_reg  <= data_i[41];
    end 
    if(N9137) begin
      \nz.mem_2760_sv2v_reg  <= data_i[40];
    end 
    if(N9136) begin
      \nz.mem_2759_sv2v_reg  <= data_i[39];
    end 
    if(N9135) begin
      \nz.mem_2758_sv2v_reg  <= data_i[38];
    end 
    if(N9134) begin
      \nz.mem_2757_sv2v_reg  <= data_i[37];
    end 
    if(N9133) begin
      \nz.mem_2756_sv2v_reg  <= data_i[36];
    end 
    if(N9132) begin
      \nz.mem_2755_sv2v_reg  <= data_i[35];
    end 
    if(N9131) begin
      \nz.mem_2754_sv2v_reg  <= data_i[34];
    end 
    if(N9130) begin
      \nz.mem_2753_sv2v_reg  <= data_i[33];
    end 
    if(N9129) begin
      \nz.mem_2752_sv2v_reg  <= data_i[32];
    end 
    if(N9128) begin
      \nz.mem_2751_sv2v_reg  <= data_i[31];
    end 
    if(N9127) begin
      \nz.mem_2750_sv2v_reg  <= data_i[30];
    end 
    if(N9126) begin
      \nz.mem_2749_sv2v_reg  <= data_i[29];
    end 
    if(N9125) begin
      \nz.mem_2748_sv2v_reg  <= data_i[28];
    end 
    if(N9124) begin
      \nz.mem_2747_sv2v_reg  <= data_i[27];
    end 
    if(N9123) begin
      \nz.mem_2746_sv2v_reg  <= data_i[26];
    end 
    if(N9122) begin
      \nz.mem_2745_sv2v_reg  <= data_i[25];
    end 
    if(N9121) begin
      \nz.mem_2744_sv2v_reg  <= data_i[24];
    end 
    if(N9120) begin
      \nz.mem_2743_sv2v_reg  <= data_i[23];
    end 
    if(N9119) begin
      \nz.mem_2742_sv2v_reg  <= data_i[22];
    end 
    if(N9118) begin
      \nz.mem_2741_sv2v_reg  <= data_i[21];
    end 
    if(N9117) begin
      \nz.mem_2740_sv2v_reg  <= data_i[20];
    end 
    if(N9116) begin
      \nz.mem_2739_sv2v_reg  <= data_i[19];
    end 
    if(N9115) begin
      \nz.mem_2738_sv2v_reg  <= data_i[18];
    end 
    if(N9114) begin
      \nz.mem_2737_sv2v_reg  <= data_i[17];
    end 
    if(N9113) begin
      \nz.mem_2736_sv2v_reg  <= data_i[16];
    end 
    if(N9112) begin
      \nz.mem_2735_sv2v_reg  <= data_i[15];
    end 
    if(N9111) begin
      \nz.mem_2734_sv2v_reg  <= data_i[14];
    end 
    if(N9110) begin
      \nz.mem_2733_sv2v_reg  <= data_i[13];
    end 
    if(N9109) begin
      \nz.mem_2732_sv2v_reg  <= data_i[12];
    end 
    if(N9108) begin
      \nz.mem_2731_sv2v_reg  <= data_i[11];
    end 
    if(N9107) begin
      \nz.mem_2730_sv2v_reg  <= data_i[10];
    end 
    if(N9106) begin
      \nz.mem_2729_sv2v_reg  <= data_i[9];
    end 
    if(N9105) begin
      \nz.mem_2728_sv2v_reg  <= data_i[8];
    end 
    if(N9104) begin
      \nz.mem_2727_sv2v_reg  <= data_i[7];
    end 
    if(N9103) begin
      \nz.mem_2726_sv2v_reg  <= data_i[6];
    end 
    if(N9102) begin
      \nz.mem_2725_sv2v_reg  <= data_i[5];
    end 
    if(N9101) begin
      \nz.mem_2724_sv2v_reg  <= data_i[4];
    end 
    if(N9100) begin
      \nz.mem_2723_sv2v_reg  <= data_i[3];
    end 
    if(N9099) begin
      \nz.mem_2722_sv2v_reg  <= data_i[2];
    end 
    if(N9098) begin
      \nz.mem_2721_sv2v_reg  <= data_i[1];
    end 
    if(N9097) begin
      \nz.mem_2720_sv2v_reg  <= data_i[0];
    end 
    if(N9096) begin
      \nz.mem_2719_sv2v_reg  <= data_i[79];
    end 
    if(N9095) begin
      \nz.mem_2718_sv2v_reg  <= data_i[78];
    end 
    if(N9094) begin
      \nz.mem_2717_sv2v_reg  <= data_i[77];
    end 
    if(N9093) begin
      \nz.mem_2716_sv2v_reg  <= data_i[76];
    end 
    if(N9092) begin
      \nz.mem_2715_sv2v_reg  <= data_i[75];
    end 
    if(N9091) begin
      \nz.mem_2714_sv2v_reg  <= data_i[74];
    end 
    if(N9090) begin
      \nz.mem_2713_sv2v_reg  <= data_i[73];
    end 
    if(N9089) begin
      \nz.mem_2712_sv2v_reg  <= data_i[72];
    end 
    if(N9088) begin
      \nz.mem_2711_sv2v_reg  <= data_i[71];
    end 
    if(N9087) begin
      \nz.mem_2710_sv2v_reg  <= data_i[70];
    end 
    if(N9086) begin
      \nz.mem_2709_sv2v_reg  <= data_i[69];
    end 
    if(N9085) begin
      \nz.mem_2708_sv2v_reg  <= data_i[68];
    end 
    if(N9084) begin
      \nz.mem_2707_sv2v_reg  <= data_i[67];
    end 
    if(N9083) begin
      \nz.mem_2706_sv2v_reg  <= data_i[66];
    end 
    if(N9082) begin
      \nz.mem_2705_sv2v_reg  <= data_i[65];
    end 
    if(N9081) begin
      \nz.mem_2704_sv2v_reg  <= data_i[64];
    end 
    if(N9080) begin
      \nz.mem_2703_sv2v_reg  <= data_i[63];
    end 
    if(N9079) begin
      \nz.mem_2702_sv2v_reg  <= data_i[62];
    end 
    if(N9078) begin
      \nz.mem_2701_sv2v_reg  <= data_i[61];
    end 
    if(N9077) begin
      \nz.mem_2700_sv2v_reg  <= data_i[60];
    end 
    if(N9076) begin
      \nz.mem_2699_sv2v_reg  <= data_i[59];
    end 
    if(N9075) begin
      \nz.mem_2698_sv2v_reg  <= data_i[58];
    end 
    if(N9074) begin
      \nz.mem_2697_sv2v_reg  <= data_i[57];
    end 
    if(N9073) begin
      \nz.mem_2696_sv2v_reg  <= data_i[56];
    end 
    if(N9072) begin
      \nz.mem_2695_sv2v_reg  <= data_i[55];
    end 
    if(N9071) begin
      \nz.mem_2694_sv2v_reg  <= data_i[54];
    end 
    if(N9070) begin
      \nz.mem_2693_sv2v_reg  <= data_i[53];
    end 
    if(N9069) begin
      \nz.mem_2692_sv2v_reg  <= data_i[52];
    end 
    if(N9068) begin
      \nz.mem_2691_sv2v_reg  <= data_i[51];
    end 
    if(N9067) begin
      \nz.mem_2690_sv2v_reg  <= data_i[50];
    end 
    if(N9066) begin
      \nz.mem_2689_sv2v_reg  <= data_i[49];
    end 
    if(N9065) begin
      \nz.mem_2688_sv2v_reg  <= data_i[48];
    end 
    if(N9064) begin
      \nz.mem_2687_sv2v_reg  <= data_i[47];
    end 
    if(N9063) begin
      \nz.mem_2686_sv2v_reg  <= data_i[46];
    end 
    if(N9062) begin
      \nz.mem_2685_sv2v_reg  <= data_i[45];
    end 
    if(N9061) begin
      \nz.mem_2684_sv2v_reg  <= data_i[44];
    end 
    if(N9060) begin
      \nz.mem_2683_sv2v_reg  <= data_i[43];
    end 
    if(N9059) begin
      \nz.mem_2682_sv2v_reg  <= data_i[42];
    end 
    if(N9058) begin
      \nz.mem_2681_sv2v_reg  <= data_i[41];
    end 
    if(N9057) begin
      \nz.mem_2680_sv2v_reg  <= data_i[40];
    end 
    if(N9056) begin
      \nz.mem_2679_sv2v_reg  <= data_i[39];
    end 
    if(N9055) begin
      \nz.mem_2678_sv2v_reg  <= data_i[38];
    end 
    if(N9054) begin
      \nz.mem_2677_sv2v_reg  <= data_i[37];
    end 
    if(N9053) begin
      \nz.mem_2676_sv2v_reg  <= data_i[36];
    end 
    if(N9052) begin
      \nz.mem_2675_sv2v_reg  <= data_i[35];
    end 
    if(N9051) begin
      \nz.mem_2674_sv2v_reg  <= data_i[34];
    end 
    if(N9050) begin
      \nz.mem_2673_sv2v_reg  <= data_i[33];
    end 
    if(N9049) begin
      \nz.mem_2672_sv2v_reg  <= data_i[32];
    end 
    if(N9048) begin
      \nz.mem_2671_sv2v_reg  <= data_i[31];
    end 
    if(N9047) begin
      \nz.mem_2670_sv2v_reg  <= data_i[30];
    end 
    if(N9046) begin
      \nz.mem_2669_sv2v_reg  <= data_i[29];
    end 
    if(N9045) begin
      \nz.mem_2668_sv2v_reg  <= data_i[28];
    end 
    if(N9044) begin
      \nz.mem_2667_sv2v_reg  <= data_i[27];
    end 
    if(N9043) begin
      \nz.mem_2666_sv2v_reg  <= data_i[26];
    end 
    if(N9042) begin
      \nz.mem_2665_sv2v_reg  <= data_i[25];
    end 
    if(N9041) begin
      \nz.mem_2664_sv2v_reg  <= data_i[24];
    end 
    if(N9040) begin
      \nz.mem_2663_sv2v_reg  <= data_i[23];
    end 
    if(N9039) begin
      \nz.mem_2662_sv2v_reg  <= data_i[22];
    end 
    if(N9038) begin
      \nz.mem_2661_sv2v_reg  <= data_i[21];
    end 
    if(N9037) begin
      \nz.mem_2660_sv2v_reg  <= data_i[20];
    end 
    if(N9036) begin
      \nz.mem_2659_sv2v_reg  <= data_i[19];
    end 
    if(N9035) begin
      \nz.mem_2658_sv2v_reg  <= data_i[18];
    end 
    if(N9034) begin
      \nz.mem_2657_sv2v_reg  <= data_i[17];
    end 
    if(N9033) begin
      \nz.mem_2656_sv2v_reg  <= data_i[16];
    end 
    if(N9032) begin
      \nz.mem_2655_sv2v_reg  <= data_i[15];
    end 
    if(N9031) begin
      \nz.mem_2654_sv2v_reg  <= data_i[14];
    end 
    if(N9030) begin
      \nz.mem_2653_sv2v_reg  <= data_i[13];
    end 
    if(N9029) begin
      \nz.mem_2652_sv2v_reg  <= data_i[12];
    end 
    if(N9028) begin
      \nz.mem_2651_sv2v_reg  <= data_i[11];
    end 
    if(N9027) begin
      \nz.mem_2650_sv2v_reg  <= data_i[10];
    end 
    if(N9026) begin
      \nz.mem_2649_sv2v_reg  <= data_i[9];
    end 
    if(N9025) begin
      \nz.mem_2648_sv2v_reg  <= data_i[8];
    end 
    if(N9024) begin
      \nz.mem_2647_sv2v_reg  <= data_i[7];
    end 
    if(N9023) begin
      \nz.mem_2646_sv2v_reg  <= data_i[6];
    end 
    if(N9022) begin
      \nz.mem_2645_sv2v_reg  <= data_i[5];
    end 
    if(N9021) begin
      \nz.mem_2644_sv2v_reg  <= data_i[4];
    end 
    if(N9020) begin
      \nz.mem_2643_sv2v_reg  <= data_i[3];
    end 
    if(N9019) begin
      \nz.mem_2642_sv2v_reg  <= data_i[2];
    end 
    if(N9018) begin
      \nz.mem_2641_sv2v_reg  <= data_i[1];
    end 
    if(N9017) begin
      \nz.mem_2640_sv2v_reg  <= data_i[0];
    end 
    if(N9016) begin
      \nz.mem_2639_sv2v_reg  <= data_i[79];
    end 
    if(N9015) begin
      \nz.mem_2638_sv2v_reg  <= data_i[78];
    end 
    if(N9014) begin
      \nz.mem_2637_sv2v_reg  <= data_i[77];
    end 
    if(N9013) begin
      \nz.mem_2636_sv2v_reg  <= data_i[76];
    end 
    if(N9012) begin
      \nz.mem_2635_sv2v_reg  <= data_i[75];
    end 
    if(N9011) begin
      \nz.mem_2634_sv2v_reg  <= data_i[74];
    end 
    if(N9010) begin
      \nz.mem_2633_sv2v_reg  <= data_i[73];
    end 
    if(N9009) begin
      \nz.mem_2632_sv2v_reg  <= data_i[72];
    end 
    if(N9008) begin
      \nz.mem_2631_sv2v_reg  <= data_i[71];
    end 
    if(N9007) begin
      \nz.mem_2630_sv2v_reg  <= data_i[70];
    end 
    if(N9006) begin
      \nz.mem_2629_sv2v_reg  <= data_i[69];
    end 
    if(N9005) begin
      \nz.mem_2628_sv2v_reg  <= data_i[68];
    end 
    if(N9004) begin
      \nz.mem_2627_sv2v_reg  <= data_i[67];
    end 
    if(N9003) begin
      \nz.mem_2626_sv2v_reg  <= data_i[66];
    end 
    if(N9002) begin
      \nz.mem_2625_sv2v_reg  <= data_i[65];
    end 
    if(N9001) begin
      \nz.mem_2624_sv2v_reg  <= data_i[64];
    end 
    if(N9000) begin
      \nz.mem_2623_sv2v_reg  <= data_i[63];
    end 
    if(N8999) begin
      \nz.mem_2622_sv2v_reg  <= data_i[62];
    end 
    if(N8998) begin
      \nz.mem_2621_sv2v_reg  <= data_i[61];
    end 
    if(N8997) begin
      \nz.mem_2620_sv2v_reg  <= data_i[60];
    end 
    if(N8996) begin
      \nz.mem_2619_sv2v_reg  <= data_i[59];
    end 
    if(N8995) begin
      \nz.mem_2618_sv2v_reg  <= data_i[58];
    end 
    if(N8994) begin
      \nz.mem_2617_sv2v_reg  <= data_i[57];
    end 
    if(N8993) begin
      \nz.mem_2616_sv2v_reg  <= data_i[56];
    end 
    if(N8992) begin
      \nz.mem_2615_sv2v_reg  <= data_i[55];
    end 
    if(N8991) begin
      \nz.mem_2614_sv2v_reg  <= data_i[54];
    end 
    if(N8990) begin
      \nz.mem_2613_sv2v_reg  <= data_i[53];
    end 
    if(N8989) begin
      \nz.mem_2612_sv2v_reg  <= data_i[52];
    end 
    if(N8988) begin
      \nz.mem_2611_sv2v_reg  <= data_i[51];
    end 
    if(N8987) begin
      \nz.mem_2610_sv2v_reg  <= data_i[50];
    end 
    if(N8986) begin
      \nz.mem_2609_sv2v_reg  <= data_i[49];
    end 
    if(N8985) begin
      \nz.mem_2608_sv2v_reg  <= data_i[48];
    end 
    if(N8984) begin
      \nz.mem_2607_sv2v_reg  <= data_i[47];
    end 
    if(N8983) begin
      \nz.mem_2606_sv2v_reg  <= data_i[46];
    end 
    if(N8982) begin
      \nz.mem_2605_sv2v_reg  <= data_i[45];
    end 
    if(N8981) begin
      \nz.mem_2604_sv2v_reg  <= data_i[44];
    end 
    if(N8980) begin
      \nz.mem_2603_sv2v_reg  <= data_i[43];
    end 
    if(N8979) begin
      \nz.mem_2602_sv2v_reg  <= data_i[42];
    end 
    if(N8978) begin
      \nz.mem_2601_sv2v_reg  <= data_i[41];
    end 
    if(N8977) begin
      \nz.mem_2600_sv2v_reg  <= data_i[40];
    end 
    if(N8976) begin
      \nz.mem_2599_sv2v_reg  <= data_i[39];
    end 
    if(N8975) begin
      \nz.mem_2598_sv2v_reg  <= data_i[38];
    end 
    if(N8974) begin
      \nz.mem_2597_sv2v_reg  <= data_i[37];
    end 
    if(N8973) begin
      \nz.mem_2596_sv2v_reg  <= data_i[36];
    end 
    if(N8972) begin
      \nz.mem_2595_sv2v_reg  <= data_i[35];
    end 
    if(N8971) begin
      \nz.mem_2594_sv2v_reg  <= data_i[34];
    end 
    if(N8970) begin
      \nz.mem_2593_sv2v_reg  <= data_i[33];
    end 
    if(N8969) begin
      \nz.mem_2592_sv2v_reg  <= data_i[32];
    end 
    if(N8968) begin
      \nz.mem_2591_sv2v_reg  <= data_i[31];
    end 
    if(N8967) begin
      \nz.mem_2590_sv2v_reg  <= data_i[30];
    end 
    if(N8966) begin
      \nz.mem_2589_sv2v_reg  <= data_i[29];
    end 
    if(N8965) begin
      \nz.mem_2588_sv2v_reg  <= data_i[28];
    end 
    if(N8964) begin
      \nz.mem_2587_sv2v_reg  <= data_i[27];
    end 
    if(N8963) begin
      \nz.mem_2586_sv2v_reg  <= data_i[26];
    end 
    if(N8962) begin
      \nz.mem_2585_sv2v_reg  <= data_i[25];
    end 
    if(N8961) begin
      \nz.mem_2584_sv2v_reg  <= data_i[24];
    end 
    if(N8960) begin
      \nz.mem_2583_sv2v_reg  <= data_i[23];
    end 
    if(N8959) begin
      \nz.mem_2582_sv2v_reg  <= data_i[22];
    end 
    if(N8958) begin
      \nz.mem_2581_sv2v_reg  <= data_i[21];
    end 
    if(N8957) begin
      \nz.mem_2580_sv2v_reg  <= data_i[20];
    end 
    if(N8956) begin
      \nz.mem_2579_sv2v_reg  <= data_i[19];
    end 
    if(N8955) begin
      \nz.mem_2578_sv2v_reg  <= data_i[18];
    end 
    if(N8954) begin
      \nz.mem_2577_sv2v_reg  <= data_i[17];
    end 
    if(N8953) begin
      \nz.mem_2576_sv2v_reg  <= data_i[16];
    end 
    if(N8952) begin
      \nz.mem_2575_sv2v_reg  <= data_i[15];
    end 
    if(N8951) begin
      \nz.mem_2574_sv2v_reg  <= data_i[14];
    end 
    if(N8950) begin
      \nz.mem_2573_sv2v_reg  <= data_i[13];
    end 
    if(N8949) begin
      \nz.mem_2572_sv2v_reg  <= data_i[12];
    end 
    if(N8948) begin
      \nz.mem_2571_sv2v_reg  <= data_i[11];
    end 
    if(N8947) begin
      \nz.mem_2570_sv2v_reg  <= data_i[10];
    end 
    if(N8946) begin
      \nz.mem_2569_sv2v_reg  <= data_i[9];
    end 
    if(N8945) begin
      \nz.mem_2568_sv2v_reg  <= data_i[8];
    end 
    if(N8944) begin
      \nz.mem_2567_sv2v_reg  <= data_i[7];
    end 
    if(N8943) begin
      \nz.mem_2566_sv2v_reg  <= data_i[6];
    end 
    if(N8942) begin
      \nz.mem_2565_sv2v_reg  <= data_i[5];
    end 
    if(N8941) begin
      \nz.mem_2564_sv2v_reg  <= data_i[4];
    end 
    if(N8940) begin
      \nz.mem_2563_sv2v_reg  <= data_i[3];
    end 
    if(N8939) begin
      \nz.mem_2562_sv2v_reg  <= data_i[2];
    end 
    if(N8938) begin
      \nz.mem_2561_sv2v_reg  <= data_i[1];
    end 
    if(N8937) begin
      \nz.mem_2560_sv2v_reg  <= data_i[0];
    end 
    if(N8936) begin
      \nz.mem_2559_sv2v_reg  <= data_i[79];
    end 
    if(N8935) begin
      \nz.mem_2558_sv2v_reg  <= data_i[78];
    end 
    if(N8934) begin
      \nz.mem_2557_sv2v_reg  <= data_i[77];
    end 
    if(N8933) begin
      \nz.mem_2556_sv2v_reg  <= data_i[76];
    end 
    if(N8932) begin
      \nz.mem_2555_sv2v_reg  <= data_i[75];
    end 
    if(N8931) begin
      \nz.mem_2554_sv2v_reg  <= data_i[74];
    end 
    if(N8930) begin
      \nz.mem_2553_sv2v_reg  <= data_i[73];
    end 
    if(N8929) begin
      \nz.mem_2552_sv2v_reg  <= data_i[72];
    end 
    if(N8928) begin
      \nz.mem_2551_sv2v_reg  <= data_i[71];
    end 
    if(N8927) begin
      \nz.mem_2550_sv2v_reg  <= data_i[70];
    end 
    if(N8926) begin
      \nz.mem_2549_sv2v_reg  <= data_i[69];
    end 
    if(N8925) begin
      \nz.mem_2548_sv2v_reg  <= data_i[68];
    end 
    if(N8924) begin
      \nz.mem_2547_sv2v_reg  <= data_i[67];
    end 
    if(N8923) begin
      \nz.mem_2546_sv2v_reg  <= data_i[66];
    end 
    if(N8922) begin
      \nz.mem_2545_sv2v_reg  <= data_i[65];
    end 
    if(N8921) begin
      \nz.mem_2544_sv2v_reg  <= data_i[64];
    end 
    if(N8920) begin
      \nz.mem_2543_sv2v_reg  <= data_i[63];
    end 
    if(N8919) begin
      \nz.mem_2542_sv2v_reg  <= data_i[62];
    end 
    if(N8918) begin
      \nz.mem_2541_sv2v_reg  <= data_i[61];
    end 
    if(N8917) begin
      \nz.mem_2540_sv2v_reg  <= data_i[60];
    end 
    if(N8916) begin
      \nz.mem_2539_sv2v_reg  <= data_i[59];
    end 
    if(N8915) begin
      \nz.mem_2538_sv2v_reg  <= data_i[58];
    end 
    if(N8914) begin
      \nz.mem_2537_sv2v_reg  <= data_i[57];
    end 
    if(N8913) begin
      \nz.mem_2536_sv2v_reg  <= data_i[56];
    end 
    if(N8912) begin
      \nz.mem_2535_sv2v_reg  <= data_i[55];
    end 
    if(N8911) begin
      \nz.mem_2534_sv2v_reg  <= data_i[54];
    end 
    if(N8910) begin
      \nz.mem_2533_sv2v_reg  <= data_i[53];
    end 
    if(N8909) begin
      \nz.mem_2532_sv2v_reg  <= data_i[52];
    end 
    if(N8908) begin
      \nz.mem_2531_sv2v_reg  <= data_i[51];
    end 
    if(N8907) begin
      \nz.mem_2530_sv2v_reg  <= data_i[50];
    end 
    if(N8906) begin
      \nz.mem_2529_sv2v_reg  <= data_i[49];
    end 
    if(N8905) begin
      \nz.mem_2528_sv2v_reg  <= data_i[48];
    end 
    if(N8904) begin
      \nz.mem_2527_sv2v_reg  <= data_i[47];
    end 
    if(N8903) begin
      \nz.mem_2526_sv2v_reg  <= data_i[46];
    end 
    if(N8902) begin
      \nz.mem_2525_sv2v_reg  <= data_i[45];
    end 
    if(N8901) begin
      \nz.mem_2524_sv2v_reg  <= data_i[44];
    end 
    if(N8900) begin
      \nz.mem_2523_sv2v_reg  <= data_i[43];
    end 
    if(N8899) begin
      \nz.mem_2522_sv2v_reg  <= data_i[42];
    end 
    if(N8898) begin
      \nz.mem_2521_sv2v_reg  <= data_i[41];
    end 
    if(N8897) begin
      \nz.mem_2520_sv2v_reg  <= data_i[40];
    end 
    if(N8896) begin
      \nz.mem_2519_sv2v_reg  <= data_i[39];
    end 
    if(N8895) begin
      \nz.mem_2518_sv2v_reg  <= data_i[38];
    end 
    if(N8894) begin
      \nz.mem_2517_sv2v_reg  <= data_i[37];
    end 
    if(N8893) begin
      \nz.mem_2516_sv2v_reg  <= data_i[36];
    end 
    if(N8892) begin
      \nz.mem_2515_sv2v_reg  <= data_i[35];
    end 
    if(N8891) begin
      \nz.mem_2514_sv2v_reg  <= data_i[34];
    end 
    if(N8890) begin
      \nz.mem_2513_sv2v_reg  <= data_i[33];
    end 
    if(N8889) begin
      \nz.mem_2512_sv2v_reg  <= data_i[32];
    end 
    if(N8888) begin
      \nz.mem_2511_sv2v_reg  <= data_i[31];
    end 
    if(N8887) begin
      \nz.mem_2510_sv2v_reg  <= data_i[30];
    end 
    if(N8886) begin
      \nz.mem_2509_sv2v_reg  <= data_i[29];
    end 
    if(N8885) begin
      \nz.mem_2508_sv2v_reg  <= data_i[28];
    end 
    if(N8884) begin
      \nz.mem_2507_sv2v_reg  <= data_i[27];
    end 
    if(N8883) begin
      \nz.mem_2506_sv2v_reg  <= data_i[26];
    end 
    if(N8882) begin
      \nz.mem_2505_sv2v_reg  <= data_i[25];
    end 
    if(N8881) begin
      \nz.mem_2504_sv2v_reg  <= data_i[24];
    end 
    if(N8880) begin
      \nz.mem_2503_sv2v_reg  <= data_i[23];
    end 
    if(N8879) begin
      \nz.mem_2502_sv2v_reg  <= data_i[22];
    end 
    if(N8878) begin
      \nz.mem_2501_sv2v_reg  <= data_i[21];
    end 
    if(N8877) begin
      \nz.mem_2500_sv2v_reg  <= data_i[20];
    end 
    if(N8876) begin
      \nz.mem_2499_sv2v_reg  <= data_i[19];
    end 
    if(N8875) begin
      \nz.mem_2498_sv2v_reg  <= data_i[18];
    end 
    if(N8874) begin
      \nz.mem_2497_sv2v_reg  <= data_i[17];
    end 
    if(N8873) begin
      \nz.mem_2496_sv2v_reg  <= data_i[16];
    end 
    if(N8872) begin
      \nz.mem_2495_sv2v_reg  <= data_i[15];
    end 
    if(N8871) begin
      \nz.mem_2494_sv2v_reg  <= data_i[14];
    end 
    if(N8870) begin
      \nz.mem_2493_sv2v_reg  <= data_i[13];
    end 
    if(N8869) begin
      \nz.mem_2492_sv2v_reg  <= data_i[12];
    end 
    if(N8868) begin
      \nz.mem_2491_sv2v_reg  <= data_i[11];
    end 
    if(N8867) begin
      \nz.mem_2490_sv2v_reg  <= data_i[10];
    end 
    if(N8866) begin
      \nz.mem_2489_sv2v_reg  <= data_i[9];
    end 
    if(N8865) begin
      \nz.mem_2488_sv2v_reg  <= data_i[8];
    end 
    if(N8864) begin
      \nz.mem_2487_sv2v_reg  <= data_i[7];
    end 
    if(N8863) begin
      \nz.mem_2486_sv2v_reg  <= data_i[6];
    end 
    if(N8862) begin
      \nz.mem_2485_sv2v_reg  <= data_i[5];
    end 
    if(N8861) begin
      \nz.mem_2484_sv2v_reg  <= data_i[4];
    end 
    if(N8860) begin
      \nz.mem_2483_sv2v_reg  <= data_i[3];
    end 
    if(N8859) begin
      \nz.mem_2482_sv2v_reg  <= data_i[2];
    end 
    if(N8858) begin
      \nz.mem_2481_sv2v_reg  <= data_i[1];
    end 
    if(N8857) begin
      \nz.mem_2480_sv2v_reg  <= data_i[0];
    end 
    if(N8856) begin
      \nz.mem_2479_sv2v_reg  <= data_i[79];
    end 
    if(N8855) begin
      \nz.mem_2478_sv2v_reg  <= data_i[78];
    end 
    if(N8854) begin
      \nz.mem_2477_sv2v_reg  <= data_i[77];
    end 
    if(N8853) begin
      \nz.mem_2476_sv2v_reg  <= data_i[76];
    end 
    if(N8852) begin
      \nz.mem_2475_sv2v_reg  <= data_i[75];
    end 
    if(N8851) begin
      \nz.mem_2474_sv2v_reg  <= data_i[74];
    end 
    if(N8850) begin
      \nz.mem_2473_sv2v_reg  <= data_i[73];
    end 
    if(N8849) begin
      \nz.mem_2472_sv2v_reg  <= data_i[72];
    end 
    if(N8848) begin
      \nz.mem_2471_sv2v_reg  <= data_i[71];
    end 
    if(N8847) begin
      \nz.mem_2470_sv2v_reg  <= data_i[70];
    end 
    if(N8846) begin
      \nz.mem_2469_sv2v_reg  <= data_i[69];
    end 
    if(N8845) begin
      \nz.mem_2468_sv2v_reg  <= data_i[68];
    end 
    if(N8844) begin
      \nz.mem_2467_sv2v_reg  <= data_i[67];
    end 
    if(N8843) begin
      \nz.mem_2466_sv2v_reg  <= data_i[66];
    end 
    if(N8842) begin
      \nz.mem_2465_sv2v_reg  <= data_i[65];
    end 
    if(N8841) begin
      \nz.mem_2464_sv2v_reg  <= data_i[64];
    end 
    if(N8840) begin
      \nz.mem_2463_sv2v_reg  <= data_i[63];
    end 
    if(N8839) begin
      \nz.mem_2462_sv2v_reg  <= data_i[62];
    end 
    if(N8838) begin
      \nz.mem_2461_sv2v_reg  <= data_i[61];
    end 
    if(N8837) begin
      \nz.mem_2460_sv2v_reg  <= data_i[60];
    end 
    if(N8836) begin
      \nz.mem_2459_sv2v_reg  <= data_i[59];
    end 
    if(N8835) begin
      \nz.mem_2458_sv2v_reg  <= data_i[58];
    end 
    if(N8834) begin
      \nz.mem_2457_sv2v_reg  <= data_i[57];
    end 
    if(N8833) begin
      \nz.mem_2456_sv2v_reg  <= data_i[56];
    end 
    if(N8832) begin
      \nz.mem_2455_sv2v_reg  <= data_i[55];
    end 
    if(N8831) begin
      \nz.mem_2454_sv2v_reg  <= data_i[54];
    end 
    if(N8830) begin
      \nz.mem_2453_sv2v_reg  <= data_i[53];
    end 
    if(N8829) begin
      \nz.mem_2452_sv2v_reg  <= data_i[52];
    end 
    if(N8828) begin
      \nz.mem_2451_sv2v_reg  <= data_i[51];
    end 
    if(N8827) begin
      \nz.mem_2450_sv2v_reg  <= data_i[50];
    end 
    if(N8826) begin
      \nz.mem_2449_sv2v_reg  <= data_i[49];
    end 
    if(N8825) begin
      \nz.mem_2448_sv2v_reg  <= data_i[48];
    end 
    if(N8824) begin
      \nz.mem_2447_sv2v_reg  <= data_i[47];
    end 
    if(N8823) begin
      \nz.mem_2446_sv2v_reg  <= data_i[46];
    end 
    if(N8822) begin
      \nz.mem_2445_sv2v_reg  <= data_i[45];
    end 
    if(N8821) begin
      \nz.mem_2444_sv2v_reg  <= data_i[44];
    end 
    if(N8820) begin
      \nz.mem_2443_sv2v_reg  <= data_i[43];
    end 
    if(N8819) begin
      \nz.mem_2442_sv2v_reg  <= data_i[42];
    end 
    if(N8818) begin
      \nz.mem_2441_sv2v_reg  <= data_i[41];
    end 
    if(N8817) begin
      \nz.mem_2440_sv2v_reg  <= data_i[40];
    end 
    if(N8816) begin
      \nz.mem_2439_sv2v_reg  <= data_i[39];
    end 
    if(N8815) begin
      \nz.mem_2438_sv2v_reg  <= data_i[38];
    end 
    if(N8814) begin
      \nz.mem_2437_sv2v_reg  <= data_i[37];
    end 
    if(N8813) begin
      \nz.mem_2436_sv2v_reg  <= data_i[36];
    end 
    if(N8812) begin
      \nz.mem_2435_sv2v_reg  <= data_i[35];
    end 
    if(N8811) begin
      \nz.mem_2434_sv2v_reg  <= data_i[34];
    end 
    if(N8810) begin
      \nz.mem_2433_sv2v_reg  <= data_i[33];
    end 
    if(N8809) begin
      \nz.mem_2432_sv2v_reg  <= data_i[32];
    end 
    if(N8808) begin
      \nz.mem_2431_sv2v_reg  <= data_i[31];
    end 
    if(N8807) begin
      \nz.mem_2430_sv2v_reg  <= data_i[30];
    end 
    if(N8806) begin
      \nz.mem_2429_sv2v_reg  <= data_i[29];
    end 
    if(N8805) begin
      \nz.mem_2428_sv2v_reg  <= data_i[28];
    end 
    if(N8804) begin
      \nz.mem_2427_sv2v_reg  <= data_i[27];
    end 
    if(N8803) begin
      \nz.mem_2426_sv2v_reg  <= data_i[26];
    end 
    if(N8802) begin
      \nz.mem_2425_sv2v_reg  <= data_i[25];
    end 
    if(N8801) begin
      \nz.mem_2424_sv2v_reg  <= data_i[24];
    end 
    if(N8800) begin
      \nz.mem_2423_sv2v_reg  <= data_i[23];
    end 
    if(N8799) begin
      \nz.mem_2422_sv2v_reg  <= data_i[22];
    end 
    if(N8798) begin
      \nz.mem_2421_sv2v_reg  <= data_i[21];
    end 
    if(N8797) begin
      \nz.mem_2420_sv2v_reg  <= data_i[20];
    end 
    if(N8796) begin
      \nz.mem_2419_sv2v_reg  <= data_i[19];
    end 
    if(N8795) begin
      \nz.mem_2418_sv2v_reg  <= data_i[18];
    end 
    if(N8794) begin
      \nz.mem_2417_sv2v_reg  <= data_i[17];
    end 
    if(N8793) begin
      \nz.mem_2416_sv2v_reg  <= data_i[16];
    end 
    if(N8792) begin
      \nz.mem_2415_sv2v_reg  <= data_i[15];
    end 
    if(N8791) begin
      \nz.mem_2414_sv2v_reg  <= data_i[14];
    end 
    if(N8790) begin
      \nz.mem_2413_sv2v_reg  <= data_i[13];
    end 
    if(N8789) begin
      \nz.mem_2412_sv2v_reg  <= data_i[12];
    end 
    if(N8788) begin
      \nz.mem_2411_sv2v_reg  <= data_i[11];
    end 
    if(N8787) begin
      \nz.mem_2410_sv2v_reg  <= data_i[10];
    end 
    if(N8786) begin
      \nz.mem_2409_sv2v_reg  <= data_i[9];
    end 
    if(N8785) begin
      \nz.mem_2408_sv2v_reg  <= data_i[8];
    end 
    if(N8784) begin
      \nz.mem_2407_sv2v_reg  <= data_i[7];
    end 
    if(N8783) begin
      \nz.mem_2406_sv2v_reg  <= data_i[6];
    end 
    if(N8782) begin
      \nz.mem_2405_sv2v_reg  <= data_i[5];
    end 
    if(N8781) begin
      \nz.mem_2404_sv2v_reg  <= data_i[4];
    end 
    if(N8780) begin
      \nz.mem_2403_sv2v_reg  <= data_i[3];
    end 
    if(N8779) begin
      \nz.mem_2402_sv2v_reg  <= data_i[2];
    end 
    if(N8778) begin
      \nz.mem_2401_sv2v_reg  <= data_i[1];
    end 
    if(N8777) begin
      \nz.mem_2400_sv2v_reg  <= data_i[0];
    end 
    if(N8776) begin
      \nz.mem_2399_sv2v_reg  <= data_i[79];
    end 
    if(N8775) begin
      \nz.mem_2398_sv2v_reg  <= data_i[78];
    end 
    if(N8774) begin
      \nz.mem_2397_sv2v_reg  <= data_i[77];
    end 
    if(N8773) begin
      \nz.mem_2396_sv2v_reg  <= data_i[76];
    end 
    if(N8772) begin
      \nz.mem_2395_sv2v_reg  <= data_i[75];
    end 
    if(N8771) begin
      \nz.mem_2394_sv2v_reg  <= data_i[74];
    end 
    if(N8770) begin
      \nz.mem_2393_sv2v_reg  <= data_i[73];
    end 
    if(N8769) begin
      \nz.mem_2392_sv2v_reg  <= data_i[72];
    end 
    if(N8768) begin
      \nz.mem_2391_sv2v_reg  <= data_i[71];
    end 
    if(N8767) begin
      \nz.mem_2390_sv2v_reg  <= data_i[70];
    end 
    if(N8766) begin
      \nz.mem_2389_sv2v_reg  <= data_i[69];
    end 
    if(N8765) begin
      \nz.mem_2388_sv2v_reg  <= data_i[68];
    end 
    if(N8764) begin
      \nz.mem_2387_sv2v_reg  <= data_i[67];
    end 
    if(N8763) begin
      \nz.mem_2386_sv2v_reg  <= data_i[66];
    end 
    if(N8762) begin
      \nz.mem_2385_sv2v_reg  <= data_i[65];
    end 
    if(N8761) begin
      \nz.mem_2384_sv2v_reg  <= data_i[64];
    end 
    if(N8760) begin
      \nz.mem_2383_sv2v_reg  <= data_i[63];
    end 
    if(N8759) begin
      \nz.mem_2382_sv2v_reg  <= data_i[62];
    end 
    if(N8758) begin
      \nz.mem_2381_sv2v_reg  <= data_i[61];
    end 
    if(N8757) begin
      \nz.mem_2380_sv2v_reg  <= data_i[60];
    end 
    if(N8756) begin
      \nz.mem_2379_sv2v_reg  <= data_i[59];
    end 
    if(N8755) begin
      \nz.mem_2378_sv2v_reg  <= data_i[58];
    end 
    if(N8754) begin
      \nz.mem_2377_sv2v_reg  <= data_i[57];
    end 
    if(N8753) begin
      \nz.mem_2376_sv2v_reg  <= data_i[56];
    end 
    if(N8752) begin
      \nz.mem_2375_sv2v_reg  <= data_i[55];
    end 
    if(N8751) begin
      \nz.mem_2374_sv2v_reg  <= data_i[54];
    end 
    if(N8750) begin
      \nz.mem_2373_sv2v_reg  <= data_i[53];
    end 
    if(N8749) begin
      \nz.mem_2372_sv2v_reg  <= data_i[52];
    end 
    if(N8748) begin
      \nz.mem_2371_sv2v_reg  <= data_i[51];
    end 
    if(N8747) begin
      \nz.mem_2370_sv2v_reg  <= data_i[50];
    end 
    if(N8746) begin
      \nz.mem_2369_sv2v_reg  <= data_i[49];
    end 
    if(N8745) begin
      \nz.mem_2368_sv2v_reg  <= data_i[48];
    end 
    if(N8744) begin
      \nz.mem_2367_sv2v_reg  <= data_i[47];
    end 
    if(N8743) begin
      \nz.mem_2366_sv2v_reg  <= data_i[46];
    end 
    if(N8742) begin
      \nz.mem_2365_sv2v_reg  <= data_i[45];
    end 
    if(N8741) begin
      \nz.mem_2364_sv2v_reg  <= data_i[44];
    end 
    if(N8740) begin
      \nz.mem_2363_sv2v_reg  <= data_i[43];
    end 
    if(N8739) begin
      \nz.mem_2362_sv2v_reg  <= data_i[42];
    end 
    if(N8738) begin
      \nz.mem_2361_sv2v_reg  <= data_i[41];
    end 
    if(N8737) begin
      \nz.mem_2360_sv2v_reg  <= data_i[40];
    end 
    if(N8736) begin
      \nz.mem_2359_sv2v_reg  <= data_i[39];
    end 
    if(N8735) begin
      \nz.mem_2358_sv2v_reg  <= data_i[38];
    end 
    if(N8734) begin
      \nz.mem_2357_sv2v_reg  <= data_i[37];
    end 
    if(N8733) begin
      \nz.mem_2356_sv2v_reg  <= data_i[36];
    end 
    if(N8732) begin
      \nz.mem_2355_sv2v_reg  <= data_i[35];
    end 
    if(N8731) begin
      \nz.mem_2354_sv2v_reg  <= data_i[34];
    end 
    if(N8730) begin
      \nz.mem_2353_sv2v_reg  <= data_i[33];
    end 
    if(N8729) begin
      \nz.mem_2352_sv2v_reg  <= data_i[32];
    end 
    if(N8728) begin
      \nz.mem_2351_sv2v_reg  <= data_i[31];
    end 
    if(N8727) begin
      \nz.mem_2350_sv2v_reg  <= data_i[30];
    end 
    if(N8726) begin
      \nz.mem_2349_sv2v_reg  <= data_i[29];
    end 
    if(N8725) begin
      \nz.mem_2348_sv2v_reg  <= data_i[28];
    end 
    if(N8724) begin
      \nz.mem_2347_sv2v_reg  <= data_i[27];
    end 
    if(N8723) begin
      \nz.mem_2346_sv2v_reg  <= data_i[26];
    end 
    if(N8722) begin
      \nz.mem_2345_sv2v_reg  <= data_i[25];
    end 
    if(N8721) begin
      \nz.mem_2344_sv2v_reg  <= data_i[24];
    end 
    if(N8720) begin
      \nz.mem_2343_sv2v_reg  <= data_i[23];
    end 
    if(N8719) begin
      \nz.mem_2342_sv2v_reg  <= data_i[22];
    end 
    if(N8718) begin
      \nz.mem_2341_sv2v_reg  <= data_i[21];
    end 
    if(N8717) begin
      \nz.mem_2340_sv2v_reg  <= data_i[20];
    end 
    if(N8716) begin
      \nz.mem_2339_sv2v_reg  <= data_i[19];
    end 
    if(N8715) begin
      \nz.mem_2338_sv2v_reg  <= data_i[18];
    end 
    if(N8714) begin
      \nz.mem_2337_sv2v_reg  <= data_i[17];
    end 
    if(N8713) begin
      \nz.mem_2336_sv2v_reg  <= data_i[16];
    end 
    if(N8712) begin
      \nz.mem_2335_sv2v_reg  <= data_i[15];
    end 
    if(N8711) begin
      \nz.mem_2334_sv2v_reg  <= data_i[14];
    end 
    if(N8710) begin
      \nz.mem_2333_sv2v_reg  <= data_i[13];
    end 
    if(N8709) begin
      \nz.mem_2332_sv2v_reg  <= data_i[12];
    end 
    if(N8708) begin
      \nz.mem_2331_sv2v_reg  <= data_i[11];
    end 
    if(N8707) begin
      \nz.mem_2330_sv2v_reg  <= data_i[10];
    end 
    if(N8706) begin
      \nz.mem_2329_sv2v_reg  <= data_i[9];
    end 
    if(N8705) begin
      \nz.mem_2328_sv2v_reg  <= data_i[8];
    end 
    if(N8704) begin
      \nz.mem_2327_sv2v_reg  <= data_i[7];
    end 
    if(N8703) begin
      \nz.mem_2326_sv2v_reg  <= data_i[6];
    end 
    if(N8702) begin
      \nz.mem_2325_sv2v_reg  <= data_i[5];
    end 
    if(N8701) begin
      \nz.mem_2324_sv2v_reg  <= data_i[4];
    end 
    if(N8700) begin
      \nz.mem_2323_sv2v_reg  <= data_i[3];
    end 
    if(N8699) begin
      \nz.mem_2322_sv2v_reg  <= data_i[2];
    end 
    if(N8698) begin
      \nz.mem_2321_sv2v_reg  <= data_i[1];
    end 
    if(N8697) begin
      \nz.mem_2320_sv2v_reg  <= data_i[0];
    end 
    if(N8696) begin
      \nz.mem_2319_sv2v_reg  <= data_i[79];
    end 
    if(N8695) begin
      \nz.mem_2318_sv2v_reg  <= data_i[78];
    end 
    if(N8694) begin
      \nz.mem_2317_sv2v_reg  <= data_i[77];
    end 
    if(N8693) begin
      \nz.mem_2316_sv2v_reg  <= data_i[76];
    end 
    if(N8692) begin
      \nz.mem_2315_sv2v_reg  <= data_i[75];
    end 
    if(N8691) begin
      \nz.mem_2314_sv2v_reg  <= data_i[74];
    end 
    if(N8690) begin
      \nz.mem_2313_sv2v_reg  <= data_i[73];
    end 
    if(N8689) begin
      \nz.mem_2312_sv2v_reg  <= data_i[72];
    end 
    if(N8688) begin
      \nz.mem_2311_sv2v_reg  <= data_i[71];
    end 
    if(N8687) begin
      \nz.mem_2310_sv2v_reg  <= data_i[70];
    end 
    if(N8686) begin
      \nz.mem_2309_sv2v_reg  <= data_i[69];
    end 
    if(N8685) begin
      \nz.mem_2308_sv2v_reg  <= data_i[68];
    end 
    if(N8684) begin
      \nz.mem_2307_sv2v_reg  <= data_i[67];
    end 
    if(N8683) begin
      \nz.mem_2306_sv2v_reg  <= data_i[66];
    end 
    if(N8682) begin
      \nz.mem_2305_sv2v_reg  <= data_i[65];
    end 
    if(N8681) begin
      \nz.mem_2304_sv2v_reg  <= data_i[64];
    end 
    if(N8680) begin
      \nz.mem_2303_sv2v_reg  <= data_i[63];
    end 
    if(N8679) begin
      \nz.mem_2302_sv2v_reg  <= data_i[62];
    end 
    if(N8678) begin
      \nz.mem_2301_sv2v_reg  <= data_i[61];
    end 
    if(N8677) begin
      \nz.mem_2300_sv2v_reg  <= data_i[60];
    end 
    if(N8676) begin
      \nz.mem_2299_sv2v_reg  <= data_i[59];
    end 
    if(N8675) begin
      \nz.mem_2298_sv2v_reg  <= data_i[58];
    end 
    if(N8674) begin
      \nz.mem_2297_sv2v_reg  <= data_i[57];
    end 
    if(N8673) begin
      \nz.mem_2296_sv2v_reg  <= data_i[56];
    end 
    if(N8672) begin
      \nz.mem_2295_sv2v_reg  <= data_i[55];
    end 
    if(N8671) begin
      \nz.mem_2294_sv2v_reg  <= data_i[54];
    end 
    if(N8670) begin
      \nz.mem_2293_sv2v_reg  <= data_i[53];
    end 
    if(N8669) begin
      \nz.mem_2292_sv2v_reg  <= data_i[52];
    end 
    if(N8668) begin
      \nz.mem_2291_sv2v_reg  <= data_i[51];
    end 
    if(N8667) begin
      \nz.mem_2290_sv2v_reg  <= data_i[50];
    end 
    if(N8666) begin
      \nz.mem_2289_sv2v_reg  <= data_i[49];
    end 
    if(N8665) begin
      \nz.mem_2288_sv2v_reg  <= data_i[48];
    end 
    if(N8664) begin
      \nz.mem_2287_sv2v_reg  <= data_i[47];
    end 
    if(N8663) begin
      \nz.mem_2286_sv2v_reg  <= data_i[46];
    end 
    if(N8662) begin
      \nz.mem_2285_sv2v_reg  <= data_i[45];
    end 
    if(N8661) begin
      \nz.mem_2284_sv2v_reg  <= data_i[44];
    end 
    if(N8660) begin
      \nz.mem_2283_sv2v_reg  <= data_i[43];
    end 
    if(N8659) begin
      \nz.mem_2282_sv2v_reg  <= data_i[42];
    end 
    if(N8658) begin
      \nz.mem_2281_sv2v_reg  <= data_i[41];
    end 
    if(N8657) begin
      \nz.mem_2280_sv2v_reg  <= data_i[40];
    end 
    if(N8656) begin
      \nz.mem_2279_sv2v_reg  <= data_i[39];
    end 
    if(N8655) begin
      \nz.mem_2278_sv2v_reg  <= data_i[38];
    end 
    if(N8654) begin
      \nz.mem_2277_sv2v_reg  <= data_i[37];
    end 
    if(N8653) begin
      \nz.mem_2276_sv2v_reg  <= data_i[36];
    end 
    if(N8652) begin
      \nz.mem_2275_sv2v_reg  <= data_i[35];
    end 
    if(N8651) begin
      \nz.mem_2274_sv2v_reg  <= data_i[34];
    end 
    if(N8650) begin
      \nz.mem_2273_sv2v_reg  <= data_i[33];
    end 
    if(N8649) begin
      \nz.mem_2272_sv2v_reg  <= data_i[32];
    end 
    if(N8648) begin
      \nz.mem_2271_sv2v_reg  <= data_i[31];
    end 
    if(N8647) begin
      \nz.mem_2270_sv2v_reg  <= data_i[30];
    end 
    if(N8646) begin
      \nz.mem_2269_sv2v_reg  <= data_i[29];
    end 
    if(N8645) begin
      \nz.mem_2268_sv2v_reg  <= data_i[28];
    end 
    if(N8644) begin
      \nz.mem_2267_sv2v_reg  <= data_i[27];
    end 
    if(N8643) begin
      \nz.mem_2266_sv2v_reg  <= data_i[26];
    end 
    if(N8642) begin
      \nz.mem_2265_sv2v_reg  <= data_i[25];
    end 
    if(N8641) begin
      \nz.mem_2264_sv2v_reg  <= data_i[24];
    end 
    if(N8640) begin
      \nz.mem_2263_sv2v_reg  <= data_i[23];
    end 
    if(N8639) begin
      \nz.mem_2262_sv2v_reg  <= data_i[22];
    end 
    if(N8638) begin
      \nz.mem_2261_sv2v_reg  <= data_i[21];
    end 
    if(N8637) begin
      \nz.mem_2260_sv2v_reg  <= data_i[20];
    end 
    if(N8636) begin
      \nz.mem_2259_sv2v_reg  <= data_i[19];
    end 
    if(N8635) begin
      \nz.mem_2258_sv2v_reg  <= data_i[18];
    end 
    if(N8634) begin
      \nz.mem_2257_sv2v_reg  <= data_i[17];
    end 
    if(N8633) begin
      \nz.mem_2256_sv2v_reg  <= data_i[16];
    end 
    if(N8632) begin
      \nz.mem_2255_sv2v_reg  <= data_i[15];
    end 
    if(N8631) begin
      \nz.mem_2254_sv2v_reg  <= data_i[14];
    end 
    if(N8630) begin
      \nz.mem_2253_sv2v_reg  <= data_i[13];
    end 
    if(N8629) begin
      \nz.mem_2252_sv2v_reg  <= data_i[12];
    end 
    if(N8628) begin
      \nz.mem_2251_sv2v_reg  <= data_i[11];
    end 
    if(N8627) begin
      \nz.mem_2250_sv2v_reg  <= data_i[10];
    end 
    if(N8626) begin
      \nz.mem_2249_sv2v_reg  <= data_i[9];
    end 
    if(N8625) begin
      \nz.mem_2248_sv2v_reg  <= data_i[8];
    end 
    if(N8624) begin
      \nz.mem_2247_sv2v_reg  <= data_i[7];
    end 
    if(N8623) begin
      \nz.mem_2246_sv2v_reg  <= data_i[6];
    end 
    if(N8622) begin
      \nz.mem_2245_sv2v_reg  <= data_i[5];
    end 
    if(N8621) begin
      \nz.mem_2244_sv2v_reg  <= data_i[4];
    end 
    if(N8620) begin
      \nz.mem_2243_sv2v_reg  <= data_i[3];
    end 
    if(N8619) begin
      \nz.mem_2242_sv2v_reg  <= data_i[2];
    end 
    if(N8618) begin
      \nz.mem_2241_sv2v_reg  <= data_i[1];
    end 
    if(N8617) begin
      \nz.mem_2240_sv2v_reg  <= data_i[0];
    end 
    if(N8616) begin
      \nz.mem_2239_sv2v_reg  <= data_i[79];
    end 
    if(N8615) begin
      \nz.mem_2238_sv2v_reg  <= data_i[78];
    end 
    if(N8614) begin
      \nz.mem_2237_sv2v_reg  <= data_i[77];
    end 
    if(N8613) begin
      \nz.mem_2236_sv2v_reg  <= data_i[76];
    end 
    if(N8612) begin
      \nz.mem_2235_sv2v_reg  <= data_i[75];
    end 
    if(N8611) begin
      \nz.mem_2234_sv2v_reg  <= data_i[74];
    end 
    if(N8610) begin
      \nz.mem_2233_sv2v_reg  <= data_i[73];
    end 
    if(N8609) begin
      \nz.mem_2232_sv2v_reg  <= data_i[72];
    end 
    if(N8608) begin
      \nz.mem_2231_sv2v_reg  <= data_i[71];
    end 
    if(N8607) begin
      \nz.mem_2230_sv2v_reg  <= data_i[70];
    end 
    if(N8606) begin
      \nz.mem_2229_sv2v_reg  <= data_i[69];
    end 
    if(N8605) begin
      \nz.mem_2228_sv2v_reg  <= data_i[68];
    end 
    if(N8604) begin
      \nz.mem_2227_sv2v_reg  <= data_i[67];
    end 
    if(N8603) begin
      \nz.mem_2226_sv2v_reg  <= data_i[66];
    end 
    if(N8602) begin
      \nz.mem_2225_sv2v_reg  <= data_i[65];
    end 
    if(N8601) begin
      \nz.mem_2224_sv2v_reg  <= data_i[64];
    end 
    if(N8600) begin
      \nz.mem_2223_sv2v_reg  <= data_i[63];
    end 
    if(N8599) begin
      \nz.mem_2222_sv2v_reg  <= data_i[62];
    end 
    if(N8598) begin
      \nz.mem_2221_sv2v_reg  <= data_i[61];
    end 
    if(N8597) begin
      \nz.mem_2220_sv2v_reg  <= data_i[60];
    end 
    if(N8596) begin
      \nz.mem_2219_sv2v_reg  <= data_i[59];
    end 
    if(N8595) begin
      \nz.mem_2218_sv2v_reg  <= data_i[58];
    end 
    if(N8594) begin
      \nz.mem_2217_sv2v_reg  <= data_i[57];
    end 
    if(N8593) begin
      \nz.mem_2216_sv2v_reg  <= data_i[56];
    end 
    if(N8592) begin
      \nz.mem_2215_sv2v_reg  <= data_i[55];
    end 
    if(N8591) begin
      \nz.mem_2214_sv2v_reg  <= data_i[54];
    end 
    if(N8590) begin
      \nz.mem_2213_sv2v_reg  <= data_i[53];
    end 
    if(N8589) begin
      \nz.mem_2212_sv2v_reg  <= data_i[52];
    end 
    if(N8588) begin
      \nz.mem_2211_sv2v_reg  <= data_i[51];
    end 
    if(N8587) begin
      \nz.mem_2210_sv2v_reg  <= data_i[50];
    end 
    if(N8586) begin
      \nz.mem_2209_sv2v_reg  <= data_i[49];
    end 
    if(N8585) begin
      \nz.mem_2208_sv2v_reg  <= data_i[48];
    end 
    if(N8584) begin
      \nz.mem_2207_sv2v_reg  <= data_i[47];
    end 
    if(N8583) begin
      \nz.mem_2206_sv2v_reg  <= data_i[46];
    end 
    if(N8582) begin
      \nz.mem_2205_sv2v_reg  <= data_i[45];
    end 
    if(N8581) begin
      \nz.mem_2204_sv2v_reg  <= data_i[44];
    end 
    if(N8580) begin
      \nz.mem_2203_sv2v_reg  <= data_i[43];
    end 
    if(N8579) begin
      \nz.mem_2202_sv2v_reg  <= data_i[42];
    end 
    if(N8578) begin
      \nz.mem_2201_sv2v_reg  <= data_i[41];
    end 
    if(N8577) begin
      \nz.mem_2200_sv2v_reg  <= data_i[40];
    end 
    if(N8576) begin
      \nz.mem_2199_sv2v_reg  <= data_i[39];
    end 
    if(N8575) begin
      \nz.mem_2198_sv2v_reg  <= data_i[38];
    end 
    if(N8574) begin
      \nz.mem_2197_sv2v_reg  <= data_i[37];
    end 
    if(N8573) begin
      \nz.mem_2196_sv2v_reg  <= data_i[36];
    end 
    if(N8572) begin
      \nz.mem_2195_sv2v_reg  <= data_i[35];
    end 
    if(N8571) begin
      \nz.mem_2194_sv2v_reg  <= data_i[34];
    end 
    if(N8570) begin
      \nz.mem_2193_sv2v_reg  <= data_i[33];
    end 
    if(N8569) begin
      \nz.mem_2192_sv2v_reg  <= data_i[32];
    end 
    if(N8568) begin
      \nz.mem_2191_sv2v_reg  <= data_i[31];
    end 
    if(N8567) begin
      \nz.mem_2190_sv2v_reg  <= data_i[30];
    end 
    if(N8566) begin
      \nz.mem_2189_sv2v_reg  <= data_i[29];
    end 
    if(N8565) begin
      \nz.mem_2188_sv2v_reg  <= data_i[28];
    end 
    if(N8564) begin
      \nz.mem_2187_sv2v_reg  <= data_i[27];
    end 
    if(N8563) begin
      \nz.mem_2186_sv2v_reg  <= data_i[26];
    end 
    if(N8562) begin
      \nz.mem_2185_sv2v_reg  <= data_i[25];
    end 
    if(N8561) begin
      \nz.mem_2184_sv2v_reg  <= data_i[24];
    end 
    if(N8560) begin
      \nz.mem_2183_sv2v_reg  <= data_i[23];
    end 
    if(N8559) begin
      \nz.mem_2182_sv2v_reg  <= data_i[22];
    end 
    if(N8558) begin
      \nz.mem_2181_sv2v_reg  <= data_i[21];
    end 
    if(N8557) begin
      \nz.mem_2180_sv2v_reg  <= data_i[20];
    end 
    if(N8556) begin
      \nz.mem_2179_sv2v_reg  <= data_i[19];
    end 
    if(N8555) begin
      \nz.mem_2178_sv2v_reg  <= data_i[18];
    end 
    if(N8554) begin
      \nz.mem_2177_sv2v_reg  <= data_i[17];
    end 
    if(N8553) begin
      \nz.mem_2176_sv2v_reg  <= data_i[16];
    end 
    if(N8552) begin
      \nz.mem_2175_sv2v_reg  <= data_i[15];
    end 
    if(N8551) begin
      \nz.mem_2174_sv2v_reg  <= data_i[14];
    end 
    if(N8550) begin
      \nz.mem_2173_sv2v_reg  <= data_i[13];
    end 
    if(N8549) begin
      \nz.mem_2172_sv2v_reg  <= data_i[12];
    end 
    if(N8548) begin
      \nz.mem_2171_sv2v_reg  <= data_i[11];
    end 
    if(N8547) begin
      \nz.mem_2170_sv2v_reg  <= data_i[10];
    end 
    if(N8546) begin
      \nz.mem_2169_sv2v_reg  <= data_i[9];
    end 
    if(N8545) begin
      \nz.mem_2168_sv2v_reg  <= data_i[8];
    end 
    if(N8544) begin
      \nz.mem_2167_sv2v_reg  <= data_i[7];
    end 
    if(N8543) begin
      \nz.mem_2166_sv2v_reg  <= data_i[6];
    end 
    if(N8542) begin
      \nz.mem_2165_sv2v_reg  <= data_i[5];
    end 
    if(N8541) begin
      \nz.mem_2164_sv2v_reg  <= data_i[4];
    end 
    if(N8540) begin
      \nz.mem_2163_sv2v_reg  <= data_i[3];
    end 
    if(N8539) begin
      \nz.mem_2162_sv2v_reg  <= data_i[2];
    end 
    if(N8538) begin
      \nz.mem_2161_sv2v_reg  <= data_i[1];
    end 
    if(N8537) begin
      \nz.mem_2160_sv2v_reg  <= data_i[0];
    end 
    if(N8536) begin
      \nz.mem_2159_sv2v_reg  <= data_i[79];
    end 
    if(N8535) begin
      \nz.mem_2158_sv2v_reg  <= data_i[78];
    end 
    if(N8534) begin
      \nz.mem_2157_sv2v_reg  <= data_i[77];
    end 
    if(N8533) begin
      \nz.mem_2156_sv2v_reg  <= data_i[76];
    end 
    if(N8532) begin
      \nz.mem_2155_sv2v_reg  <= data_i[75];
    end 
    if(N8531) begin
      \nz.mem_2154_sv2v_reg  <= data_i[74];
    end 
    if(N8530) begin
      \nz.mem_2153_sv2v_reg  <= data_i[73];
    end 
    if(N8529) begin
      \nz.mem_2152_sv2v_reg  <= data_i[72];
    end 
    if(N8528) begin
      \nz.mem_2151_sv2v_reg  <= data_i[71];
    end 
    if(N8527) begin
      \nz.mem_2150_sv2v_reg  <= data_i[70];
    end 
    if(N8526) begin
      \nz.mem_2149_sv2v_reg  <= data_i[69];
    end 
    if(N8525) begin
      \nz.mem_2148_sv2v_reg  <= data_i[68];
    end 
    if(N8524) begin
      \nz.mem_2147_sv2v_reg  <= data_i[67];
    end 
    if(N8523) begin
      \nz.mem_2146_sv2v_reg  <= data_i[66];
    end 
    if(N8522) begin
      \nz.mem_2145_sv2v_reg  <= data_i[65];
    end 
    if(N8521) begin
      \nz.mem_2144_sv2v_reg  <= data_i[64];
    end 
    if(N8520) begin
      \nz.mem_2143_sv2v_reg  <= data_i[63];
    end 
    if(N8519) begin
      \nz.mem_2142_sv2v_reg  <= data_i[62];
    end 
    if(N8518) begin
      \nz.mem_2141_sv2v_reg  <= data_i[61];
    end 
    if(N8517) begin
      \nz.mem_2140_sv2v_reg  <= data_i[60];
    end 
    if(N8516) begin
      \nz.mem_2139_sv2v_reg  <= data_i[59];
    end 
    if(N8515) begin
      \nz.mem_2138_sv2v_reg  <= data_i[58];
    end 
    if(N8514) begin
      \nz.mem_2137_sv2v_reg  <= data_i[57];
    end 
    if(N8513) begin
      \nz.mem_2136_sv2v_reg  <= data_i[56];
    end 
    if(N8512) begin
      \nz.mem_2135_sv2v_reg  <= data_i[55];
    end 
    if(N8511) begin
      \nz.mem_2134_sv2v_reg  <= data_i[54];
    end 
    if(N8510) begin
      \nz.mem_2133_sv2v_reg  <= data_i[53];
    end 
    if(N8509) begin
      \nz.mem_2132_sv2v_reg  <= data_i[52];
    end 
    if(N8508) begin
      \nz.mem_2131_sv2v_reg  <= data_i[51];
    end 
    if(N8507) begin
      \nz.mem_2130_sv2v_reg  <= data_i[50];
    end 
    if(N8506) begin
      \nz.mem_2129_sv2v_reg  <= data_i[49];
    end 
    if(N8505) begin
      \nz.mem_2128_sv2v_reg  <= data_i[48];
    end 
    if(N8504) begin
      \nz.mem_2127_sv2v_reg  <= data_i[47];
    end 
    if(N8503) begin
      \nz.mem_2126_sv2v_reg  <= data_i[46];
    end 
    if(N8502) begin
      \nz.mem_2125_sv2v_reg  <= data_i[45];
    end 
    if(N8501) begin
      \nz.mem_2124_sv2v_reg  <= data_i[44];
    end 
    if(N8500) begin
      \nz.mem_2123_sv2v_reg  <= data_i[43];
    end 
    if(N8499) begin
      \nz.mem_2122_sv2v_reg  <= data_i[42];
    end 
    if(N8498) begin
      \nz.mem_2121_sv2v_reg  <= data_i[41];
    end 
    if(N8497) begin
      \nz.mem_2120_sv2v_reg  <= data_i[40];
    end 
    if(N8496) begin
      \nz.mem_2119_sv2v_reg  <= data_i[39];
    end 
    if(N8495) begin
      \nz.mem_2118_sv2v_reg  <= data_i[38];
    end 
    if(N8494) begin
      \nz.mem_2117_sv2v_reg  <= data_i[37];
    end 
    if(N8493) begin
      \nz.mem_2116_sv2v_reg  <= data_i[36];
    end 
    if(N8492) begin
      \nz.mem_2115_sv2v_reg  <= data_i[35];
    end 
    if(N8491) begin
      \nz.mem_2114_sv2v_reg  <= data_i[34];
    end 
    if(N8490) begin
      \nz.mem_2113_sv2v_reg  <= data_i[33];
    end 
    if(N8489) begin
      \nz.mem_2112_sv2v_reg  <= data_i[32];
    end 
    if(N8488) begin
      \nz.mem_2111_sv2v_reg  <= data_i[31];
    end 
    if(N8487) begin
      \nz.mem_2110_sv2v_reg  <= data_i[30];
    end 
    if(N8486) begin
      \nz.mem_2109_sv2v_reg  <= data_i[29];
    end 
    if(N8485) begin
      \nz.mem_2108_sv2v_reg  <= data_i[28];
    end 
    if(N8484) begin
      \nz.mem_2107_sv2v_reg  <= data_i[27];
    end 
    if(N8483) begin
      \nz.mem_2106_sv2v_reg  <= data_i[26];
    end 
    if(N8482) begin
      \nz.mem_2105_sv2v_reg  <= data_i[25];
    end 
    if(N8481) begin
      \nz.mem_2104_sv2v_reg  <= data_i[24];
    end 
    if(N8480) begin
      \nz.mem_2103_sv2v_reg  <= data_i[23];
    end 
    if(N8479) begin
      \nz.mem_2102_sv2v_reg  <= data_i[22];
    end 
    if(N8478) begin
      \nz.mem_2101_sv2v_reg  <= data_i[21];
    end 
    if(N8477) begin
      \nz.mem_2100_sv2v_reg  <= data_i[20];
    end 
    if(N8476) begin
      \nz.mem_2099_sv2v_reg  <= data_i[19];
    end 
    if(N8475) begin
      \nz.mem_2098_sv2v_reg  <= data_i[18];
    end 
    if(N8474) begin
      \nz.mem_2097_sv2v_reg  <= data_i[17];
    end 
    if(N8473) begin
      \nz.mem_2096_sv2v_reg  <= data_i[16];
    end 
    if(N8472) begin
      \nz.mem_2095_sv2v_reg  <= data_i[15];
    end 
    if(N8471) begin
      \nz.mem_2094_sv2v_reg  <= data_i[14];
    end 
    if(N8470) begin
      \nz.mem_2093_sv2v_reg  <= data_i[13];
    end 
    if(N8469) begin
      \nz.mem_2092_sv2v_reg  <= data_i[12];
    end 
    if(N8468) begin
      \nz.mem_2091_sv2v_reg  <= data_i[11];
    end 
    if(N8467) begin
      \nz.mem_2090_sv2v_reg  <= data_i[10];
    end 
    if(N8466) begin
      \nz.mem_2089_sv2v_reg  <= data_i[9];
    end 
    if(N8465) begin
      \nz.mem_2088_sv2v_reg  <= data_i[8];
    end 
    if(N8464) begin
      \nz.mem_2087_sv2v_reg  <= data_i[7];
    end 
    if(N8463) begin
      \nz.mem_2086_sv2v_reg  <= data_i[6];
    end 
    if(N8462) begin
      \nz.mem_2085_sv2v_reg  <= data_i[5];
    end 
    if(N8461) begin
      \nz.mem_2084_sv2v_reg  <= data_i[4];
    end 
    if(N8460) begin
      \nz.mem_2083_sv2v_reg  <= data_i[3];
    end 
    if(N8459) begin
      \nz.mem_2082_sv2v_reg  <= data_i[2];
    end 
    if(N8458) begin
      \nz.mem_2081_sv2v_reg  <= data_i[1];
    end 
    if(N8457) begin
      \nz.mem_2080_sv2v_reg  <= data_i[0];
    end 
    if(N8456) begin
      \nz.mem_2079_sv2v_reg  <= data_i[79];
    end 
    if(N8455) begin
      \nz.mem_2078_sv2v_reg  <= data_i[78];
    end 
    if(N8454) begin
      \nz.mem_2077_sv2v_reg  <= data_i[77];
    end 
    if(N8453) begin
      \nz.mem_2076_sv2v_reg  <= data_i[76];
    end 
    if(N8452) begin
      \nz.mem_2075_sv2v_reg  <= data_i[75];
    end 
    if(N8451) begin
      \nz.mem_2074_sv2v_reg  <= data_i[74];
    end 
    if(N8450) begin
      \nz.mem_2073_sv2v_reg  <= data_i[73];
    end 
    if(N8449) begin
      \nz.mem_2072_sv2v_reg  <= data_i[72];
    end 
    if(N8448) begin
      \nz.mem_2071_sv2v_reg  <= data_i[71];
    end 
    if(N8447) begin
      \nz.mem_2070_sv2v_reg  <= data_i[70];
    end 
    if(N8446) begin
      \nz.mem_2069_sv2v_reg  <= data_i[69];
    end 
    if(N8445) begin
      \nz.mem_2068_sv2v_reg  <= data_i[68];
    end 
    if(N8444) begin
      \nz.mem_2067_sv2v_reg  <= data_i[67];
    end 
    if(N8443) begin
      \nz.mem_2066_sv2v_reg  <= data_i[66];
    end 
    if(N8442) begin
      \nz.mem_2065_sv2v_reg  <= data_i[65];
    end 
    if(N8441) begin
      \nz.mem_2064_sv2v_reg  <= data_i[64];
    end 
    if(N8440) begin
      \nz.mem_2063_sv2v_reg  <= data_i[63];
    end 
    if(N8439) begin
      \nz.mem_2062_sv2v_reg  <= data_i[62];
    end 
    if(N8438) begin
      \nz.mem_2061_sv2v_reg  <= data_i[61];
    end 
    if(N8437) begin
      \nz.mem_2060_sv2v_reg  <= data_i[60];
    end 
    if(N8436) begin
      \nz.mem_2059_sv2v_reg  <= data_i[59];
    end 
    if(N8435) begin
      \nz.mem_2058_sv2v_reg  <= data_i[58];
    end 
    if(N8434) begin
      \nz.mem_2057_sv2v_reg  <= data_i[57];
    end 
    if(N8433) begin
      \nz.mem_2056_sv2v_reg  <= data_i[56];
    end 
    if(N8432) begin
      \nz.mem_2055_sv2v_reg  <= data_i[55];
    end 
    if(N8431) begin
      \nz.mem_2054_sv2v_reg  <= data_i[54];
    end 
    if(N8430) begin
      \nz.mem_2053_sv2v_reg  <= data_i[53];
    end 
    if(N8429) begin
      \nz.mem_2052_sv2v_reg  <= data_i[52];
    end 
    if(N8428) begin
      \nz.mem_2051_sv2v_reg  <= data_i[51];
    end 
    if(N8427) begin
      \nz.mem_2050_sv2v_reg  <= data_i[50];
    end 
    if(N8426) begin
      \nz.mem_2049_sv2v_reg  <= data_i[49];
    end 
    if(N8425) begin
      \nz.mem_2048_sv2v_reg  <= data_i[48];
    end 
    if(N8424) begin
      \nz.mem_2047_sv2v_reg  <= data_i[47];
    end 
    if(N8423) begin
      \nz.mem_2046_sv2v_reg  <= data_i[46];
    end 
    if(N8422) begin
      \nz.mem_2045_sv2v_reg  <= data_i[45];
    end 
    if(N8421) begin
      \nz.mem_2044_sv2v_reg  <= data_i[44];
    end 
    if(N8420) begin
      \nz.mem_2043_sv2v_reg  <= data_i[43];
    end 
    if(N8419) begin
      \nz.mem_2042_sv2v_reg  <= data_i[42];
    end 
    if(N8418) begin
      \nz.mem_2041_sv2v_reg  <= data_i[41];
    end 
    if(N8417) begin
      \nz.mem_2040_sv2v_reg  <= data_i[40];
    end 
    if(N8416) begin
      \nz.mem_2039_sv2v_reg  <= data_i[39];
    end 
    if(N8415) begin
      \nz.mem_2038_sv2v_reg  <= data_i[38];
    end 
    if(N8414) begin
      \nz.mem_2037_sv2v_reg  <= data_i[37];
    end 
    if(N8413) begin
      \nz.mem_2036_sv2v_reg  <= data_i[36];
    end 
    if(N8412) begin
      \nz.mem_2035_sv2v_reg  <= data_i[35];
    end 
    if(N8411) begin
      \nz.mem_2034_sv2v_reg  <= data_i[34];
    end 
    if(N8410) begin
      \nz.mem_2033_sv2v_reg  <= data_i[33];
    end 
    if(N8409) begin
      \nz.mem_2032_sv2v_reg  <= data_i[32];
    end 
    if(N8408) begin
      \nz.mem_2031_sv2v_reg  <= data_i[31];
    end 
    if(N8407) begin
      \nz.mem_2030_sv2v_reg  <= data_i[30];
    end 
    if(N8406) begin
      \nz.mem_2029_sv2v_reg  <= data_i[29];
    end 
    if(N8405) begin
      \nz.mem_2028_sv2v_reg  <= data_i[28];
    end 
    if(N8404) begin
      \nz.mem_2027_sv2v_reg  <= data_i[27];
    end 
    if(N8403) begin
      \nz.mem_2026_sv2v_reg  <= data_i[26];
    end 
    if(N8402) begin
      \nz.mem_2025_sv2v_reg  <= data_i[25];
    end 
    if(N8401) begin
      \nz.mem_2024_sv2v_reg  <= data_i[24];
    end 
    if(N8400) begin
      \nz.mem_2023_sv2v_reg  <= data_i[23];
    end 
    if(N8399) begin
      \nz.mem_2022_sv2v_reg  <= data_i[22];
    end 
    if(N8398) begin
      \nz.mem_2021_sv2v_reg  <= data_i[21];
    end 
    if(N8397) begin
      \nz.mem_2020_sv2v_reg  <= data_i[20];
    end 
    if(N8396) begin
      \nz.mem_2019_sv2v_reg  <= data_i[19];
    end 
    if(N8395) begin
      \nz.mem_2018_sv2v_reg  <= data_i[18];
    end 
    if(N8394) begin
      \nz.mem_2017_sv2v_reg  <= data_i[17];
    end 
    if(N8393) begin
      \nz.mem_2016_sv2v_reg  <= data_i[16];
    end 
    if(N8392) begin
      \nz.mem_2015_sv2v_reg  <= data_i[15];
    end 
    if(N8391) begin
      \nz.mem_2014_sv2v_reg  <= data_i[14];
    end 
    if(N8390) begin
      \nz.mem_2013_sv2v_reg  <= data_i[13];
    end 
    if(N8389) begin
      \nz.mem_2012_sv2v_reg  <= data_i[12];
    end 
    if(N8388) begin
      \nz.mem_2011_sv2v_reg  <= data_i[11];
    end 
    if(N8387) begin
      \nz.mem_2010_sv2v_reg  <= data_i[10];
    end 
    if(N8386) begin
      \nz.mem_2009_sv2v_reg  <= data_i[9];
    end 
    if(N8385) begin
      \nz.mem_2008_sv2v_reg  <= data_i[8];
    end 
    if(N8384) begin
      \nz.mem_2007_sv2v_reg  <= data_i[7];
    end 
    if(N8383) begin
      \nz.mem_2006_sv2v_reg  <= data_i[6];
    end 
    if(N8382) begin
      \nz.mem_2005_sv2v_reg  <= data_i[5];
    end 
    if(N8381) begin
      \nz.mem_2004_sv2v_reg  <= data_i[4];
    end 
    if(N8380) begin
      \nz.mem_2003_sv2v_reg  <= data_i[3];
    end 
    if(N8379) begin
      \nz.mem_2002_sv2v_reg  <= data_i[2];
    end 
    if(N8378) begin
      \nz.mem_2001_sv2v_reg  <= data_i[1];
    end 
    if(N8377) begin
      \nz.mem_2000_sv2v_reg  <= data_i[0];
    end 
    if(N8376) begin
      \nz.mem_1999_sv2v_reg  <= data_i[79];
    end 
    if(N8375) begin
      \nz.mem_1998_sv2v_reg  <= data_i[78];
    end 
    if(N8374) begin
      \nz.mem_1997_sv2v_reg  <= data_i[77];
    end 
    if(N8373) begin
      \nz.mem_1996_sv2v_reg  <= data_i[76];
    end 
    if(N8372) begin
      \nz.mem_1995_sv2v_reg  <= data_i[75];
    end 
    if(N8371) begin
      \nz.mem_1994_sv2v_reg  <= data_i[74];
    end 
    if(N8370) begin
      \nz.mem_1993_sv2v_reg  <= data_i[73];
    end 
    if(N8369) begin
      \nz.mem_1992_sv2v_reg  <= data_i[72];
    end 
    if(N8368) begin
      \nz.mem_1991_sv2v_reg  <= data_i[71];
    end 
    if(N8367) begin
      \nz.mem_1990_sv2v_reg  <= data_i[70];
    end 
    if(N8366) begin
      \nz.mem_1989_sv2v_reg  <= data_i[69];
    end 
    if(N8365) begin
      \nz.mem_1988_sv2v_reg  <= data_i[68];
    end 
    if(N8364) begin
      \nz.mem_1987_sv2v_reg  <= data_i[67];
    end 
    if(N8363) begin
      \nz.mem_1986_sv2v_reg  <= data_i[66];
    end 
    if(N8362) begin
      \nz.mem_1985_sv2v_reg  <= data_i[65];
    end 
    if(N8361) begin
      \nz.mem_1984_sv2v_reg  <= data_i[64];
    end 
    if(N8360) begin
      \nz.mem_1983_sv2v_reg  <= data_i[63];
    end 
    if(N8359) begin
      \nz.mem_1982_sv2v_reg  <= data_i[62];
    end 
    if(N8358) begin
      \nz.mem_1981_sv2v_reg  <= data_i[61];
    end 
    if(N8357) begin
      \nz.mem_1980_sv2v_reg  <= data_i[60];
    end 
    if(N8356) begin
      \nz.mem_1979_sv2v_reg  <= data_i[59];
    end 
    if(N8355) begin
      \nz.mem_1978_sv2v_reg  <= data_i[58];
    end 
    if(N8354) begin
      \nz.mem_1977_sv2v_reg  <= data_i[57];
    end 
    if(N8353) begin
      \nz.mem_1976_sv2v_reg  <= data_i[56];
    end 
    if(N8352) begin
      \nz.mem_1975_sv2v_reg  <= data_i[55];
    end 
    if(N8351) begin
      \nz.mem_1974_sv2v_reg  <= data_i[54];
    end 
    if(N8350) begin
      \nz.mem_1973_sv2v_reg  <= data_i[53];
    end 
    if(N8349) begin
      \nz.mem_1972_sv2v_reg  <= data_i[52];
    end 
    if(N8348) begin
      \nz.mem_1971_sv2v_reg  <= data_i[51];
    end 
    if(N8347) begin
      \nz.mem_1970_sv2v_reg  <= data_i[50];
    end 
    if(N8346) begin
      \nz.mem_1969_sv2v_reg  <= data_i[49];
    end 
    if(N8345) begin
      \nz.mem_1968_sv2v_reg  <= data_i[48];
    end 
    if(N8344) begin
      \nz.mem_1967_sv2v_reg  <= data_i[47];
    end 
    if(N8343) begin
      \nz.mem_1966_sv2v_reg  <= data_i[46];
    end 
    if(N8342) begin
      \nz.mem_1965_sv2v_reg  <= data_i[45];
    end 
    if(N8341) begin
      \nz.mem_1964_sv2v_reg  <= data_i[44];
    end 
    if(N8340) begin
      \nz.mem_1963_sv2v_reg  <= data_i[43];
    end 
    if(N8339) begin
      \nz.mem_1962_sv2v_reg  <= data_i[42];
    end 
    if(N8338) begin
      \nz.mem_1961_sv2v_reg  <= data_i[41];
    end 
    if(N8337) begin
      \nz.mem_1960_sv2v_reg  <= data_i[40];
    end 
    if(N8336) begin
      \nz.mem_1959_sv2v_reg  <= data_i[39];
    end 
    if(N8335) begin
      \nz.mem_1958_sv2v_reg  <= data_i[38];
    end 
    if(N8334) begin
      \nz.mem_1957_sv2v_reg  <= data_i[37];
    end 
    if(N8333) begin
      \nz.mem_1956_sv2v_reg  <= data_i[36];
    end 
    if(N8332) begin
      \nz.mem_1955_sv2v_reg  <= data_i[35];
    end 
    if(N8331) begin
      \nz.mem_1954_sv2v_reg  <= data_i[34];
    end 
    if(N8330) begin
      \nz.mem_1953_sv2v_reg  <= data_i[33];
    end 
    if(N8329) begin
      \nz.mem_1952_sv2v_reg  <= data_i[32];
    end 
    if(N8328) begin
      \nz.mem_1951_sv2v_reg  <= data_i[31];
    end 
    if(N8327) begin
      \nz.mem_1950_sv2v_reg  <= data_i[30];
    end 
    if(N8326) begin
      \nz.mem_1949_sv2v_reg  <= data_i[29];
    end 
    if(N8325) begin
      \nz.mem_1948_sv2v_reg  <= data_i[28];
    end 
    if(N8324) begin
      \nz.mem_1947_sv2v_reg  <= data_i[27];
    end 
    if(N8323) begin
      \nz.mem_1946_sv2v_reg  <= data_i[26];
    end 
    if(N8322) begin
      \nz.mem_1945_sv2v_reg  <= data_i[25];
    end 
    if(N8321) begin
      \nz.mem_1944_sv2v_reg  <= data_i[24];
    end 
    if(N8320) begin
      \nz.mem_1943_sv2v_reg  <= data_i[23];
    end 
    if(N8319) begin
      \nz.mem_1942_sv2v_reg  <= data_i[22];
    end 
    if(N8318) begin
      \nz.mem_1941_sv2v_reg  <= data_i[21];
    end 
    if(N8317) begin
      \nz.mem_1940_sv2v_reg  <= data_i[20];
    end 
    if(N8316) begin
      \nz.mem_1939_sv2v_reg  <= data_i[19];
    end 
    if(N8315) begin
      \nz.mem_1938_sv2v_reg  <= data_i[18];
    end 
    if(N8314) begin
      \nz.mem_1937_sv2v_reg  <= data_i[17];
    end 
    if(N8313) begin
      \nz.mem_1936_sv2v_reg  <= data_i[16];
    end 
    if(N8312) begin
      \nz.mem_1935_sv2v_reg  <= data_i[15];
    end 
    if(N8311) begin
      \nz.mem_1934_sv2v_reg  <= data_i[14];
    end 
    if(N8310) begin
      \nz.mem_1933_sv2v_reg  <= data_i[13];
    end 
    if(N8309) begin
      \nz.mem_1932_sv2v_reg  <= data_i[12];
    end 
    if(N8308) begin
      \nz.mem_1931_sv2v_reg  <= data_i[11];
    end 
    if(N8307) begin
      \nz.mem_1930_sv2v_reg  <= data_i[10];
    end 
    if(N8306) begin
      \nz.mem_1929_sv2v_reg  <= data_i[9];
    end 
    if(N8305) begin
      \nz.mem_1928_sv2v_reg  <= data_i[8];
    end 
    if(N8304) begin
      \nz.mem_1927_sv2v_reg  <= data_i[7];
    end 
    if(N8303) begin
      \nz.mem_1926_sv2v_reg  <= data_i[6];
    end 
    if(N8302) begin
      \nz.mem_1925_sv2v_reg  <= data_i[5];
    end 
    if(N8301) begin
      \nz.mem_1924_sv2v_reg  <= data_i[4];
    end 
    if(N8300) begin
      \nz.mem_1923_sv2v_reg  <= data_i[3];
    end 
    if(N8299) begin
      \nz.mem_1922_sv2v_reg  <= data_i[2];
    end 
    if(N8298) begin
      \nz.mem_1921_sv2v_reg  <= data_i[1];
    end 
    if(N8297) begin
      \nz.mem_1920_sv2v_reg  <= data_i[0];
    end 
    if(N8296) begin
      \nz.mem_1919_sv2v_reg  <= data_i[79];
    end 
    if(N8295) begin
      \nz.mem_1918_sv2v_reg  <= data_i[78];
    end 
    if(N8294) begin
      \nz.mem_1917_sv2v_reg  <= data_i[77];
    end 
    if(N8293) begin
      \nz.mem_1916_sv2v_reg  <= data_i[76];
    end 
    if(N8292) begin
      \nz.mem_1915_sv2v_reg  <= data_i[75];
    end 
    if(N8291) begin
      \nz.mem_1914_sv2v_reg  <= data_i[74];
    end 
    if(N8290) begin
      \nz.mem_1913_sv2v_reg  <= data_i[73];
    end 
    if(N8289) begin
      \nz.mem_1912_sv2v_reg  <= data_i[72];
    end 
    if(N8288) begin
      \nz.mem_1911_sv2v_reg  <= data_i[71];
    end 
    if(N8287) begin
      \nz.mem_1910_sv2v_reg  <= data_i[70];
    end 
    if(N8286) begin
      \nz.mem_1909_sv2v_reg  <= data_i[69];
    end 
    if(N8285) begin
      \nz.mem_1908_sv2v_reg  <= data_i[68];
    end 
    if(N8284) begin
      \nz.mem_1907_sv2v_reg  <= data_i[67];
    end 
    if(N8283) begin
      \nz.mem_1906_sv2v_reg  <= data_i[66];
    end 
    if(N8282) begin
      \nz.mem_1905_sv2v_reg  <= data_i[65];
    end 
    if(N8281) begin
      \nz.mem_1904_sv2v_reg  <= data_i[64];
    end 
    if(N8280) begin
      \nz.mem_1903_sv2v_reg  <= data_i[63];
    end 
    if(N8279) begin
      \nz.mem_1902_sv2v_reg  <= data_i[62];
    end 
    if(N8278) begin
      \nz.mem_1901_sv2v_reg  <= data_i[61];
    end 
    if(N8277) begin
      \nz.mem_1900_sv2v_reg  <= data_i[60];
    end 
    if(N8276) begin
      \nz.mem_1899_sv2v_reg  <= data_i[59];
    end 
    if(N8275) begin
      \nz.mem_1898_sv2v_reg  <= data_i[58];
    end 
    if(N8274) begin
      \nz.mem_1897_sv2v_reg  <= data_i[57];
    end 
    if(N8273) begin
      \nz.mem_1896_sv2v_reg  <= data_i[56];
    end 
    if(N8272) begin
      \nz.mem_1895_sv2v_reg  <= data_i[55];
    end 
    if(N8271) begin
      \nz.mem_1894_sv2v_reg  <= data_i[54];
    end 
    if(N8270) begin
      \nz.mem_1893_sv2v_reg  <= data_i[53];
    end 
    if(N8269) begin
      \nz.mem_1892_sv2v_reg  <= data_i[52];
    end 
    if(N8268) begin
      \nz.mem_1891_sv2v_reg  <= data_i[51];
    end 
    if(N8267) begin
      \nz.mem_1890_sv2v_reg  <= data_i[50];
    end 
    if(N8266) begin
      \nz.mem_1889_sv2v_reg  <= data_i[49];
    end 
    if(N8265) begin
      \nz.mem_1888_sv2v_reg  <= data_i[48];
    end 
    if(N8264) begin
      \nz.mem_1887_sv2v_reg  <= data_i[47];
    end 
    if(N8263) begin
      \nz.mem_1886_sv2v_reg  <= data_i[46];
    end 
    if(N8262) begin
      \nz.mem_1885_sv2v_reg  <= data_i[45];
    end 
    if(N8261) begin
      \nz.mem_1884_sv2v_reg  <= data_i[44];
    end 
    if(N8260) begin
      \nz.mem_1883_sv2v_reg  <= data_i[43];
    end 
    if(N8259) begin
      \nz.mem_1882_sv2v_reg  <= data_i[42];
    end 
    if(N8258) begin
      \nz.mem_1881_sv2v_reg  <= data_i[41];
    end 
    if(N8257) begin
      \nz.mem_1880_sv2v_reg  <= data_i[40];
    end 
    if(N8256) begin
      \nz.mem_1879_sv2v_reg  <= data_i[39];
    end 
    if(N8255) begin
      \nz.mem_1878_sv2v_reg  <= data_i[38];
    end 
    if(N8254) begin
      \nz.mem_1877_sv2v_reg  <= data_i[37];
    end 
    if(N8253) begin
      \nz.mem_1876_sv2v_reg  <= data_i[36];
    end 
    if(N8252) begin
      \nz.mem_1875_sv2v_reg  <= data_i[35];
    end 
    if(N8251) begin
      \nz.mem_1874_sv2v_reg  <= data_i[34];
    end 
    if(N8250) begin
      \nz.mem_1873_sv2v_reg  <= data_i[33];
    end 
    if(N8249) begin
      \nz.mem_1872_sv2v_reg  <= data_i[32];
    end 
    if(N8248) begin
      \nz.mem_1871_sv2v_reg  <= data_i[31];
    end 
    if(N8247) begin
      \nz.mem_1870_sv2v_reg  <= data_i[30];
    end 
    if(N8246) begin
      \nz.mem_1869_sv2v_reg  <= data_i[29];
    end 
    if(N8245) begin
      \nz.mem_1868_sv2v_reg  <= data_i[28];
    end 
    if(N8244) begin
      \nz.mem_1867_sv2v_reg  <= data_i[27];
    end 
    if(N8243) begin
      \nz.mem_1866_sv2v_reg  <= data_i[26];
    end 
    if(N8242) begin
      \nz.mem_1865_sv2v_reg  <= data_i[25];
    end 
    if(N8241) begin
      \nz.mem_1864_sv2v_reg  <= data_i[24];
    end 
    if(N8240) begin
      \nz.mem_1863_sv2v_reg  <= data_i[23];
    end 
    if(N8239) begin
      \nz.mem_1862_sv2v_reg  <= data_i[22];
    end 
    if(N8238) begin
      \nz.mem_1861_sv2v_reg  <= data_i[21];
    end 
    if(N8237) begin
      \nz.mem_1860_sv2v_reg  <= data_i[20];
    end 
    if(N8236) begin
      \nz.mem_1859_sv2v_reg  <= data_i[19];
    end 
    if(N8235) begin
      \nz.mem_1858_sv2v_reg  <= data_i[18];
    end 
    if(N8234) begin
      \nz.mem_1857_sv2v_reg  <= data_i[17];
    end 
    if(N8233) begin
      \nz.mem_1856_sv2v_reg  <= data_i[16];
    end 
    if(N8232) begin
      \nz.mem_1855_sv2v_reg  <= data_i[15];
    end 
    if(N8231) begin
      \nz.mem_1854_sv2v_reg  <= data_i[14];
    end 
    if(N8230) begin
      \nz.mem_1853_sv2v_reg  <= data_i[13];
    end 
    if(N8229) begin
      \nz.mem_1852_sv2v_reg  <= data_i[12];
    end 
    if(N8228) begin
      \nz.mem_1851_sv2v_reg  <= data_i[11];
    end 
    if(N8227) begin
      \nz.mem_1850_sv2v_reg  <= data_i[10];
    end 
    if(N8226) begin
      \nz.mem_1849_sv2v_reg  <= data_i[9];
    end 
    if(N8225) begin
      \nz.mem_1848_sv2v_reg  <= data_i[8];
    end 
    if(N8224) begin
      \nz.mem_1847_sv2v_reg  <= data_i[7];
    end 
    if(N8223) begin
      \nz.mem_1846_sv2v_reg  <= data_i[6];
    end 
    if(N8222) begin
      \nz.mem_1845_sv2v_reg  <= data_i[5];
    end 
    if(N8221) begin
      \nz.mem_1844_sv2v_reg  <= data_i[4];
    end 
    if(N8220) begin
      \nz.mem_1843_sv2v_reg  <= data_i[3];
    end 
    if(N8219) begin
      \nz.mem_1842_sv2v_reg  <= data_i[2];
    end 
    if(N8218) begin
      \nz.mem_1841_sv2v_reg  <= data_i[1];
    end 
    if(N8217) begin
      \nz.mem_1840_sv2v_reg  <= data_i[0];
    end 
    if(N8216) begin
      \nz.mem_1839_sv2v_reg  <= data_i[79];
    end 
    if(N8215) begin
      \nz.mem_1838_sv2v_reg  <= data_i[78];
    end 
    if(N8214) begin
      \nz.mem_1837_sv2v_reg  <= data_i[77];
    end 
    if(N8213) begin
      \nz.mem_1836_sv2v_reg  <= data_i[76];
    end 
    if(N8212) begin
      \nz.mem_1835_sv2v_reg  <= data_i[75];
    end 
    if(N8211) begin
      \nz.mem_1834_sv2v_reg  <= data_i[74];
    end 
    if(N8210) begin
      \nz.mem_1833_sv2v_reg  <= data_i[73];
    end 
    if(N8209) begin
      \nz.mem_1832_sv2v_reg  <= data_i[72];
    end 
    if(N8208) begin
      \nz.mem_1831_sv2v_reg  <= data_i[71];
    end 
    if(N8207) begin
      \nz.mem_1830_sv2v_reg  <= data_i[70];
    end 
    if(N8206) begin
      \nz.mem_1829_sv2v_reg  <= data_i[69];
    end 
    if(N8205) begin
      \nz.mem_1828_sv2v_reg  <= data_i[68];
    end 
    if(N8204) begin
      \nz.mem_1827_sv2v_reg  <= data_i[67];
    end 
    if(N8203) begin
      \nz.mem_1826_sv2v_reg  <= data_i[66];
    end 
    if(N8202) begin
      \nz.mem_1825_sv2v_reg  <= data_i[65];
    end 
    if(N8201) begin
      \nz.mem_1824_sv2v_reg  <= data_i[64];
    end 
    if(N8200) begin
      \nz.mem_1823_sv2v_reg  <= data_i[63];
    end 
    if(N8199) begin
      \nz.mem_1822_sv2v_reg  <= data_i[62];
    end 
    if(N8198) begin
      \nz.mem_1821_sv2v_reg  <= data_i[61];
    end 
    if(N8197) begin
      \nz.mem_1820_sv2v_reg  <= data_i[60];
    end 
    if(N8196) begin
      \nz.mem_1819_sv2v_reg  <= data_i[59];
    end 
    if(N8195) begin
      \nz.mem_1818_sv2v_reg  <= data_i[58];
    end 
    if(N8194) begin
      \nz.mem_1817_sv2v_reg  <= data_i[57];
    end 
    if(N8193) begin
      \nz.mem_1816_sv2v_reg  <= data_i[56];
    end 
    if(N8192) begin
      \nz.mem_1815_sv2v_reg  <= data_i[55];
    end 
    if(N8191) begin
      \nz.mem_1814_sv2v_reg  <= data_i[54];
    end 
    if(N8190) begin
      \nz.mem_1813_sv2v_reg  <= data_i[53];
    end 
    if(N8189) begin
      \nz.mem_1812_sv2v_reg  <= data_i[52];
    end 
    if(N8188) begin
      \nz.mem_1811_sv2v_reg  <= data_i[51];
    end 
    if(N8187) begin
      \nz.mem_1810_sv2v_reg  <= data_i[50];
    end 
    if(N8186) begin
      \nz.mem_1809_sv2v_reg  <= data_i[49];
    end 
    if(N8185) begin
      \nz.mem_1808_sv2v_reg  <= data_i[48];
    end 
    if(N8184) begin
      \nz.mem_1807_sv2v_reg  <= data_i[47];
    end 
    if(N8183) begin
      \nz.mem_1806_sv2v_reg  <= data_i[46];
    end 
    if(N8182) begin
      \nz.mem_1805_sv2v_reg  <= data_i[45];
    end 
    if(N8181) begin
      \nz.mem_1804_sv2v_reg  <= data_i[44];
    end 
    if(N8180) begin
      \nz.mem_1803_sv2v_reg  <= data_i[43];
    end 
    if(N8179) begin
      \nz.mem_1802_sv2v_reg  <= data_i[42];
    end 
    if(N8178) begin
      \nz.mem_1801_sv2v_reg  <= data_i[41];
    end 
    if(N8177) begin
      \nz.mem_1800_sv2v_reg  <= data_i[40];
    end 
    if(N8176) begin
      \nz.mem_1799_sv2v_reg  <= data_i[39];
    end 
    if(N8175) begin
      \nz.mem_1798_sv2v_reg  <= data_i[38];
    end 
    if(N8174) begin
      \nz.mem_1797_sv2v_reg  <= data_i[37];
    end 
    if(N8173) begin
      \nz.mem_1796_sv2v_reg  <= data_i[36];
    end 
    if(N8172) begin
      \nz.mem_1795_sv2v_reg  <= data_i[35];
    end 
    if(N8171) begin
      \nz.mem_1794_sv2v_reg  <= data_i[34];
    end 
    if(N8170) begin
      \nz.mem_1793_sv2v_reg  <= data_i[33];
    end 
    if(N8169) begin
      \nz.mem_1792_sv2v_reg  <= data_i[32];
    end 
    if(N8168) begin
      \nz.mem_1791_sv2v_reg  <= data_i[31];
    end 
    if(N8167) begin
      \nz.mem_1790_sv2v_reg  <= data_i[30];
    end 
    if(N8166) begin
      \nz.mem_1789_sv2v_reg  <= data_i[29];
    end 
    if(N8165) begin
      \nz.mem_1788_sv2v_reg  <= data_i[28];
    end 
    if(N8164) begin
      \nz.mem_1787_sv2v_reg  <= data_i[27];
    end 
    if(N8163) begin
      \nz.mem_1786_sv2v_reg  <= data_i[26];
    end 
    if(N8162) begin
      \nz.mem_1785_sv2v_reg  <= data_i[25];
    end 
    if(N8161) begin
      \nz.mem_1784_sv2v_reg  <= data_i[24];
    end 
    if(N8160) begin
      \nz.mem_1783_sv2v_reg  <= data_i[23];
    end 
    if(N8159) begin
      \nz.mem_1782_sv2v_reg  <= data_i[22];
    end 
    if(N8158) begin
      \nz.mem_1781_sv2v_reg  <= data_i[21];
    end 
    if(N8157) begin
      \nz.mem_1780_sv2v_reg  <= data_i[20];
    end 
    if(N8156) begin
      \nz.mem_1779_sv2v_reg  <= data_i[19];
    end 
    if(N8155) begin
      \nz.mem_1778_sv2v_reg  <= data_i[18];
    end 
    if(N8154) begin
      \nz.mem_1777_sv2v_reg  <= data_i[17];
    end 
    if(N8153) begin
      \nz.mem_1776_sv2v_reg  <= data_i[16];
    end 
    if(N8152) begin
      \nz.mem_1775_sv2v_reg  <= data_i[15];
    end 
    if(N8151) begin
      \nz.mem_1774_sv2v_reg  <= data_i[14];
    end 
    if(N8150) begin
      \nz.mem_1773_sv2v_reg  <= data_i[13];
    end 
    if(N8149) begin
      \nz.mem_1772_sv2v_reg  <= data_i[12];
    end 
    if(N8148) begin
      \nz.mem_1771_sv2v_reg  <= data_i[11];
    end 
    if(N8147) begin
      \nz.mem_1770_sv2v_reg  <= data_i[10];
    end 
    if(N8146) begin
      \nz.mem_1769_sv2v_reg  <= data_i[9];
    end 
    if(N8145) begin
      \nz.mem_1768_sv2v_reg  <= data_i[8];
    end 
    if(N8144) begin
      \nz.mem_1767_sv2v_reg  <= data_i[7];
    end 
    if(N8143) begin
      \nz.mem_1766_sv2v_reg  <= data_i[6];
    end 
    if(N8142) begin
      \nz.mem_1765_sv2v_reg  <= data_i[5];
    end 
    if(N8141) begin
      \nz.mem_1764_sv2v_reg  <= data_i[4];
    end 
    if(N8140) begin
      \nz.mem_1763_sv2v_reg  <= data_i[3];
    end 
    if(N8139) begin
      \nz.mem_1762_sv2v_reg  <= data_i[2];
    end 
    if(N8138) begin
      \nz.mem_1761_sv2v_reg  <= data_i[1];
    end 
    if(N8137) begin
      \nz.mem_1760_sv2v_reg  <= data_i[0];
    end 
    if(N8136) begin
      \nz.mem_1759_sv2v_reg  <= data_i[79];
    end 
    if(N8135) begin
      \nz.mem_1758_sv2v_reg  <= data_i[78];
    end 
    if(N8134) begin
      \nz.mem_1757_sv2v_reg  <= data_i[77];
    end 
    if(N8133) begin
      \nz.mem_1756_sv2v_reg  <= data_i[76];
    end 
    if(N8132) begin
      \nz.mem_1755_sv2v_reg  <= data_i[75];
    end 
    if(N8131) begin
      \nz.mem_1754_sv2v_reg  <= data_i[74];
    end 
    if(N8130) begin
      \nz.mem_1753_sv2v_reg  <= data_i[73];
    end 
    if(N8129) begin
      \nz.mem_1752_sv2v_reg  <= data_i[72];
    end 
    if(N8128) begin
      \nz.mem_1751_sv2v_reg  <= data_i[71];
    end 
    if(N8127) begin
      \nz.mem_1750_sv2v_reg  <= data_i[70];
    end 
    if(N8126) begin
      \nz.mem_1749_sv2v_reg  <= data_i[69];
    end 
    if(N8125) begin
      \nz.mem_1748_sv2v_reg  <= data_i[68];
    end 
    if(N8124) begin
      \nz.mem_1747_sv2v_reg  <= data_i[67];
    end 
    if(N8123) begin
      \nz.mem_1746_sv2v_reg  <= data_i[66];
    end 
    if(N8122) begin
      \nz.mem_1745_sv2v_reg  <= data_i[65];
    end 
    if(N8121) begin
      \nz.mem_1744_sv2v_reg  <= data_i[64];
    end 
    if(N8120) begin
      \nz.mem_1743_sv2v_reg  <= data_i[63];
    end 
    if(N8119) begin
      \nz.mem_1742_sv2v_reg  <= data_i[62];
    end 
    if(N8118) begin
      \nz.mem_1741_sv2v_reg  <= data_i[61];
    end 
    if(N8117) begin
      \nz.mem_1740_sv2v_reg  <= data_i[60];
    end 
    if(N8116) begin
      \nz.mem_1739_sv2v_reg  <= data_i[59];
    end 
    if(N8115) begin
      \nz.mem_1738_sv2v_reg  <= data_i[58];
    end 
    if(N8114) begin
      \nz.mem_1737_sv2v_reg  <= data_i[57];
    end 
    if(N8113) begin
      \nz.mem_1736_sv2v_reg  <= data_i[56];
    end 
    if(N8112) begin
      \nz.mem_1735_sv2v_reg  <= data_i[55];
    end 
    if(N8111) begin
      \nz.mem_1734_sv2v_reg  <= data_i[54];
    end 
    if(N8110) begin
      \nz.mem_1733_sv2v_reg  <= data_i[53];
    end 
    if(N8109) begin
      \nz.mem_1732_sv2v_reg  <= data_i[52];
    end 
    if(N8108) begin
      \nz.mem_1731_sv2v_reg  <= data_i[51];
    end 
    if(N8107) begin
      \nz.mem_1730_sv2v_reg  <= data_i[50];
    end 
    if(N8106) begin
      \nz.mem_1729_sv2v_reg  <= data_i[49];
    end 
    if(N8105) begin
      \nz.mem_1728_sv2v_reg  <= data_i[48];
    end 
    if(N8104) begin
      \nz.mem_1727_sv2v_reg  <= data_i[47];
    end 
    if(N8103) begin
      \nz.mem_1726_sv2v_reg  <= data_i[46];
    end 
    if(N8102) begin
      \nz.mem_1725_sv2v_reg  <= data_i[45];
    end 
    if(N8101) begin
      \nz.mem_1724_sv2v_reg  <= data_i[44];
    end 
    if(N8100) begin
      \nz.mem_1723_sv2v_reg  <= data_i[43];
    end 
    if(N8099) begin
      \nz.mem_1722_sv2v_reg  <= data_i[42];
    end 
    if(N8098) begin
      \nz.mem_1721_sv2v_reg  <= data_i[41];
    end 
    if(N8097) begin
      \nz.mem_1720_sv2v_reg  <= data_i[40];
    end 
    if(N8096) begin
      \nz.mem_1719_sv2v_reg  <= data_i[39];
    end 
    if(N8095) begin
      \nz.mem_1718_sv2v_reg  <= data_i[38];
    end 
    if(N8094) begin
      \nz.mem_1717_sv2v_reg  <= data_i[37];
    end 
    if(N8093) begin
      \nz.mem_1716_sv2v_reg  <= data_i[36];
    end 
    if(N8092) begin
      \nz.mem_1715_sv2v_reg  <= data_i[35];
    end 
    if(N8091) begin
      \nz.mem_1714_sv2v_reg  <= data_i[34];
    end 
    if(N8090) begin
      \nz.mem_1713_sv2v_reg  <= data_i[33];
    end 
    if(N8089) begin
      \nz.mem_1712_sv2v_reg  <= data_i[32];
    end 
    if(N8088) begin
      \nz.mem_1711_sv2v_reg  <= data_i[31];
    end 
    if(N8087) begin
      \nz.mem_1710_sv2v_reg  <= data_i[30];
    end 
    if(N8086) begin
      \nz.mem_1709_sv2v_reg  <= data_i[29];
    end 
    if(N8085) begin
      \nz.mem_1708_sv2v_reg  <= data_i[28];
    end 
    if(N8084) begin
      \nz.mem_1707_sv2v_reg  <= data_i[27];
    end 
    if(N8083) begin
      \nz.mem_1706_sv2v_reg  <= data_i[26];
    end 
    if(N8082) begin
      \nz.mem_1705_sv2v_reg  <= data_i[25];
    end 
    if(N8081) begin
      \nz.mem_1704_sv2v_reg  <= data_i[24];
    end 
    if(N8080) begin
      \nz.mem_1703_sv2v_reg  <= data_i[23];
    end 
    if(N8079) begin
      \nz.mem_1702_sv2v_reg  <= data_i[22];
    end 
    if(N8078) begin
      \nz.mem_1701_sv2v_reg  <= data_i[21];
    end 
    if(N8077) begin
      \nz.mem_1700_sv2v_reg  <= data_i[20];
    end 
    if(N8076) begin
      \nz.mem_1699_sv2v_reg  <= data_i[19];
    end 
    if(N8075) begin
      \nz.mem_1698_sv2v_reg  <= data_i[18];
    end 
    if(N8074) begin
      \nz.mem_1697_sv2v_reg  <= data_i[17];
    end 
    if(N8073) begin
      \nz.mem_1696_sv2v_reg  <= data_i[16];
    end 
    if(N8072) begin
      \nz.mem_1695_sv2v_reg  <= data_i[15];
    end 
    if(N8071) begin
      \nz.mem_1694_sv2v_reg  <= data_i[14];
    end 
    if(N8070) begin
      \nz.mem_1693_sv2v_reg  <= data_i[13];
    end 
    if(N8069) begin
      \nz.mem_1692_sv2v_reg  <= data_i[12];
    end 
    if(N8068) begin
      \nz.mem_1691_sv2v_reg  <= data_i[11];
    end 
    if(N8067) begin
      \nz.mem_1690_sv2v_reg  <= data_i[10];
    end 
    if(N8066) begin
      \nz.mem_1689_sv2v_reg  <= data_i[9];
    end 
    if(N8065) begin
      \nz.mem_1688_sv2v_reg  <= data_i[8];
    end 
    if(N8064) begin
      \nz.mem_1687_sv2v_reg  <= data_i[7];
    end 
    if(N8063) begin
      \nz.mem_1686_sv2v_reg  <= data_i[6];
    end 
    if(N8062) begin
      \nz.mem_1685_sv2v_reg  <= data_i[5];
    end 
    if(N8061) begin
      \nz.mem_1684_sv2v_reg  <= data_i[4];
    end 
    if(N8060) begin
      \nz.mem_1683_sv2v_reg  <= data_i[3];
    end 
    if(N8059) begin
      \nz.mem_1682_sv2v_reg  <= data_i[2];
    end 
    if(N8058) begin
      \nz.mem_1681_sv2v_reg  <= data_i[1];
    end 
    if(N8057) begin
      \nz.mem_1680_sv2v_reg  <= data_i[0];
    end 
    if(N8056) begin
      \nz.mem_1679_sv2v_reg  <= data_i[79];
    end 
    if(N8055) begin
      \nz.mem_1678_sv2v_reg  <= data_i[78];
    end 
    if(N8054) begin
      \nz.mem_1677_sv2v_reg  <= data_i[77];
    end 
    if(N8053) begin
      \nz.mem_1676_sv2v_reg  <= data_i[76];
    end 
    if(N8052) begin
      \nz.mem_1675_sv2v_reg  <= data_i[75];
    end 
    if(N8051) begin
      \nz.mem_1674_sv2v_reg  <= data_i[74];
    end 
    if(N8050) begin
      \nz.mem_1673_sv2v_reg  <= data_i[73];
    end 
    if(N8049) begin
      \nz.mem_1672_sv2v_reg  <= data_i[72];
    end 
    if(N8048) begin
      \nz.mem_1671_sv2v_reg  <= data_i[71];
    end 
    if(N8047) begin
      \nz.mem_1670_sv2v_reg  <= data_i[70];
    end 
    if(N8046) begin
      \nz.mem_1669_sv2v_reg  <= data_i[69];
    end 
    if(N8045) begin
      \nz.mem_1668_sv2v_reg  <= data_i[68];
    end 
    if(N8044) begin
      \nz.mem_1667_sv2v_reg  <= data_i[67];
    end 
    if(N8043) begin
      \nz.mem_1666_sv2v_reg  <= data_i[66];
    end 
    if(N8042) begin
      \nz.mem_1665_sv2v_reg  <= data_i[65];
    end 
    if(N8041) begin
      \nz.mem_1664_sv2v_reg  <= data_i[64];
    end 
    if(N8040) begin
      \nz.mem_1663_sv2v_reg  <= data_i[63];
    end 
    if(N8039) begin
      \nz.mem_1662_sv2v_reg  <= data_i[62];
    end 
    if(N8038) begin
      \nz.mem_1661_sv2v_reg  <= data_i[61];
    end 
    if(N8037) begin
      \nz.mem_1660_sv2v_reg  <= data_i[60];
    end 
    if(N8036) begin
      \nz.mem_1659_sv2v_reg  <= data_i[59];
    end 
    if(N8035) begin
      \nz.mem_1658_sv2v_reg  <= data_i[58];
    end 
    if(N8034) begin
      \nz.mem_1657_sv2v_reg  <= data_i[57];
    end 
    if(N8033) begin
      \nz.mem_1656_sv2v_reg  <= data_i[56];
    end 
    if(N8032) begin
      \nz.mem_1655_sv2v_reg  <= data_i[55];
    end 
    if(N8031) begin
      \nz.mem_1654_sv2v_reg  <= data_i[54];
    end 
    if(N8030) begin
      \nz.mem_1653_sv2v_reg  <= data_i[53];
    end 
    if(N8029) begin
      \nz.mem_1652_sv2v_reg  <= data_i[52];
    end 
    if(N8028) begin
      \nz.mem_1651_sv2v_reg  <= data_i[51];
    end 
    if(N8027) begin
      \nz.mem_1650_sv2v_reg  <= data_i[50];
    end 
    if(N8026) begin
      \nz.mem_1649_sv2v_reg  <= data_i[49];
    end 
    if(N8025) begin
      \nz.mem_1648_sv2v_reg  <= data_i[48];
    end 
    if(N8024) begin
      \nz.mem_1647_sv2v_reg  <= data_i[47];
    end 
    if(N8023) begin
      \nz.mem_1646_sv2v_reg  <= data_i[46];
    end 
    if(N8022) begin
      \nz.mem_1645_sv2v_reg  <= data_i[45];
    end 
    if(N8021) begin
      \nz.mem_1644_sv2v_reg  <= data_i[44];
    end 
    if(N8020) begin
      \nz.mem_1643_sv2v_reg  <= data_i[43];
    end 
    if(N8019) begin
      \nz.mem_1642_sv2v_reg  <= data_i[42];
    end 
    if(N8018) begin
      \nz.mem_1641_sv2v_reg  <= data_i[41];
    end 
    if(N8017) begin
      \nz.mem_1640_sv2v_reg  <= data_i[40];
    end 
    if(N8016) begin
      \nz.mem_1639_sv2v_reg  <= data_i[39];
    end 
    if(N8015) begin
      \nz.mem_1638_sv2v_reg  <= data_i[38];
    end 
    if(N8014) begin
      \nz.mem_1637_sv2v_reg  <= data_i[37];
    end 
    if(N8013) begin
      \nz.mem_1636_sv2v_reg  <= data_i[36];
    end 
    if(N8012) begin
      \nz.mem_1635_sv2v_reg  <= data_i[35];
    end 
    if(N8011) begin
      \nz.mem_1634_sv2v_reg  <= data_i[34];
    end 
    if(N8010) begin
      \nz.mem_1633_sv2v_reg  <= data_i[33];
    end 
    if(N8009) begin
      \nz.mem_1632_sv2v_reg  <= data_i[32];
    end 
    if(N8008) begin
      \nz.mem_1631_sv2v_reg  <= data_i[31];
    end 
    if(N8007) begin
      \nz.mem_1630_sv2v_reg  <= data_i[30];
    end 
    if(N8006) begin
      \nz.mem_1629_sv2v_reg  <= data_i[29];
    end 
    if(N8005) begin
      \nz.mem_1628_sv2v_reg  <= data_i[28];
    end 
    if(N8004) begin
      \nz.mem_1627_sv2v_reg  <= data_i[27];
    end 
    if(N8003) begin
      \nz.mem_1626_sv2v_reg  <= data_i[26];
    end 
    if(N8002) begin
      \nz.mem_1625_sv2v_reg  <= data_i[25];
    end 
    if(N8001) begin
      \nz.mem_1624_sv2v_reg  <= data_i[24];
    end 
    if(N8000) begin
      \nz.mem_1623_sv2v_reg  <= data_i[23];
    end 
    if(N7999) begin
      \nz.mem_1622_sv2v_reg  <= data_i[22];
    end 
    if(N7998) begin
      \nz.mem_1621_sv2v_reg  <= data_i[21];
    end 
    if(N7997) begin
      \nz.mem_1620_sv2v_reg  <= data_i[20];
    end 
    if(N7996) begin
      \nz.mem_1619_sv2v_reg  <= data_i[19];
    end 
    if(N7995) begin
      \nz.mem_1618_sv2v_reg  <= data_i[18];
    end 
    if(N7994) begin
      \nz.mem_1617_sv2v_reg  <= data_i[17];
    end 
    if(N7993) begin
      \nz.mem_1616_sv2v_reg  <= data_i[16];
    end 
    if(N7992) begin
      \nz.mem_1615_sv2v_reg  <= data_i[15];
    end 
    if(N7991) begin
      \nz.mem_1614_sv2v_reg  <= data_i[14];
    end 
    if(N7990) begin
      \nz.mem_1613_sv2v_reg  <= data_i[13];
    end 
    if(N7989) begin
      \nz.mem_1612_sv2v_reg  <= data_i[12];
    end 
    if(N7988) begin
      \nz.mem_1611_sv2v_reg  <= data_i[11];
    end 
    if(N7987) begin
      \nz.mem_1610_sv2v_reg  <= data_i[10];
    end 
    if(N7986) begin
      \nz.mem_1609_sv2v_reg  <= data_i[9];
    end 
    if(N7985) begin
      \nz.mem_1608_sv2v_reg  <= data_i[8];
    end 
    if(N7984) begin
      \nz.mem_1607_sv2v_reg  <= data_i[7];
    end 
    if(N7983) begin
      \nz.mem_1606_sv2v_reg  <= data_i[6];
    end 
    if(N7982) begin
      \nz.mem_1605_sv2v_reg  <= data_i[5];
    end 
    if(N7981) begin
      \nz.mem_1604_sv2v_reg  <= data_i[4];
    end 
    if(N7980) begin
      \nz.mem_1603_sv2v_reg  <= data_i[3];
    end 
    if(N7979) begin
      \nz.mem_1602_sv2v_reg  <= data_i[2];
    end 
    if(N7978) begin
      \nz.mem_1601_sv2v_reg  <= data_i[1];
    end 
    if(N7977) begin
      \nz.mem_1600_sv2v_reg  <= data_i[0];
    end 
    if(N7976) begin
      \nz.mem_1599_sv2v_reg  <= data_i[79];
    end 
    if(N7975) begin
      \nz.mem_1598_sv2v_reg  <= data_i[78];
    end 
    if(N7974) begin
      \nz.mem_1597_sv2v_reg  <= data_i[77];
    end 
    if(N7973) begin
      \nz.mem_1596_sv2v_reg  <= data_i[76];
    end 
    if(N7972) begin
      \nz.mem_1595_sv2v_reg  <= data_i[75];
    end 
    if(N7971) begin
      \nz.mem_1594_sv2v_reg  <= data_i[74];
    end 
    if(N7970) begin
      \nz.mem_1593_sv2v_reg  <= data_i[73];
    end 
    if(N7969) begin
      \nz.mem_1592_sv2v_reg  <= data_i[72];
    end 
    if(N7968) begin
      \nz.mem_1591_sv2v_reg  <= data_i[71];
    end 
    if(N7967) begin
      \nz.mem_1590_sv2v_reg  <= data_i[70];
    end 
    if(N7966) begin
      \nz.mem_1589_sv2v_reg  <= data_i[69];
    end 
    if(N7965) begin
      \nz.mem_1588_sv2v_reg  <= data_i[68];
    end 
    if(N7964) begin
      \nz.mem_1587_sv2v_reg  <= data_i[67];
    end 
    if(N7963) begin
      \nz.mem_1586_sv2v_reg  <= data_i[66];
    end 
    if(N7962) begin
      \nz.mem_1585_sv2v_reg  <= data_i[65];
    end 
    if(N7961) begin
      \nz.mem_1584_sv2v_reg  <= data_i[64];
    end 
    if(N7960) begin
      \nz.mem_1583_sv2v_reg  <= data_i[63];
    end 
    if(N7959) begin
      \nz.mem_1582_sv2v_reg  <= data_i[62];
    end 
    if(N7958) begin
      \nz.mem_1581_sv2v_reg  <= data_i[61];
    end 
    if(N7957) begin
      \nz.mem_1580_sv2v_reg  <= data_i[60];
    end 
    if(N7956) begin
      \nz.mem_1579_sv2v_reg  <= data_i[59];
    end 
    if(N7955) begin
      \nz.mem_1578_sv2v_reg  <= data_i[58];
    end 
    if(N7954) begin
      \nz.mem_1577_sv2v_reg  <= data_i[57];
    end 
    if(N7953) begin
      \nz.mem_1576_sv2v_reg  <= data_i[56];
    end 
    if(N7952) begin
      \nz.mem_1575_sv2v_reg  <= data_i[55];
    end 
    if(N7951) begin
      \nz.mem_1574_sv2v_reg  <= data_i[54];
    end 
    if(N7950) begin
      \nz.mem_1573_sv2v_reg  <= data_i[53];
    end 
    if(N7949) begin
      \nz.mem_1572_sv2v_reg  <= data_i[52];
    end 
    if(N7948) begin
      \nz.mem_1571_sv2v_reg  <= data_i[51];
    end 
    if(N7947) begin
      \nz.mem_1570_sv2v_reg  <= data_i[50];
    end 
    if(N7946) begin
      \nz.mem_1569_sv2v_reg  <= data_i[49];
    end 
    if(N7945) begin
      \nz.mem_1568_sv2v_reg  <= data_i[48];
    end 
    if(N7944) begin
      \nz.mem_1567_sv2v_reg  <= data_i[47];
    end 
    if(N7943) begin
      \nz.mem_1566_sv2v_reg  <= data_i[46];
    end 
    if(N7942) begin
      \nz.mem_1565_sv2v_reg  <= data_i[45];
    end 
    if(N7941) begin
      \nz.mem_1564_sv2v_reg  <= data_i[44];
    end 
    if(N7940) begin
      \nz.mem_1563_sv2v_reg  <= data_i[43];
    end 
    if(N7939) begin
      \nz.mem_1562_sv2v_reg  <= data_i[42];
    end 
    if(N7938) begin
      \nz.mem_1561_sv2v_reg  <= data_i[41];
    end 
    if(N7937) begin
      \nz.mem_1560_sv2v_reg  <= data_i[40];
    end 
    if(N7936) begin
      \nz.mem_1559_sv2v_reg  <= data_i[39];
    end 
    if(N7935) begin
      \nz.mem_1558_sv2v_reg  <= data_i[38];
    end 
    if(N7934) begin
      \nz.mem_1557_sv2v_reg  <= data_i[37];
    end 
    if(N7933) begin
      \nz.mem_1556_sv2v_reg  <= data_i[36];
    end 
    if(N7932) begin
      \nz.mem_1555_sv2v_reg  <= data_i[35];
    end 
    if(N7931) begin
      \nz.mem_1554_sv2v_reg  <= data_i[34];
    end 
    if(N7930) begin
      \nz.mem_1553_sv2v_reg  <= data_i[33];
    end 
    if(N7929) begin
      \nz.mem_1552_sv2v_reg  <= data_i[32];
    end 
    if(N7928) begin
      \nz.mem_1551_sv2v_reg  <= data_i[31];
    end 
    if(N7927) begin
      \nz.mem_1550_sv2v_reg  <= data_i[30];
    end 
    if(N7926) begin
      \nz.mem_1549_sv2v_reg  <= data_i[29];
    end 
    if(N7925) begin
      \nz.mem_1548_sv2v_reg  <= data_i[28];
    end 
    if(N7924) begin
      \nz.mem_1547_sv2v_reg  <= data_i[27];
    end 
    if(N7923) begin
      \nz.mem_1546_sv2v_reg  <= data_i[26];
    end 
    if(N7922) begin
      \nz.mem_1545_sv2v_reg  <= data_i[25];
    end 
    if(N7921) begin
      \nz.mem_1544_sv2v_reg  <= data_i[24];
    end 
    if(N7920) begin
      \nz.mem_1543_sv2v_reg  <= data_i[23];
    end 
    if(N7919) begin
      \nz.mem_1542_sv2v_reg  <= data_i[22];
    end 
    if(N7918) begin
      \nz.mem_1541_sv2v_reg  <= data_i[21];
    end 
    if(N7917) begin
      \nz.mem_1540_sv2v_reg  <= data_i[20];
    end 
    if(N7916) begin
      \nz.mem_1539_sv2v_reg  <= data_i[19];
    end 
    if(N7915) begin
      \nz.mem_1538_sv2v_reg  <= data_i[18];
    end 
    if(N7914) begin
      \nz.mem_1537_sv2v_reg  <= data_i[17];
    end 
    if(N7913) begin
      \nz.mem_1536_sv2v_reg  <= data_i[16];
    end 
    if(N7912) begin
      \nz.mem_1535_sv2v_reg  <= data_i[15];
    end 
    if(N7911) begin
      \nz.mem_1534_sv2v_reg  <= data_i[14];
    end 
    if(N7910) begin
      \nz.mem_1533_sv2v_reg  <= data_i[13];
    end 
    if(N7909) begin
      \nz.mem_1532_sv2v_reg  <= data_i[12];
    end 
    if(N7908) begin
      \nz.mem_1531_sv2v_reg  <= data_i[11];
    end 
    if(N7907) begin
      \nz.mem_1530_sv2v_reg  <= data_i[10];
    end 
    if(N7906) begin
      \nz.mem_1529_sv2v_reg  <= data_i[9];
    end 
    if(N7905) begin
      \nz.mem_1528_sv2v_reg  <= data_i[8];
    end 
    if(N7904) begin
      \nz.mem_1527_sv2v_reg  <= data_i[7];
    end 
    if(N7903) begin
      \nz.mem_1526_sv2v_reg  <= data_i[6];
    end 
    if(N7902) begin
      \nz.mem_1525_sv2v_reg  <= data_i[5];
    end 
    if(N7901) begin
      \nz.mem_1524_sv2v_reg  <= data_i[4];
    end 
    if(N7900) begin
      \nz.mem_1523_sv2v_reg  <= data_i[3];
    end 
    if(N7899) begin
      \nz.mem_1522_sv2v_reg  <= data_i[2];
    end 
    if(N7898) begin
      \nz.mem_1521_sv2v_reg  <= data_i[1];
    end 
    if(N7897) begin
      \nz.mem_1520_sv2v_reg  <= data_i[0];
    end 
    if(N7896) begin
      \nz.mem_1519_sv2v_reg  <= data_i[79];
    end 
    if(N7895) begin
      \nz.mem_1518_sv2v_reg  <= data_i[78];
    end 
    if(N7894) begin
      \nz.mem_1517_sv2v_reg  <= data_i[77];
    end 
    if(N7893) begin
      \nz.mem_1516_sv2v_reg  <= data_i[76];
    end 
    if(N7892) begin
      \nz.mem_1515_sv2v_reg  <= data_i[75];
    end 
    if(N7891) begin
      \nz.mem_1514_sv2v_reg  <= data_i[74];
    end 
    if(N7890) begin
      \nz.mem_1513_sv2v_reg  <= data_i[73];
    end 
    if(N7889) begin
      \nz.mem_1512_sv2v_reg  <= data_i[72];
    end 
    if(N7888) begin
      \nz.mem_1511_sv2v_reg  <= data_i[71];
    end 
    if(N7887) begin
      \nz.mem_1510_sv2v_reg  <= data_i[70];
    end 
    if(N7886) begin
      \nz.mem_1509_sv2v_reg  <= data_i[69];
    end 
    if(N7885) begin
      \nz.mem_1508_sv2v_reg  <= data_i[68];
    end 
    if(N7884) begin
      \nz.mem_1507_sv2v_reg  <= data_i[67];
    end 
    if(N7883) begin
      \nz.mem_1506_sv2v_reg  <= data_i[66];
    end 
    if(N7882) begin
      \nz.mem_1505_sv2v_reg  <= data_i[65];
    end 
    if(N7881) begin
      \nz.mem_1504_sv2v_reg  <= data_i[64];
    end 
    if(N7880) begin
      \nz.mem_1503_sv2v_reg  <= data_i[63];
    end 
    if(N7879) begin
      \nz.mem_1502_sv2v_reg  <= data_i[62];
    end 
    if(N7878) begin
      \nz.mem_1501_sv2v_reg  <= data_i[61];
    end 
    if(N7877) begin
      \nz.mem_1500_sv2v_reg  <= data_i[60];
    end 
    if(N7876) begin
      \nz.mem_1499_sv2v_reg  <= data_i[59];
    end 
    if(N7875) begin
      \nz.mem_1498_sv2v_reg  <= data_i[58];
    end 
    if(N7874) begin
      \nz.mem_1497_sv2v_reg  <= data_i[57];
    end 
    if(N7873) begin
      \nz.mem_1496_sv2v_reg  <= data_i[56];
    end 
    if(N7872) begin
      \nz.mem_1495_sv2v_reg  <= data_i[55];
    end 
    if(N7871) begin
      \nz.mem_1494_sv2v_reg  <= data_i[54];
    end 
    if(N7870) begin
      \nz.mem_1493_sv2v_reg  <= data_i[53];
    end 
    if(N7869) begin
      \nz.mem_1492_sv2v_reg  <= data_i[52];
    end 
    if(N7868) begin
      \nz.mem_1491_sv2v_reg  <= data_i[51];
    end 
    if(N7867) begin
      \nz.mem_1490_sv2v_reg  <= data_i[50];
    end 
    if(N7866) begin
      \nz.mem_1489_sv2v_reg  <= data_i[49];
    end 
    if(N7865) begin
      \nz.mem_1488_sv2v_reg  <= data_i[48];
    end 
    if(N7864) begin
      \nz.mem_1487_sv2v_reg  <= data_i[47];
    end 
    if(N7863) begin
      \nz.mem_1486_sv2v_reg  <= data_i[46];
    end 
    if(N7862) begin
      \nz.mem_1485_sv2v_reg  <= data_i[45];
    end 
    if(N7861) begin
      \nz.mem_1484_sv2v_reg  <= data_i[44];
    end 
    if(N7860) begin
      \nz.mem_1483_sv2v_reg  <= data_i[43];
    end 
    if(N7859) begin
      \nz.mem_1482_sv2v_reg  <= data_i[42];
    end 
    if(N7858) begin
      \nz.mem_1481_sv2v_reg  <= data_i[41];
    end 
    if(N7857) begin
      \nz.mem_1480_sv2v_reg  <= data_i[40];
    end 
    if(N7856) begin
      \nz.mem_1479_sv2v_reg  <= data_i[39];
    end 
    if(N7855) begin
      \nz.mem_1478_sv2v_reg  <= data_i[38];
    end 
    if(N7854) begin
      \nz.mem_1477_sv2v_reg  <= data_i[37];
    end 
    if(N7853) begin
      \nz.mem_1476_sv2v_reg  <= data_i[36];
    end 
    if(N7852) begin
      \nz.mem_1475_sv2v_reg  <= data_i[35];
    end 
    if(N7851) begin
      \nz.mem_1474_sv2v_reg  <= data_i[34];
    end 
    if(N7850) begin
      \nz.mem_1473_sv2v_reg  <= data_i[33];
    end 
    if(N7849) begin
      \nz.mem_1472_sv2v_reg  <= data_i[32];
    end 
    if(N7848) begin
      \nz.mem_1471_sv2v_reg  <= data_i[31];
    end 
    if(N7847) begin
      \nz.mem_1470_sv2v_reg  <= data_i[30];
    end 
    if(N7846) begin
      \nz.mem_1469_sv2v_reg  <= data_i[29];
    end 
    if(N7845) begin
      \nz.mem_1468_sv2v_reg  <= data_i[28];
    end 
    if(N7844) begin
      \nz.mem_1467_sv2v_reg  <= data_i[27];
    end 
    if(N7843) begin
      \nz.mem_1466_sv2v_reg  <= data_i[26];
    end 
    if(N7842) begin
      \nz.mem_1465_sv2v_reg  <= data_i[25];
    end 
    if(N7841) begin
      \nz.mem_1464_sv2v_reg  <= data_i[24];
    end 
    if(N7840) begin
      \nz.mem_1463_sv2v_reg  <= data_i[23];
    end 
    if(N7839) begin
      \nz.mem_1462_sv2v_reg  <= data_i[22];
    end 
    if(N7838) begin
      \nz.mem_1461_sv2v_reg  <= data_i[21];
    end 
    if(N7837) begin
      \nz.mem_1460_sv2v_reg  <= data_i[20];
    end 
    if(N7836) begin
      \nz.mem_1459_sv2v_reg  <= data_i[19];
    end 
    if(N7835) begin
      \nz.mem_1458_sv2v_reg  <= data_i[18];
    end 
    if(N7834) begin
      \nz.mem_1457_sv2v_reg  <= data_i[17];
    end 
    if(N7833) begin
      \nz.mem_1456_sv2v_reg  <= data_i[16];
    end 
    if(N7832) begin
      \nz.mem_1455_sv2v_reg  <= data_i[15];
    end 
    if(N7831) begin
      \nz.mem_1454_sv2v_reg  <= data_i[14];
    end 
    if(N7830) begin
      \nz.mem_1453_sv2v_reg  <= data_i[13];
    end 
    if(N7829) begin
      \nz.mem_1452_sv2v_reg  <= data_i[12];
    end 
    if(N7828) begin
      \nz.mem_1451_sv2v_reg  <= data_i[11];
    end 
    if(N7827) begin
      \nz.mem_1450_sv2v_reg  <= data_i[10];
    end 
    if(N7826) begin
      \nz.mem_1449_sv2v_reg  <= data_i[9];
    end 
    if(N7825) begin
      \nz.mem_1448_sv2v_reg  <= data_i[8];
    end 
    if(N7824) begin
      \nz.mem_1447_sv2v_reg  <= data_i[7];
    end 
    if(N7823) begin
      \nz.mem_1446_sv2v_reg  <= data_i[6];
    end 
    if(N7822) begin
      \nz.mem_1445_sv2v_reg  <= data_i[5];
    end 
    if(N7821) begin
      \nz.mem_1444_sv2v_reg  <= data_i[4];
    end 
    if(N7820) begin
      \nz.mem_1443_sv2v_reg  <= data_i[3];
    end 
    if(N7819) begin
      \nz.mem_1442_sv2v_reg  <= data_i[2];
    end 
    if(N7818) begin
      \nz.mem_1441_sv2v_reg  <= data_i[1];
    end 
    if(N7817) begin
      \nz.mem_1440_sv2v_reg  <= data_i[0];
    end 
    if(N7816) begin
      \nz.mem_1439_sv2v_reg  <= data_i[79];
    end 
    if(N7815) begin
      \nz.mem_1438_sv2v_reg  <= data_i[78];
    end 
    if(N7814) begin
      \nz.mem_1437_sv2v_reg  <= data_i[77];
    end 
    if(N7813) begin
      \nz.mem_1436_sv2v_reg  <= data_i[76];
    end 
    if(N7812) begin
      \nz.mem_1435_sv2v_reg  <= data_i[75];
    end 
    if(N7811) begin
      \nz.mem_1434_sv2v_reg  <= data_i[74];
    end 
    if(N7810) begin
      \nz.mem_1433_sv2v_reg  <= data_i[73];
    end 
    if(N7809) begin
      \nz.mem_1432_sv2v_reg  <= data_i[72];
    end 
    if(N7808) begin
      \nz.mem_1431_sv2v_reg  <= data_i[71];
    end 
    if(N7807) begin
      \nz.mem_1430_sv2v_reg  <= data_i[70];
    end 
    if(N7806) begin
      \nz.mem_1429_sv2v_reg  <= data_i[69];
    end 
    if(N7805) begin
      \nz.mem_1428_sv2v_reg  <= data_i[68];
    end 
    if(N7804) begin
      \nz.mem_1427_sv2v_reg  <= data_i[67];
    end 
    if(N7803) begin
      \nz.mem_1426_sv2v_reg  <= data_i[66];
    end 
    if(N7802) begin
      \nz.mem_1425_sv2v_reg  <= data_i[65];
    end 
    if(N7801) begin
      \nz.mem_1424_sv2v_reg  <= data_i[64];
    end 
    if(N7800) begin
      \nz.mem_1423_sv2v_reg  <= data_i[63];
    end 
    if(N7799) begin
      \nz.mem_1422_sv2v_reg  <= data_i[62];
    end 
    if(N7798) begin
      \nz.mem_1421_sv2v_reg  <= data_i[61];
    end 
    if(N7797) begin
      \nz.mem_1420_sv2v_reg  <= data_i[60];
    end 
    if(N7796) begin
      \nz.mem_1419_sv2v_reg  <= data_i[59];
    end 
    if(N7795) begin
      \nz.mem_1418_sv2v_reg  <= data_i[58];
    end 
    if(N7794) begin
      \nz.mem_1417_sv2v_reg  <= data_i[57];
    end 
    if(N7793) begin
      \nz.mem_1416_sv2v_reg  <= data_i[56];
    end 
    if(N7792) begin
      \nz.mem_1415_sv2v_reg  <= data_i[55];
    end 
    if(N7791) begin
      \nz.mem_1414_sv2v_reg  <= data_i[54];
    end 
    if(N7790) begin
      \nz.mem_1413_sv2v_reg  <= data_i[53];
    end 
    if(N7789) begin
      \nz.mem_1412_sv2v_reg  <= data_i[52];
    end 
    if(N7788) begin
      \nz.mem_1411_sv2v_reg  <= data_i[51];
    end 
    if(N7787) begin
      \nz.mem_1410_sv2v_reg  <= data_i[50];
    end 
    if(N7786) begin
      \nz.mem_1409_sv2v_reg  <= data_i[49];
    end 
    if(N7785) begin
      \nz.mem_1408_sv2v_reg  <= data_i[48];
    end 
    if(N7784) begin
      \nz.mem_1407_sv2v_reg  <= data_i[47];
    end 
    if(N7783) begin
      \nz.mem_1406_sv2v_reg  <= data_i[46];
    end 
    if(N7782) begin
      \nz.mem_1405_sv2v_reg  <= data_i[45];
    end 
    if(N7781) begin
      \nz.mem_1404_sv2v_reg  <= data_i[44];
    end 
    if(N7780) begin
      \nz.mem_1403_sv2v_reg  <= data_i[43];
    end 
    if(N7779) begin
      \nz.mem_1402_sv2v_reg  <= data_i[42];
    end 
    if(N7778) begin
      \nz.mem_1401_sv2v_reg  <= data_i[41];
    end 
    if(N7777) begin
      \nz.mem_1400_sv2v_reg  <= data_i[40];
    end 
    if(N7776) begin
      \nz.mem_1399_sv2v_reg  <= data_i[39];
    end 
    if(N7775) begin
      \nz.mem_1398_sv2v_reg  <= data_i[38];
    end 
    if(N7774) begin
      \nz.mem_1397_sv2v_reg  <= data_i[37];
    end 
    if(N7773) begin
      \nz.mem_1396_sv2v_reg  <= data_i[36];
    end 
    if(N7772) begin
      \nz.mem_1395_sv2v_reg  <= data_i[35];
    end 
    if(N7771) begin
      \nz.mem_1394_sv2v_reg  <= data_i[34];
    end 
    if(N7770) begin
      \nz.mem_1393_sv2v_reg  <= data_i[33];
    end 
    if(N7769) begin
      \nz.mem_1392_sv2v_reg  <= data_i[32];
    end 
    if(N7768) begin
      \nz.mem_1391_sv2v_reg  <= data_i[31];
    end 
    if(N7767) begin
      \nz.mem_1390_sv2v_reg  <= data_i[30];
    end 
    if(N7766) begin
      \nz.mem_1389_sv2v_reg  <= data_i[29];
    end 
    if(N7765) begin
      \nz.mem_1388_sv2v_reg  <= data_i[28];
    end 
    if(N7764) begin
      \nz.mem_1387_sv2v_reg  <= data_i[27];
    end 
    if(N7763) begin
      \nz.mem_1386_sv2v_reg  <= data_i[26];
    end 
    if(N7762) begin
      \nz.mem_1385_sv2v_reg  <= data_i[25];
    end 
    if(N7761) begin
      \nz.mem_1384_sv2v_reg  <= data_i[24];
    end 
    if(N7760) begin
      \nz.mem_1383_sv2v_reg  <= data_i[23];
    end 
    if(N7759) begin
      \nz.mem_1382_sv2v_reg  <= data_i[22];
    end 
    if(N7758) begin
      \nz.mem_1381_sv2v_reg  <= data_i[21];
    end 
    if(N7757) begin
      \nz.mem_1380_sv2v_reg  <= data_i[20];
    end 
    if(N7756) begin
      \nz.mem_1379_sv2v_reg  <= data_i[19];
    end 
    if(N7755) begin
      \nz.mem_1378_sv2v_reg  <= data_i[18];
    end 
    if(N7754) begin
      \nz.mem_1377_sv2v_reg  <= data_i[17];
    end 
    if(N7753) begin
      \nz.mem_1376_sv2v_reg  <= data_i[16];
    end 
    if(N7752) begin
      \nz.mem_1375_sv2v_reg  <= data_i[15];
    end 
    if(N7751) begin
      \nz.mem_1374_sv2v_reg  <= data_i[14];
    end 
    if(N7750) begin
      \nz.mem_1373_sv2v_reg  <= data_i[13];
    end 
    if(N7749) begin
      \nz.mem_1372_sv2v_reg  <= data_i[12];
    end 
    if(N7748) begin
      \nz.mem_1371_sv2v_reg  <= data_i[11];
    end 
    if(N7747) begin
      \nz.mem_1370_sv2v_reg  <= data_i[10];
    end 
    if(N7746) begin
      \nz.mem_1369_sv2v_reg  <= data_i[9];
    end 
    if(N7745) begin
      \nz.mem_1368_sv2v_reg  <= data_i[8];
    end 
    if(N7744) begin
      \nz.mem_1367_sv2v_reg  <= data_i[7];
    end 
    if(N7743) begin
      \nz.mem_1366_sv2v_reg  <= data_i[6];
    end 
    if(N7742) begin
      \nz.mem_1365_sv2v_reg  <= data_i[5];
    end 
    if(N7741) begin
      \nz.mem_1364_sv2v_reg  <= data_i[4];
    end 
    if(N7740) begin
      \nz.mem_1363_sv2v_reg  <= data_i[3];
    end 
    if(N7739) begin
      \nz.mem_1362_sv2v_reg  <= data_i[2];
    end 
    if(N7738) begin
      \nz.mem_1361_sv2v_reg  <= data_i[1];
    end 
    if(N7737) begin
      \nz.mem_1360_sv2v_reg  <= data_i[0];
    end 
    if(N7736) begin
      \nz.mem_1359_sv2v_reg  <= data_i[79];
    end 
    if(N7735) begin
      \nz.mem_1358_sv2v_reg  <= data_i[78];
    end 
    if(N7734) begin
      \nz.mem_1357_sv2v_reg  <= data_i[77];
    end 
    if(N7733) begin
      \nz.mem_1356_sv2v_reg  <= data_i[76];
    end 
    if(N7732) begin
      \nz.mem_1355_sv2v_reg  <= data_i[75];
    end 
    if(N7731) begin
      \nz.mem_1354_sv2v_reg  <= data_i[74];
    end 
    if(N7730) begin
      \nz.mem_1353_sv2v_reg  <= data_i[73];
    end 
    if(N7729) begin
      \nz.mem_1352_sv2v_reg  <= data_i[72];
    end 
    if(N7728) begin
      \nz.mem_1351_sv2v_reg  <= data_i[71];
    end 
    if(N7727) begin
      \nz.mem_1350_sv2v_reg  <= data_i[70];
    end 
    if(N7726) begin
      \nz.mem_1349_sv2v_reg  <= data_i[69];
    end 
    if(N7725) begin
      \nz.mem_1348_sv2v_reg  <= data_i[68];
    end 
    if(N7724) begin
      \nz.mem_1347_sv2v_reg  <= data_i[67];
    end 
    if(N7723) begin
      \nz.mem_1346_sv2v_reg  <= data_i[66];
    end 
    if(N7722) begin
      \nz.mem_1345_sv2v_reg  <= data_i[65];
    end 
    if(N7721) begin
      \nz.mem_1344_sv2v_reg  <= data_i[64];
    end 
    if(N7720) begin
      \nz.mem_1343_sv2v_reg  <= data_i[63];
    end 
    if(N7719) begin
      \nz.mem_1342_sv2v_reg  <= data_i[62];
    end 
    if(N7718) begin
      \nz.mem_1341_sv2v_reg  <= data_i[61];
    end 
    if(N7717) begin
      \nz.mem_1340_sv2v_reg  <= data_i[60];
    end 
    if(N7716) begin
      \nz.mem_1339_sv2v_reg  <= data_i[59];
    end 
    if(N7715) begin
      \nz.mem_1338_sv2v_reg  <= data_i[58];
    end 
    if(N7714) begin
      \nz.mem_1337_sv2v_reg  <= data_i[57];
    end 
    if(N7713) begin
      \nz.mem_1336_sv2v_reg  <= data_i[56];
    end 
    if(N7712) begin
      \nz.mem_1335_sv2v_reg  <= data_i[55];
    end 
    if(N7711) begin
      \nz.mem_1334_sv2v_reg  <= data_i[54];
    end 
    if(N7710) begin
      \nz.mem_1333_sv2v_reg  <= data_i[53];
    end 
    if(N7709) begin
      \nz.mem_1332_sv2v_reg  <= data_i[52];
    end 
    if(N7708) begin
      \nz.mem_1331_sv2v_reg  <= data_i[51];
    end 
    if(N7707) begin
      \nz.mem_1330_sv2v_reg  <= data_i[50];
    end 
    if(N7706) begin
      \nz.mem_1329_sv2v_reg  <= data_i[49];
    end 
    if(N7705) begin
      \nz.mem_1328_sv2v_reg  <= data_i[48];
    end 
    if(N7704) begin
      \nz.mem_1327_sv2v_reg  <= data_i[47];
    end 
    if(N7703) begin
      \nz.mem_1326_sv2v_reg  <= data_i[46];
    end 
    if(N7702) begin
      \nz.mem_1325_sv2v_reg  <= data_i[45];
    end 
    if(N7701) begin
      \nz.mem_1324_sv2v_reg  <= data_i[44];
    end 
    if(N7700) begin
      \nz.mem_1323_sv2v_reg  <= data_i[43];
    end 
    if(N7699) begin
      \nz.mem_1322_sv2v_reg  <= data_i[42];
    end 
    if(N7698) begin
      \nz.mem_1321_sv2v_reg  <= data_i[41];
    end 
    if(N7697) begin
      \nz.mem_1320_sv2v_reg  <= data_i[40];
    end 
    if(N7696) begin
      \nz.mem_1319_sv2v_reg  <= data_i[39];
    end 
    if(N7695) begin
      \nz.mem_1318_sv2v_reg  <= data_i[38];
    end 
    if(N7694) begin
      \nz.mem_1317_sv2v_reg  <= data_i[37];
    end 
    if(N7693) begin
      \nz.mem_1316_sv2v_reg  <= data_i[36];
    end 
    if(N7692) begin
      \nz.mem_1315_sv2v_reg  <= data_i[35];
    end 
    if(N7691) begin
      \nz.mem_1314_sv2v_reg  <= data_i[34];
    end 
    if(N7690) begin
      \nz.mem_1313_sv2v_reg  <= data_i[33];
    end 
    if(N7689) begin
      \nz.mem_1312_sv2v_reg  <= data_i[32];
    end 
    if(N7688) begin
      \nz.mem_1311_sv2v_reg  <= data_i[31];
    end 
    if(N7687) begin
      \nz.mem_1310_sv2v_reg  <= data_i[30];
    end 
    if(N7686) begin
      \nz.mem_1309_sv2v_reg  <= data_i[29];
    end 
    if(N7685) begin
      \nz.mem_1308_sv2v_reg  <= data_i[28];
    end 
    if(N7684) begin
      \nz.mem_1307_sv2v_reg  <= data_i[27];
    end 
    if(N7683) begin
      \nz.mem_1306_sv2v_reg  <= data_i[26];
    end 
    if(N7682) begin
      \nz.mem_1305_sv2v_reg  <= data_i[25];
    end 
    if(N7681) begin
      \nz.mem_1304_sv2v_reg  <= data_i[24];
    end 
    if(N7680) begin
      \nz.mem_1303_sv2v_reg  <= data_i[23];
    end 
    if(N7679) begin
      \nz.mem_1302_sv2v_reg  <= data_i[22];
    end 
    if(N7678) begin
      \nz.mem_1301_sv2v_reg  <= data_i[21];
    end 
    if(N7677) begin
      \nz.mem_1300_sv2v_reg  <= data_i[20];
    end 
    if(N7676) begin
      \nz.mem_1299_sv2v_reg  <= data_i[19];
    end 
    if(N7675) begin
      \nz.mem_1298_sv2v_reg  <= data_i[18];
    end 
    if(N7674) begin
      \nz.mem_1297_sv2v_reg  <= data_i[17];
    end 
    if(N7673) begin
      \nz.mem_1296_sv2v_reg  <= data_i[16];
    end 
    if(N7672) begin
      \nz.mem_1295_sv2v_reg  <= data_i[15];
    end 
    if(N7671) begin
      \nz.mem_1294_sv2v_reg  <= data_i[14];
    end 
    if(N7670) begin
      \nz.mem_1293_sv2v_reg  <= data_i[13];
    end 
    if(N7669) begin
      \nz.mem_1292_sv2v_reg  <= data_i[12];
    end 
    if(N7668) begin
      \nz.mem_1291_sv2v_reg  <= data_i[11];
    end 
    if(N7667) begin
      \nz.mem_1290_sv2v_reg  <= data_i[10];
    end 
    if(N7666) begin
      \nz.mem_1289_sv2v_reg  <= data_i[9];
    end 
    if(N7665) begin
      \nz.mem_1288_sv2v_reg  <= data_i[8];
    end 
    if(N7664) begin
      \nz.mem_1287_sv2v_reg  <= data_i[7];
    end 
    if(N7663) begin
      \nz.mem_1286_sv2v_reg  <= data_i[6];
    end 
    if(N7662) begin
      \nz.mem_1285_sv2v_reg  <= data_i[5];
    end 
    if(N7661) begin
      \nz.mem_1284_sv2v_reg  <= data_i[4];
    end 
    if(N7660) begin
      \nz.mem_1283_sv2v_reg  <= data_i[3];
    end 
    if(N7659) begin
      \nz.mem_1282_sv2v_reg  <= data_i[2];
    end 
    if(N7658) begin
      \nz.mem_1281_sv2v_reg  <= data_i[1];
    end 
    if(N7657) begin
      \nz.mem_1280_sv2v_reg  <= data_i[0];
    end 
    if(N7656) begin
      \nz.mem_1279_sv2v_reg  <= data_i[79];
    end 
    if(N7655) begin
      \nz.mem_1278_sv2v_reg  <= data_i[78];
    end 
    if(N7654) begin
      \nz.mem_1277_sv2v_reg  <= data_i[77];
    end 
    if(N7653) begin
      \nz.mem_1276_sv2v_reg  <= data_i[76];
    end 
    if(N7652) begin
      \nz.mem_1275_sv2v_reg  <= data_i[75];
    end 
    if(N7651) begin
      \nz.mem_1274_sv2v_reg  <= data_i[74];
    end 
    if(N7650) begin
      \nz.mem_1273_sv2v_reg  <= data_i[73];
    end 
    if(N7649) begin
      \nz.mem_1272_sv2v_reg  <= data_i[72];
    end 
    if(N7648) begin
      \nz.mem_1271_sv2v_reg  <= data_i[71];
    end 
    if(N7647) begin
      \nz.mem_1270_sv2v_reg  <= data_i[70];
    end 
    if(N7646) begin
      \nz.mem_1269_sv2v_reg  <= data_i[69];
    end 
    if(N7645) begin
      \nz.mem_1268_sv2v_reg  <= data_i[68];
    end 
    if(N7644) begin
      \nz.mem_1267_sv2v_reg  <= data_i[67];
    end 
    if(N7643) begin
      \nz.mem_1266_sv2v_reg  <= data_i[66];
    end 
    if(N7642) begin
      \nz.mem_1265_sv2v_reg  <= data_i[65];
    end 
    if(N7641) begin
      \nz.mem_1264_sv2v_reg  <= data_i[64];
    end 
    if(N7640) begin
      \nz.mem_1263_sv2v_reg  <= data_i[63];
    end 
    if(N7639) begin
      \nz.mem_1262_sv2v_reg  <= data_i[62];
    end 
    if(N7638) begin
      \nz.mem_1261_sv2v_reg  <= data_i[61];
    end 
    if(N7637) begin
      \nz.mem_1260_sv2v_reg  <= data_i[60];
    end 
    if(N7636) begin
      \nz.mem_1259_sv2v_reg  <= data_i[59];
    end 
    if(N7635) begin
      \nz.mem_1258_sv2v_reg  <= data_i[58];
    end 
    if(N7634) begin
      \nz.mem_1257_sv2v_reg  <= data_i[57];
    end 
    if(N7633) begin
      \nz.mem_1256_sv2v_reg  <= data_i[56];
    end 
    if(N7632) begin
      \nz.mem_1255_sv2v_reg  <= data_i[55];
    end 
    if(N7631) begin
      \nz.mem_1254_sv2v_reg  <= data_i[54];
    end 
    if(N7630) begin
      \nz.mem_1253_sv2v_reg  <= data_i[53];
    end 
    if(N7629) begin
      \nz.mem_1252_sv2v_reg  <= data_i[52];
    end 
    if(N7628) begin
      \nz.mem_1251_sv2v_reg  <= data_i[51];
    end 
    if(N7627) begin
      \nz.mem_1250_sv2v_reg  <= data_i[50];
    end 
    if(N7626) begin
      \nz.mem_1249_sv2v_reg  <= data_i[49];
    end 
    if(N7625) begin
      \nz.mem_1248_sv2v_reg  <= data_i[48];
    end 
    if(N7624) begin
      \nz.mem_1247_sv2v_reg  <= data_i[47];
    end 
    if(N7623) begin
      \nz.mem_1246_sv2v_reg  <= data_i[46];
    end 
    if(N7622) begin
      \nz.mem_1245_sv2v_reg  <= data_i[45];
    end 
    if(N7621) begin
      \nz.mem_1244_sv2v_reg  <= data_i[44];
    end 
    if(N7620) begin
      \nz.mem_1243_sv2v_reg  <= data_i[43];
    end 
    if(N7619) begin
      \nz.mem_1242_sv2v_reg  <= data_i[42];
    end 
    if(N7618) begin
      \nz.mem_1241_sv2v_reg  <= data_i[41];
    end 
    if(N7617) begin
      \nz.mem_1240_sv2v_reg  <= data_i[40];
    end 
    if(N7616) begin
      \nz.mem_1239_sv2v_reg  <= data_i[39];
    end 
    if(N7615) begin
      \nz.mem_1238_sv2v_reg  <= data_i[38];
    end 
    if(N7614) begin
      \nz.mem_1237_sv2v_reg  <= data_i[37];
    end 
    if(N7613) begin
      \nz.mem_1236_sv2v_reg  <= data_i[36];
    end 
    if(N7612) begin
      \nz.mem_1235_sv2v_reg  <= data_i[35];
    end 
    if(N7611) begin
      \nz.mem_1234_sv2v_reg  <= data_i[34];
    end 
    if(N7610) begin
      \nz.mem_1233_sv2v_reg  <= data_i[33];
    end 
    if(N7609) begin
      \nz.mem_1232_sv2v_reg  <= data_i[32];
    end 
    if(N7608) begin
      \nz.mem_1231_sv2v_reg  <= data_i[31];
    end 
    if(N7607) begin
      \nz.mem_1230_sv2v_reg  <= data_i[30];
    end 
    if(N7606) begin
      \nz.mem_1229_sv2v_reg  <= data_i[29];
    end 
    if(N7605) begin
      \nz.mem_1228_sv2v_reg  <= data_i[28];
    end 
    if(N7604) begin
      \nz.mem_1227_sv2v_reg  <= data_i[27];
    end 
    if(N7603) begin
      \nz.mem_1226_sv2v_reg  <= data_i[26];
    end 
    if(N7602) begin
      \nz.mem_1225_sv2v_reg  <= data_i[25];
    end 
    if(N7601) begin
      \nz.mem_1224_sv2v_reg  <= data_i[24];
    end 
    if(N7600) begin
      \nz.mem_1223_sv2v_reg  <= data_i[23];
    end 
    if(N7599) begin
      \nz.mem_1222_sv2v_reg  <= data_i[22];
    end 
    if(N7598) begin
      \nz.mem_1221_sv2v_reg  <= data_i[21];
    end 
    if(N7597) begin
      \nz.mem_1220_sv2v_reg  <= data_i[20];
    end 
    if(N7596) begin
      \nz.mem_1219_sv2v_reg  <= data_i[19];
    end 
    if(N7595) begin
      \nz.mem_1218_sv2v_reg  <= data_i[18];
    end 
    if(N7594) begin
      \nz.mem_1217_sv2v_reg  <= data_i[17];
    end 
    if(N7593) begin
      \nz.mem_1216_sv2v_reg  <= data_i[16];
    end 
    if(N7592) begin
      \nz.mem_1215_sv2v_reg  <= data_i[15];
    end 
    if(N7591) begin
      \nz.mem_1214_sv2v_reg  <= data_i[14];
    end 
    if(N7590) begin
      \nz.mem_1213_sv2v_reg  <= data_i[13];
    end 
    if(N7589) begin
      \nz.mem_1212_sv2v_reg  <= data_i[12];
    end 
    if(N7588) begin
      \nz.mem_1211_sv2v_reg  <= data_i[11];
    end 
    if(N7587) begin
      \nz.mem_1210_sv2v_reg  <= data_i[10];
    end 
    if(N7586) begin
      \nz.mem_1209_sv2v_reg  <= data_i[9];
    end 
    if(N7585) begin
      \nz.mem_1208_sv2v_reg  <= data_i[8];
    end 
    if(N7584) begin
      \nz.mem_1207_sv2v_reg  <= data_i[7];
    end 
    if(N7583) begin
      \nz.mem_1206_sv2v_reg  <= data_i[6];
    end 
    if(N7582) begin
      \nz.mem_1205_sv2v_reg  <= data_i[5];
    end 
    if(N7581) begin
      \nz.mem_1204_sv2v_reg  <= data_i[4];
    end 
    if(N7580) begin
      \nz.mem_1203_sv2v_reg  <= data_i[3];
    end 
    if(N7579) begin
      \nz.mem_1202_sv2v_reg  <= data_i[2];
    end 
    if(N7578) begin
      \nz.mem_1201_sv2v_reg  <= data_i[1];
    end 
    if(N7577) begin
      \nz.mem_1200_sv2v_reg  <= data_i[0];
    end 
    if(N7576) begin
      \nz.mem_1199_sv2v_reg  <= data_i[79];
    end 
    if(N7575) begin
      \nz.mem_1198_sv2v_reg  <= data_i[78];
    end 
    if(N7574) begin
      \nz.mem_1197_sv2v_reg  <= data_i[77];
    end 
    if(N7573) begin
      \nz.mem_1196_sv2v_reg  <= data_i[76];
    end 
    if(N7572) begin
      \nz.mem_1195_sv2v_reg  <= data_i[75];
    end 
    if(N7571) begin
      \nz.mem_1194_sv2v_reg  <= data_i[74];
    end 
    if(N7570) begin
      \nz.mem_1193_sv2v_reg  <= data_i[73];
    end 
    if(N7569) begin
      \nz.mem_1192_sv2v_reg  <= data_i[72];
    end 
    if(N7568) begin
      \nz.mem_1191_sv2v_reg  <= data_i[71];
    end 
    if(N7567) begin
      \nz.mem_1190_sv2v_reg  <= data_i[70];
    end 
    if(N7566) begin
      \nz.mem_1189_sv2v_reg  <= data_i[69];
    end 
    if(N7565) begin
      \nz.mem_1188_sv2v_reg  <= data_i[68];
    end 
    if(N7564) begin
      \nz.mem_1187_sv2v_reg  <= data_i[67];
    end 
    if(N7563) begin
      \nz.mem_1186_sv2v_reg  <= data_i[66];
    end 
    if(N7562) begin
      \nz.mem_1185_sv2v_reg  <= data_i[65];
    end 
    if(N7561) begin
      \nz.mem_1184_sv2v_reg  <= data_i[64];
    end 
    if(N7560) begin
      \nz.mem_1183_sv2v_reg  <= data_i[63];
    end 
    if(N7559) begin
      \nz.mem_1182_sv2v_reg  <= data_i[62];
    end 
    if(N7558) begin
      \nz.mem_1181_sv2v_reg  <= data_i[61];
    end 
    if(N7557) begin
      \nz.mem_1180_sv2v_reg  <= data_i[60];
    end 
    if(N7556) begin
      \nz.mem_1179_sv2v_reg  <= data_i[59];
    end 
    if(N7555) begin
      \nz.mem_1178_sv2v_reg  <= data_i[58];
    end 
    if(N7554) begin
      \nz.mem_1177_sv2v_reg  <= data_i[57];
    end 
    if(N7553) begin
      \nz.mem_1176_sv2v_reg  <= data_i[56];
    end 
    if(N7552) begin
      \nz.mem_1175_sv2v_reg  <= data_i[55];
    end 
    if(N7551) begin
      \nz.mem_1174_sv2v_reg  <= data_i[54];
    end 
    if(N7550) begin
      \nz.mem_1173_sv2v_reg  <= data_i[53];
    end 
    if(N7549) begin
      \nz.mem_1172_sv2v_reg  <= data_i[52];
    end 
    if(N7548) begin
      \nz.mem_1171_sv2v_reg  <= data_i[51];
    end 
    if(N7547) begin
      \nz.mem_1170_sv2v_reg  <= data_i[50];
    end 
    if(N7546) begin
      \nz.mem_1169_sv2v_reg  <= data_i[49];
    end 
    if(N7545) begin
      \nz.mem_1168_sv2v_reg  <= data_i[48];
    end 
    if(N7544) begin
      \nz.mem_1167_sv2v_reg  <= data_i[47];
    end 
    if(N7543) begin
      \nz.mem_1166_sv2v_reg  <= data_i[46];
    end 
    if(N7542) begin
      \nz.mem_1165_sv2v_reg  <= data_i[45];
    end 
    if(N7541) begin
      \nz.mem_1164_sv2v_reg  <= data_i[44];
    end 
    if(N7540) begin
      \nz.mem_1163_sv2v_reg  <= data_i[43];
    end 
    if(N7539) begin
      \nz.mem_1162_sv2v_reg  <= data_i[42];
    end 
    if(N7538) begin
      \nz.mem_1161_sv2v_reg  <= data_i[41];
    end 
    if(N7537) begin
      \nz.mem_1160_sv2v_reg  <= data_i[40];
    end 
    if(N7536) begin
      \nz.mem_1159_sv2v_reg  <= data_i[39];
    end 
    if(N7535) begin
      \nz.mem_1158_sv2v_reg  <= data_i[38];
    end 
    if(N7534) begin
      \nz.mem_1157_sv2v_reg  <= data_i[37];
    end 
    if(N7533) begin
      \nz.mem_1156_sv2v_reg  <= data_i[36];
    end 
    if(N7532) begin
      \nz.mem_1155_sv2v_reg  <= data_i[35];
    end 
    if(N7531) begin
      \nz.mem_1154_sv2v_reg  <= data_i[34];
    end 
    if(N7530) begin
      \nz.mem_1153_sv2v_reg  <= data_i[33];
    end 
    if(N7529) begin
      \nz.mem_1152_sv2v_reg  <= data_i[32];
    end 
    if(N7528) begin
      \nz.mem_1151_sv2v_reg  <= data_i[31];
    end 
    if(N7527) begin
      \nz.mem_1150_sv2v_reg  <= data_i[30];
    end 
    if(N7526) begin
      \nz.mem_1149_sv2v_reg  <= data_i[29];
    end 
    if(N7525) begin
      \nz.mem_1148_sv2v_reg  <= data_i[28];
    end 
    if(N7524) begin
      \nz.mem_1147_sv2v_reg  <= data_i[27];
    end 
    if(N7523) begin
      \nz.mem_1146_sv2v_reg  <= data_i[26];
    end 
    if(N7522) begin
      \nz.mem_1145_sv2v_reg  <= data_i[25];
    end 
    if(N7521) begin
      \nz.mem_1144_sv2v_reg  <= data_i[24];
    end 
    if(N7520) begin
      \nz.mem_1143_sv2v_reg  <= data_i[23];
    end 
    if(N7519) begin
      \nz.mem_1142_sv2v_reg  <= data_i[22];
    end 
    if(N7518) begin
      \nz.mem_1141_sv2v_reg  <= data_i[21];
    end 
    if(N7517) begin
      \nz.mem_1140_sv2v_reg  <= data_i[20];
    end 
    if(N7516) begin
      \nz.mem_1139_sv2v_reg  <= data_i[19];
    end 
    if(N7515) begin
      \nz.mem_1138_sv2v_reg  <= data_i[18];
    end 
    if(N7514) begin
      \nz.mem_1137_sv2v_reg  <= data_i[17];
    end 
    if(N7513) begin
      \nz.mem_1136_sv2v_reg  <= data_i[16];
    end 
    if(N7512) begin
      \nz.mem_1135_sv2v_reg  <= data_i[15];
    end 
    if(N7511) begin
      \nz.mem_1134_sv2v_reg  <= data_i[14];
    end 
    if(N7510) begin
      \nz.mem_1133_sv2v_reg  <= data_i[13];
    end 
    if(N7509) begin
      \nz.mem_1132_sv2v_reg  <= data_i[12];
    end 
    if(N7508) begin
      \nz.mem_1131_sv2v_reg  <= data_i[11];
    end 
    if(N7507) begin
      \nz.mem_1130_sv2v_reg  <= data_i[10];
    end 
    if(N7506) begin
      \nz.mem_1129_sv2v_reg  <= data_i[9];
    end 
    if(N7505) begin
      \nz.mem_1128_sv2v_reg  <= data_i[8];
    end 
    if(N7504) begin
      \nz.mem_1127_sv2v_reg  <= data_i[7];
    end 
    if(N7503) begin
      \nz.mem_1126_sv2v_reg  <= data_i[6];
    end 
    if(N7502) begin
      \nz.mem_1125_sv2v_reg  <= data_i[5];
    end 
    if(N7501) begin
      \nz.mem_1124_sv2v_reg  <= data_i[4];
    end 
    if(N7500) begin
      \nz.mem_1123_sv2v_reg  <= data_i[3];
    end 
    if(N7499) begin
      \nz.mem_1122_sv2v_reg  <= data_i[2];
    end 
    if(N7498) begin
      \nz.mem_1121_sv2v_reg  <= data_i[1];
    end 
    if(N7497) begin
      \nz.mem_1120_sv2v_reg  <= data_i[0];
    end 
    if(N7496) begin
      \nz.mem_1119_sv2v_reg  <= data_i[79];
    end 
    if(N7495) begin
      \nz.mem_1118_sv2v_reg  <= data_i[78];
    end 
    if(N7494) begin
      \nz.mem_1117_sv2v_reg  <= data_i[77];
    end 
    if(N7493) begin
      \nz.mem_1116_sv2v_reg  <= data_i[76];
    end 
    if(N7492) begin
      \nz.mem_1115_sv2v_reg  <= data_i[75];
    end 
    if(N7491) begin
      \nz.mem_1114_sv2v_reg  <= data_i[74];
    end 
    if(N7490) begin
      \nz.mem_1113_sv2v_reg  <= data_i[73];
    end 
    if(N7489) begin
      \nz.mem_1112_sv2v_reg  <= data_i[72];
    end 
    if(N7488) begin
      \nz.mem_1111_sv2v_reg  <= data_i[71];
    end 
    if(N7487) begin
      \nz.mem_1110_sv2v_reg  <= data_i[70];
    end 
    if(N7486) begin
      \nz.mem_1109_sv2v_reg  <= data_i[69];
    end 
    if(N7485) begin
      \nz.mem_1108_sv2v_reg  <= data_i[68];
    end 
    if(N7484) begin
      \nz.mem_1107_sv2v_reg  <= data_i[67];
    end 
    if(N7483) begin
      \nz.mem_1106_sv2v_reg  <= data_i[66];
    end 
    if(N7482) begin
      \nz.mem_1105_sv2v_reg  <= data_i[65];
    end 
    if(N7481) begin
      \nz.mem_1104_sv2v_reg  <= data_i[64];
    end 
    if(N7480) begin
      \nz.mem_1103_sv2v_reg  <= data_i[63];
    end 
    if(N7479) begin
      \nz.mem_1102_sv2v_reg  <= data_i[62];
    end 
    if(N7478) begin
      \nz.mem_1101_sv2v_reg  <= data_i[61];
    end 
    if(N7477) begin
      \nz.mem_1100_sv2v_reg  <= data_i[60];
    end 
    if(N7476) begin
      \nz.mem_1099_sv2v_reg  <= data_i[59];
    end 
    if(N7475) begin
      \nz.mem_1098_sv2v_reg  <= data_i[58];
    end 
    if(N7474) begin
      \nz.mem_1097_sv2v_reg  <= data_i[57];
    end 
    if(N7473) begin
      \nz.mem_1096_sv2v_reg  <= data_i[56];
    end 
    if(N7472) begin
      \nz.mem_1095_sv2v_reg  <= data_i[55];
    end 
    if(N7471) begin
      \nz.mem_1094_sv2v_reg  <= data_i[54];
    end 
    if(N7470) begin
      \nz.mem_1093_sv2v_reg  <= data_i[53];
    end 
    if(N7469) begin
      \nz.mem_1092_sv2v_reg  <= data_i[52];
    end 
    if(N7468) begin
      \nz.mem_1091_sv2v_reg  <= data_i[51];
    end 
    if(N7467) begin
      \nz.mem_1090_sv2v_reg  <= data_i[50];
    end 
    if(N7466) begin
      \nz.mem_1089_sv2v_reg  <= data_i[49];
    end 
    if(N7465) begin
      \nz.mem_1088_sv2v_reg  <= data_i[48];
    end 
    if(N7464) begin
      \nz.mem_1087_sv2v_reg  <= data_i[47];
    end 
    if(N7463) begin
      \nz.mem_1086_sv2v_reg  <= data_i[46];
    end 
    if(N7462) begin
      \nz.mem_1085_sv2v_reg  <= data_i[45];
    end 
    if(N7461) begin
      \nz.mem_1084_sv2v_reg  <= data_i[44];
    end 
    if(N7460) begin
      \nz.mem_1083_sv2v_reg  <= data_i[43];
    end 
    if(N7459) begin
      \nz.mem_1082_sv2v_reg  <= data_i[42];
    end 
    if(N7458) begin
      \nz.mem_1081_sv2v_reg  <= data_i[41];
    end 
    if(N7457) begin
      \nz.mem_1080_sv2v_reg  <= data_i[40];
    end 
    if(N7456) begin
      \nz.mem_1079_sv2v_reg  <= data_i[39];
    end 
    if(N7455) begin
      \nz.mem_1078_sv2v_reg  <= data_i[38];
    end 
    if(N7454) begin
      \nz.mem_1077_sv2v_reg  <= data_i[37];
    end 
    if(N7453) begin
      \nz.mem_1076_sv2v_reg  <= data_i[36];
    end 
    if(N7452) begin
      \nz.mem_1075_sv2v_reg  <= data_i[35];
    end 
    if(N7451) begin
      \nz.mem_1074_sv2v_reg  <= data_i[34];
    end 
    if(N7450) begin
      \nz.mem_1073_sv2v_reg  <= data_i[33];
    end 
    if(N7449) begin
      \nz.mem_1072_sv2v_reg  <= data_i[32];
    end 
    if(N7448) begin
      \nz.mem_1071_sv2v_reg  <= data_i[31];
    end 
    if(N7447) begin
      \nz.mem_1070_sv2v_reg  <= data_i[30];
    end 
    if(N7446) begin
      \nz.mem_1069_sv2v_reg  <= data_i[29];
    end 
    if(N7445) begin
      \nz.mem_1068_sv2v_reg  <= data_i[28];
    end 
    if(N7444) begin
      \nz.mem_1067_sv2v_reg  <= data_i[27];
    end 
    if(N7443) begin
      \nz.mem_1066_sv2v_reg  <= data_i[26];
    end 
    if(N7442) begin
      \nz.mem_1065_sv2v_reg  <= data_i[25];
    end 
    if(N7441) begin
      \nz.mem_1064_sv2v_reg  <= data_i[24];
    end 
    if(N7440) begin
      \nz.mem_1063_sv2v_reg  <= data_i[23];
    end 
    if(N7439) begin
      \nz.mem_1062_sv2v_reg  <= data_i[22];
    end 
    if(N7438) begin
      \nz.mem_1061_sv2v_reg  <= data_i[21];
    end 
    if(N7437) begin
      \nz.mem_1060_sv2v_reg  <= data_i[20];
    end 
    if(N7436) begin
      \nz.mem_1059_sv2v_reg  <= data_i[19];
    end 
    if(N7435) begin
      \nz.mem_1058_sv2v_reg  <= data_i[18];
    end 
    if(N7434) begin
      \nz.mem_1057_sv2v_reg  <= data_i[17];
    end 
    if(N7433) begin
      \nz.mem_1056_sv2v_reg  <= data_i[16];
    end 
    if(N7432) begin
      \nz.mem_1055_sv2v_reg  <= data_i[15];
    end 
    if(N7431) begin
      \nz.mem_1054_sv2v_reg  <= data_i[14];
    end 
    if(N7430) begin
      \nz.mem_1053_sv2v_reg  <= data_i[13];
    end 
    if(N7429) begin
      \nz.mem_1052_sv2v_reg  <= data_i[12];
    end 
    if(N7428) begin
      \nz.mem_1051_sv2v_reg  <= data_i[11];
    end 
    if(N7427) begin
      \nz.mem_1050_sv2v_reg  <= data_i[10];
    end 
    if(N7426) begin
      \nz.mem_1049_sv2v_reg  <= data_i[9];
    end 
    if(N7425) begin
      \nz.mem_1048_sv2v_reg  <= data_i[8];
    end 
    if(N7424) begin
      \nz.mem_1047_sv2v_reg  <= data_i[7];
    end 
    if(N7423) begin
      \nz.mem_1046_sv2v_reg  <= data_i[6];
    end 
    if(N7422) begin
      \nz.mem_1045_sv2v_reg  <= data_i[5];
    end 
    if(N7421) begin
      \nz.mem_1044_sv2v_reg  <= data_i[4];
    end 
    if(N7420) begin
      \nz.mem_1043_sv2v_reg  <= data_i[3];
    end 
    if(N7419) begin
      \nz.mem_1042_sv2v_reg  <= data_i[2];
    end 
    if(N7418) begin
      \nz.mem_1041_sv2v_reg  <= data_i[1];
    end 
    if(N7417) begin
      \nz.mem_1040_sv2v_reg  <= data_i[0];
    end 
    if(N7416) begin
      \nz.mem_1039_sv2v_reg  <= data_i[79];
    end 
    if(N7415) begin
      \nz.mem_1038_sv2v_reg  <= data_i[78];
    end 
    if(N7414) begin
      \nz.mem_1037_sv2v_reg  <= data_i[77];
    end 
    if(N7413) begin
      \nz.mem_1036_sv2v_reg  <= data_i[76];
    end 
    if(N7412) begin
      \nz.mem_1035_sv2v_reg  <= data_i[75];
    end 
    if(N7411) begin
      \nz.mem_1034_sv2v_reg  <= data_i[74];
    end 
    if(N7410) begin
      \nz.mem_1033_sv2v_reg  <= data_i[73];
    end 
    if(N7409) begin
      \nz.mem_1032_sv2v_reg  <= data_i[72];
    end 
    if(N7408) begin
      \nz.mem_1031_sv2v_reg  <= data_i[71];
    end 
    if(N7407) begin
      \nz.mem_1030_sv2v_reg  <= data_i[70];
    end 
    if(N7406) begin
      \nz.mem_1029_sv2v_reg  <= data_i[69];
    end 
    if(N7405) begin
      \nz.mem_1028_sv2v_reg  <= data_i[68];
    end 
    if(N7404) begin
      \nz.mem_1027_sv2v_reg  <= data_i[67];
    end 
    if(N7403) begin
      \nz.mem_1026_sv2v_reg  <= data_i[66];
    end 
    if(N7402) begin
      \nz.mem_1025_sv2v_reg  <= data_i[65];
    end 
    if(N7401) begin
      \nz.mem_1024_sv2v_reg  <= data_i[64];
    end 
    if(N7400) begin
      \nz.mem_1023_sv2v_reg  <= data_i[63];
    end 
    if(N7399) begin
      \nz.mem_1022_sv2v_reg  <= data_i[62];
    end 
    if(N7398) begin
      \nz.mem_1021_sv2v_reg  <= data_i[61];
    end 
    if(N7397) begin
      \nz.mem_1020_sv2v_reg  <= data_i[60];
    end 
    if(N7396) begin
      \nz.mem_1019_sv2v_reg  <= data_i[59];
    end 
    if(N7395) begin
      \nz.mem_1018_sv2v_reg  <= data_i[58];
    end 
    if(N7394) begin
      \nz.mem_1017_sv2v_reg  <= data_i[57];
    end 
    if(N7393) begin
      \nz.mem_1016_sv2v_reg  <= data_i[56];
    end 
    if(N7392) begin
      \nz.mem_1015_sv2v_reg  <= data_i[55];
    end 
    if(N7391) begin
      \nz.mem_1014_sv2v_reg  <= data_i[54];
    end 
    if(N7390) begin
      \nz.mem_1013_sv2v_reg  <= data_i[53];
    end 
    if(N7389) begin
      \nz.mem_1012_sv2v_reg  <= data_i[52];
    end 
    if(N7388) begin
      \nz.mem_1011_sv2v_reg  <= data_i[51];
    end 
    if(N7387) begin
      \nz.mem_1010_sv2v_reg  <= data_i[50];
    end 
    if(N7386) begin
      \nz.mem_1009_sv2v_reg  <= data_i[49];
    end 
    if(N7385) begin
      \nz.mem_1008_sv2v_reg  <= data_i[48];
    end 
    if(N7384) begin
      \nz.mem_1007_sv2v_reg  <= data_i[47];
    end 
    if(N7383) begin
      \nz.mem_1006_sv2v_reg  <= data_i[46];
    end 
    if(N7382) begin
      \nz.mem_1005_sv2v_reg  <= data_i[45];
    end 
    if(N7381) begin
      \nz.mem_1004_sv2v_reg  <= data_i[44];
    end 
    if(N7380) begin
      \nz.mem_1003_sv2v_reg  <= data_i[43];
    end 
    if(N7379) begin
      \nz.mem_1002_sv2v_reg  <= data_i[42];
    end 
    if(N7378) begin
      \nz.mem_1001_sv2v_reg  <= data_i[41];
    end 
    if(N7377) begin
      \nz.mem_1000_sv2v_reg  <= data_i[40];
    end 
    if(N7376) begin
      \nz.mem_999_sv2v_reg  <= data_i[39];
    end 
    if(N7375) begin
      \nz.mem_998_sv2v_reg  <= data_i[38];
    end 
    if(N7374) begin
      \nz.mem_997_sv2v_reg  <= data_i[37];
    end 
    if(N7373) begin
      \nz.mem_996_sv2v_reg  <= data_i[36];
    end 
    if(N7372) begin
      \nz.mem_995_sv2v_reg  <= data_i[35];
    end 
    if(N7371) begin
      \nz.mem_994_sv2v_reg  <= data_i[34];
    end 
    if(N7370) begin
      \nz.mem_993_sv2v_reg  <= data_i[33];
    end 
    if(N7369) begin
      \nz.mem_992_sv2v_reg  <= data_i[32];
    end 
    if(N7368) begin
      \nz.mem_991_sv2v_reg  <= data_i[31];
    end 
    if(N7367) begin
      \nz.mem_990_sv2v_reg  <= data_i[30];
    end 
    if(N7366) begin
      \nz.mem_989_sv2v_reg  <= data_i[29];
    end 
    if(N7365) begin
      \nz.mem_988_sv2v_reg  <= data_i[28];
    end 
    if(N7364) begin
      \nz.mem_987_sv2v_reg  <= data_i[27];
    end 
    if(N7363) begin
      \nz.mem_986_sv2v_reg  <= data_i[26];
    end 
    if(N7362) begin
      \nz.mem_985_sv2v_reg  <= data_i[25];
    end 
    if(N7361) begin
      \nz.mem_984_sv2v_reg  <= data_i[24];
    end 
    if(N7360) begin
      \nz.mem_983_sv2v_reg  <= data_i[23];
    end 
    if(N7359) begin
      \nz.mem_982_sv2v_reg  <= data_i[22];
    end 
    if(N7358) begin
      \nz.mem_981_sv2v_reg  <= data_i[21];
    end 
    if(N7357) begin
      \nz.mem_980_sv2v_reg  <= data_i[20];
    end 
    if(N7356) begin
      \nz.mem_979_sv2v_reg  <= data_i[19];
    end 
    if(N7355) begin
      \nz.mem_978_sv2v_reg  <= data_i[18];
    end 
    if(N7354) begin
      \nz.mem_977_sv2v_reg  <= data_i[17];
    end 
    if(N7353) begin
      \nz.mem_976_sv2v_reg  <= data_i[16];
    end 
    if(N7352) begin
      \nz.mem_975_sv2v_reg  <= data_i[15];
    end 
    if(N7351) begin
      \nz.mem_974_sv2v_reg  <= data_i[14];
    end 
    if(N7350) begin
      \nz.mem_973_sv2v_reg  <= data_i[13];
    end 
    if(N7349) begin
      \nz.mem_972_sv2v_reg  <= data_i[12];
    end 
    if(N7348) begin
      \nz.mem_971_sv2v_reg  <= data_i[11];
    end 
    if(N7347) begin
      \nz.mem_970_sv2v_reg  <= data_i[10];
    end 
    if(N7346) begin
      \nz.mem_969_sv2v_reg  <= data_i[9];
    end 
    if(N7345) begin
      \nz.mem_968_sv2v_reg  <= data_i[8];
    end 
    if(N7344) begin
      \nz.mem_967_sv2v_reg  <= data_i[7];
    end 
    if(N7343) begin
      \nz.mem_966_sv2v_reg  <= data_i[6];
    end 
    if(N7342) begin
      \nz.mem_965_sv2v_reg  <= data_i[5];
    end 
    if(N7341) begin
      \nz.mem_964_sv2v_reg  <= data_i[4];
    end 
    if(N7340) begin
      \nz.mem_963_sv2v_reg  <= data_i[3];
    end 
    if(N7339) begin
      \nz.mem_962_sv2v_reg  <= data_i[2];
    end 
    if(N7338) begin
      \nz.mem_961_sv2v_reg  <= data_i[1];
    end 
    if(N7337) begin
      \nz.mem_960_sv2v_reg  <= data_i[0];
    end 
    if(N7336) begin
      \nz.mem_959_sv2v_reg  <= data_i[79];
    end 
    if(N7335) begin
      \nz.mem_958_sv2v_reg  <= data_i[78];
    end 
    if(N7334) begin
      \nz.mem_957_sv2v_reg  <= data_i[77];
    end 
    if(N7333) begin
      \nz.mem_956_sv2v_reg  <= data_i[76];
    end 
    if(N7332) begin
      \nz.mem_955_sv2v_reg  <= data_i[75];
    end 
    if(N7331) begin
      \nz.mem_954_sv2v_reg  <= data_i[74];
    end 
    if(N7330) begin
      \nz.mem_953_sv2v_reg  <= data_i[73];
    end 
    if(N7329) begin
      \nz.mem_952_sv2v_reg  <= data_i[72];
    end 
    if(N7328) begin
      \nz.mem_951_sv2v_reg  <= data_i[71];
    end 
    if(N7327) begin
      \nz.mem_950_sv2v_reg  <= data_i[70];
    end 
    if(N7326) begin
      \nz.mem_949_sv2v_reg  <= data_i[69];
    end 
    if(N7325) begin
      \nz.mem_948_sv2v_reg  <= data_i[68];
    end 
    if(N7324) begin
      \nz.mem_947_sv2v_reg  <= data_i[67];
    end 
    if(N7323) begin
      \nz.mem_946_sv2v_reg  <= data_i[66];
    end 
    if(N7322) begin
      \nz.mem_945_sv2v_reg  <= data_i[65];
    end 
    if(N7321) begin
      \nz.mem_944_sv2v_reg  <= data_i[64];
    end 
    if(N7320) begin
      \nz.mem_943_sv2v_reg  <= data_i[63];
    end 
    if(N7319) begin
      \nz.mem_942_sv2v_reg  <= data_i[62];
    end 
    if(N7318) begin
      \nz.mem_941_sv2v_reg  <= data_i[61];
    end 
    if(N7317) begin
      \nz.mem_940_sv2v_reg  <= data_i[60];
    end 
    if(N7316) begin
      \nz.mem_939_sv2v_reg  <= data_i[59];
    end 
    if(N7315) begin
      \nz.mem_938_sv2v_reg  <= data_i[58];
    end 
    if(N7314) begin
      \nz.mem_937_sv2v_reg  <= data_i[57];
    end 
    if(N7313) begin
      \nz.mem_936_sv2v_reg  <= data_i[56];
    end 
    if(N7312) begin
      \nz.mem_935_sv2v_reg  <= data_i[55];
    end 
    if(N7311) begin
      \nz.mem_934_sv2v_reg  <= data_i[54];
    end 
    if(N7310) begin
      \nz.mem_933_sv2v_reg  <= data_i[53];
    end 
    if(N7309) begin
      \nz.mem_932_sv2v_reg  <= data_i[52];
    end 
    if(N7308) begin
      \nz.mem_931_sv2v_reg  <= data_i[51];
    end 
    if(N7307) begin
      \nz.mem_930_sv2v_reg  <= data_i[50];
    end 
    if(N7306) begin
      \nz.mem_929_sv2v_reg  <= data_i[49];
    end 
    if(N7305) begin
      \nz.mem_928_sv2v_reg  <= data_i[48];
    end 
    if(N7304) begin
      \nz.mem_927_sv2v_reg  <= data_i[47];
    end 
    if(N7303) begin
      \nz.mem_926_sv2v_reg  <= data_i[46];
    end 
    if(N7302) begin
      \nz.mem_925_sv2v_reg  <= data_i[45];
    end 
    if(N7301) begin
      \nz.mem_924_sv2v_reg  <= data_i[44];
    end 
    if(N7300) begin
      \nz.mem_923_sv2v_reg  <= data_i[43];
    end 
    if(N7299) begin
      \nz.mem_922_sv2v_reg  <= data_i[42];
    end 
    if(N7298) begin
      \nz.mem_921_sv2v_reg  <= data_i[41];
    end 
    if(N7297) begin
      \nz.mem_920_sv2v_reg  <= data_i[40];
    end 
    if(N7296) begin
      \nz.mem_919_sv2v_reg  <= data_i[39];
    end 
    if(N7295) begin
      \nz.mem_918_sv2v_reg  <= data_i[38];
    end 
    if(N7294) begin
      \nz.mem_917_sv2v_reg  <= data_i[37];
    end 
    if(N7293) begin
      \nz.mem_916_sv2v_reg  <= data_i[36];
    end 
    if(N7292) begin
      \nz.mem_915_sv2v_reg  <= data_i[35];
    end 
    if(N7291) begin
      \nz.mem_914_sv2v_reg  <= data_i[34];
    end 
    if(N7290) begin
      \nz.mem_913_sv2v_reg  <= data_i[33];
    end 
    if(N7289) begin
      \nz.mem_912_sv2v_reg  <= data_i[32];
    end 
    if(N7288) begin
      \nz.mem_911_sv2v_reg  <= data_i[31];
    end 
    if(N7287) begin
      \nz.mem_910_sv2v_reg  <= data_i[30];
    end 
    if(N7286) begin
      \nz.mem_909_sv2v_reg  <= data_i[29];
    end 
    if(N7285) begin
      \nz.mem_908_sv2v_reg  <= data_i[28];
    end 
    if(N7284) begin
      \nz.mem_907_sv2v_reg  <= data_i[27];
    end 
    if(N7283) begin
      \nz.mem_906_sv2v_reg  <= data_i[26];
    end 
    if(N7282) begin
      \nz.mem_905_sv2v_reg  <= data_i[25];
    end 
    if(N7281) begin
      \nz.mem_904_sv2v_reg  <= data_i[24];
    end 
    if(N7280) begin
      \nz.mem_903_sv2v_reg  <= data_i[23];
    end 
    if(N7279) begin
      \nz.mem_902_sv2v_reg  <= data_i[22];
    end 
    if(N7278) begin
      \nz.mem_901_sv2v_reg  <= data_i[21];
    end 
    if(N7277) begin
      \nz.mem_900_sv2v_reg  <= data_i[20];
    end 
    if(N7276) begin
      \nz.mem_899_sv2v_reg  <= data_i[19];
    end 
    if(N7275) begin
      \nz.mem_898_sv2v_reg  <= data_i[18];
    end 
    if(N7274) begin
      \nz.mem_897_sv2v_reg  <= data_i[17];
    end 
    if(N7273) begin
      \nz.mem_896_sv2v_reg  <= data_i[16];
    end 
    if(N7272) begin
      \nz.mem_895_sv2v_reg  <= data_i[15];
    end 
    if(N7271) begin
      \nz.mem_894_sv2v_reg  <= data_i[14];
    end 
    if(N7270) begin
      \nz.mem_893_sv2v_reg  <= data_i[13];
    end 
    if(N7269) begin
      \nz.mem_892_sv2v_reg  <= data_i[12];
    end 
    if(N7268) begin
      \nz.mem_891_sv2v_reg  <= data_i[11];
    end 
    if(N7267) begin
      \nz.mem_890_sv2v_reg  <= data_i[10];
    end 
    if(N7266) begin
      \nz.mem_889_sv2v_reg  <= data_i[9];
    end 
    if(N7265) begin
      \nz.mem_888_sv2v_reg  <= data_i[8];
    end 
    if(N7264) begin
      \nz.mem_887_sv2v_reg  <= data_i[7];
    end 
    if(N7263) begin
      \nz.mem_886_sv2v_reg  <= data_i[6];
    end 
    if(N7262) begin
      \nz.mem_885_sv2v_reg  <= data_i[5];
    end 
    if(N7261) begin
      \nz.mem_884_sv2v_reg  <= data_i[4];
    end 
    if(N7260) begin
      \nz.mem_883_sv2v_reg  <= data_i[3];
    end 
    if(N7259) begin
      \nz.mem_882_sv2v_reg  <= data_i[2];
    end 
    if(N7258) begin
      \nz.mem_881_sv2v_reg  <= data_i[1];
    end 
    if(N7257) begin
      \nz.mem_880_sv2v_reg  <= data_i[0];
    end 
    if(N7256) begin
      \nz.mem_879_sv2v_reg  <= data_i[79];
    end 
    if(N7255) begin
      \nz.mem_878_sv2v_reg  <= data_i[78];
    end 
    if(N7254) begin
      \nz.mem_877_sv2v_reg  <= data_i[77];
    end 
    if(N7253) begin
      \nz.mem_876_sv2v_reg  <= data_i[76];
    end 
    if(N7252) begin
      \nz.mem_875_sv2v_reg  <= data_i[75];
    end 
    if(N7251) begin
      \nz.mem_874_sv2v_reg  <= data_i[74];
    end 
    if(N7250) begin
      \nz.mem_873_sv2v_reg  <= data_i[73];
    end 
    if(N7249) begin
      \nz.mem_872_sv2v_reg  <= data_i[72];
    end 
    if(N7248) begin
      \nz.mem_871_sv2v_reg  <= data_i[71];
    end 
    if(N7247) begin
      \nz.mem_870_sv2v_reg  <= data_i[70];
    end 
    if(N7246) begin
      \nz.mem_869_sv2v_reg  <= data_i[69];
    end 
    if(N7245) begin
      \nz.mem_868_sv2v_reg  <= data_i[68];
    end 
    if(N7244) begin
      \nz.mem_867_sv2v_reg  <= data_i[67];
    end 
    if(N7243) begin
      \nz.mem_866_sv2v_reg  <= data_i[66];
    end 
    if(N7242) begin
      \nz.mem_865_sv2v_reg  <= data_i[65];
    end 
    if(N7241) begin
      \nz.mem_864_sv2v_reg  <= data_i[64];
    end 
    if(N7240) begin
      \nz.mem_863_sv2v_reg  <= data_i[63];
    end 
    if(N7239) begin
      \nz.mem_862_sv2v_reg  <= data_i[62];
    end 
    if(N7238) begin
      \nz.mem_861_sv2v_reg  <= data_i[61];
    end 
    if(N7237) begin
      \nz.mem_860_sv2v_reg  <= data_i[60];
    end 
    if(N7236) begin
      \nz.mem_859_sv2v_reg  <= data_i[59];
    end 
    if(N7235) begin
      \nz.mem_858_sv2v_reg  <= data_i[58];
    end 
    if(N7234) begin
      \nz.mem_857_sv2v_reg  <= data_i[57];
    end 
    if(N7233) begin
      \nz.mem_856_sv2v_reg  <= data_i[56];
    end 
    if(N7232) begin
      \nz.mem_855_sv2v_reg  <= data_i[55];
    end 
    if(N7231) begin
      \nz.mem_854_sv2v_reg  <= data_i[54];
    end 
    if(N7230) begin
      \nz.mem_853_sv2v_reg  <= data_i[53];
    end 
    if(N7229) begin
      \nz.mem_852_sv2v_reg  <= data_i[52];
    end 
    if(N7228) begin
      \nz.mem_851_sv2v_reg  <= data_i[51];
    end 
    if(N7227) begin
      \nz.mem_850_sv2v_reg  <= data_i[50];
    end 
    if(N7226) begin
      \nz.mem_849_sv2v_reg  <= data_i[49];
    end 
    if(N7225) begin
      \nz.mem_848_sv2v_reg  <= data_i[48];
    end 
    if(N7224) begin
      \nz.mem_847_sv2v_reg  <= data_i[47];
    end 
    if(N7223) begin
      \nz.mem_846_sv2v_reg  <= data_i[46];
    end 
    if(N7222) begin
      \nz.mem_845_sv2v_reg  <= data_i[45];
    end 
    if(N7221) begin
      \nz.mem_844_sv2v_reg  <= data_i[44];
    end 
    if(N7220) begin
      \nz.mem_843_sv2v_reg  <= data_i[43];
    end 
    if(N7219) begin
      \nz.mem_842_sv2v_reg  <= data_i[42];
    end 
    if(N7218) begin
      \nz.mem_841_sv2v_reg  <= data_i[41];
    end 
    if(N7217) begin
      \nz.mem_840_sv2v_reg  <= data_i[40];
    end 
    if(N7216) begin
      \nz.mem_839_sv2v_reg  <= data_i[39];
    end 
    if(N7215) begin
      \nz.mem_838_sv2v_reg  <= data_i[38];
    end 
    if(N7214) begin
      \nz.mem_837_sv2v_reg  <= data_i[37];
    end 
    if(N7213) begin
      \nz.mem_836_sv2v_reg  <= data_i[36];
    end 
    if(N7212) begin
      \nz.mem_835_sv2v_reg  <= data_i[35];
    end 
    if(N7211) begin
      \nz.mem_834_sv2v_reg  <= data_i[34];
    end 
    if(N7210) begin
      \nz.mem_833_sv2v_reg  <= data_i[33];
    end 
    if(N7209) begin
      \nz.mem_832_sv2v_reg  <= data_i[32];
    end 
    if(N7208) begin
      \nz.mem_831_sv2v_reg  <= data_i[31];
    end 
    if(N7207) begin
      \nz.mem_830_sv2v_reg  <= data_i[30];
    end 
    if(N7206) begin
      \nz.mem_829_sv2v_reg  <= data_i[29];
    end 
    if(N7205) begin
      \nz.mem_828_sv2v_reg  <= data_i[28];
    end 
    if(N7204) begin
      \nz.mem_827_sv2v_reg  <= data_i[27];
    end 
    if(N7203) begin
      \nz.mem_826_sv2v_reg  <= data_i[26];
    end 
    if(N7202) begin
      \nz.mem_825_sv2v_reg  <= data_i[25];
    end 
    if(N7201) begin
      \nz.mem_824_sv2v_reg  <= data_i[24];
    end 
    if(N7200) begin
      \nz.mem_823_sv2v_reg  <= data_i[23];
    end 
    if(N7199) begin
      \nz.mem_822_sv2v_reg  <= data_i[22];
    end 
    if(N7198) begin
      \nz.mem_821_sv2v_reg  <= data_i[21];
    end 
    if(N7197) begin
      \nz.mem_820_sv2v_reg  <= data_i[20];
    end 
    if(N7196) begin
      \nz.mem_819_sv2v_reg  <= data_i[19];
    end 
    if(N7195) begin
      \nz.mem_818_sv2v_reg  <= data_i[18];
    end 
    if(N7194) begin
      \nz.mem_817_sv2v_reg  <= data_i[17];
    end 
    if(N7193) begin
      \nz.mem_816_sv2v_reg  <= data_i[16];
    end 
    if(N7192) begin
      \nz.mem_815_sv2v_reg  <= data_i[15];
    end 
    if(N7191) begin
      \nz.mem_814_sv2v_reg  <= data_i[14];
    end 
    if(N7190) begin
      \nz.mem_813_sv2v_reg  <= data_i[13];
    end 
    if(N7189) begin
      \nz.mem_812_sv2v_reg  <= data_i[12];
    end 
    if(N7188) begin
      \nz.mem_811_sv2v_reg  <= data_i[11];
    end 
    if(N7187) begin
      \nz.mem_810_sv2v_reg  <= data_i[10];
    end 
    if(N7186) begin
      \nz.mem_809_sv2v_reg  <= data_i[9];
    end 
    if(N7185) begin
      \nz.mem_808_sv2v_reg  <= data_i[8];
    end 
    if(N7184) begin
      \nz.mem_807_sv2v_reg  <= data_i[7];
    end 
    if(N7183) begin
      \nz.mem_806_sv2v_reg  <= data_i[6];
    end 
    if(N7182) begin
      \nz.mem_805_sv2v_reg  <= data_i[5];
    end 
    if(N7181) begin
      \nz.mem_804_sv2v_reg  <= data_i[4];
    end 
    if(N7180) begin
      \nz.mem_803_sv2v_reg  <= data_i[3];
    end 
    if(N7179) begin
      \nz.mem_802_sv2v_reg  <= data_i[2];
    end 
    if(N7178) begin
      \nz.mem_801_sv2v_reg  <= data_i[1];
    end 
    if(N7177) begin
      \nz.mem_800_sv2v_reg  <= data_i[0];
    end 
    if(N7176) begin
      \nz.mem_799_sv2v_reg  <= data_i[79];
    end 
    if(N7175) begin
      \nz.mem_798_sv2v_reg  <= data_i[78];
    end 
    if(N7174) begin
      \nz.mem_797_sv2v_reg  <= data_i[77];
    end 
    if(N7173) begin
      \nz.mem_796_sv2v_reg  <= data_i[76];
    end 
    if(N7172) begin
      \nz.mem_795_sv2v_reg  <= data_i[75];
    end 
    if(N7171) begin
      \nz.mem_794_sv2v_reg  <= data_i[74];
    end 
    if(N7170) begin
      \nz.mem_793_sv2v_reg  <= data_i[73];
    end 
    if(N7169) begin
      \nz.mem_792_sv2v_reg  <= data_i[72];
    end 
    if(N7168) begin
      \nz.mem_791_sv2v_reg  <= data_i[71];
    end 
    if(N7167) begin
      \nz.mem_790_sv2v_reg  <= data_i[70];
    end 
    if(N7166) begin
      \nz.mem_789_sv2v_reg  <= data_i[69];
    end 
    if(N7165) begin
      \nz.mem_788_sv2v_reg  <= data_i[68];
    end 
    if(N7164) begin
      \nz.mem_787_sv2v_reg  <= data_i[67];
    end 
    if(N7163) begin
      \nz.mem_786_sv2v_reg  <= data_i[66];
    end 
    if(N7162) begin
      \nz.mem_785_sv2v_reg  <= data_i[65];
    end 
    if(N7161) begin
      \nz.mem_784_sv2v_reg  <= data_i[64];
    end 
    if(N7160) begin
      \nz.mem_783_sv2v_reg  <= data_i[63];
    end 
    if(N7159) begin
      \nz.mem_782_sv2v_reg  <= data_i[62];
    end 
    if(N7158) begin
      \nz.mem_781_sv2v_reg  <= data_i[61];
    end 
    if(N7157) begin
      \nz.mem_780_sv2v_reg  <= data_i[60];
    end 
    if(N7156) begin
      \nz.mem_779_sv2v_reg  <= data_i[59];
    end 
    if(N7155) begin
      \nz.mem_778_sv2v_reg  <= data_i[58];
    end 
    if(N7154) begin
      \nz.mem_777_sv2v_reg  <= data_i[57];
    end 
    if(N7153) begin
      \nz.mem_776_sv2v_reg  <= data_i[56];
    end 
    if(N7152) begin
      \nz.mem_775_sv2v_reg  <= data_i[55];
    end 
    if(N7151) begin
      \nz.mem_774_sv2v_reg  <= data_i[54];
    end 
    if(N7150) begin
      \nz.mem_773_sv2v_reg  <= data_i[53];
    end 
    if(N7149) begin
      \nz.mem_772_sv2v_reg  <= data_i[52];
    end 
    if(N7148) begin
      \nz.mem_771_sv2v_reg  <= data_i[51];
    end 
    if(N7147) begin
      \nz.mem_770_sv2v_reg  <= data_i[50];
    end 
    if(N7146) begin
      \nz.mem_769_sv2v_reg  <= data_i[49];
    end 
    if(N7145) begin
      \nz.mem_768_sv2v_reg  <= data_i[48];
    end 
    if(N7144) begin
      \nz.mem_767_sv2v_reg  <= data_i[47];
    end 
    if(N7143) begin
      \nz.mem_766_sv2v_reg  <= data_i[46];
    end 
    if(N7142) begin
      \nz.mem_765_sv2v_reg  <= data_i[45];
    end 
    if(N7141) begin
      \nz.mem_764_sv2v_reg  <= data_i[44];
    end 
    if(N7140) begin
      \nz.mem_763_sv2v_reg  <= data_i[43];
    end 
    if(N7139) begin
      \nz.mem_762_sv2v_reg  <= data_i[42];
    end 
    if(N7138) begin
      \nz.mem_761_sv2v_reg  <= data_i[41];
    end 
    if(N7137) begin
      \nz.mem_760_sv2v_reg  <= data_i[40];
    end 
    if(N7136) begin
      \nz.mem_759_sv2v_reg  <= data_i[39];
    end 
    if(N7135) begin
      \nz.mem_758_sv2v_reg  <= data_i[38];
    end 
    if(N7134) begin
      \nz.mem_757_sv2v_reg  <= data_i[37];
    end 
    if(N7133) begin
      \nz.mem_756_sv2v_reg  <= data_i[36];
    end 
    if(N7132) begin
      \nz.mem_755_sv2v_reg  <= data_i[35];
    end 
    if(N7131) begin
      \nz.mem_754_sv2v_reg  <= data_i[34];
    end 
    if(N7130) begin
      \nz.mem_753_sv2v_reg  <= data_i[33];
    end 
    if(N7129) begin
      \nz.mem_752_sv2v_reg  <= data_i[32];
    end 
    if(N7128) begin
      \nz.mem_751_sv2v_reg  <= data_i[31];
    end 
    if(N7127) begin
      \nz.mem_750_sv2v_reg  <= data_i[30];
    end 
    if(N7126) begin
      \nz.mem_749_sv2v_reg  <= data_i[29];
    end 
    if(N7125) begin
      \nz.mem_748_sv2v_reg  <= data_i[28];
    end 
    if(N7124) begin
      \nz.mem_747_sv2v_reg  <= data_i[27];
    end 
    if(N7123) begin
      \nz.mem_746_sv2v_reg  <= data_i[26];
    end 
    if(N7122) begin
      \nz.mem_745_sv2v_reg  <= data_i[25];
    end 
    if(N7121) begin
      \nz.mem_744_sv2v_reg  <= data_i[24];
    end 
    if(N7120) begin
      \nz.mem_743_sv2v_reg  <= data_i[23];
    end 
    if(N7119) begin
      \nz.mem_742_sv2v_reg  <= data_i[22];
    end 
    if(N7118) begin
      \nz.mem_741_sv2v_reg  <= data_i[21];
    end 
    if(N7117) begin
      \nz.mem_740_sv2v_reg  <= data_i[20];
    end 
    if(N7116) begin
      \nz.mem_739_sv2v_reg  <= data_i[19];
    end 
    if(N7115) begin
      \nz.mem_738_sv2v_reg  <= data_i[18];
    end 
    if(N7114) begin
      \nz.mem_737_sv2v_reg  <= data_i[17];
    end 
    if(N7113) begin
      \nz.mem_736_sv2v_reg  <= data_i[16];
    end 
    if(N7112) begin
      \nz.mem_735_sv2v_reg  <= data_i[15];
    end 
    if(N7111) begin
      \nz.mem_734_sv2v_reg  <= data_i[14];
    end 
    if(N7110) begin
      \nz.mem_733_sv2v_reg  <= data_i[13];
    end 
    if(N7109) begin
      \nz.mem_732_sv2v_reg  <= data_i[12];
    end 
    if(N7108) begin
      \nz.mem_731_sv2v_reg  <= data_i[11];
    end 
    if(N7107) begin
      \nz.mem_730_sv2v_reg  <= data_i[10];
    end 
    if(N7106) begin
      \nz.mem_729_sv2v_reg  <= data_i[9];
    end 
    if(N7105) begin
      \nz.mem_728_sv2v_reg  <= data_i[8];
    end 
    if(N7104) begin
      \nz.mem_727_sv2v_reg  <= data_i[7];
    end 
    if(N7103) begin
      \nz.mem_726_sv2v_reg  <= data_i[6];
    end 
    if(N7102) begin
      \nz.mem_725_sv2v_reg  <= data_i[5];
    end 
    if(N7101) begin
      \nz.mem_724_sv2v_reg  <= data_i[4];
    end 
    if(N7100) begin
      \nz.mem_723_sv2v_reg  <= data_i[3];
    end 
    if(N7099) begin
      \nz.mem_722_sv2v_reg  <= data_i[2];
    end 
    if(N7098) begin
      \nz.mem_721_sv2v_reg  <= data_i[1];
    end 
    if(N7097) begin
      \nz.mem_720_sv2v_reg  <= data_i[0];
    end 
    if(N7096) begin
      \nz.mem_719_sv2v_reg  <= data_i[79];
    end 
    if(N7095) begin
      \nz.mem_718_sv2v_reg  <= data_i[78];
    end 
    if(N7094) begin
      \nz.mem_717_sv2v_reg  <= data_i[77];
    end 
    if(N7093) begin
      \nz.mem_716_sv2v_reg  <= data_i[76];
    end 
    if(N7092) begin
      \nz.mem_715_sv2v_reg  <= data_i[75];
    end 
    if(N7091) begin
      \nz.mem_714_sv2v_reg  <= data_i[74];
    end 
    if(N7090) begin
      \nz.mem_713_sv2v_reg  <= data_i[73];
    end 
    if(N7089) begin
      \nz.mem_712_sv2v_reg  <= data_i[72];
    end 
    if(N7088) begin
      \nz.mem_711_sv2v_reg  <= data_i[71];
    end 
    if(N7087) begin
      \nz.mem_710_sv2v_reg  <= data_i[70];
    end 
    if(N7086) begin
      \nz.mem_709_sv2v_reg  <= data_i[69];
    end 
    if(N7085) begin
      \nz.mem_708_sv2v_reg  <= data_i[68];
    end 
    if(N7084) begin
      \nz.mem_707_sv2v_reg  <= data_i[67];
    end 
    if(N7083) begin
      \nz.mem_706_sv2v_reg  <= data_i[66];
    end 
    if(N7082) begin
      \nz.mem_705_sv2v_reg  <= data_i[65];
    end 
    if(N7081) begin
      \nz.mem_704_sv2v_reg  <= data_i[64];
    end 
    if(N7080) begin
      \nz.mem_703_sv2v_reg  <= data_i[63];
    end 
    if(N7079) begin
      \nz.mem_702_sv2v_reg  <= data_i[62];
    end 
    if(N7078) begin
      \nz.mem_701_sv2v_reg  <= data_i[61];
    end 
    if(N7077) begin
      \nz.mem_700_sv2v_reg  <= data_i[60];
    end 
    if(N7076) begin
      \nz.mem_699_sv2v_reg  <= data_i[59];
    end 
    if(N7075) begin
      \nz.mem_698_sv2v_reg  <= data_i[58];
    end 
    if(N7074) begin
      \nz.mem_697_sv2v_reg  <= data_i[57];
    end 
    if(N7073) begin
      \nz.mem_696_sv2v_reg  <= data_i[56];
    end 
    if(N7072) begin
      \nz.mem_695_sv2v_reg  <= data_i[55];
    end 
    if(N7071) begin
      \nz.mem_694_sv2v_reg  <= data_i[54];
    end 
    if(N7070) begin
      \nz.mem_693_sv2v_reg  <= data_i[53];
    end 
    if(N7069) begin
      \nz.mem_692_sv2v_reg  <= data_i[52];
    end 
    if(N7068) begin
      \nz.mem_691_sv2v_reg  <= data_i[51];
    end 
    if(N7067) begin
      \nz.mem_690_sv2v_reg  <= data_i[50];
    end 
    if(N7066) begin
      \nz.mem_689_sv2v_reg  <= data_i[49];
    end 
    if(N7065) begin
      \nz.mem_688_sv2v_reg  <= data_i[48];
    end 
    if(N7064) begin
      \nz.mem_687_sv2v_reg  <= data_i[47];
    end 
    if(N7063) begin
      \nz.mem_686_sv2v_reg  <= data_i[46];
    end 
    if(N7062) begin
      \nz.mem_685_sv2v_reg  <= data_i[45];
    end 
    if(N7061) begin
      \nz.mem_684_sv2v_reg  <= data_i[44];
    end 
    if(N7060) begin
      \nz.mem_683_sv2v_reg  <= data_i[43];
    end 
    if(N7059) begin
      \nz.mem_682_sv2v_reg  <= data_i[42];
    end 
    if(N7058) begin
      \nz.mem_681_sv2v_reg  <= data_i[41];
    end 
    if(N7057) begin
      \nz.mem_680_sv2v_reg  <= data_i[40];
    end 
    if(N7056) begin
      \nz.mem_679_sv2v_reg  <= data_i[39];
    end 
    if(N7055) begin
      \nz.mem_678_sv2v_reg  <= data_i[38];
    end 
    if(N7054) begin
      \nz.mem_677_sv2v_reg  <= data_i[37];
    end 
    if(N7053) begin
      \nz.mem_676_sv2v_reg  <= data_i[36];
    end 
    if(N7052) begin
      \nz.mem_675_sv2v_reg  <= data_i[35];
    end 
    if(N7051) begin
      \nz.mem_674_sv2v_reg  <= data_i[34];
    end 
    if(N7050) begin
      \nz.mem_673_sv2v_reg  <= data_i[33];
    end 
    if(N7049) begin
      \nz.mem_672_sv2v_reg  <= data_i[32];
    end 
    if(N7048) begin
      \nz.mem_671_sv2v_reg  <= data_i[31];
    end 
    if(N7047) begin
      \nz.mem_670_sv2v_reg  <= data_i[30];
    end 
    if(N7046) begin
      \nz.mem_669_sv2v_reg  <= data_i[29];
    end 
    if(N7045) begin
      \nz.mem_668_sv2v_reg  <= data_i[28];
    end 
    if(N7044) begin
      \nz.mem_667_sv2v_reg  <= data_i[27];
    end 
    if(N7043) begin
      \nz.mem_666_sv2v_reg  <= data_i[26];
    end 
    if(N7042) begin
      \nz.mem_665_sv2v_reg  <= data_i[25];
    end 
    if(N7041) begin
      \nz.mem_664_sv2v_reg  <= data_i[24];
    end 
    if(N7040) begin
      \nz.mem_663_sv2v_reg  <= data_i[23];
    end 
    if(N7039) begin
      \nz.mem_662_sv2v_reg  <= data_i[22];
    end 
    if(N7038) begin
      \nz.mem_661_sv2v_reg  <= data_i[21];
    end 
    if(N7037) begin
      \nz.mem_660_sv2v_reg  <= data_i[20];
    end 
    if(N7036) begin
      \nz.mem_659_sv2v_reg  <= data_i[19];
    end 
    if(N7035) begin
      \nz.mem_658_sv2v_reg  <= data_i[18];
    end 
    if(N7034) begin
      \nz.mem_657_sv2v_reg  <= data_i[17];
    end 
    if(N7033) begin
      \nz.mem_656_sv2v_reg  <= data_i[16];
    end 
    if(N7032) begin
      \nz.mem_655_sv2v_reg  <= data_i[15];
    end 
    if(N7031) begin
      \nz.mem_654_sv2v_reg  <= data_i[14];
    end 
    if(N7030) begin
      \nz.mem_653_sv2v_reg  <= data_i[13];
    end 
    if(N7029) begin
      \nz.mem_652_sv2v_reg  <= data_i[12];
    end 
    if(N7028) begin
      \nz.mem_651_sv2v_reg  <= data_i[11];
    end 
    if(N7027) begin
      \nz.mem_650_sv2v_reg  <= data_i[10];
    end 
    if(N7026) begin
      \nz.mem_649_sv2v_reg  <= data_i[9];
    end 
    if(N7025) begin
      \nz.mem_648_sv2v_reg  <= data_i[8];
    end 
    if(N7024) begin
      \nz.mem_647_sv2v_reg  <= data_i[7];
    end 
    if(N7023) begin
      \nz.mem_646_sv2v_reg  <= data_i[6];
    end 
    if(N7022) begin
      \nz.mem_645_sv2v_reg  <= data_i[5];
    end 
    if(N7021) begin
      \nz.mem_644_sv2v_reg  <= data_i[4];
    end 
    if(N7020) begin
      \nz.mem_643_sv2v_reg  <= data_i[3];
    end 
    if(N7019) begin
      \nz.mem_642_sv2v_reg  <= data_i[2];
    end 
    if(N7018) begin
      \nz.mem_641_sv2v_reg  <= data_i[1];
    end 
    if(N7017) begin
      \nz.mem_640_sv2v_reg  <= data_i[0];
    end 
    if(N7016) begin
      \nz.mem_639_sv2v_reg  <= data_i[79];
    end 
    if(N7015) begin
      \nz.mem_638_sv2v_reg  <= data_i[78];
    end 
    if(N7014) begin
      \nz.mem_637_sv2v_reg  <= data_i[77];
    end 
    if(N7013) begin
      \nz.mem_636_sv2v_reg  <= data_i[76];
    end 
    if(N7012) begin
      \nz.mem_635_sv2v_reg  <= data_i[75];
    end 
    if(N7011) begin
      \nz.mem_634_sv2v_reg  <= data_i[74];
    end 
    if(N7010) begin
      \nz.mem_633_sv2v_reg  <= data_i[73];
    end 
    if(N7009) begin
      \nz.mem_632_sv2v_reg  <= data_i[72];
    end 
    if(N7008) begin
      \nz.mem_631_sv2v_reg  <= data_i[71];
    end 
    if(N7007) begin
      \nz.mem_630_sv2v_reg  <= data_i[70];
    end 
    if(N7006) begin
      \nz.mem_629_sv2v_reg  <= data_i[69];
    end 
    if(N7005) begin
      \nz.mem_628_sv2v_reg  <= data_i[68];
    end 
    if(N7004) begin
      \nz.mem_627_sv2v_reg  <= data_i[67];
    end 
    if(N7003) begin
      \nz.mem_626_sv2v_reg  <= data_i[66];
    end 
    if(N7002) begin
      \nz.mem_625_sv2v_reg  <= data_i[65];
    end 
    if(N7001) begin
      \nz.mem_624_sv2v_reg  <= data_i[64];
    end 
    if(N7000) begin
      \nz.mem_623_sv2v_reg  <= data_i[63];
    end 
    if(N6999) begin
      \nz.mem_622_sv2v_reg  <= data_i[62];
    end 
    if(N6998) begin
      \nz.mem_621_sv2v_reg  <= data_i[61];
    end 
    if(N6997) begin
      \nz.mem_620_sv2v_reg  <= data_i[60];
    end 
    if(N6996) begin
      \nz.mem_619_sv2v_reg  <= data_i[59];
    end 
    if(N6995) begin
      \nz.mem_618_sv2v_reg  <= data_i[58];
    end 
    if(N6994) begin
      \nz.mem_617_sv2v_reg  <= data_i[57];
    end 
    if(N6993) begin
      \nz.mem_616_sv2v_reg  <= data_i[56];
    end 
    if(N6992) begin
      \nz.mem_615_sv2v_reg  <= data_i[55];
    end 
    if(N6991) begin
      \nz.mem_614_sv2v_reg  <= data_i[54];
    end 
    if(N6990) begin
      \nz.mem_613_sv2v_reg  <= data_i[53];
    end 
    if(N6989) begin
      \nz.mem_612_sv2v_reg  <= data_i[52];
    end 
    if(N6988) begin
      \nz.mem_611_sv2v_reg  <= data_i[51];
    end 
    if(N6987) begin
      \nz.mem_610_sv2v_reg  <= data_i[50];
    end 
    if(N6986) begin
      \nz.mem_609_sv2v_reg  <= data_i[49];
    end 
    if(N6985) begin
      \nz.mem_608_sv2v_reg  <= data_i[48];
    end 
    if(N6984) begin
      \nz.mem_607_sv2v_reg  <= data_i[47];
    end 
    if(N6983) begin
      \nz.mem_606_sv2v_reg  <= data_i[46];
    end 
    if(N6982) begin
      \nz.mem_605_sv2v_reg  <= data_i[45];
    end 
    if(N6981) begin
      \nz.mem_604_sv2v_reg  <= data_i[44];
    end 
    if(N6980) begin
      \nz.mem_603_sv2v_reg  <= data_i[43];
    end 
    if(N6979) begin
      \nz.mem_602_sv2v_reg  <= data_i[42];
    end 
    if(N6978) begin
      \nz.mem_601_sv2v_reg  <= data_i[41];
    end 
    if(N6977) begin
      \nz.mem_600_sv2v_reg  <= data_i[40];
    end 
    if(N6976) begin
      \nz.mem_599_sv2v_reg  <= data_i[39];
    end 
    if(N6975) begin
      \nz.mem_598_sv2v_reg  <= data_i[38];
    end 
    if(N6974) begin
      \nz.mem_597_sv2v_reg  <= data_i[37];
    end 
    if(N6973) begin
      \nz.mem_596_sv2v_reg  <= data_i[36];
    end 
    if(N6972) begin
      \nz.mem_595_sv2v_reg  <= data_i[35];
    end 
    if(N6971) begin
      \nz.mem_594_sv2v_reg  <= data_i[34];
    end 
    if(N6970) begin
      \nz.mem_593_sv2v_reg  <= data_i[33];
    end 
    if(N6969) begin
      \nz.mem_592_sv2v_reg  <= data_i[32];
    end 
    if(N6968) begin
      \nz.mem_591_sv2v_reg  <= data_i[31];
    end 
    if(N6967) begin
      \nz.mem_590_sv2v_reg  <= data_i[30];
    end 
    if(N6966) begin
      \nz.mem_589_sv2v_reg  <= data_i[29];
    end 
    if(N6965) begin
      \nz.mem_588_sv2v_reg  <= data_i[28];
    end 
    if(N6964) begin
      \nz.mem_587_sv2v_reg  <= data_i[27];
    end 
    if(N6963) begin
      \nz.mem_586_sv2v_reg  <= data_i[26];
    end 
    if(N6962) begin
      \nz.mem_585_sv2v_reg  <= data_i[25];
    end 
    if(N6961) begin
      \nz.mem_584_sv2v_reg  <= data_i[24];
    end 
    if(N6960) begin
      \nz.mem_583_sv2v_reg  <= data_i[23];
    end 
    if(N6959) begin
      \nz.mem_582_sv2v_reg  <= data_i[22];
    end 
    if(N6958) begin
      \nz.mem_581_sv2v_reg  <= data_i[21];
    end 
    if(N6957) begin
      \nz.mem_580_sv2v_reg  <= data_i[20];
    end 
    if(N6956) begin
      \nz.mem_579_sv2v_reg  <= data_i[19];
    end 
    if(N6955) begin
      \nz.mem_578_sv2v_reg  <= data_i[18];
    end 
    if(N6954) begin
      \nz.mem_577_sv2v_reg  <= data_i[17];
    end 
    if(N6953) begin
      \nz.mem_576_sv2v_reg  <= data_i[16];
    end 
    if(N6952) begin
      \nz.mem_575_sv2v_reg  <= data_i[15];
    end 
    if(N6951) begin
      \nz.mem_574_sv2v_reg  <= data_i[14];
    end 
    if(N6950) begin
      \nz.mem_573_sv2v_reg  <= data_i[13];
    end 
    if(N6949) begin
      \nz.mem_572_sv2v_reg  <= data_i[12];
    end 
    if(N6948) begin
      \nz.mem_571_sv2v_reg  <= data_i[11];
    end 
    if(N6947) begin
      \nz.mem_570_sv2v_reg  <= data_i[10];
    end 
    if(N6946) begin
      \nz.mem_569_sv2v_reg  <= data_i[9];
    end 
    if(N6945) begin
      \nz.mem_568_sv2v_reg  <= data_i[8];
    end 
    if(N6944) begin
      \nz.mem_567_sv2v_reg  <= data_i[7];
    end 
    if(N6943) begin
      \nz.mem_566_sv2v_reg  <= data_i[6];
    end 
    if(N6942) begin
      \nz.mem_565_sv2v_reg  <= data_i[5];
    end 
    if(N6941) begin
      \nz.mem_564_sv2v_reg  <= data_i[4];
    end 
    if(N6940) begin
      \nz.mem_563_sv2v_reg  <= data_i[3];
    end 
    if(N6939) begin
      \nz.mem_562_sv2v_reg  <= data_i[2];
    end 
    if(N6938) begin
      \nz.mem_561_sv2v_reg  <= data_i[1];
    end 
    if(N6937) begin
      \nz.mem_560_sv2v_reg  <= data_i[0];
    end 
    if(N6936) begin
      \nz.mem_559_sv2v_reg  <= data_i[79];
    end 
    if(N6935) begin
      \nz.mem_558_sv2v_reg  <= data_i[78];
    end 
    if(N6934) begin
      \nz.mem_557_sv2v_reg  <= data_i[77];
    end 
    if(N6933) begin
      \nz.mem_556_sv2v_reg  <= data_i[76];
    end 
    if(N6932) begin
      \nz.mem_555_sv2v_reg  <= data_i[75];
    end 
    if(N6931) begin
      \nz.mem_554_sv2v_reg  <= data_i[74];
    end 
    if(N6930) begin
      \nz.mem_553_sv2v_reg  <= data_i[73];
    end 
    if(N6929) begin
      \nz.mem_552_sv2v_reg  <= data_i[72];
    end 
    if(N6928) begin
      \nz.mem_551_sv2v_reg  <= data_i[71];
    end 
    if(N6927) begin
      \nz.mem_550_sv2v_reg  <= data_i[70];
    end 
    if(N6926) begin
      \nz.mem_549_sv2v_reg  <= data_i[69];
    end 
    if(N6925) begin
      \nz.mem_548_sv2v_reg  <= data_i[68];
    end 
    if(N6924) begin
      \nz.mem_547_sv2v_reg  <= data_i[67];
    end 
    if(N6923) begin
      \nz.mem_546_sv2v_reg  <= data_i[66];
    end 
    if(N6922) begin
      \nz.mem_545_sv2v_reg  <= data_i[65];
    end 
    if(N6921) begin
      \nz.mem_544_sv2v_reg  <= data_i[64];
    end 
    if(N6920) begin
      \nz.mem_543_sv2v_reg  <= data_i[63];
    end 
    if(N6919) begin
      \nz.mem_542_sv2v_reg  <= data_i[62];
    end 
    if(N6918) begin
      \nz.mem_541_sv2v_reg  <= data_i[61];
    end 
    if(N6917) begin
      \nz.mem_540_sv2v_reg  <= data_i[60];
    end 
    if(N6916) begin
      \nz.mem_539_sv2v_reg  <= data_i[59];
    end 
    if(N6915) begin
      \nz.mem_538_sv2v_reg  <= data_i[58];
    end 
    if(N6914) begin
      \nz.mem_537_sv2v_reg  <= data_i[57];
    end 
    if(N6913) begin
      \nz.mem_536_sv2v_reg  <= data_i[56];
    end 
    if(N6912) begin
      \nz.mem_535_sv2v_reg  <= data_i[55];
    end 
    if(N6911) begin
      \nz.mem_534_sv2v_reg  <= data_i[54];
    end 
    if(N6910) begin
      \nz.mem_533_sv2v_reg  <= data_i[53];
    end 
    if(N6909) begin
      \nz.mem_532_sv2v_reg  <= data_i[52];
    end 
    if(N6908) begin
      \nz.mem_531_sv2v_reg  <= data_i[51];
    end 
    if(N6907) begin
      \nz.mem_530_sv2v_reg  <= data_i[50];
    end 
    if(N6906) begin
      \nz.mem_529_sv2v_reg  <= data_i[49];
    end 
    if(N6905) begin
      \nz.mem_528_sv2v_reg  <= data_i[48];
    end 
    if(N6904) begin
      \nz.mem_527_sv2v_reg  <= data_i[47];
    end 
    if(N6903) begin
      \nz.mem_526_sv2v_reg  <= data_i[46];
    end 
    if(N6902) begin
      \nz.mem_525_sv2v_reg  <= data_i[45];
    end 
    if(N6901) begin
      \nz.mem_524_sv2v_reg  <= data_i[44];
    end 
    if(N6900) begin
      \nz.mem_523_sv2v_reg  <= data_i[43];
    end 
    if(N6899) begin
      \nz.mem_522_sv2v_reg  <= data_i[42];
    end 
    if(N6898) begin
      \nz.mem_521_sv2v_reg  <= data_i[41];
    end 
    if(N6897) begin
      \nz.mem_520_sv2v_reg  <= data_i[40];
    end 
    if(N6896) begin
      \nz.mem_519_sv2v_reg  <= data_i[39];
    end 
    if(N6895) begin
      \nz.mem_518_sv2v_reg  <= data_i[38];
    end 
    if(N6894) begin
      \nz.mem_517_sv2v_reg  <= data_i[37];
    end 
    if(N6893) begin
      \nz.mem_516_sv2v_reg  <= data_i[36];
    end 
    if(N6892) begin
      \nz.mem_515_sv2v_reg  <= data_i[35];
    end 
    if(N6891) begin
      \nz.mem_514_sv2v_reg  <= data_i[34];
    end 
    if(N6890) begin
      \nz.mem_513_sv2v_reg  <= data_i[33];
    end 
    if(N6889) begin
      \nz.mem_512_sv2v_reg  <= data_i[32];
    end 
    if(N6888) begin
      \nz.mem_511_sv2v_reg  <= data_i[31];
    end 
    if(N6887) begin
      \nz.mem_510_sv2v_reg  <= data_i[30];
    end 
    if(N6886) begin
      \nz.mem_509_sv2v_reg  <= data_i[29];
    end 
    if(N6885) begin
      \nz.mem_508_sv2v_reg  <= data_i[28];
    end 
    if(N6884) begin
      \nz.mem_507_sv2v_reg  <= data_i[27];
    end 
    if(N6883) begin
      \nz.mem_506_sv2v_reg  <= data_i[26];
    end 
    if(N6882) begin
      \nz.mem_505_sv2v_reg  <= data_i[25];
    end 
    if(N6881) begin
      \nz.mem_504_sv2v_reg  <= data_i[24];
    end 
    if(N6880) begin
      \nz.mem_503_sv2v_reg  <= data_i[23];
    end 
    if(N6879) begin
      \nz.mem_502_sv2v_reg  <= data_i[22];
    end 
    if(N6878) begin
      \nz.mem_501_sv2v_reg  <= data_i[21];
    end 
    if(N6877) begin
      \nz.mem_500_sv2v_reg  <= data_i[20];
    end 
    if(N6876) begin
      \nz.mem_499_sv2v_reg  <= data_i[19];
    end 
    if(N6875) begin
      \nz.mem_498_sv2v_reg  <= data_i[18];
    end 
    if(N6874) begin
      \nz.mem_497_sv2v_reg  <= data_i[17];
    end 
    if(N6873) begin
      \nz.mem_496_sv2v_reg  <= data_i[16];
    end 
    if(N6872) begin
      \nz.mem_495_sv2v_reg  <= data_i[15];
    end 
    if(N6871) begin
      \nz.mem_494_sv2v_reg  <= data_i[14];
    end 
    if(N6870) begin
      \nz.mem_493_sv2v_reg  <= data_i[13];
    end 
    if(N6869) begin
      \nz.mem_492_sv2v_reg  <= data_i[12];
    end 
    if(N6868) begin
      \nz.mem_491_sv2v_reg  <= data_i[11];
    end 
    if(N6867) begin
      \nz.mem_490_sv2v_reg  <= data_i[10];
    end 
    if(N6866) begin
      \nz.mem_489_sv2v_reg  <= data_i[9];
    end 
    if(N6865) begin
      \nz.mem_488_sv2v_reg  <= data_i[8];
    end 
    if(N6864) begin
      \nz.mem_487_sv2v_reg  <= data_i[7];
    end 
    if(N6863) begin
      \nz.mem_486_sv2v_reg  <= data_i[6];
    end 
    if(N6862) begin
      \nz.mem_485_sv2v_reg  <= data_i[5];
    end 
    if(N6861) begin
      \nz.mem_484_sv2v_reg  <= data_i[4];
    end 
    if(N6860) begin
      \nz.mem_483_sv2v_reg  <= data_i[3];
    end 
    if(N6859) begin
      \nz.mem_482_sv2v_reg  <= data_i[2];
    end 
    if(N6858) begin
      \nz.mem_481_sv2v_reg  <= data_i[1];
    end 
    if(N6857) begin
      \nz.mem_480_sv2v_reg  <= data_i[0];
    end 
    if(N6856) begin
      \nz.mem_479_sv2v_reg  <= data_i[79];
    end 
    if(N6855) begin
      \nz.mem_478_sv2v_reg  <= data_i[78];
    end 
    if(N6854) begin
      \nz.mem_477_sv2v_reg  <= data_i[77];
    end 
    if(N6853) begin
      \nz.mem_476_sv2v_reg  <= data_i[76];
    end 
    if(N6852) begin
      \nz.mem_475_sv2v_reg  <= data_i[75];
    end 
    if(N6851) begin
      \nz.mem_474_sv2v_reg  <= data_i[74];
    end 
    if(N6850) begin
      \nz.mem_473_sv2v_reg  <= data_i[73];
    end 
    if(N6849) begin
      \nz.mem_472_sv2v_reg  <= data_i[72];
    end 
    if(N6848) begin
      \nz.mem_471_sv2v_reg  <= data_i[71];
    end 
    if(N6847) begin
      \nz.mem_470_sv2v_reg  <= data_i[70];
    end 
    if(N6846) begin
      \nz.mem_469_sv2v_reg  <= data_i[69];
    end 
    if(N6845) begin
      \nz.mem_468_sv2v_reg  <= data_i[68];
    end 
    if(N6844) begin
      \nz.mem_467_sv2v_reg  <= data_i[67];
    end 
    if(N6843) begin
      \nz.mem_466_sv2v_reg  <= data_i[66];
    end 
    if(N6842) begin
      \nz.mem_465_sv2v_reg  <= data_i[65];
    end 
    if(N6841) begin
      \nz.mem_464_sv2v_reg  <= data_i[64];
    end 
    if(N6840) begin
      \nz.mem_463_sv2v_reg  <= data_i[63];
    end 
    if(N6839) begin
      \nz.mem_462_sv2v_reg  <= data_i[62];
    end 
    if(N6838) begin
      \nz.mem_461_sv2v_reg  <= data_i[61];
    end 
    if(N6837) begin
      \nz.mem_460_sv2v_reg  <= data_i[60];
    end 
    if(N6836) begin
      \nz.mem_459_sv2v_reg  <= data_i[59];
    end 
    if(N6835) begin
      \nz.mem_458_sv2v_reg  <= data_i[58];
    end 
    if(N6834) begin
      \nz.mem_457_sv2v_reg  <= data_i[57];
    end 
    if(N6833) begin
      \nz.mem_456_sv2v_reg  <= data_i[56];
    end 
    if(N6832) begin
      \nz.mem_455_sv2v_reg  <= data_i[55];
    end 
    if(N6831) begin
      \nz.mem_454_sv2v_reg  <= data_i[54];
    end 
    if(N6830) begin
      \nz.mem_453_sv2v_reg  <= data_i[53];
    end 
    if(N6829) begin
      \nz.mem_452_sv2v_reg  <= data_i[52];
    end 
    if(N6828) begin
      \nz.mem_451_sv2v_reg  <= data_i[51];
    end 
    if(N6827) begin
      \nz.mem_450_sv2v_reg  <= data_i[50];
    end 
    if(N6826) begin
      \nz.mem_449_sv2v_reg  <= data_i[49];
    end 
    if(N6825) begin
      \nz.mem_448_sv2v_reg  <= data_i[48];
    end 
    if(N6824) begin
      \nz.mem_447_sv2v_reg  <= data_i[47];
    end 
    if(N6823) begin
      \nz.mem_446_sv2v_reg  <= data_i[46];
    end 
    if(N6822) begin
      \nz.mem_445_sv2v_reg  <= data_i[45];
    end 
    if(N6821) begin
      \nz.mem_444_sv2v_reg  <= data_i[44];
    end 
    if(N6820) begin
      \nz.mem_443_sv2v_reg  <= data_i[43];
    end 
    if(N6819) begin
      \nz.mem_442_sv2v_reg  <= data_i[42];
    end 
    if(N6818) begin
      \nz.mem_441_sv2v_reg  <= data_i[41];
    end 
    if(N6817) begin
      \nz.mem_440_sv2v_reg  <= data_i[40];
    end 
    if(N6816) begin
      \nz.mem_439_sv2v_reg  <= data_i[39];
    end 
    if(N6815) begin
      \nz.mem_438_sv2v_reg  <= data_i[38];
    end 
    if(N6814) begin
      \nz.mem_437_sv2v_reg  <= data_i[37];
    end 
    if(N6813) begin
      \nz.mem_436_sv2v_reg  <= data_i[36];
    end 
    if(N6812) begin
      \nz.mem_435_sv2v_reg  <= data_i[35];
    end 
    if(N6811) begin
      \nz.mem_434_sv2v_reg  <= data_i[34];
    end 
    if(N6810) begin
      \nz.mem_433_sv2v_reg  <= data_i[33];
    end 
    if(N6809) begin
      \nz.mem_432_sv2v_reg  <= data_i[32];
    end 
    if(N6808) begin
      \nz.mem_431_sv2v_reg  <= data_i[31];
    end 
    if(N6807) begin
      \nz.mem_430_sv2v_reg  <= data_i[30];
    end 
    if(N6806) begin
      \nz.mem_429_sv2v_reg  <= data_i[29];
    end 
    if(N6805) begin
      \nz.mem_428_sv2v_reg  <= data_i[28];
    end 
    if(N6804) begin
      \nz.mem_427_sv2v_reg  <= data_i[27];
    end 
    if(N6803) begin
      \nz.mem_426_sv2v_reg  <= data_i[26];
    end 
    if(N6802) begin
      \nz.mem_425_sv2v_reg  <= data_i[25];
    end 
    if(N6801) begin
      \nz.mem_424_sv2v_reg  <= data_i[24];
    end 
    if(N6800) begin
      \nz.mem_423_sv2v_reg  <= data_i[23];
    end 
    if(N6799) begin
      \nz.mem_422_sv2v_reg  <= data_i[22];
    end 
    if(N6798) begin
      \nz.mem_421_sv2v_reg  <= data_i[21];
    end 
    if(N6797) begin
      \nz.mem_420_sv2v_reg  <= data_i[20];
    end 
    if(N6796) begin
      \nz.mem_419_sv2v_reg  <= data_i[19];
    end 
    if(N6795) begin
      \nz.mem_418_sv2v_reg  <= data_i[18];
    end 
    if(N6794) begin
      \nz.mem_417_sv2v_reg  <= data_i[17];
    end 
    if(N6793) begin
      \nz.mem_416_sv2v_reg  <= data_i[16];
    end 
    if(N6792) begin
      \nz.mem_415_sv2v_reg  <= data_i[15];
    end 
    if(N6791) begin
      \nz.mem_414_sv2v_reg  <= data_i[14];
    end 
    if(N6790) begin
      \nz.mem_413_sv2v_reg  <= data_i[13];
    end 
    if(N6789) begin
      \nz.mem_412_sv2v_reg  <= data_i[12];
    end 
    if(N6788) begin
      \nz.mem_411_sv2v_reg  <= data_i[11];
    end 
    if(N6787) begin
      \nz.mem_410_sv2v_reg  <= data_i[10];
    end 
    if(N6786) begin
      \nz.mem_409_sv2v_reg  <= data_i[9];
    end 
    if(N6785) begin
      \nz.mem_408_sv2v_reg  <= data_i[8];
    end 
    if(N6784) begin
      \nz.mem_407_sv2v_reg  <= data_i[7];
    end 
    if(N6783) begin
      \nz.mem_406_sv2v_reg  <= data_i[6];
    end 
    if(N6782) begin
      \nz.mem_405_sv2v_reg  <= data_i[5];
    end 
    if(N6781) begin
      \nz.mem_404_sv2v_reg  <= data_i[4];
    end 
    if(N6780) begin
      \nz.mem_403_sv2v_reg  <= data_i[3];
    end 
    if(N6779) begin
      \nz.mem_402_sv2v_reg  <= data_i[2];
    end 
    if(N6778) begin
      \nz.mem_401_sv2v_reg  <= data_i[1];
    end 
    if(N6777) begin
      \nz.mem_400_sv2v_reg  <= data_i[0];
    end 
    if(N6776) begin
      \nz.mem_399_sv2v_reg  <= data_i[79];
    end 
    if(N6775) begin
      \nz.mem_398_sv2v_reg  <= data_i[78];
    end 
    if(N6774) begin
      \nz.mem_397_sv2v_reg  <= data_i[77];
    end 
    if(N6773) begin
      \nz.mem_396_sv2v_reg  <= data_i[76];
    end 
    if(N6772) begin
      \nz.mem_395_sv2v_reg  <= data_i[75];
    end 
    if(N6771) begin
      \nz.mem_394_sv2v_reg  <= data_i[74];
    end 
    if(N6770) begin
      \nz.mem_393_sv2v_reg  <= data_i[73];
    end 
    if(N6769) begin
      \nz.mem_392_sv2v_reg  <= data_i[72];
    end 
    if(N6768) begin
      \nz.mem_391_sv2v_reg  <= data_i[71];
    end 
    if(N6767) begin
      \nz.mem_390_sv2v_reg  <= data_i[70];
    end 
    if(N6766) begin
      \nz.mem_389_sv2v_reg  <= data_i[69];
    end 
    if(N6765) begin
      \nz.mem_388_sv2v_reg  <= data_i[68];
    end 
    if(N6764) begin
      \nz.mem_387_sv2v_reg  <= data_i[67];
    end 
    if(N6763) begin
      \nz.mem_386_sv2v_reg  <= data_i[66];
    end 
    if(N6762) begin
      \nz.mem_385_sv2v_reg  <= data_i[65];
    end 
    if(N6761) begin
      \nz.mem_384_sv2v_reg  <= data_i[64];
    end 
    if(N6760) begin
      \nz.mem_383_sv2v_reg  <= data_i[63];
    end 
    if(N6759) begin
      \nz.mem_382_sv2v_reg  <= data_i[62];
    end 
    if(N6758) begin
      \nz.mem_381_sv2v_reg  <= data_i[61];
    end 
    if(N6757) begin
      \nz.mem_380_sv2v_reg  <= data_i[60];
    end 
    if(N6756) begin
      \nz.mem_379_sv2v_reg  <= data_i[59];
    end 
    if(N6755) begin
      \nz.mem_378_sv2v_reg  <= data_i[58];
    end 
    if(N6754) begin
      \nz.mem_377_sv2v_reg  <= data_i[57];
    end 
    if(N6753) begin
      \nz.mem_376_sv2v_reg  <= data_i[56];
    end 
    if(N6752) begin
      \nz.mem_375_sv2v_reg  <= data_i[55];
    end 
    if(N6751) begin
      \nz.mem_374_sv2v_reg  <= data_i[54];
    end 
    if(N6750) begin
      \nz.mem_373_sv2v_reg  <= data_i[53];
    end 
    if(N6749) begin
      \nz.mem_372_sv2v_reg  <= data_i[52];
    end 
    if(N6748) begin
      \nz.mem_371_sv2v_reg  <= data_i[51];
    end 
    if(N6747) begin
      \nz.mem_370_sv2v_reg  <= data_i[50];
    end 
    if(N6746) begin
      \nz.mem_369_sv2v_reg  <= data_i[49];
    end 
    if(N6745) begin
      \nz.mem_368_sv2v_reg  <= data_i[48];
    end 
    if(N6744) begin
      \nz.mem_367_sv2v_reg  <= data_i[47];
    end 
    if(N6743) begin
      \nz.mem_366_sv2v_reg  <= data_i[46];
    end 
    if(N6742) begin
      \nz.mem_365_sv2v_reg  <= data_i[45];
    end 
    if(N6741) begin
      \nz.mem_364_sv2v_reg  <= data_i[44];
    end 
    if(N6740) begin
      \nz.mem_363_sv2v_reg  <= data_i[43];
    end 
    if(N6739) begin
      \nz.mem_362_sv2v_reg  <= data_i[42];
    end 
    if(N6738) begin
      \nz.mem_361_sv2v_reg  <= data_i[41];
    end 
    if(N6737) begin
      \nz.mem_360_sv2v_reg  <= data_i[40];
    end 
    if(N6736) begin
      \nz.mem_359_sv2v_reg  <= data_i[39];
    end 
    if(N6735) begin
      \nz.mem_358_sv2v_reg  <= data_i[38];
    end 
    if(N6734) begin
      \nz.mem_357_sv2v_reg  <= data_i[37];
    end 
    if(N6733) begin
      \nz.mem_356_sv2v_reg  <= data_i[36];
    end 
    if(N6732) begin
      \nz.mem_355_sv2v_reg  <= data_i[35];
    end 
    if(N6731) begin
      \nz.mem_354_sv2v_reg  <= data_i[34];
    end 
    if(N6730) begin
      \nz.mem_353_sv2v_reg  <= data_i[33];
    end 
    if(N6729) begin
      \nz.mem_352_sv2v_reg  <= data_i[32];
    end 
    if(N6728) begin
      \nz.mem_351_sv2v_reg  <= data_i[31];
    end 
    if(N6727) begin
      \nz.mem_350_sv2v_reg  <= data_i[30];
    end 
    if(N6726) begin
      \nz.mem_349_sv2v_reg  <= data_i[29];
    end 
    if(N6725) begin
      \nz.mem_348_sv2v_reg  <= data_i[28];
    end 
    if(N6724) begin
      \nz.mem_347_sv2v_reg  <= data_i[27];
    end 
    if(N6723) begin
      \nz.mem_346_sv2v_reg  <= data_i[26];
    end 
    if(N6722) begin
      \nz.mem_345_sv2v_reg  <= data_i[25];
    end 
    if(N6721) begin
      \nz.mem_344_sv2v_reg  <= data_i[24];
    end 
    if(N6720) begin
      \nz.mem_343_sv2v_reg  <= data_i[23];
    end 
    if(N6719) begin
      \nz.mem_342_sv2v_reg  <= data_i[22];
    end 
    if(N6718) begin
      \nz.mem_341_sv2v_reg  <= data_i[21];
    end 
    if(N6717) begin
      \nz.mem_340_sv2v_reg  <= data_i[20];
    end 
    if(N6716) begin
      \nz.mem_339_sv2v_reg  <= data_i[19];
    end 
    if(N6715) begin
      \nz.mem_338_sv2v_reg  <= data_i[18];
    end 
    if(N6714) begin
      \nz.mem_337_sv2v_reg  <= data_i[17];
    end 
    if(N6713) begin
      \nz.mem_336_sv2v_reg  <= data_i[16];
    end 
    if(N6712) begin
      \nz.mem_335_sv2v_reg  <= data_i[15];
    end 
    if(N6711) begin
      \nz.mem_334_sv2v_reg  <= data_i[14];
    end 
    if(N6710) begin
      \nz.mem_333_sv2v_reg  <= data_i[13];
    end 
    if(N6709) begin
      \nz.mem_332_sv2v_reg  <= data_i[12];
    end 
    if(N6708) begin
      \nz.mem_331_sv2v_reg  <= data_i[11];
    end 
    if(N6707) begin
      \nz.mem_330_sv2v_reg  <= data_i[10];
    end 
    if(N6706) begin
      \nz.mem_329_sv2v_reg  <= data_i[9];
    end 
    if(N6705) begin
      \nz.mem_328_sv2v_reg  <= data_i[8];
    end 
    if(N6704) begin
      \nz.mem_327_sv2v_reg  <= data_i[7];
    end 
    if(N6703) begin
      \nz.mem_326_sv2v_reg  <= data_i[6];
    end 
    if(N6702) begin
      \nz.mem_325_sv2v_reg  <= data_i[5];
    end 
    if(N6701) begin
      \nz.mem_324_sv2v_reg  <= data_i[4];
    end 
    if(N6700) begin
      \nz.mem_323_sv2v_reg  <= data_i[3];
    end 
    if(N6699) begin
      \nz.mem_322_sv2v_reg  <= data_i[2];
    end 
    if(N6698) begin
      \nz.mem_321_sv2v_reg  <= data_i[1];
    end 
    if(N6697) begin
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N6696) begin
      \nz.mem_319_sv2v_reg  <= data_i[79];
    end 
    if(N6695) begin
      \nz.mem_318_sv2v_reg  <= data_i[78];
    end 
    if(N6694) begin
      \nz.mem_317_sv2v_reg  <= data_i[77];
    end 
    if(N6693) begin
      \nz.mem_316_sv2v_reg  <= data_i[76];
    end 
    if(N6692) begin
      \nz.mem_315_sv2v_reg  <= data_i[75];
    end 
    if(N6691) begin
      \nz.mem_314_sv2v_reg  <= data_i[74];
    end 
    if(N6690) begin
      \nz.mem_313_sv2v_reg  <= data_i[73];
    end 
    if(N6689) begin
      \nz.mem_312_sv2v_reg  <= data_i[72];
    end 
    if(N6688) begin
      \nz.mem_311_sv2v_reg  <= data_i[71];
    end 
    if(N6687) begin
      \nz.mem_310_sv2v_reg  <= data_i[70];
    end 
    if(N6686) begin
      \nz.mem_309_sv2v_reg  <= data_i[69];
    end 
    if(N6685) begin
      \nz.mem_308_sv2v_reg  <= data_i[68];
    end 
    if(N6684) begin
      \nz.mem_307_sv2v_reg  <= data_i[67];
    end 
    if(N6683) begin
      \nz.mem_306_sv2v_reg  <= data_i[66];
    end 
    if(N6682) begin
      \nz.mem_305_sv2v_reg  <= data_i[65];
    end 
    if(N6681) begin
      \nz.mem_304_sv2v_reg  <= data_i[64];
    end 
    if(N6680) begin
      \nz.mem_303_sv2v_reg  <= data_i[63];
    end 
    if(N6679) begin
      \nz.mem_302_sv2v_reg  <= data_i[62];
    end 
    if(N6678) begin
      \nz.mem_301_sv2v_reg  <= data_i[61];
    end 
    if(N6677) begin
      \nz.mem_300_sv2v_reg  <= data_i[60];
    end 
    if(N6676) begin
      \nz.mem_299_sv2v_reg  <= data_i[59];
    end 
    if(N6675) begin
      \nz.mem_298_sv2v_reg  <= data_i[58];
    end 
    if(N6674) begin
      \nz.mem_297_sv2v_reg  <= data_i[57];
    end 
    if(N6673) begin
      \nz.mem_296_sv2v_reg  <= data_i[56];
    end 
    if(N6672) begin
      \nz.mem_295_sv2v_reg  <= data_i[55];
    end 
    if(N6671) begin
      \nz.mem_294_sv2v_reg  <= data_i[54];
    end 
    if(N6670) begin
      \nz.mem_293_sv2v_reg  <= data_i[53];
    end 
    if(N6669) begin
      \nz.mem_292_sv2v_reg  <= data_i[52];
    end 
    if(N6668) begin
      \nz.mem_291_sv2v_reg  <= data_i[51];
    end 
    if(N6667) begin
      \nz.mem_290_sv2v_reg  <= data_i[50];
    end 
    if(N6666) begin
      \nz.mem_289_sv2v_reg  <= data_i[49];
    end 
    if(N6665) begin
      \nz.mem_288_sv2v_reg  <= data_i[48];
    end 
    if(N6664) begin
      \nz.mem_287_sv2v_reg  <= data_i[47];
    end 
    if(N6663) begin
      \nz.mem_286_sv2v_reg  <= data_i[46];
    end 
    if(N6662) begin
      \nz.mem_285_sv2v_reg  <= data_i[45];
    end 
    if(N6661) begin
      \nz.mem_284_sv2v_reg  <= data_i[44];
    end 
    if(N6660) begin
      \nz.mem_283_sv2v_reg  <= data_i[43];
    end 
    if(N6659) begin
      \nz.mem_282_sv2v_reg  <= data_i[42];
    end 
    if(N6658) begin
      \nz.mem_281_sv2v_reg  <= data_i[41];
    end 
    if(N6657) begin
      \nz.mem_280_sv2v_reg  <= data_i[40];
    end 
    if(N6656) begin
      \nz.mem_279_sv2v_reg  <= data_i[39];
    end 
    if(N6655) begin
      \nz.mem_278_sv2v_reg  <= data_i[38];
    end 
    if(N6654) begin
      \nz.mem_277_sv2v_reg  <= data_i[37];
    end 
    if(N6653) begin
      \nz.mem_276_sv2v_reg  <= data_i[36];
    end 
    if(N6652) begin
      \nz.mem_275_sv2v_reg  <= data_i[35];
    end 
    if(N6651) begin
      \nz.mem_274_sv2v_reg  <= data_i[34];
    end 
    if(N6650) begin
      \nz.mem_273_sv2v_reg  <= data_i[33];
    end 
    if(N6649) begin
      \nz.mem_272_sv2v_reg  <= data_i[32];
    end 
    if(N6648) begin
      \nz.mem_271_sv2v_reg  <= data_i[31];
    end 
    if(N6647) begin
      \nz.mem_270_sv2v_reg  <= data_i[30];
    end 
    if(N6646) begin
      \nz.mem_269_sv2v_reg  <= data_i[29];
    end 
    if(N6645) begin
      \nz.mem_268_sv2v_reg  <= data_i[28];
    end 
    if(N6644) begin
      \nz.mem_267_sv2v_reg  <= data_i[27];
    end 
    if(N6643) begin
      \nz.mem_266_sv2v_reg  <= data_i[26];
    end 
    if(N6642) begin
      \nz.mem_265_sv2v_reg  <= data_i[25];
    end 
    if(N6641) begin
      \nz.mem_264_sv2v_reg  <= data_i[24];
    end 
    if(N6640) begin
      \nz.mem_263_sv2v_reg  <= data_i[23];
    end 
    if(N6639) begin
      \nz.mem_262_sv2v_reg  <= data_i[22];
    end 
    if(N6638) begin
      \nz.mem_261_sv2v_reg  <= data_i[21];
    end 
    if(N6637) begin
      \nz.mem_260_sv2v_reg  <= data_i[20];
    end 
    if(N6636) begin
      \nz.mem_259_sv2v_reg  <= data_i[19];
    end 
    if(N6635) begin
      \nz.mem_258_sv2v_reg  <= data_i[18];
    end 
    if(N6634) begin
      \nz.mem_257_sv2v_reg  <= data_i[17];
    end 
    if(N6633) begin
      \nz.mem_256_sv2v_reg  <= data_i[16];
    end 
    if(N6632) begin
      \nz.mem_255_sv2v_reg  <= data_i[15];
    end 
    if(N6631) begin
      \nz.mem_254_sv2v_reg  <= data_i[14];
    end 
    if(N6630) begin
      \nz.mem_253_sv2v_reg  <= data_i[13];
    end 
    if(N6629) begin
      \nz.mem_252_sv2v_reg  <= data_i[12];
    end 
    if(N6628) begin
      \nz.mem_251_sv2v_reg  <= data_i[11];
    end 
    if(N6627) begin
      \nz.mem_250_sv2v_reg  <= data_i[10];
    end 
    if(N6626) begin
      \nz.mem_249_sv2v_reg  <= data_i[9];
    end 
    if(N6625) begin
      \nz.mem_248_sv2v_reg  <= data_i[8];
    end 
    if(N6624) begin
      \nz.mem_247_sv2v_reg  <= data_i[7];
    end 
    if(N6623) begin
      \nz.mem_246_sv2v_reg  <= data_i[6];
    end 
    if(N6622) begin
      \nz.mem_245_sv2v_reg  <= data_i[5];
    end 
    if(N6621) begin
      \nz.mem_244_sv2v_reg  <= data_i[4];
    end 
    if(N6620) begin
      \nz.mem_243_sv2v_reg  <= data_i[3];
    end 
    if(N6619) begin
      \nz.mem_242_sv2v_reg  <= data_i[2];
    end 
    if(N6618) begin
      \nz.mem_241_sv2v_reg  <= data_i[1];
    end 
    if(N6617) begin
      \nz.mem_240_sv2v_reg  <= data_i[0];
    end 
    if(N6616) begin
      \nz.mem_239_sv2v_reg  <= data_i[79];
    end 
    if(N6615) begin
      \nz.mem_238_sv2v_reg  <= data_i[78];
    end 
    if(N6614) begin
      \nz.mem_237_sv2v_reg  <= data_i[77];
    end 
    if(N6613) begin
      \nz.mem_236_sv2v_reg  <= data_i[76];
    end 
    if(N6612) begin
      \nz.mem_235_sv2v_reg  <= data_i[75];
    end 
    if(N6611) begin
      \nz.mem_234_sv2v_reg  <= data_i[74];
    end 
    if(N6610) begin
      \nz.mem_233_sv2v_reg  <= data_i[73];
    end 
    if(N6609) begin
      \nz.mem_232_sv2v_reg  <= data_i[72];
    end 
    if(N6608) begin
      \nz.mem_231_sv2v_reg  <= data_i[71];
    end 
    if(N6607) begin
      \nz.mem_230_sv2v_reg  <= data_i[70];
    end 
    if(N6606) begin
      \nz.mem_229_sv2v_reg  <= data_i[69];
    end 
    if(N6605) begin
      \nz.mem_228_sv2v_reg  <= data_i[68];
    end 
    if(N6604) begin
      \nz.mem_227_sv2v_reg  <= data_i[67];
    end 
    if(N6603) begin
      \nz.mem_226_sv2v_reg  <= data_i[66];
    end 
    if(N6602) begin
      \nz.mem_225_sv2v_reg  <= data_i[65];
    end 
    if(N6601) begin
      \nz.mem_224_sv2v_reg  <= data_i[64];
    end 
    if(N6600) begin
      \nz.mem_223_sv2v_reg  <= data_i[63];
    end 
    if(N6599) begin
      \nz.mem_222_sv2v_reg  <= data_i[62];
    end 
    if(N6598) begin
      \nz.mem_221_sv2v_reg  <= data_i[61];
    end 
    if(N6597) begin
      \nz.mem_220_sv2v_reg  <= data_i[60];
    end 
    if(N6596) begin
      \nz.mem_219_sv2v_reg  <= data_i[59];
    end 
    if(N6595) begin
      \nz.mem_218_sv2v_reg  <= data_i[58];
    end 
    if(N6594) begin
      \nz.mem_217_sv2v_reg  <= data_i[57];
    end 
    if(N6593) begin
      \nz.mem_216_sv2v_reg  <= data_i[56];
    end 
    if(N6592) begin
      \nz.mem_215_sv2v_reg  <= data_i[55];
    end 
    if(N6591) begin
      \nz.mem_214_sv2v_reg  <= data_i[54];
    end 
    if(N6590) begin
      \nz.mem_213_sv2v_reg  <= data_i[53];
    end 
    if(N6589) begin
      \nz.mem_212_sv2v_reg  <= data_i[52];
    end 
    if(N6588) begin
      \nz.mem_211_sv2v_reg  <= data_i[51];
    end 
    if(N6587) begin
      \nz.mem_210_sv2v_reg  <= data_i[50];
    end 
    if(N6586) begin
      \nz.mem_209_sv2v_reg  <= data_i[49];
    end 
    if(N6585) begin
      \nz.mem_208_sv2v_reg  <= data_i[48];
    end 
    if(N6584) begin
      \nz.mem_207_sv2v_reg  <= data_i[47];
    end 
    if(N6583) begin
      \nz.mem_206_sv2v_reg  <= data_i[46];
    end 
    if(N6582) begin
      \nz.mem_205_sv2v_reg  <= data_i[45];
    end 
    if(N6581) begin
      \nz.mem_204_sv2v_reg  <= data_i[44];
    end 
    if(N6580) begin
      \nz.mem_203_sv2v_reg  <= data_i[43];
    end 
    if(N6579) begin
      \nz.mem_202_sv2v_reg  <= data_i[42];
    end 
    if(N6578) begin
      \nz.mem_201_sv2v_reg  <= data_i[41];
    end 
    if(N6577) begin
      \nz.mem_200_sv2v_reg  <= data_i[40];
    end 
    if(N6576) begin
      \nz.mem_199_sv2v_reg  <= data_i[39];
    end 
    if(N6575) begin
      \nz.mem_198_sv2v_reg  <= data_i[38];
    end 
    if(N6574) begin
      \nz.mem_197_sv2v_reg  <= data_i[37];
    end 
    if(N6573) begin
      \nz.mem_196_sv2v_reg  <= data_i[36];
    end 
    if(N6572) begin
      \nz.mem_195_sv2v_reg  <= data_i[35];
    end 
    if(N6571) begin
      \nz.mem_194_sv2v_reg  <= data_i[34];
    end 
    if(N6570) begin
      \nz.mem_193_sv2v_reg  <= data_i[33];
    end 
    if(N6569) begin
      \nz.mem_192_sv2v_reg  <= data_i[32];
    end 
    if(N6568) begin
      \nz.mem_191_sv2v_reg  <= data_i[31];
    end 
    if(N6567) begin
      \nz.mem_190_sv2v_reg  <= data_i[30];
    end 
    if(N6566) begin
      \nz.mem_189_sv2v_reg  <= data_i[29];
    end 
    if(N6565) begin
      \nz.mem_188_sv2v_reg  <= data_i[28];
    end 
    if(N6564) begin
      \nz.mem_187_sv2v_reg  <= data_i[27];
    end 
    if(N6563) begin
      \nz.mem_186_sv2v_reg  <= data_i[26];
    end 
    if(N6562) begin
      \nz.mem_185_sv2v_reg  <= data_i[25];
    end 
    if(N6561) begin
      \nz.mem_184_sv2v_reg  <= data_i[24];
    end 
    if(N6560) begin
      \nz.mem_183_sv2v_reg  <= data_i[23];
    end 
    if(N6559) begin
      \nz.mem_182_sv2v_reg  <= data_i[22];
    end 
    if(N6558) begin
      \nz.mem_181_sv2v_reg  <= data_i[21];
    end 
    if(N6557) begin
      \nz.mem_180_sv2v_reg  <= data_i[20];
    end 
    if(N6556) begin
      \nz.mem_179_sv2v_reg  <= data_i[19];
    end 
    if(N6555) begin
      \nz.mem_178_sv2v_reg  <= data_i[18];
    end 
    if(N6554) begin
      \nz.mem_177_sv2v_reg  <= data_i[17];
    end 
    if(N6553) begin
      \nz.mem_176_sv2v_reg  <= data_i[16];
    end 
    if(N6552) begin
      \nz.mem_175_sv2v_reg  <= data_i[15];
    end 
    if(N6551) begin
      \nz.mem_174_sv2v_reg  <= data_i[14];
    end 
    if(N6550) begin
      \nz.mem_173_sv2v_reg  <= data_i[13];
    end 
    if(N6549) begin
      \nz.mem_172_sv2v_reg  <= data_i[12];
    end 
    if(N6548) begin
      \nz.mem_171_sv2v_reg  <= data_i[11];
    end 
    if(N6547) begin
      \nz.mem_170_sv2v_reg  <= data_i[10];
    end 
    if(N6546) begin
      \nz.mem_169_sv2v_reg  <= data_i[9];
    end 
    if(N6545) begin
      \nz.mem_168_sv2v_reg  <= data_i[8];
    end 
    if(N6544) begin
      \nz.mem_167_sv2v_reg  <= data_i[7];
    end 
    if(N6543) begin
      \nz.mem_166_sv2v_reg  <= data_i[6];
    end 
    if(N6542) begin
      \nz.mem_165_sv2v_reg  <= data_i[5];
    end 
    if(N6541) begin
      \nz.mem_164_sv2v_reg  <= data_i[4];
    end 
    if(N6540) begin
      \nz.mem_163_sv2v_reg  <= data_i[3];
    end 
    if(N6539) begin
      \nz.mem_162_sv2v_reg  <= data_i[2];
    end 
    if(N6538) begin
      \nz.mem_161_sv2v_reg  <= data_i[1];
    end 
    if(N6537) begin
      \nz.mem_160_sv2v_reg  <= data_i[0];
    end 
    if(N6536) begin
      \nz.mem_159_sv2v_reg  <= data_i[79];
    end 
    if(N6535) begin
      \nz.mem_158_sv2v_reg  <= data_i[78];
    end 
    if(N6534) begin
      \nz.mem_157_sv2v_reg  <= data_i[77];
    end 
    if(N6533) begin
      \nz.mem_156_sv2v_reg  <= data_i[76];
    end 
    if(N6532) begin
      \nz.mem_155_sv2v_reg  <= data_i[75];
    end 
    if(N6531) begin
      \nz.mem_154_sv2v_reg  <= data_i[74];
    end 
    if(N6530) begin
      \nz.mem_153_sv2v_reg  <= data_i[73];
    end 
    if(N6529) begin
      \nz.mem_152_sv2v_reg  <= data_i[72];
    end 
    if(N6528) begin
      \nz.mem_151_sv2v_reg  <= data_i[71];
    end 
    if(N6527) begin
      \nz.mem_150_sv2v_reg  <= data_i[70];
    end 
    if(N6526) begin
      \nz.mem_149_sv2v_reg  <= data_i[69];
    end 
    if(N6525) begin
      \nz.mem_148_sv2v_reg  <= data_i[68];
    end 
    if(N6524) begin
      \nz.mem_147_sv2v_reg  <= data_i[67];
    end 
    if(N6523) begin
      \nz.mem_146_sv2v_reg  <= data_i[66];
    end 
    if(N6522) begin
      \nz.mem_145_sv2v_reg  <= data_i[65];
    end 
    if(N6521) begin
      \nz.mem_144_sv2v_reg  <= data_i[64];
    end 
    if(N6520) begin
      \nz.mem_143_sv2v_reg  <= data_i[63];
    end 
    if(N6519) begin
      \nz.mem_142_sv2v_reg  <= data_i[62];
    end 
    if(N6518) begin
      \nz.mem_141_sv2v_reg  <= data_i[61];
    end 
    if(N6517) begin
      \nz.mem_140_sv2v_reg  <= data_i[60];
    end 
    if(N6516) begin
      \nz.mem_139_sv2v_reg  <= data_i[59];
    end 
    if(N6515) begin
      \nz.mem_138_sv2v_reg  <= data_i[58];
    end 
    if(N6514) begin
      \nz.mem_137_sv2v_reg  <= data_i[57];
    end 
    if(N6513) begin
      \nz.mem_136_sv2v_reg  <= data_i[56];
    end 
    if(N6512) begin
      \nz.mem_135_sv2v_reg  <= data_i[55];
    end 
    if(N6511) begin
      \nz.mem_134_sv2v_reg  <= data_i[54];
    end 
    if(N6510) begin
      \nz.mem_133_sv2v_reg  <= data_i[53];
    end 
    if(N6509) begin
      \nz.mem_132_sv2v_reg  <= data_i[52];
    end 
    if(N6508) begin
      \nz.mem_131_sv2v_reg  <= data_i[51];
    end 
    if(N6507) begin
      \nz.mem_130_sv2v_reg  <= data_i[50];
    end 
    if(N6506) begin
      \nz.mem_129_sv2v_reg  <= data_i[49];
    end 
    if(N6505) begin
      \nz.mem_128_sv2v_reg  <= data_i[48];
    end 
    if(N6504) begin
      \nz.mem_127_sv2v_reg  <= data_i[47];
    end 
    if(N6503) begin
      \nz.mem_126_sv2v_reg  <= data_i[46];
    end 
    if(N6502) begin
      \nz.mem_125_sv2v_reg  <= data_i[45];
    end 
    if(N6501) begin
      \nz.mem_124_sv2v_reg  <= data_i[44];
    end 
    if(N6500) begin
      \nz.mem_123_sv2v_reg  <= data_i[43];
    end 
    if(N6499) begin
      \nz.mem_122_sv2v_reg  <= data_i[42];
    end 
    if(N6498) begin
      \nz.mem_121_sv2v_reg  <= data_i[41];
    end 
    if(N6497) begin
      \nz.mem_120_sv2v_reg  <= data_i[40];
    end 
    if(N6496) begin
      \nz.mem_119_sv2v_reg  <= data_i[39];
    end 
    if(N6495) begin
      \nz.mem_118_sv2v_reg  <= data_i[38];
    end 
    if(N6494) begin
      \nz.mem_117_sv2v_reg  <= data_i[37];
    end 
    if(N6493) begin
      \nz.mem_116_sv2v_reg  <= data_i[36];
    end 
    if(N6492) begin
      \nz.mem_115_sv2v_reg  <= data_i[35];
    end 
    if(N6491) begin
      \nz.mem_114_sv2v_reg  <= data_i[34];
    end 
    if(N6490) begin
      \nz.mem_113_sv2v_reg  <= data_i[33];
    end 
    if(N6489) begin
      \nz.mem_112_sv2v_reg  <= data_i[32];
    end 
    if(N6488) begin
      \nz.mem_111_sv2v_reg  <= data_i[31];
    end 
    if(N6487) begin
      \nz.mem_110_sv2v_reg  <= data_i[30];
    end 
    if(N6486) begin
      \nz.mem_109_sv2v_reg  <= data_i[29];
    end 
    if(N6485) begin
      \nz.mem_108_sv2v_reg  <= data_i[28];
    end 
    if(N6484) begin
      \nz.mem_107_sv2v_reg  <= data_i[27];
    end 
    if(N6483) begin
      \nz.mem_106_sv2v_reg  <= data_i[26];
    end 
    if(N6482) begin
      \nz.mem_105_sv2v_reg  <= data_i[25];
    end 
    if(N6481) begin
      \nz.mem_104_sv2v_reg  <= data_i[24];
    end 
    if(N6480) begin
      \nz.mem_103_sv2v_reg  <= data_i[23];
    end 
    if(N6479) begin
      \nz.mem_102_sv2v_reg  <= data_i[22];
    end 
    if(N6478) begin
      \nz.mem_101_sv2v_reg  <= data_i[21];
    end 
    if(N6477) begin
      \nz.mem_100_sv2v_reg  <= data_i[20];
    end 
    if(N6476) begin
      \nz.mem_99_sv2v_reg  <= data_i[19];
    end 
    if(N6475) begin
      \nz.mem_98_sv2v_reg  <= data_i[18];
    end 
    if(N6474) begin
      \nz.mem_97_sv2v_reg  <= data_i[17];
    end 
    if(N6473) begin
      \nz.mem_96_sv2v_reg  <= data_i[16];
    end 
    if(N6472) begin
      \nz.mem_95_sv2v_reg  <= data_i[15];
    end 
    if(N6471) begin
      \nz.mem_94_sv2v_reg  <= data_i[14];
    end 
    if(N6470) begin
      \nz.mem_93_sv2v_reg  <= data_i[13];
    end 
    if(N6469) begin
      \nz.mem_92_sv2v_reg  <= data_i[12];
    end 
    if(N6468) begin
      \nz.mem_91_sv2v_reg  <= data_i[11];
    end 
    if(N6467) begin
      \nz.mem_90_sv2v_reg  <= data_i[10];
    end 
    if(N6466) begin
      \nz.mem_89_sv2v_reg  <= data_i[9];
    end 
    if(N6465) begin
      \nz.mem_88_sv2v_reg  <= data_i[8];
    end 
    if(N6464) begin
      \nz.mem_87_sv2v_reg  <= data_i[7];
    end 
    if(N6463) begin
      \nz.mem_86_sv2v_reg  <= data_i[6];
    end 
    if(N6462) begin
      \nz.mem_85_sv2v_reg  <= data_i[5];
    end 
    if(N6461) begin
      \nz.mem_84_sv2v_reg  <= data_i[4];
    end 
    if(N6460) begin
      \nz.mem_83_sv2v_reg  <= data_i[3];
    end 
    if(N6459) begin
      \nz.mem_82_sv2v_reg  <= data_i[2];
    end 
    if(N6458) begin
      \nz.mem_81_sv2v_reg  <= data_i[1];
    end 
    if(N6457) begin
      \nz.mem_80_sv2v_reg  <= data_i[0];
    end 
    if(N6456) begin
      \nz.mem_79_sv2v_reg  <= data_i[79];
    end 
    if(N6455) begin
      \nz.mem_78_sv2v_reg  <= data_i[78];
    end 
    if(N6454) begin
      \nz.mem_77_sv2v_reg  <= data_i[77];
    end 
    if(N6453) begin
      \nz.mem_76_sv2v_reg  <= data_i[76];
    end 
    if(N6452) begin
      \nz.mem_75_sv2v_reg  <= data_i[75];
    end 
    if(N6451) begin
      \nz.mem_74_sv2v_reg  <= data_i[74];
    end 
    if(N6450) begin
      \nz.mem_73_sv2v_reg  <= data_i[73];
    end 
    if(N6449) begin
      \nz.mem_72_sv2v_reg  <= data_i[72];
    end 
    if(N6448) begin
      \nz.mem_71_sv2v_reg  <= data_i[71];
    end 
    if(N6447) begin
      \nz.mem_70_sv2v_reg  <= data_i[70];
    end 
    if(N6446) begin
      \nz.mem_69_sv2v_reg  <= data_i[69];
    end 
    if(N6445) begin
      \nz.mem_68_sv2v_reg  <= data_i[68];
    end 
    if(N6444) begin
      \nz.mem_67_sv2v_reg  <= data_i[67];
    end 
    if(N6443) begin
      \nz.mem_66_sv2v_reg  <= data_i[66];
    end 
    if(N6442) begin
      \nz.mem_65_sv2v_reg  <= data_i[65];
    end 
    if(N6441) begin
      \nz.mem_64_sv2v_reg  <= data_i[64];
    end 
    if(N6440) begin
      \nz.mem_63_sv2v_reg  <= data_i[63];
    end 
    if(N6439) begin
      \nz.mem_62_sv2v_reg  <= data_i[62];
    end 
    if(N6438) begin
      \nz.mem_61_sv2v_reg  <= data_i[61];
    end 
    if(N6437) begin
      \nz.mem_60_sv2v_reg  <= data_i[60];
    end 
    if(N6436) begin
      \nz.mem_59_sv2v_reg  <= data_i[59];
    end 
    if(N6435) begin
      \nz.mem_58_sv2v_reg  <= data_i[58];
    end 
    if(N6434) begin
      \nz.mem_57_sv2v_reg  <= data_i[57];
    end 
    if(N6433) begin
      \nz.mem_56_sv2v_reg  <= data_i[56];
    end 
    if(N6432) begin
      \nz.mem_55_sv2v_reg  <= data_i[55];
    end 
    if(N6431) begin
      \nz.mem_54_sv2v_reg  <= data_i[54];
    end 
    if(N6430) begin
      \nz.mem_53_sv2v_reg  <= data_i[53];
    end 
    if(N6429) begin
      \nz.mem_52_sv2v_reg  <= data_i[52];
    end 
    if(N6428) begin
      \nz.mem_51_sv2v_reg  <= data_i[51];
    end 
    if(N6427) begin
      \nz.mem_50_sv2v_reg  <= data_i[50];
    end 
    if(N6426) begin
      \nz.mem_49_sv2v_reg  <= data_i[49];
    end 
    if(N6425) begin
      \nz.mem_48_sv2v_reg  <= data_i[48];
    end 
    if(N6424) begin
      \nz.mem_47_sv2v_reg  <= data_i[47];
    end 
    if(N6423) begin
      \nz.mem_46_sv2v_reg  <= data_i[46];
    end 
    if(N6422) begin
      \nz.mem_45_sv2v_reg  <= data_i[45];
    end 
    if(N6421) begin
      \nz.mem_44_sv2v_reg  <= data_i[44];
    end 
    if(N6420) begin
      \nz.mem_43_sv2v_reg  <= data_i[43];
    end 
    if(N6419) begin
      \nz.mem_42_sv2v_reg  <= data_i[42];
    end 
    if(N6418) begin
      \nz.mem_41_sv2v_reg  <= data_i[41];
    end 
    if(N6417) begin
      \nz.mem_40_sv2v_reg  <= data_i[40];
    end 
    if(N6416) begin
      \nz.mem_39_sv2v_reg  <= data_i[39];
    end 
    if(N6415) begin
      \nz.mem_38_sv2v_reg  <= data_i[38];
    end 
    if(N6414) begin
      \nz.mem_37_sv2v_reg  <= data_i[37];
    end 
    if(N6413) begin
      \nz.mem_36_sv2v_reg  <= data_i[36];
    end 
    if(N6412) begin
      \nz.mem_35_sv2v_reg  <= data_i[35];
    end 
    if(N6411) begin
      \nz.mem_34_sv2v_reg  <= data_i[34];
    end 
    if(N6410) begin
      \nz.mem_33_sv2v_reg  <= data_i[33];
    end 
    if(N6409) begin
      \nz.mem_32_sv2v_reg  <= data_i[32];
    end 
    if(N6408) begin
      \nz.mem_31_sv2v_reg  <= data_i[31];
    end 
    if(N6407) begin
      \nz.mem_30_sv2v_reg  <= data_i[30];
    end 
    if(N6406) begin
      \nz.mem_29_sv2v_reg  <= data_i[29];
    end 
    if(N6405) begin
      \nz.mem_28_sv2v_reg  <= data_i[28];
    end 
    if(N6404) begin
      \nz.mem_27_sv2v_reg  <= data_i[27];
    end 
    if(N6403) begin
      \nz.mem_26_sv2v_reg  <= data_i[26];
    end 
    if(N6402) begin
      \nz.mem_25_sv2v_reg  <= data_i[25];
    end 
    if(N6401) begin
      \nz.mem_24_sv2v_reg  <= data_i[24];
    end 
    if(N6400) begin
      \nz.mem_23_sv2v_reg  <= data_i[23];
    end 
    if(N6399) begin
      \nz.mem_22_sv2v_reg  <= data_i[22];
    end 
    if(N6398) begin
      \nz.mem_21_sv2v_reg  <= data_i[21];
    end 
    if(N6397) begin
      \nz.mem_20_sv2v_reg  <= data_i[20];
    end 
    if(N6396) begin
      \nz.mem_19_sv2v_reg  <= data_i[19];
    end 
    if(N6395) begin
      \nz.mem_18_sv2v_reg  <= data_i[18];
    end 
    if(N6394) begin
      \nz.mem_17_sv2v_reg  <= data_i[17];
    end 
    if(N6393) begin
      \nz.mem_16_sv2v_reg  <= data_i[16];
    end 
    if(N6392) begin
      \nz.mem_15_sv2v_reg  <= data_i[15];
    end 
    if(N6391) begin
      \nz.mem_14_sv2v_reg  <= data_i[14];
    end 
    if(N6390) begin
      \nz.mem_13_sv2v_reg  <= data_i[13];
    end 
    if(N6389) begin
      \nz.mem_12_sv2v_reg  <= data_i[12];
    end 
    if(N6388) begin
      \nz.mem_11_sv2v_reg  <= data_i[11];
    end 
    if(N6387) begin
      \nz.mem_10_sv2v_reg  <= data_i[10];
    end 
    if(N6386) begin
      \nz.mem_9_sv2v_reg  <= data_i[9];
    end 
    if(N6385) begin
      \nz.mem_8_sv2v_reg  <= data_i[8];
    end 
    if(N6384) begin
      \nz.mem_7_sv2v_reg  <= data_i[7];
    end 
    if(N6383) begin
      \nz.mem_6_sv2v_reg  <= data_i[6];
    end 
    if(N6382) begin
      \nz.mem_5_sv2v_reg  <= data_i[5];
    end 
    if(N6381) begin
      \nz.mem_4_sv2v_reg  <= data_i[4];
    end 
    if(N6380) begin
      \nz.mem_3_sv2v_reg  <= data_i[3];
    end 
    if(N6379) begin
      \nz.mem_2_sv2v_reg  <= data_i[2];
    end 
    if(N6378) begin
      \nz.mem_1_sv2v_reg  <= data_i[1];
    end 
    if(N6377) begin
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p80_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [79:0] data_i;
  input [5:0] addr_i;
  input [79:0] w_mask_i;
  output [79:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [79:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p80_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_en_width_p8_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  wire [7:0] data_o;
  reg data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p8
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  wire [7:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p8_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1_verbose_p0
(
  clk_i,
  v_i,
  reset_i,
  data_i,
  addr_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input v_i;
  input reset_i;
  input w_i;
  wire [7:0] data_o,\nz.addr_r ,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,\nz.read_en ,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,\nz.llr.read_en_r ,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095;
  wire [2047:0] \nz.mem ;
  reg \nz.addr_r_7_sv2v_reg ,\nz.addr_r_6_sv2v_reg ,\nz.addr_r_5_sv2v_reg ,
  \nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,\nz.addr_r_2_sv2v_reg ,
  \nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,\nz.mem_2047_sv2v_reg ,\nz.mem_2046_sv2v_reg ,
  \nz.mem_2045_sv2v_reg ,\nz.mem_2044_sv2v_reg ,\nz.mem_2043_sv2v_reg ,
  \nz.mem_2042_sv2v_reg ,\nz.mem_2041_sv2v_reg ,\nz.mem_2040_sv2v_reg ,\nz.mem_2039_sv2v_reg ,
  \nz.mem_2038_sv2v_reg ,\nz.mem_2037_sv2v_reg ,\nz.mem_2036_sv2v_reg ,
  \nz.mem_2035_sv2v_reg ,\nz.mem_2034_sv2v_reg ,\nz.mem_2033_sv2v_reg ,\nz.mem_2032_sv2v_reg ,
  \nz.mem_2031_sv2v_reg ,\nz.mem_2030_sv2v_reg ,\nz.mem_2029_sv2v_reg ,
  \nz.mem_2028_sv2v_reg ,\nz.mem_2027_sv2v_reg ,\nz.mem_2026_sv2v_reg ,\nz.mem_2025_sv2v_reg ,
  \nz.mem_2024_sv2v_reg ,\nz.mem_2023_sv2v_reg ,\nz.mem_2022_sv2v_reg ,
  \nz.mem_2021_sv2v_reg ,\nz.mem_2020_sv2v_reg ,\nz.mem_2019_sv2v_reg ,\nz.mem_2018_sv2v_reg ,
  \nz.mem_2017_sv2v_reg ,\nz.mem_2016_sv2v_reg ,\nz.mem_2015_sv2v_reg ,
  \nz.mem_2014_sv2v_reg ,\nz.mem_2013_sv2v_reg ,\nz.mem_2012_sv2v_reg ,\nz.mem_2011_sv2v_reg ,
  \nz.mem_2010_sv2v_reg ,\nz.mem_2009_sv2v_reg ,\nz.mem_2008_sv2v_reg ,
  \nz.mem_2007_sv2v_reg ,\nz.mem_2006_sv2v_reg ,\nz.mem_2005_sv2v_reg ,\nz.mem_2004_sv2v_reg ,
  \nz.mem_2003_sv2v_reg ,\nz.mem_2002_sv2v_reg ,\nz.mem_2001_sv2v_reg ,
  \nz.mem_2000_sv2v_reg ,\nz.mem_1999_sv2v_reg ,\nz.mem_1998_sv2v_reg ,\nz.mem_1997_sv2v_reg ,
  \nz.mem_1996_sv2v_reg ,\nz.mem_1995_sv2v_reg ,\nz.mem_1994_sv2v_reg ,
  \nz.mem_1993_sv2v_reg ,\nz.mem_1992_sv2v_reg ,\nz.mem_1991_sv2v_reg ,\nz.mem_1990_sv2v_reg ,
  \nz.mem_1989_sv2v_reg ,\nz.mem_1988_sv2v_reg ,\nz.mem_1987_sv2v_reg ,
  \nz.mem_1986_sv2v_reg ,\nz.mem_1985_sv2v_reg ,\nz.mem_1984_sv2v_reg ,\nz.mem_1983_sv2v_reg ,
  \nz.mem_1982_sv2v_reg ,\nz.mem_1981_sv2v_reg ,\nz.mem_1980_sv2v_reg ,
  \nz.mem_1979_sv2v_reg ,\nz.mem_1978_sv2v_reg ,\nz.mem_1977_sv2v_reg ,\nz.mem_1976_sv2v_reg ,
  \nz.mem_1975_sv2v_reg ,\nz.mem_1974_sv2v_reg ,\nz.mem_1973_sv2v_reg ,
  \nz.mem_1972_sv2v_reg ,\nz.mem_1971_sv2v_reg ,\nz.mem_1970_sv2v_reg ,
  \nz.mem_1969_sv2v_reg ,\nz.mem_1968_sv2v_reg ,\nz.mem_1967_sv2v_reg ,\nz.mem_1966_sv2v_reg ,
  \nz.mem_1965_sv2v_reg ,\nz.mem_1964_sv2v_reg ,\nz.mem_1963_sv2v_reg ,
  \nz.mem_1962_sv2v_reg ,\nz.mem_1961_sv2v_reg ,\nz.mem_1960_sv2v_reg ,\nz.mem_1959_sv2v_reg ,
  \nz.mem_1958_sv2v_reg ,\nz.mem_1957_sv2v_reg ,\nz.mem_1956_sv2v_reg ,
  \nz.mem_1955_sv2v_reg ,\nz.mem_1954_sv2v_reg ,\nz.mem_1953_sv2v_reg ,\nz.mem_1952_sv2v_reg ,
  \nz.mem_1951_sv2v_reg ,\nz.mem_1950_sv2v_reg ,\nz.mem_1949_sv2v_reg ,
  \nz.mem_1948_sv2v_reg ,\nz.mem_1947_sv2v_reg ,\nz.mem_1946_sv2v_reg ,\nz.mem_1945_sv2v_reg ,
  \nz.mem_1944_sv2v_reg ,\nz.mem_1943_sv2v_reg ,\nz.mem_1942_sv2v_reg ,
  \nz.mem_1941_sv2v_reg ,\nz.mem_1940_sv2v_reg ,\nz.mem_1939_sv2v_reg ,\nz.mem_1938_sv2v_reg ,
  \nz.mem_1937_sv2v_reg ,\nz.mem_1936_sv2v_reg ,\nz.mem_1935_sv2v_reg ,
  \nz.mem_1934_sv2v_reg ,\nz.mem_1933_sv2v_reg ,\nz.mem_1932_sv2v_reg ,\nz.mem_1931_sv2v_reg ,
  \nz.mem_1930_sv2v_reg ,\nz.mem_1929_sv2v_reg ,\nz.mem_1928_sv2v_reg ,
  \nz.mem_1927_sv2v_reg ,\nz.mem_1926_sv2v_reg ,\nz.mem_1925_sv2v_reg ,\nz.mem_1924_sv2v_reg ,
  \nz.mem_1923_sv2v_reg ,\nz.mem_1922_sv2v_reg ,\nz.mem_1921_sv2v_reg ,
  \nz.mem_1920_sv2v_reg ,\nz.mem_1919_sv2v_reg ,\nz.mem_1918_sv2v_reg ,\nz.mem_1917_sv2v_reg ,
  \nz.mem_1916_sv2v_reg ,\nz.mem_1915_sv2v_reg ,\nz.mem_1914_sv2v_reg ,
  \nz.mem_1913_sv2v_reg ,\nz.mem_1912_sv2v_reg ,\nz.mem_1911_sv2v_reg ,\nz.mem_1910_sv2v_reg ,
  \nz.mem_1909_sv2v_reg ,\nz.mem_1908_sv2v_reg ,\nz.mem_1907_sv2v_reg ,
  \nz.mem_1906_sv2v_reg ,\nz.mem_1905_sv2v_reg ,\nz.mem_1904_sv2v_reg ,\nz.mem_1903_sv2v_reg ,
  \nz.mem_1902_sv2v_reg ,\nz.mem_1901_sv2v_reg ,\nz.mem_1900_sv2v_reg ,
  \nz.mem_1899_sv2v_reg ,\nz.mem_1898_sv2v_reg ,\nz.mem_1897_sv2v_reg ,\nz.mem_1896_sv2v_reg ,
  \nz.mem_1895_sv2v_reg ,\nz.mem_1894_sv2v_reg ,\nz.mem_1893_sv2v_reg ,
  \nz.mem_1892_sv2v_reg ,\nz.mem_1891_sv2v_reg ,\nz.mem_1890_sv2v_reg ,
  \nz.mem_1889_sv2v_reg ,\nz.mem_1888_sv2v_reg ,\nz.mem_1887_sv2v_reg ,\nz.mem_1886_sv2v_reg ,
  \nz.mem_1885_sv2v_reg ,\nz.mem_1884_sv2v_reg ,\nz.mem_1883_sv2v_reg ,
  \nz.mem_1882_sv2v_reg ,\nz.mem_1881_sv2v_reg ,\nz.mem_1880_sv2v_reg ,\nz.mem_1879_sv2v_reg ,
  \nz.mem_1878_sv2v_reg ,\nz.mem_1877_sv2v_reg ,\nz.mem_1876_sv2v_reg ,
  \nz.mem_1875_sv2v_reg ,\nz.mem_1874_sv2v_reg ,\nz.mem_1873_sv2v_reg ,\nz.mem_1872_sv2v_reg ,
  \nz.mem_1871_sv2v_reg ,\nz.mem_1870_sv2v_reg ,\nz.mem_1869_sv2v_reg ,
  \nz.mem_1868_sv2v_reg ,\nz.mem_1867_sv2v_reg ,\nz.mem_1866_sv2v_reg ,\nz.mem_1865_sv2v_reg ,
  \nz.mem_1864_sv2v_reg ,\nz.mem_1863_sv2v_reg ,\nz.mem_1862_sv2v_reg ,
  \nz.mem_1861_sv2v_reg ,\nz.mem_1860_sv2v_reg ,\nz.mem_1859_sv2v_reg ,\nz.mem_1858_sv2v_reg ,
  \nz.mem_1857_sv2v_reg ,\nz.mem_1856_sv2v_reg ,\nz.mem_1855_sv2v_reg ,
  \nz.mem_1854_sv2v_reg ,\nz.mem_1853_sv2v_reg ,\nz.mem_1852_sv2v_reg ,\nz.mem_1851_sv2v_reg ,
  \nz.mem_1850_sv2v_reg ,\nz.mem_1849_sv2v_reg ,\nz.mem_1848_sv2v_reg ,
  \nz.mem_1847_sv2v_reg ,\nz.mem_1846_sv2v_reg ,\nz.mem_1845_sv2v_reg ,\nz.mem_1844_sv2v_reg ,
  \nz.mem_1843_sv2v_reg ,\nz.mem_1842_sv2v_reg ,\nz.mem_1841_sv2v_reg ,
  \nz.mem_1840_sv2v_reg ,\nz.mem_1839_sv2v_reg ,\nz.mem_1838_sv2v_reg ,\nz.mem_1837_sv2v_reg ,
  \nz.mem_1836_sv2v_reg ,\nz.mem_1835_sv2v_reg ,\nz.mem_1834_sv2v_reg ,
  \nz.mem_1833_sv2v_reg ,\nz.mem_1832_sv2v_reg ,\nz.mem_1831_sv2v_reg ,\nz.mem_1830_sv2v_reg ,
  \nz.mem_1829_sv2v_reg ,\nz.mem_1828_sv2v_reg ,\nz.mem_1827_sv2v_reg ,
  \nz.mem_1826_sv2v_reg ,\nz.mem_1825_sv2v_reg ,\nz.mem_1824_sv2v_reg ,\nz.mem_1823_sv2v_reg ,
  \nz.mem_1822_sv2v_reg ,\nz.mem_1821_sv2v_reg ,\nz.mem_1820_sv2v_reg ,
  \nz.mem_1819_sv2v_reg ,\nz.mem_1818_sv2v_reg ,\nz.mem_1817_sv2v_reg ,\nz.mem_1816_sv2v_reg ,
  \nz.mem_1815_sv2v_reg ,\nz.mem_1814_sv2v_reg ,\nz.mem_1813_sv2v_reg ,
  \nz.mem_1812_sv2v_reg ,\nz.mem_1811_sv2v_reg ,\nz.mem_1810_sv2v_reg ,
  \nz.mem_1809_sv2v_reg ,\nz.mem_1808_sv2v_reg ,\nz.mem_1807_sv2v_reg ,\nz.mem_1806_sv2v_reg ,
  \nz.mem_1805_sv2v_reg ,\nz.mem_1804_sv2v_reg ,\nz.mem_1803_sv2v_reg ,
  \nz.mem_1802_sv2v_reg ,\nz.mem_1801_sv2v_reg ,\nz.mem_1800_sv2v_reg ,\nz.mem_1799_sv2v_reg ,
  \nz.mem_1798_sv2v_reg ,\nz.mem_1797_sv2v_reg ,\nz.mem_1796_sv2v_reg ,
  \nz.mem_1795_sv2v_reg ,\nz.mem_1794_sv2v_reg ,\nz.mem_1793_sv2v_reg ,\nz.mem_1792_sv2v_reg ,
  \nz.mem_1791_sv2v_reg ,\nz.mem_1790_sv2v_reg ,\nz.mem_1789_sv2v_reg ,
  \nz.mem_1788_sv2v_reg ,\nz.mem_1787_sv2v_reg ,\nz.mem_1786_sv2v_reg ,\nz.mem_1785_sv2v_reg ,
  \nz.mem_1784_sv2v_reg ,\nz.mem_1783_sv2v_reg ,\nz.mem_1782_sv2v_reg ,
  \nz.mem_1781_sv2v_reg ,\nz.mem_1780_sv2v_reg ,\nz.mem_1779_sv2v_reg ,\nz.mem_1778_sv2v_reg ,
  \nz.mem_1777_sv2v_reg ,\nz.mem_1776_sv2v_reg ,\nz.mem_1775_sv2v_reg ,
  \nz.mem_1774_sv2v_reg ,\nz.mem_1773_sv2v_reg ,\nz.mem_1772_sv2v_reg ,\nz.mem_1771_sv2v_reg ,
  \nz.mem_1770_sv2v_reg ,\nz.mem_1769_sv2v_reg ,\nz.mem_1768_sv2v_reg ,
  \nz.mem_1767_sv2v_reg ,\nz.mem_1766_sv2v_reg ,\nz.mem_1765_sv2v_reg ,\nz.mem_1764_sv2v_reg ,
  \nz.mem_1763_sv2v_reg ,\nz.mem_1762_sv2v_reg ,\nz.mem_1761_sv2v_reg ,
  \nz.mem_1760_sv2v_reg ,\nz.mem_1759_sv2v_reg ,\nz.mem_1758_sv2v_reg ,\nz.mem_1757_sv2v_reg ,
  \nz.mem_1756_sv2v_reg ,\nz.mem_1755_sv2v_reg ,\nz.mem_1754_sv2v_reg ,
  \nz.mem_1753_sv2v_reg ,\nz.mem_1752_sv2v_reg ,\nz.mem_1751_sv2v_reg ,\nz.mem_1750_sv2v_reg ,
  \nz.mem_1749_sv2v_reg ,\nz.mem_1748_sv2v_reg ,\nz.mem_1747_sv2v_reg ,
  \nz.mem_1746_sv2v_reg ,\nz.mem_1745_sv2v_reg ,\nz.mem_1744_sv2v_reg ,\nz.mem_1743_sv2v_reg ,
  \nz.mem_1742_sv2v_reg ,\nz.mem_1741_sv2v_reg ,\nz.mem_1740_sv2v_reg ,
  \nz.mem_1739_sv2v_reg ,\nz.mem_1738_sv2v_reg ,\nz.mem_1737_sv2v_reg ,\nz.mem_1736_sv2v_reg ,
  \nz.mem_1735_sv2v_reg ,\nz.mem_1734_sv2v_reg ,\nz.mem_1733_sv2v_reg ,
  \nz.mem_1732_sv2v_reg ,\nz.mem_1731_sv2v_reg ,\nz.mem_1730_sv2v_reg ,
  \nz.mem_1729_sv2v_reg ,\nz.mem_1728_sv2v_reg ,\nz.mem_1727_sv2v_reg ,\nz.mem_1726_sv2v_reg ,
  \nz.mem_1725_sv2v_reg ,\nz.mem_1724_sv2v_reg ,\nz.mem_1723_sv2v_reg ,
  \nz.mem_1722_sv2v_reg ,\nz.mem_1721_sv2v_reg ,\nz.mem_1720_sv2v_reg ,\nz.mem_1719_sv2v_reg ,
  \nz.mem_1718_sv2v_reg ,\nz.mem_1717_sv2v_reg ,\nz.mem_1716_sv2v_reg ,
  \nz.mem_1715_sv2v_reg ,\nz.mem_1714_sv2v_reg ,\nz.mem_1713_sv2v_reg ,\nz.mem_1712_sv2v_reg ,
  \nz.mem_1711_sv2v_reg ,\nz.mem_1710_sv2v_reg ,\nz.mem_1709_sv2v_reg ,
  \nz.mem_1708_sv2v_reg ,\nz.mem_1707_sv2v_reg ,\nz.mem_1706_sv2v_reg ,\nz.mem_1705_sv2v_reg ,
  \nz.mem_1704_sv2v_reg ,\nz.mem_1703_sv2v_reg ,\nz.mem_1702_sv2v_reg ,
  \nz.mem_1701_sv2v_reg ,\nz.mem_1700_sv2v_reg ,\nz.mem_1699_sv2v_reg ,\nz.mem_1698_sv2v_reg ,
  \nz.mem_1697_sv2v_reg ,\nz.mem_1696_sv2v_reg ,\nz.mem_1695_sv2v_reg ,
  \nz.mem_1694_sv2v_reg ,\nz.mem_1693_sv2v_reg ,\nz.mem_1692_sv2v_reg ,\nz.mem_1691_sv2v_reg ,
  \nz.mem_1690_sv2v_reg ,\nz.mem_1689_sv2v_reg ,\nz.mem_1688_sv2v_reg ,
  \nz.mem_1687_sv2v_reg ,\nz.mem_1686_sv2v_reg ,\nz.mem_1685_sv2v_reg ,\nz.mem_1684_sv2v_reg ,
  \nz.mem_1683_sv2v_reg ,\nz.mem_1682_sv2v_reg ,\nz.mem_1681_sv2v_reg ,
  \nz.mem_1680_sv2v_reg ,\nz.mem_1679_sv2v_reg ,\nz.mem_1678_sv2v_reg ,\nz.mem_1677_sv2v_reg ,
  \nz.mem_1676_sv2v_reg ,\nz.mem_1675_sv2v_reg ,\nz.mem_1674_sv2v_reg ,
  \nz.mem_1673_sv2v_reg ,\nz.mem_1672_sv2v_reg ,\nz.mem_1671_sv2v_reg ,\nz.mem_1670_sv2v_reg ,
  \nz.mem_1669_sv2v_reg ,\nz.mem_1668_sv2v_reg ,\nz.mem_1667_sv2v_reg ,
  \nz.mem_1666_sv2v_reg ,\nz.mem_1665_sv2v_reg ,\nz.mem_1664_sv2v_reg ,\nz.mem_1663_sv2v_reg ,
  \nz.mem_1662_sv2v_reg ,\nz.mem_1661_sv2v_reg ,\nz.mem_1660_sv2v_reg ,
  \nz.mem_1659_sv2v_reg ,\nz.mem_1658_sv2v_reg ,\nz.mem_1657_sv2v_reg ,\nz.mem_1656_sv2v_reg ,
  \nz.mem_1655_sv2v_reg ,\nz.mem_1654_sv2v_reg ,\nz.mem_1653_sv2v_reg ,
  \nz.mem_1652_sv2v_reg ,\nz.mem_1651_sv2v_reg ,\nz.mem_1650_sv2v_reg ,
  \nz.mem_1649_sv2v_reg ,\nz.mem_1648_sv2v_reg ,\nz.mem_1647_sv2v_reg ,\nz.mem_1646_sv2v_reg ,
  \nz.mem_1645_sv2v_reg ,\nz.mem_1644_sv2v_reg ,\nz.mem_1643_sv2v_reg ,
  \nz.mem_1642_sv2v_reg ,\nz.mem_1641_sv2v_reg ,\nz.mem_1640_sv2v_reg ,\nz.mem_1639_sv2v_reg ,
  \nz.mem_1638_sv2v_reg ,\nz.mem_1637_sv2v_reg ,\nz.mem_1636_sv2v_reg ,
  \nz.mem_1635_sv2v_reg ,\nz.mem_1634_sv2v_reg ,\nz.mem_1633_sv2v_reg ,\nz.mem_1632_sv2v_reg ,
  \nz.mem_1631_sv2v_reg ,\nz.mem_1630_sv2v_reg ,\nz.mem_1629_sv2v_reg ,
  \nz.mem_1628_sv2v_reg ,\nz.mem_1627_sv2v_reg ,\nz.mem_1626_sv2v_reg ,\nz.mem_1625_sv2v_reg ,
  \nz.mem_1624_sv2v_reg ,\nz.mem_1623_sv2v_reg ,\nz.mem_1622_sv2v_reg ,
  \nz.mem_1621_sv2v_reg ,\nz.mem_1620_sv2v_reg ,\nz.mem_1619_sv2v_reg ,\nz.mem_1618_sv2v_reg ,
  \nz.mem_1617_sv2v_reg ,\nz.mem_1616_sv2v_reg ,\nz.mem_1615_sv2v_reg ,
  \nz.mem_1614_sv2v_reg ,\nz.mem_1613_sv2v_reg ,\nz.mem_1612_sv2v_reg ,\nz.mem_1611_sv2v_reg ,
  \nz.mem_1610_sv2v_reg ,\nz.mem_1609_sv2v_reg ,\nz.mem_1608_sv2v_reg ,
  \nz.mem_1607_sv2v_reg ,\nz.mem_1606_sv2v_reg ,\nz.mem_1605_sv2v_reg ,\nz.mem_1604_sv2v_reg ,
  \nz.mem_1603_sv2v_reg ,\nz.mem_1602_sv2v_reg ,\nz.mem_1601_sv2v_reg ,
  \nz.mem_1600_sv2v_reg ,\nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,
  \nz.mem_1596_sv2v_reg ,\nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,
  \nz.mem_1593_sv2v_reg ,\nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,
  \nz.mem_1589_sv2v_reg ,\nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,
  \nz.mem_1586_sv2v_reg ,\nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,
  \nz.mem_1582_sv2v_reg ,\nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,
  \nz.mem_1579_sv2v_reg ,\nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,
  \nz.mem_1575_sv2v_reg ,\nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,
  \nz.mem_1572_sv2v_reg ,\nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,
  \nz.mem_1569_sv2v_reg ,\nz.mem_1568_sv2v_reg ,\nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,
  \nz.mem_1565_sv2v_reg ,\nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,
  \nz.mem_1562_sv2v_reg ,\nz.mem_1561_sv2v_reg ,\nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,
  \nz.mem_1558_sv2v_reg ,\nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,
  \nz.mem_1555_sv2v_reg ,\nz.mem_1554_sv2v_reg ,\nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,
  \nz.mem_1551_sv2v_reg ,\nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,
  \nz.mem_1548_sv2v_reg ,\nz.mem_1547_sv2v_reg ,\nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,
  \nz.mem_1544_sv2v_reg ,\nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,
  \nz.mem_1541_sv2v_reg ,\nz.mem_1540_sv2v_reg ,\nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,
  \nz.mem_1537_sv2v_reg ,\nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,
  \nz.mem_1534_sv2v_reg ,\nz.mem_1533_sv2v_reg ,\nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,
  \nz.mem_1530_sv2v_reg ,\nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,
  \nz.mem_1527_sv2v_reg ,\nz.mem_1526_sv2v_reg ,\nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,
  \nz.mem_1523_sv2v_reg ,\nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,
  \nz.mem_1520_sv2v_reg ,\nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,
  \nz.mem_1516_sv2v_reg ,\nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,
  \nz.mem_1513_sv2v_reg ,\nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,
  \nz.mem_1509_sv2v_reg ,\nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,
  \nz.mem_1506_sv2v_reg ,\nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,
  \nz.mem_1502_sv2v_reg ,\nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,
  \nz.mem_1499_sv2v_reg ,\nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,
  \nz.mem_1495_sv2v_reg ,\nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,
  \nz.mem_1492_sv2v_reg ,\nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,
  \nz.mem_1489_sv2v_reg ,\nz.mem_1488_sv2v_reg ,\nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,
  \nz.mem_1485_sv2v_reg ,\nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,
  \nz.mem_1482_sv2v_reg ,\nz.mem_1481_sv2v_reg ,\nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,
  \nz.mem_1478_sv2v_reg ,\nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,
  \nz.mem_1475_sv2v_reg ,\nz.mem_1474_sv2v_reg ,\nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,
  \nz.mem_1471_sv2v_reg ,\nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,
  \nz.mem_1468_sv2v_reg ,\nz.mem_1467_sv2v_reg ,\nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,
  \nz.mem_1464_sv2v_reg ,\nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,
  \nz.mem_1461_sv2v_reg ,\nz.mem_1460_sv2v_reg ,\nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,
  \nz.mem_1457_sv2v_reg ,\nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,
  \nz.mem_1454_sv2v_reg ,\nz.mem_1453_sv2v_reg ,\nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,
  \nz.mem_1450_sv2v_reg ,\nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,
  \nz.mem_1447_sv2v_reg ,\nz.mem_1446_sv2v_reg ,\nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,
  \nz.mem_1443_sv2v_reg ,\nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,
  \nz.mem_1440_sv2v_reg ,\nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,
  \nz.mem_1436_sv2v_reg ,\nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,
  \nz.mem_1433_sv2v_reg ,\nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,
  \nz.mem_1429_sv2v_reg ,\nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,
  \nz.mem_1426_sv2v_reg ,\nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,
  \nz.mem_1422_sv2v_reg ,\nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,
  \nz.mem_1419_sv2v_reg ,\nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,
  \nz.mem_1415_sv2v_reg ,\nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,
  \nz.mem_1412_sv2v_reg ,\nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,
  \nz.mem_1409_sv2v_reg ,\nz.mem_1408_sv2v_reg ,\nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,
  \nz.mem_1405_sv2v_reg ,\nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,
  \nz.mem_1402_sv2v_reg ,\nz.mem_1401_sv2v_reg ,\nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,
  \nz.mem_1398_sv2v_reg ,\nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,
  \nz.mem_1395_sv2v_reg ,\nz.mem_1394_sv2v_reg ,\nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,
  \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,
  \nz.mem_1388_sv2v_reg ,\nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,
  \nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,
  \nz.mem_1381_sv2v_reg ,\nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,
  \nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,
  \nz.mem_1374_sv2v_reg ,\nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,
  \nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,
  \nz.mem_1367_sv2v_reg ,\nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,
  \nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,
  \nz.mem_1360_sv2v_reg ,\nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,
  \nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,
  \nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,
  \nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,
  \nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,
  \nz.mem_1329_sv2v_reg ,\nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,
  \nz.mem_1322_sv2v_reg ,\nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,
  \nz.mem_1315_sv2v_reg ,\nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,
  \nz.mem_1308_sv2v_reg ,\nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,
  \nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,
  \nz.mem_1301_sv2v_reg ,\nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,
  \nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,
  \nz.mem_1294_sv2v_reg ,\nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,
  \nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,
  \nz.mem_1287_sv2v_reg ,\nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,
  \nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,
  \nz.mem_1280_sv2v_reg ,\nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,
  \nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,
  \nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,
  \nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,
  \nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,
  \nz.mem_1249_sv2v_reg ,\nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,
  \nz.mem_1242_sv2v_reg ,\nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,
  \nz.mem_1235_sv2v_reg ,\nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,
  \nz.mem_1228_sv2v_reg ,\nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,
  \nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,
  \nz.mem_1221_sv2v_reg ,\nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,
  \nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,
  \nz.mem_1214_sv2v_reg ,\nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,
  \nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,
  \nz.mem_1207_sv2v_reg ,\nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,
  \nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,
  \nz.mem_1200_sv2v_reg ,\nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,
  \nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,
  \nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,
  \nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,
  \nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,
  \nz.mem_1169_sv2v_reg ,\nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,
  \nz.mem_1162_sv2v_reg ,\nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,
  \nz.mem_1155_sv2v_reg ,\nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,
  \nz.mem_1148_sv2v_reg ,\nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,
  \nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,
  \nz.mem_1141_sv2v_reg ,\nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,
  \nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,
  \nz.mem_1134_sv2v_reg ,\nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,
  \nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,
  \nz.mem_1127_sv2v_reg ,\nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,
  \nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,
  \nz.mem_1120_sv2v_reg ,\nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,
  \nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,
  \nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,
  \nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,
  \nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,
  \nz.mem_1089_sv2v_reg ,\nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,
  \nz.mem_1082_sv2v_reg ,\nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,
  \nz.mem_1075_sv2v_reg ,\nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,
  \nz.mem_1068_sv2v_reg ,\nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,
  \nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,
  \nz.mem_1061_sv2v_reg ,\nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,
  \nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,
  \nz.mem_1054_sv2v_reg ,\nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,
  \nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,
  \nz.mem_1047_sv2v_reg ,\nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,
  \nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,
  \nz.mem_1040_sv2v_reg ,\nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,
  \nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,
  \nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,
  \nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,
  \nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,
  \nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,
  \nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,
  \nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,
  \nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,
  \nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,
  \nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,
  \nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,
  \nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,
  \nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,
  \nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,
  \nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,
  \nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,
  \nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,
  \nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,
  \nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,
  \nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,
  \nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,
  \nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,
  \nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,
  \nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,
  \nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,
  \nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,
  \nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,
  \nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,
  \nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,
  \nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,
  \nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,
  \nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,
  \nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,
  \nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,
  \nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,
  \nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,
  \nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,
  \nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,
  \nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,
  \nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,
  \nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,
  \nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,
  \nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,
  \nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,
  \nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,
  \nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,
  \nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,
  \nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,
  \nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,
  \nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,
  \nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,
  \nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,
  \nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,
  \nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,
  \nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,
  \nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,
  \nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,
  \nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,
  \nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,
  \nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,
  \nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,
  \nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,
  \nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,
  \nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,
  \nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,
  \nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,
  \nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,
  \nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,
  \nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,
  \nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,
  \nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,
  \nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,
  \nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,
  \nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,
  \nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,
  \nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,
  \nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,
  \nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,
  \nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,
  \nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,
  \nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,
  \nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,
  \nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,
  \nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,
  \nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,
  \nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,
  \nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,
  \nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,
  \nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,
  \nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,
  \nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,
  \nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,
  \nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,
  \nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,
  \nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,
  \nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,
  \nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,
  \nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,
  \nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,
  \nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,
  \nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,
  \nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,
  \nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,
  \nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,
  \nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,
  \nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,
  \nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,
  \nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,
  \nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,
  \nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,
  \nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,
  \nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,
  \nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,
  \nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,
  \nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,
  \nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,
  \nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,
  \nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,
  \nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,
  \nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,
  \nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,
  \nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,
  \nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,
  \nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,
  \nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,
  \nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,
  \nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,
  \nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,
  \nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,
  \nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,
  \nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,
  \nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,
  \nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,
  \nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,
  \nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,
  \nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,
  \nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,
  \nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,
  \nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,
  \nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,
  \nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,
  \nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,
  \nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,
  \nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,
  \nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [7] = \nz.addr_r_7_sv2v_reg ;
  assign \nz.addr_r [6] = \nz.addr_r_6_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [2047] = \nz.mem_2047_sv2v_reg ;
  assign \nz.mem [2046] = \nz.mem_2046_sv2v_reg ;
  assign \nz.mem [2045] = \nz.mem_2045_sv2v_reg ;
  assign \nz.mem [2044] = \nz.mem_2044_sv2v_reg ;
  assign \nz.mem [2043] = \nz.mem_2043_sv2v_reg ;
  assign \nz.mem [2042] = \nz.mem_2042_sv2v_reg ;
  assign \nz.mem [2041] = \nz.mem_2041_sv2v_reg ;
  assign \nz.mem [2040] = \nz.mem_2040_sv2v_reg ;
  assign \nz.mem [2039] = \nz.mem_2039_sv2v_reg ;
  assign \nz.mem [2038] = \nz.mem_2038_sv2v_reg ;
  assign \nz.mem [2037] = \nz.mem_2037_sv2v_reg ;
  assign \nz.mem [2036] = \nz.mem_2036_sv2v_reg ;
  assign \nz.mem [2035] = \nz.mem_2035_sv2v_reg ;
  assign \nz.mem [2034] = \nz.mem_2034_sv2v_reg ;
  assign \nz.mem [2033] = \nz.mem_2033_sv2v_reg ;
  assign \nz.mem [2032] = \nz.mem_2032_sv2v_reg ;
  assign \nz.mem [2031] = \nz.mem_2031_sv2v_reg ;
  assign \nz.mem [2030] = \nz.mem_2030_sv2v_reg ;
  assign \nz.mem [2029] = \nz.mem_2029_sv2v_reg ;
  assign \nz.mem [2028] = \nz.mem_2028_sv2v_reg ;
  assign \nz.mem [2027] = \nz.mem_2027_sv2v_reg ;
  assign \nz.mem [2026] = \nz.mem_2026_sv2v_reg ;
  assign \nz.mem [2025] = \nz.mem_2025_sv2v_reg ;
  assign \nz.mem [2024] = \nz.mem_2024_sv2v_reg ;
  assign \nz.mem [2023] = \nz.mem_2023_sv2v_reg ;
  assign \nz.mem [2022] = \nz.mem_2022_sv2v_reg ;
  assign \nz.mem [2021] = \nz.mem_2021_sv2v_reg ;
  assign \nz.mem [2020] = \nz.mem_2020_sv2v_reg ;
  assign \nz.mem [2019] = \nz.mem_2019_sv2v_reg ;
  assign \nz.mem [2018] = \nz.mem_2018_sv2v_reg ;
  assign \nz.mem [2017] = \nz.mem_2017_sv2v_reg ;
  assign \nz.mem [2016] = \nz.mem_2016_sv2v_reg ;
  assign \nz.mem [2015] = \nz.mem_2015_sv2v_reg ;
  assign \nz.mem [2014] = \nz.mem_2014_sv2v_reg ;
  assign \nz.mem [2013] = \nz.mem_2013_sv2v_reg ;
  assign \nz.mem [2012] = \nz.mem_2012_sv2v_reg ;
  assign \nz.mem [2011] = \nz.mem_2011_sv2v_reg ;
  assign \nz.mem [2010] = \nz.mem_2010_sv2v_reg ;
  assign \nz.mem [2009] = \nz.mem_2009_sv2v_reg ;
  assign \nz.mem [2008] = \nz.mem_2008_sv2v_reg ;
  assign \nz.mem [2007] = \nz.mem_2007_sv2v_reg ;
  assign \nz.mem [2006] = \nz.mem_2006_sv2v_reg ;
  assign \nz.mem [2005] = \nz.mem_2005_sv2v_reg ;
  assign \nz.mem [2004] = \nz.mem_2004_sv2v_reg ;
  assign \nz.mem [2003] = \nz.mem_2003_sv2v_reg ;
  assign \nz.mem [2002] = \nz.mem_2002_sv2v_reg ;
  assign \nz.mem [2001] = \nz.mem_2001_sv2v_reg ;
  assign \nz.mem [2000] = \nz.mem_2000_sv2v_reg ;
  assign \nz.mem [1999] = \nz.mem_1999_sv2v_reg ;
  assign \nz.mem [1998] = \nz.mem_1998_sv2v_reg ;
  assign \nz.mem [1997] = \nz.mem_1997_sv2v_reg ;
  assign \nz.mem [1996] = \nz.mem_1996_sv2v_reg ;
  assign \nz.mem [1995] = \nz.mem_1995_sv2v_reg ;
  assign \nz.mem [1994] = \nz.mem_1994_sv2v_reg ;
  assign \nz.mem [1993] = \nz.mem_1993_sv2v_reg ;
  assign \nz.mem [1992] = \nz.mem_1992_sv2v_reg ;
  assign \nz.mem [1991] = \nz.mem_1991_sv2v_reg ;
  assign \nz.mem [1990] = \nz.mem_1990_sv2v_reg ;
  assign \nz.mem [1989] = \nz.mem_1989_sv2v_reg ;
  assign \nz.mem [1988] = \nz.mem_1988_sv2v_reg ;
  assign \nz.mem [1987] = \nz.mem_1987_sv2v_reg ;
  assign \nz.mem [1986] = \nz.mem_1986_sv2v_reg ;
  assign \nz.mem [1985] = \nz.mem_1985_sv2v_reg ;
  assign \nz.mem [1984] = \nz.mem_1984_sv2v_reg ;
  assign \nz.mem [1983] = \nz.mem_1983_sv2v_reg ;
  assign \nz.mem [1982] = \nz.mem_1982_sv2v_reg ;
  assign \nz.mem [1981] = \nz.mem_1981_sv2v_reg ;
  assign \nz.mem [1980] = \nz.mem_1980_sv2v_reg ;
  assign \nz.mem [1979] = \nz.mem_1979_sv2v_reg ;
  assign \nz.mem [1978] = \nz.mem_1978_sv2v_reg ;
  assign \nz.mem [1977] = \nz.mem_1977_sv2v_reg ;
  assign \nz.mem [1976] = \nz.mem_1976_sv2v_reg ;
  assign \nz.mem [1975] = \nz.mem_1975_sv2v_reg ;
  assign \nz.mem [1974] = \nz.mem_1974_sv2v_reg ;
  assign \nz.mem [1973] = \nz.mem_1973_sv2v_reg ;
  assign \nz.mem [1972] = \nz.mem_1972_sv2v_reg ;
  assign \nz.mem [1971] = \nz.mem_1971_sv2v_reg ;
  assign \nz.mem [1970] = \nz.mem_1970_sv2v_reg ;
  assign \nz.mem [1969] = \nz.mem_1969_sv2v_reg ;
  assign \nz.mem [1968] = \nz.mem_1968_sv2v_reg ;
  assign \nz.mem [1967] = \nz.mem_1967_sv2v_reg ;
  assign \nz.mem [1966] = \nz.mem_1966_sv2v_reg ;
  assign \nz.mem [1965] = \nz.mem_1965_sv2v_reg ;
  assign \nz.mem [1964] = \nz.mem_1964_sv2v_reg ;
  assign \nz.mem [1963] = \nz.mem_1963_sv2v_reg ;
  assign \nz.mem [1962] = \nz.mem_1962_sv2v_reg ;
  assign \nz.mem [1961] = \nz.mem_1961_sv2v_reg ;
  assign \nz.mem [1960] = \nz.mem_1960_sv2v_reg ;
  assign \nz.mem [1959] = \nz.mem_1959_sv2v_reg ;
  assign \nz.mem [1958] = \nz.mem_1958_sv2v_reg ;
  assign \nz.mem [1957] = \nz.mem_1957_sv2v_reg ;
  assign \nz.mem [1956] = \nz.mem_1956_sv2v_reg ;
  assign \nz.mem [1955] = \nz.mem_1955_sv2v_reg ;
  assign \nz.mem [1954] = \nz.mem_1954_sv2v_reg ;
  assign \nz.mem [1953] = \nz.mem_1953_sv2v_reg ;
  assign \nz.mem [1952] = \nz.mem_1952_sv2v_reg ;
  assign \nz.mem [1951] = \nz.mem_1951_sv2v_reg ;
  assign \nz.mem [1950] = \nz.mem_1950_sv2v_reg ;
  assign \nz.mem [1949] = \nz.mem_1949_sv2v_reg ;
  assign \nz.mem [1948] = \nz.mem_1948_sv2v_reg ;
  assign \nz.mem [1947] = \nz.mem_1947_sv2v_reg ;
  assign \nz.mem [1946] = \nz.mem_1946_sv2v_reg ;
  assign \nz.mem [1945] = \nz.mem_1945_sv2v_reg ;
  assign \nz.mem [1944] = \nz.mem_1944_sv2v_reg ;
  assign \nz.mem [1943] = \nz.mem_1943_sv2v_reg ;
  assign \nz.mem [1942] = \nz.mem_1942_sv2v_reg ;
  assign \nz.mem [1941] = \nz.mem_1941_sv2v_reg ;
  assign \nz.mem [1940] = \nz.mem_1940_sv2v_reg ;
  assign \nz.mem [1939] = \nz.mem_1939_sv2v_reg ;
  assign \nz.mem [1938] = \nz.mem_1938_sv2v_reg ;
  assign \nz.mem [1937] = \nz.mem_1937_sv2v_reg ;
  assign \nz.mem [1936] = \nz.mem_1936_sv2v_reg ;
  assign \nz.mem [1935] = \nz.mem_1935_sv2v_reg ;
  assign \nz.mem [1934] = \nz.mem_1934_sv2v_reg ;
  assign \nz.mem [1933] = \nz.mem_1933_sv2v_reg ;
  assign \nz.mem [1932] = \nz.mem_1932_sv2v_reg ;
  assign \nz.mem [1931] = \nz.mem_1931_sv2v_reg ;
  assign \nz.mem [1930] = \nz.mem_1930_sv2v_reg ;
  assign \nz.mem [1929] = \nz.mem_1929_sv2v_reg ;
  assign \nz.mem [1928] = \nz.mem_1928_sv2v_reg ;
  assign \nz.mem [1927] = \nz.mem_1927_sv2v_reg ;
  assign \nz.mem [1926] = \nz.mem_1926_sv2v_reg ;
  assign \nz.mem [1925] = \nz.mem_1925_sv2v_reg ;
  assign \nz.mem [1924] = \nz.mem_1924_sv2v_reg ;
  assign \nz.mem [1923] = \nz.mem_1923_sv2v_reg ;
  assign \nz.mem [1922] = \nz.mem_1922_sv2v_reg ;
  assign \nz.mem [1921] = \nz.mem_1921_sv2v_reg ;
  assign \nz.mem [1920] = \nz.mem_1920_sv2v_reg ;
  assign \nz.mem [1919] = \nz.mem_1919_sv2v_reg ;
  assign \nz.mem [1918] = \nz.mem_1918_sv2v_reg ;
  assign \nz.mem [1917] = \nz.mem_1917_sv2v_reg ;
  assign \nz.mem [1916] = \nz.mem_1916_sv2v_reg ;
  assign \nz.mem [1915] = \nz.mem_1915_sv2v_reg ;
  assign \nz.mem [1914] = \nz.mem_1914_sv2v_reg ;
  assign \nz.mem [1913] = \nz.mem_1913_sv2v_reg ;
  assign \nz.mem [1912] = \nz.mem_1912_sv2v_reg ;
  assign \nz.mem [1911] = \nz.mem_1911_sv2v_reg ;
  assign \nz.mem [1910] = \nz.mem_1910_sv2v_reg ;
  assign \nz.mem [1909] = \nz.mem_1909_sv2v_reg ;
  assign \nz.mem [1908] = \nz.mem_1908_sv2v_reg ;
  assign \nz.mem [1907] = \nz.mem_1907_sv2v_reg ;
  assign \nz.mem [1906] = \nz.mem_1906_sv2v_reg ;
  assign \nz.mem [1905] = \nz.mem_1905_sv2v_reg ;
  assign \nz.mem [1904] = \nz.mem_1904_sv2v_reg ;
  assign \nz.mem [1903] = \nz.mem_1903_sv2v_reg ;
  assign \nz.mem [1902] = \nz.mem_1902_sv2v_reg ;
  assign \nz.mem [1901] = \nz.mem_1901_sv2v_reg ;
  assign \nz.mem [1900] = \nz.mem_1900_sv2v_reg ;
  assign \nz.mem [1899] = \nz.mem_1899_sv2v_reg ;
  assign \nz.mem [1898] = \nz.mem_1898_sv2v_reg ;
  assign \nz.mem [1897] = \nz.mem_1897_sv2v_reg ;
  assign \nz.mem [1896] = \nz.mem_1896_sv2v_reg ;
  assign \nz.mem [1895] = \nz.mem_1895_sv2v_reg ;
  assign \nz.mem [1894] = \nz.mem_1894_sv2v_reg ;
  assign \nz.mem [1893] = \nz.mem_1893_sv2v_reg ;
  assign \nz.mem [1892] = \nz.mem_1892_sv2v_reg ;
  assign \nz.mem [1891] = \nz.mem_1891_sv2v_reg ;
  assign \nz.mem [1890] = \nz.mem_1890_sv2v_reg ;
  assign \nz.mem [1889] = \nz.mem_1889_sv2v_reg ;
  assign \nz.mem [1888] = \nz.mem_1888_sv2v_reg ;
  assign \nz.mem [1887] = \nz.mem_1887_sv2v_reg ;
  assign \nz.mem [1886] = \nz.mem_1886_sv2v_reg ;
  assign \nz.mem [1885] = \nz.mem_1885_sv2v_reg ;
  assign \nz.mem [1884] = \nz.mem_1884_sv2v_reg ;
  assign \nz.mem [1883] = \nz.mem_1883_sv2v_reg ;
  assign \nz.mem [1882] = \nz.mem_1882_sv2v_reg ;
  assign \nz.mem [1881] = \nz.mem_1881_sv2v_reg ;
  assign \nz.mem [1880] = \nz.mem_1880_sv2v_reg ;
  assign \nz.mem [1879] = \nz.mem_1879_sv2v_reg ;
  assign \nz.mem [1878] = \nz.mem_1878_sv2v_reg ;
  assign \nz.mem [1877] = \nz.mem_1877_sv2v_reg ;
  assign \nz.mem [1876] = \nz.mem_1876_sv2v_reg ;
  assign \nz.mem [1875] = \nz.mem_1875_sv2v_reg ;
  assign \nz.mem [1874] = \nz.mem_1874_sv2v_reg ;
  assign \nz.mem [1873] = \nz.mem_1873_sv2v_reg ;
  assign \nz.mem [1872] = \nz.mem_1872_sv2v_reg ;
  assign \nz.mem [1871] = \nz.mem_1871_sv2v_reg ;
  assign \nz.mem [1870] = \nz.mem_1870_sv2v_reg ;
  assign \nz.mem [1869] = \nz.mem_1869_sv2v_reg ;
  assign \nz.mem [1868] = \nz.mem_1868_sv2v_reg ;
  assign \nz.mem [1867] = \nz.mem_1867_sv2v_reg ;
  assign \nz.mem [1866] = \nz.mem_1866_sv2v_reg ;
  assign \nz.mem [1865] = \nz.mem_1865_sv2v_reg ;
  assign \nz.mem [1864] = \nz.mem_1864_sv2v_reg ;
  assign \nz.mem [1863] = \nz.mem_1863_sv2v_reg ;
  assign \nz.mem [1862] = \nz.mem_1862_sv2v_reg ;
  assign \nz.mem [1861] = \nz.mem_1861_sv2v_reg ;
  assign \nz.mem [1860] = \nz.mem_1860_sv2v_reg ;
  assign \nz.mem [1859] = \nz.mem_1859_sv2v_reg ;
  assign \nz.mem [1858] = \nz.mem_1858_sv2v_reg ;
  assign \nz.mem [1857] = \nz.mem_1857_sv2v_reg ;
  assign \nz.mem [1856] = \nz.mem_1856_sv2v_reg ;
  assign \nz.mem [1855] = \nz.mem_1855_sv2v_reg ;
  assign \nz.mem [1854] = \nz.mem_1854_sv2v_reg ;
  assign \nz.mem [1853] = \nz.mem_1853_sv2v_reg ;
  assign \nz.mem [1852] = \nz.mem_1852_sv2v_reg ;
  assign \nz.mem [1851] = \nz.mem_1851_sv2v_reg ;
  assign \nz.mem [1850] = \nz.mem_1850_sv2v_reg ;
  assign \nz.mem [1849] = \nz.mem_1849_sv2v_reg ;
  assign \nz.mem [1848] = \nz.mem_1848_sv2v_reg ;
  assign \nz.mem [1847] = \nz.mem_1847_sv2v_reg ;
  assign \nz.mem [1846] = \nz.mem_1846_sv2v_reg ;
  assign \nz.mem [1845] = \nz.mem_1845_sv2v_reg ;
  assign \nz.mem [1844] = \nz.mem_1844_sv2v_reg ;
  assign \nz.mem [1843] = \nz.mem_1843_sv2v_reg ;
  assign \nz.mem [1842] = \nz.mem_1842_sv2v_reg ;
  assign \nz.mem [1841] = \nz.mem_1841_sv2v_reg ;
  assign \nz.mem [1840] = \nz.mem_1840_sv2v_reg ;
  assign \nz.mem [1839] = \nz.mem_1839_sv2v_reg ;
  assign \nz.mem [1838] = \nz.mem_1838_sv2v_reg ;
  assign \nz.mem [1837] = \nz.mem_1837_sv2v_reg ;
  assign \nz.mem [1836] = \nz.mem_1836_sv2v_reg ;
  assign \nz.mem [1835] = \nz.mem_1835_sv2v_reg ;
  assign \nz.mem [1834] = \nz.mem_1834_sv2v_reg ;
  assign \nz.mem [1833] = \nz.mem_1833_sv2v_reg ;
  assign \nz.mem [1832] = \nz.mem_1832_sv2v_reg ;
  assign \nz.mem [1831] = \nz.mem_1831_sv2v_reg ;
  assign \nz.mem [1830] = \nz.mem_1830_sv2v_reg ;
  assign \nz.mem [1829] = \nz.mem_1829_sv2v_reg ;
  assign \nz.mem [1828] = \nz.mem_1828_sv2v_reg ;
  assign \nz.mem [1827] = \nz.mem_1827_sv2v_reg ;
  assign \nz.mem [1826] = \nz.mem_1826_sv2v_reg ;
  assign \nz.mem [1825] = \nz.mem_1825_sv2v_reg ;
  assign \nz.mem [1824] = \nz.mem_1824_sv2v_reg ;
  assign \nz.mem [1823] = \nz.mem_1823_sv2v_reg ;
  assign \nz.mem [1822] = \nz.mem_1822_sv2v_reg ;
  assign \nz.mem [1821] = \nz.mem_1821_sv2v_reg ;
  assign \nz.mem [1820] = \nz.mem_1820_sv2v_reg ;
  assign \nz.mem [1819] = \nz.mem_1819_sv2v_reg ;
  assign \nz.mem [1818] = \nz.mem_1818_sv2v_reg ;
  assign \nz.mem [1817] = \nz.mem_1817_sv2v_reg ;
  assign \nz.mem [1816] = \nz.mem_1816_sv2v_reg ;
  assign \nz.mem [1815] = \nz.mem_1815_sv2v_reg ;
  assign \nz.mem [1814] = \nz.mem_1814_sv2v_reg ;
  assign \nz.mem [1813] = \nz.mem_1813_sv2v_reg ;
  assign \nz.mem [1812] = \nz.mem_1812_sv2v_reg ;
  assign \nz.mem [1811] = \nz.mem_1811_sv2v_reg ;
  assign \nz.mem [1810] = \nz.mem_1810_sv2v_reg ;
  assign \nz.mem [1809] = \nz.mem_1809_sv2v_reg ;
  assign \nz.mem [1808] = \nz.mem_1808_sv2v_reg ;
  assign \nz.mem [1807] = \nz.mem_1807_sv2v_reg ;
  assign \nz.mem [1806] = \nz.mem_1806_sv2v_reg ;
  assign \nz.mem [1805] = \nz.mem_1805_sv2v_reg ;
  assign \nz.mem [1804] = \nz.mem_1804_sv2v_reg ;
  assign \nz.mem [1803] = \nz.mem_1803_sv2v_reg ;
  assign \nz.mem [1802] = \nz.mem_1802_sv2v_reg ;
  assign \nz.mem [1801] = \nz.mem_1801_sv2v_reg ;
  assign \nz.mem [1800] = \nz.mem_1800_sv2v_reg ;
  assign \nz.mem [1799] = \nz.mem_1799_sv2v_reg ;
  assign \nz.mem [1798] = \nz.mem_1798_sv2v_reg ;
  assign \nz.mem [1797] = \nz.mem_1797_sv2v_reg ;
  assign \nz.mem [1796] = \nz.mem_1796_sv2v_reg ;
  assign \nz.mem [1795] = \nz.mem_1795_sv2v_reg ;
  assign \nz.mem [1794] = \nz.mem_1794_sv2v_reg ;
  assign \nz.mem [1793] = \nz.mem_1793_sv2v_reg ;
  assign \nz.mem [1792] = \nz.mem_1792_sv2v_reg ;
  assign \nz.mem [1791] = \nz.mem_1791_sv2v_reg ;
  assign \nz.mem [1790] = \nz.mem_1790_sv2v_reg ;
  assign \nz.mem [1789] = \nz.mem_1789_sv2v_reg ;
  assign \nz.mem [1788] = \nz.mem_1788_sv2v_reg ;
  assign \nz.mem [1787] = \nz.mem_1787_sv2v_reg ;
  assign \nz.mem [1786] = \nz.mem_1786_sv2v_reg ;
  assign \nz.mem [1785] = \nz.mem_1785_sv2v_reg ;
  assign \nz.mem [1784] = \nz.mem_1784_sv2v_reg ;
  assign \nz.mem [1783] = \nz.mem_1783_sv2v_reg ;
  assign \nz.mem [1782] = \nz.mem_1782_sv2v_reg ;
  assign \nz.mem [1781] = \nz.mem_1781_sv2v_reg ;
  assign \nz.mem [1780] = \nz.mem_1780_sv2v_reg ;
  assign \nz.mem [1779] = \nz.mem_1779_sv2v_reg ;
  assign \nz.mem [1778] = \nz.mem_1778_sv2v_reg ;
  assign \nz.mem [1777] = \nz.mem_1777_sv2v_reg ;
  assign \nz.mem [1776] = \nz.mem_1776_sv2v_reg ;
  assign \nz.mem [1775] = \nz.mem_1775_sv2v_reg ;
  assign \nz.mem [1774] = \nz.mem_1774_sv2v_reg ;
  assign \nz.mem [1773] = \nz.mem_1773_sv2v_reg ;
  assign \nz.mem [1772] = \nz.mem_1772_sv2v_reg ;
  assign \nz.mem [1771] = \nz.mem_1771_sv2v_reg ;
  assign \nz.mem [1770] = \nz.mem_1770_sv2v_reg ;
  assign \nz.mem [1769] = \nz.mem_1769_sv2v_reg ;
  assign \nz.mem [1768] = \nz.mem_1768_sv2v_reg ;
  assign \nz.mem [1767] = \nz.mem_1767_sv2v_reg ;
  assign \nz.mem [1766] = \nz.mem_1766_sv2v_reg ;
  assign \nz.mem [1765] = \nz.mem_1765_sv2v_reg ;
  assign \nz.mem [1764] = \nz.mem_1764_sv2v_reg ;
  assign \nz.mem [1763] = \nz.mem_1763_sv2v_reg ;
  assign \nz.mem [1762] = \nz.mem_1762_sv2v_reg ;
  assign \nz.mem [1761] = \nz.mem_1761_sv2v_reg ;
  assign \nz.mem [1760] = \nz.mem_1760_sv2v_reg ;
  assign \nz.mem [1759] = \nz.mem_1759_sv2v_reg ;
  assign \nz.mem [1758] = \nz.mem_1758_sv2v_reg ;
  assign \nz.mem [1757] = \nz.mem_1757_sv2v_reg ;
  assign \nz.mem [1756] = \nz.mem_1756_sv2v_reg ;
  assign \nz.mem [1755] = \nz.mem_1755_sv2v_reg ;
  assign \nz.mem [1754] = \nz.mem_1754_sv2v_reg ;
  assign \nz.mem [1753] = \nz.mem_1753_sv2v_reg ;
  assign \nz.mem [1752] = \nz.mem_1752_sv2v_reg ;
  assign \nz.mem [1751] = \nz.mem_1751_sv2v_reg ;
  assign \nz.mem [1750] = \nz.mem_1750_sv2v_reg ;
  assign \nz.mem [1749] = \nz.mem_1749_sv2v_reg ;
  assign \nz.mem [1748] = \nz.mem_1748_sv2v_reg ;
  assign \nz.mem [1747] = \nz.mem_1747_sv2v_reg ;
  assign \nz.mem [1746] = \nz.mem_1746_sv2v_reg ;
  assign \nz.mem [1745] = \nz.mem_1745_sv2v_reg ;
  assign \nz.mem [1744] = \nz.mem_1744_sv2v_reg ;
  assign \nz.mem [1743] = \nz.mem_1743_sv2v_reg ;
  assign \nz.mem [1742] = \nz.mem_1742_sv2v_reg ;
  assign \nz.mem [1741] = \nz.mem_1741_sv2v_reg ;
  assign \nz.mem [1740] = \nz.mem_1740_sv2v_reg ;
  assign \nz.mem [1739] = \nz.mem_1739_sv2v_reg ;
  assign \nz.mem [1738] = \nz.mem_1738_sv2v_reg ;
  assign \nz.mem [1737] = \nz.mem_1737_sv2v_reg ;
  assign \nz.mem [1736] = \nz.mem_1736_sv2v_reg ;
  assign \nz.mem [1735] = \nz.mem_1735_sv2v_reg ;
  assign \nz.mem [1734] = \nz.mem_1734_sv2v_reg ;
  assign \nz.mem [1733] = \nz.mem_1733_sv2v_reg ;
  assign \nz.mem [1732] = \nz.mem_1732_sv2v_reg ;
  assign \nz.mem [1731] = \nz.mem_1731_sv2v_reg ;
  assign \nz.mem [1730] = \nz.mem_1730_sv2v_reg ;
  assign \nz.mem [1729] = \nz.mem_1729_sv2v_reg ;
  assign \nz.mem [1728] = \nz.mem_1728_sv2v_reg ;
  assign \nz.mem [1727] = \nz.mem_1727_sv2v_reg ;
  assign \nz.mem [1726] = \nz.mem_1726_sv2v_reg ;
  assign \nz.mem [1725] = \nz.mem_1725_sv2v_reg ;
  assign \nz.mem [1724] = \nz.mem_1724_sv2v_reg ;
  assign \nz.mem [1723] = \nz.mem_1723_sv2v_reg ;
  assign \nz.mem [1722] = \nz.mem_1722_sv2v_reg ;
  assign \nz.mem [1721] = \nz.mem_1721_sv2v_reg ;
  assign \nz.mem [1720] = \nz.mem_1720_sv2v_reg ;
  assign \nz.mem [1719] = \nz.mem_1719_sv2v_reg ;
  assign \nz.mem [1718] = \nz.mem_1718_sv2v_reg ;
  assign \nz.mem [1717] = \nz.mem_1717_sv2v_reg ;
  assign \nz.mem [1716] = \nz.mem_1716_sv2v_reg ;
  assign \nz.mem [1715] = \nz.mem_1715_sv2v_reg ;
  assign \nz.mem [1714] = \nz.mem_1714_sv2v_reg ;
  assign \nz.mem [1713] = \nz.mem_1713_sv2v_reg ;
  assign \nz.mem [1712] = \nz.mem_1712_sv2v_reg ;
  assign \nz.mem [1711] = \nz.mem_1711_sv2v_reg ;
  assign \nz.mem [1710] = \nz.mem_1710_sv2v_reg ;
  assign \nz.mem [1709] = \nz.mem_1709_sv2v_reg ;
  assign \nz.mem [1708] = \nz.mem_1708_sv2v_reg ;
  assign \nz.mem [1707] = \nz.mem_1707_sv2v_reg ;
  assign \nz.mem [1706] = \nz.mem_1706_sv2v_reg ;
  assign \nz.mem [1705] = \nz.mem_1705_sv2v_reg ;
  assign \nz.mem [1704] = \nz.mem_1704_sv2v_reg ;
  assign \nz.mem [1703] = \nz.mem_1703_sv2v_reg ;
  assign \nz.mem [1702] = \nz.mem_1702_sv2v_reg ;
  assign \nz.mem [1701] = \nz.mem_1701_sv2v_reg ;
  assign \nz.mem [1700] = \nz.mem_1700_sv2v_reg ;
  assign \nz.mem [1699] = \nz.mem_1699_sv2v_reg ;
  assign \nz.mem [1698] = \nz.mem_1698_sv2v_reg ;
  assign \nz.mem [1697] = \nz.mem_1697_sv2v_reg ;
  assign \nz.mem [1696] = \nz.mem_1696_sv2v_reg ;
  assign \nz.mem [1695] = \nz.mem_1695_sv2v_reg ;
  assign \nz.mem [1694] = \nz.mem_1694_sv2v_reg ;
  assign \nz.mem [1693] = \nz.mem_1693_sv2v_reg ;
  assign \nz.mem [1692] = \nz.mem_1692_sv2v_reg ;
  assign \nz.mem [1691] = \nz.mem_1691_sv2v_reg ;
  assign \nz.mem [1690] = \nz.mem_1690_sv2v_reg ;
  assign \nz.mem [1689] = \nz.mem_1689_sv2v_reg ;
  assign \nz.mem [1688] = \nz.mem_1688_sv2v_reg ;
  assign \nz.mem [1687] = \nz.mem_1687_sv2v_reg ;
  assign \nz.mem [1686] = \nz.mem_1686_sv2v_reg ;
  assign \nz.mem [1685] = \nz.mem_1685_sv2v_reg ;
  assign \nz.mem [1684] = \nz.mem_1684_sv2v_reg ;
  assign \nz.mem [1683] = \nz.mem_1683_sv2v_reg ;
  assign \nz.mem [1682] = \nz.mem_1682_sv2v_reg ;
  assign \nz.mem [1681] = \nz.mem_1681_sv2v_reg ;
  assign \nz.mem [1680] = \nz.mem_1680_sv2v_reg ;
  assign \nz.mem [1679] = \nz.mem_1679_sv2v_reg ;
  assign \nz.mem [1678] = \nz.mem_1678_sv2v_reg ;
  assign \nz.mem [1677] = \nz.mem_1677_sv2v_reg ;
  assign \nz.mem [1676] = \nz.mem_1676_sv2v_reg ;
  assign \nz.mem [1675] = \nz.mem_1675_sv2v_reg ;
  assign \nz.mem [1674] = \nz.mem_1674_sv2v_reg ;
  assign \nz.mem [1673] = \nz.mem_1673_sv2v_reg ;
  assign \nz.mem [1672] = \nz.mem_1672_sv2v_reg ;
  assign \nz.mem [1671] = \nz.mem_1671_sv2v_reg ;
  assign \nz.mem [1670] = \nz.mem_1670_sv2v_reg ;
  assign \nz.mem [1669] = \nz.mem_1669_sv2v_reg ;
  assign \nz.mem [1668] = \nz.mem_1668_sv2v_reg ;
  assign \nz.mem [1667] = \nz.mem_1667_sv2v_reg ;
  assign \nz.mem [1666] = \nz.mem_1666_sv2v_reg ;
  assign \nz.mem [1665] = \nz.mem_1665_sv2v_reg ;
  assign \nz.mem [1664] = \nz.mem_1664_sv2v_reg ;
  assign \nz.mem [1663] = \nz.mem_1663_sv2v_reg ;
  assign \nz.mem [1662] = \nz.mem_1662_sv2v_reg ;
  assign \nz.mem [1661] = \nz.mem_1661_sv2v_reg ;
  assign \nz.mem [1660] = \nz.mem_1660_sv2v_reg ;
  assign \nz.mem [1659] = \nz.mem_1659_sv2v_reg ;
  assign \nz.mem [1658] = \nz.mem_1658_sv2v_reg ;
  assign \nz.mem [1657] = \nz.mem_1657_sv2v_reg ;
  assign \nz.mem [1656] = \nz.mem_1656_sv2v_reg ;
  assign \nz.mem [1655] = \nz.mem_1655_sv2v_reg ;
  assign \nz.mem [1654] = \nz.mem_1654_sv2v_reg ;
  assign \nz.mem [1653] = \nz.mem_1653_sv2v_reg ;
  assign \nz.mem [1652] = \nz.mem_1652_sv2v_reg ;
  assign \nz.mem [1651] = \nz.mem_1651_sv2v_reg ;
  assign \nz.mem [1650] = \nz.mem_1650_sv2v_reg ;
  assign \nz.mem [1649] = \nz.mem_1649_sv2v_reg ;
  assign \nz.mem [1648] = \nz.mem_1648_sv2v_reg ;
  assign \nz.mem [1647] = \nz.mem_1647_sv2v_reg ;
  assign \nz.mem [1646] = \nz.mem_1646_sv2v_reg ;
  assign \nz.mem [1645] = \nz.mem_1645_sv2v_reg ;
  assign \nz.mem [1644] = \nz.mem_1644_sv2v_reg ;
  assign \nz.mem [1643] = \nz.mem_1643_sv2v_reg ;
  assign \nz.mem [1642] = \nz.mem_1642_sv2v_reg ;
  assign \nz.mem [1641] = \nz.mem_1641_sv2v_reg ;
  assign \nz.mem [1640] = \nz.mem_1640_sv2v_reg ;
  assign \nz.mem [1639] = \nz.mem_1639_sv2v_reg ;
  assign \nz.mem [1638] = \nz.mem_1638_sv2v_reg ;
  assign \nz.mem [1637] = \nz.mem_1637_sv2v_reg ;
  assign \nz.mem [1636] = \nz.mem_1636_sv2v_reg ;
  assign \nz.mem [1635] = \nz.mem_1635_sv2v_reg ;
  assign \nz.mem [1634] = \nz.mem_1634_sv2v_reg ;
  assign \nz.mem [1633] = \nz.mem_1633_sv2v_reg ;
  assign \nz.mem [1632] = \nz.mem_1632_sv2v_reg ;
  assign \nz.mem [1631] = \nz.mem_1631_sv2v_reg ;
  assign \nz.mem [1630] = \nz.mem_1630_sv2v_reg ;
  assign \nz.mem [1629] = \nz.mem_1629_sv2v_reg ;
  assign \nz.mem [1628] = \nz.mem_1628_sv2v_reg ;
  assign \nz.mem [1627] = \nz.mem_1627_sv2v_reg ;
  assign \nz.mem [1626] = \nz.mem_1626_sv2v_reg ;
  assign \nz.mem [1625] = \nz.mem_1625_sv2v_reg ;
  assign \nz.mem [1624] = \nz.mem_1624_sv2v_reg ;
  assign \nz.mem [1623] = \nz.mem_1623_sv2v_reg ;
  assign \nz.mem [1622] = \nz.mem_1622_sv2v_reg ;
  assign \nz.mem [1621] = \nz.mem_1621_sv2v_reg ;
  assign \nz.mem [1620] = \nz.mem_1620_sv2v_reg ;
  assign \nz.mem [1619] = \nz.mem_1619_sv2v_reg ;
  assign \nz.mem [1618] = \nz.mem_1618_sv2v_reg ;
  assign \nz.mem [1617] = \nz.mem_1617_sv2v_reg ;
  assign \nz.mem [1616] = \nz.mem_1616_sv2v_reg ;
  assign \nz.mem [1615] = \nz.mem_1615_sv2v_reg ;
  assign \nz.mem [1614] = \nz.mem_1614_sv2v_reg ;
  assign \nz.mem [1613] = \nz.mem_1613_sv2v_reg ;
  assign \nz.mem [1612] = \nz.mem_1612_sv2v_reg ;
  assign \nz.mem [1611] = \nz.mem_1611_sv2v_reg ;
  assign \nz.mem [1610] = \nz.mem_1610_sv2v_reg ;
  assign \nz.mem [1609] = \nz.mem_1609_sv2v_reg ;
  assign \nz.mem [1608] = \nz.mem_1608_sv2v_reg ;
  assign \nz.mem [1607] = \nz.mem_1607_sv2v_reg ;
  assign \nz.mem [1606] = \nz.mem_1606_sv2v_reg ;
  assign \nz.mem [1605] = \nz.mem_1605_sv2v_reg ;
  assign \nz.mem [1604] = \nz.mem_1604_sv2v_reg ;
  assign \nz.mem [1603] = \nz.mem_1603_sv2v_reg ;
  assign \nz.mem [1602] = \nz.mem_1602_sv2v_reg ;
  assign \nz.mem [1601] = \nz.mem_1601_sv2v_reg ;
  assign \nz.mem [1600] = \nz.mem_1600_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [7] = (N277)? \nz.mem [7] : 
                            (N279)? \nz.mem [15] : 
                            (N281)? \nz.mem [23] : 
                            (N283)? \nz.mem [31] : 
                            (N285)? \nz.mem [39] : 
                            (N287)? \nz.mem [47] : 
                            (N289)? \nz.mem [55] : 
                            (N291)? \nz.mem [63] : 
                            (N293)? \nz.mem [71] : 
                            (N295)? \nz.mem [79] : 
                            (N297)? \nz.mem [87] : 
                            (N299)? \nz.mem [95] : 
                            (N301)? \nz.mem [103] : 
                            (N303)? \nz.mem [111] : 
                            (N305)? \nz.mem [119] : 
                            (N307)? \nz.mem [127] : 
                            (N309)? \nz.mem [135] : 
                            (N311)? \nz.mem [143] : 
                            (N313)? \nz.mem [151] : 
                            (N315)? \nz.mem [159] : 
                            (N317)? \nz.mem [167] : 
                            (N319)? \nz.mem [175] : 
                            (N321)? \nz.mem [183] : 
                            (N323)? \nz.mem [191] : 
                            (N325)? \nz.mem [199] : 
                            (N327)? \nz.mem [207] : 
                            (N329)? \nz.mem [215] : 
                            (N331)? \nz.mem [223] : 
                            (N333)? \nz.mem [231] : 
                            (N335)? \nz.mem [239] : 
                            (N337)? \nz.mem [247] : 
                            (N339)? \nz.mem [255] : 
                            (N341)? \nz.mem [263] : 
                            (N343)? \nz.mem [271] : 
                            (N345)? \nz.mem [279] : 
                            (N347)? \nz.mem [287] : 
                            (N349)? \nz.mem [295] : 
                            (N351)? \nz.mem [303] : 
                            (N353)? \nz.mem [311] : 
                            (N355)? \nz.mem [319] : 
                            (N357)? \nz.mem [327] : 
                            (N359)? \nz.mem [335] : 
                            (N361)? \nz.mem [343] : 
                            (N363)? \nz.mem [351] : 
                            (N365)? \nz.mem [359] : 
                            (N367)? \nz.mem [367] : 
                            (N369)? \nz.mem [375] : 
                            (N371)? \nz.mem [383] : 
                            (N373)? \nz.mem [391] : 
                            (N375)? \nz.mem [399] : 
                            (N377)? \nz.mem [407] : 
                            (N379)? \nz.mem [415] : 
                            (N381)? \nz.mem [423] : 
                            (N383)? \nz.mem [431] : 
                            (N385)? \nz.mem [439] : 
                            (N387)? \nz.mem [447] : 
                            (N389)? \nz.mem [455] : 
                            (N391)? \nz.mem [463] : 
                            (N393)? \nz.mem [471] : 
                            (N395)? \nz.mem [479] : 
                            (N397)? \nz.mem [487] : 
                            (N399)? \nz.mem [495] : 
                            (N401)? \nz.mem [503] : 
                            (N403)? \nz.mem [511] : 
                            (N405)? \nz.mem [519] : 
                            (N407)? \nz.mem [527] : 
                            (N409)? \nz.mem [535] : 
                            (N411)? \nz.mem [543] : 
                            (N413)? \nz.mem [551] : 
                            (N415)? \nz.mem [559] : 
                            (N417)? \nz.mem [567] : 
                            (N419)? \nz.mem [575] : 
                            (N421)? \nz.mem [583] : 
                            (N423)? \nz.mem [591] : 
                            (N425)? \nz.mem [599] : 
                            (N427)? \nz.mem [607] : 
                            (N429)? \nz.mem [615] : 
                            (N431)? \nz.mem [623] : 
                            (N433)? \nz.mem [631] : 
                            (N435)? \nz.mem [639] : 
                            (N437)? \nz.mem [647] : 
                            (N439)? \nz.mem [655] : 
                            (N441)? \nz.mem [663] : 
                            (N443)? \nz.mem [671] : 
                            (N445)? \nz.mem [679] : 
                            (N447)? \nz.mem [687] : 
                            (N449)? \nz.mem [695] : 
                            (N451)? \nz.mem [703] : 
                            (N453)? \nz.mem [711] : 
                            (N455)? \nz.mem [719] : 
                            (N457)? \nz.mem [727] : 
                            (N459)? \nz.mem [735] : 
                            (N461)? \nz.mem [743] : 
                            (N463)? \nz.mem [751] : 
                            (N465)? \nz.mem [759] : 
                            (N467)? \nz.mem [767] : 
                            (N469)? \nz.mem [775] : 
                            (N471)? \nz.mem [783] : 
                            (N473)? \nz.mem [791] : 
                            (N475)? \nz.mem [799] : 
                            (N477)? \nz.mem [807] : 
                            (N479)? \nz.mem [815] : 
                            (N481)? \nz.mem [823] : 
                            (N483)? \nz.mem [831] : 
                            (N485)? \nz.mem [839] : 
                            (N487)? \nz.mem [847] : 
                            (N489)? \nz.mem [855] : 
                            (N491)? \nz.mem [863] : 
                            (N493)? \nz.mem [871] : 
                            (N495)? \nz.mem [879] : 
                            (N497)? \nz.mem [887] : 
                            (N499)? \nz.mem [895] : 
                            (N501)? \nz.mem [903] : 
                            (N503)? \nz.mem [911] : 
                            (N505)? \nz.mem [919] : 
                            (N507)? \nz.mem [927] : 
                            (N509)? \nz.mem [935] : 
                            (N511)? \nz.mem [943] : 
                            (N513)? \nz.mem [951] : 
                            (N515)? \nz.mem [959] : 
                            (N517)? \nz.mem [967] : 
                            (N519)? \nz.mem [975] : 
                            (N521)? \nz.mem [983] : 
                            (N523)? \nz.mem [991] : 
                            (N525)? \nz.mem [999] : 
                            (N527)? \nz.mem [1007] : 
                            (N529)? \nz.mem [1015] : 
                            (N531)? \nz.mem [1023] : 
                            (N278)? \nz.mem [1031] : 
                            (N280)? \nz.mem [1039] : 
                            (N282)? \nz.mem [1047] : 
                            (N284)? \nz.mem [1055] : 
                            (N286)? \nz.mem [1063] : 
                            (N288)? \nz.mem [1071] : 
                            (N290)? \nz.mem [1079] : 
                            (N292)? \nz.mem [1087] : 
                            (N294)? \nz.mem [1095] : 
                            (N296)? \nz.mem [1103] : 
                            (N298)? \nz.mem [1111] : 
                            (N300)? \nz.mem [1119] : 
                            (N302)? \nz.mem [1127] : 
                            (N304)? \nz.mem [1135] : 
                            (N306)? \nz.mem [1143] : 
                            (N308)? \nz.mem [1151] : 
                            (N310)? \nz.mem [1159] : 
                            (N312)? \nz.mem [1167] : 
                            (N314)? \nz.mem [1175] : 
                            (N316)? \nz.mem [1183] : 
                            (N318)? \nz.mem [1191] : 
                            (N320)? \nz.mem [1199] : 
                            (N322)? \nz.mem [1207] : 
                            (N324)? \nz.mem [1215] : 
                            (N326)? \nz.mem [1223] : 
                            (N328)? \nz.mem [1231] : 
                            (N330)? \nz.mem [1239] : 
                            (N332)? \nz.mem [1247] : 
                            (N334)? \nz.mem [1255] : 
                            (N336)? \nz.mem [1263] : 
                            (N338)? \nz.mem [1271] : 
                            (N340)? \nz.mem [1279] : 
                            (N342)? \nz.mem [1287] : 
                            (N344)? \nz.mem [1295] : 
                            (N346)? \nz.mem [1303] : 
                            (N348)? \nz.mem [1311] : 
                            (N350)? \nz.mem [1319] : 
                            (N352)? \nz.mem [1327] : 
                            (N354)? \nz.mem [1335] : 
                            (N356)? \nz.mem [1343] : 
                            (N358)? \nz.mem [1351] : 
                            (N360)? \nz.mem [1359] : 
                            (N362)? \nz.mem [1367] : 
                            (N364)? \nz.mem [1375] : 
                            (N366)? \nz.mem [1383] : 
                            (N368)? \nz.mem [1391] : 
                            (N370)? \nz.mem [1399] : 
                            (N372)? \nz.mem [1407] : 
                            (N374)? \nz.mem [1415] : 
                            (N376)? \nz.mem [1423] : 
                            (N378)? \nz.mem [1431] : 
                            (N380)? \nz.mem [1439] : 
                            (N382)? \nz.mem [1447] : 
                            (N384)? \nz.mem [1455] : 
                            (N386)? \nz.mem [1463] : 
                            (N388)? \nz.mem [1471] : 
                            (N390)? \nz.mem [1479] : 
                            (N392)? \nz.mem [1487] : 
                            (N394)? \nz.mem [1495] : 
                            (N396)? \nz.mem [1503] : 
                            (N398)? \nz.mem [1511] : 
                            (N400)? \nz.mem [1519] : 
                            (N402)? \nz.mem [1527] : 
                            (N404)? \nz.mem [1535] : 
                            (N406)? \nz.mem [1543] : 
                            (N408)? \nz.mem [1551] : 
                            (N410)? \nz.mem [1559] : 
                            (N412)? \nz.mem [1567] : 
                            (N414)? \nz.mem [1575] : 
                            (N416)? \nz.mem [1583] : 
                            (N418)? \nz.mem [1591] : 
                            (N420)? \nz.mem [1599] : 
                            (N422)? \nz.mem [1607] : 
                            (N424)? \nz.mem [1615] : 
                            (N426)? \nz.mem [1623] : 
                            (N428)? \nz.mem [1631] : 
                            (N430)? \nz.mem [1639] : 
                            (N432)? \nz.mem [1647] : 
                            (N434)? \nz.mem [1655] : 
                            (N436)? \nz.mem [1663] : 
                            (N438)? \nz.mem [1671] : 
                            (N440)? \nz.mem [1679] : 
                            (N442)? \nz.mem [1687] : 
                            (N444)? \nz.mem [1695] : 
                            (N446)? \nz.mem [1703] : 
                            (N448)? \nz.mem [1711] : 
                            (N450)? \nz.mem [1719] : 
                            (N452)? \nz.mem [1727] : 
                            (N454)? \nz.mem [1735] : 
                            (N456)? \nz.mem [1743] : 
                            (N458)? \nz.mem [1751] : 
                            (N460)? \nz.mem [1759] : 
                            (N462)? \nz.mem [1767] : 
                            (N464)? \nz.mem [1775] : 
                            (N466)? \nz.mem [1783] : 
                            (N468)? \nz.mem [1791] : 
                            (N470)? \nz.mem [1799] : 
                            (N472)? \nz.mem [1807] : 
                            (N474)? \nz.mem [1815] : 
                            (N476)? \nz.mem [1823] : 
                            (N478)? \nz.mem [1831] : 
                            (N480)? \nz.mem [1839] : 
                            (N482)? \nz.mem [1847] : 
                            (N484)? \nz.mem [1855] : 
                            (N486)? \nz.mem [1863] : 
                            (N488)? \nz.mem [1871] : 
                            (N490)? \nz.mem [1879] : 
                            (N492)? \nz.mem [1887] : 
                            (N494)? \nz.mem [1895] : 
                            (N496)? \nz.mem [1903] : 
                            (N498)? \nz.mem [1911] : 
                            (N500)? \nz.mem [1919] : 
                            (N502)? \nz.mem [1927] : 
                            (N504)? \nz.mem [1935] : 
                            (N506)? \nz.mem [1943] : 
                            (N508)? \nz.mem [1951] : 
                            (N510)? \nz.mem [1959] : 
                            (N512)? \nz.mem [1967] : 
                            (N514)? \nz.mem [1975] : 
                            (N516)? \nz.mem [1983] : 
                            (N518)? \nz.mem [1991] : 
                            (N520)? \nz.mem [1999] : 
                            (N522)? \nz.mem [2007] : 
                            (N524)? \nz.mem [2015] : 
                            (N526)? \nz.mem [2023] : 
                            (N528)? \nz.mem [2031] : 
                            (N530)? \nz.mem [2039] : 
                            (N532)? \nz.mem [2047] : 1'b0;
  assign \nz.data_out [6] = (N277)? \nz.mem [6] : 
                            (N279)? \nz.mem [14] : 
                            (N281)? \nz.mem [22] : 
                            (N283)? \nz.mem [30] : 
                            (N285)? \nz.mem [38] : 
                            (N287)? \nz.mem [46] : 
                            (N289)? \nz.mem [54] : 
                            (N291)? \nz.mem [62] : 
                            (N293)? \nz.mem [70] : 
                            (N295)? \nz.mem [78] : 
                            (N297)? \nz.mem [86] : 
                            (N299)? \nz.mem [94] : 
                            (N301)? \nz.mem [102] : 
                            (N303)? \nz.mem [110] : 
                            (N305)? \nz.mem [118] : 
                            (N307)? \nz.mem [126] : 
                            (N309)? \nz.mem [134] : 
                            (N311)? \nz.mem [142] : 
                            (N313)? \nz.mem [150] : 
                            (N315)? \nz.mem [158] : 
                            (N317)? \nz.mem [166] : 
                            (N319)? \nz.mem [174] : 
                            (N321)? \nz.mem [182] : 
                            (N323)? \nz.mem [190] : 
                            (N325)? \nz.mem [198] : 
                            (N327)? \nz.mem [206] : 
                            (N329)? \nz.mem [214] : 
                            (N331)? \nz.mem [222] : 
                            (N333)? \nz.mem [230] : 
                            (N335)? \nz.mem [238] : 
                            (N337)? \nz.mem [246] : 
                            (N339)? \nz.mem [254] : 
                            (N341)? \nz.mem [262] : 
                            (N343)? \nz.mem [270] : 
                            (N345)? \nz.mem [278] : 
                            (N347)? \nz.mem [286] : 
                            (N349)? \nz.mem [294] : 
                            (N351)? \nz.mem [302] : 
                            (N353)? \nz.mem [310] : 
                            (N355)? \nz.mem [318] : 
                            (N357)? \nz.mem [326] : 
                            (N359)? \nz.mem [334] : 
                            (N361)? \nz.mem [342] : 
                            (N363)? \nz.mem [350] : 
                            (N365)? \nz.mem [358] : 
                            (N367)? \nz.mem [366] : 
                            (N369)? \nz.mem [374] : 
                            (N371)? \nz.mem [382] : 
                            (N373)? \nz.mem [390] : 
                            (N375)? \nz.mem [398] : 
                            (N377)? \nz.mem [406] : 
                            (N379)? \nz.mem [414] : 
                            (N381)? \nz.mem [422] : 
                            (N383)? \nz.mem [430] : 
                            (N385)? \nz.mem [438] : 
                            (N387)? \nz.mem [446] : 
                            (N389)? \nz.mem [454] : 
                            (N391)? \nz.mem [462] : 
                            (N393)? \nz.mem [470] : 
                            (N395)? \nz.mem [478] : 
                            (N397)? \nz.mem [486] : 
                            (N399)? \nz.mem [494] : 
                            (N401)? \nz.mem [502] : 
                            (N403)? \nz.mem [510] : 
                            (N405)? \nz.mem [518] : 
                            (N407)? \nz.mem [526] : 
                            (N409)? \nz.mem [534] : 
                            (N411)? \nz.mem [542] : 
                            (N413)? \nz.mem [550] : 
                            (N415)? \nz.mem [558] : 
                            (N417)? \nz.mem [566] : 
                            (N419)? \nz.mem [574] : 
                            (N421)? \nz.mem [582] : 
                            (N423)? \nz.mem [590] : 
                            (N425)? \nz.mem [598] : 
                            (N427)? \nz.mem [606] : 
                            (N429)? \nz.mem [614] : 
                            (N431)? \nz.mem [622] : 
                            (N433)? \nz.mem [630] : 
                            (N435)? \nz.mem [638] : 
                            (N437)? \nz.mem [646] : 
                            (N439)? \nz.mem [654] : 
                            (N441)? \nz.mem [662] : 
                            (N443)? \nz.mem [670] : 
                            (N445)? \nz.mem [678] : 
                            (N447)? \nz.mem [686] : 
                            (N449)? \nz.mem [694] : 
                            (N451)? \nz.mem [702] : 
                            (N453)? \nz.mem [710] : 
                            (N455)? \nz.mem [718] : 
                            (N457)? \nz.mem [726] : 
                            (N459)? \nz.mem [734] : 
                            (N461)? \nz.mem [742] : 
                            (N463)? \nz.mem [750] : 
                            (N465)? \nz.mem [758] : 
                            (N467)? \nz.mem [766] : 
                            (N469)? \nz.mem [774] : 
                            (N471)? \nz.mem [782] : 
                            (N473)? \nz.mem [790] : 
                            (N475)? \nz.mem [798] : 
                            (N477)? \nz.mem [806] : 
                            (N479)? \nz.mem [814] : 
                            (N481)? \nz.mem [822] : 
                            (N483)? \nz.mem [830] : 
                            (N485)? \nz.mem [838] : 
                            (N487)? \nz.mem [846] : 
                            (N489)? \nz.mem [854] : 
                            (N491)? \nz.mem [862] : 
                            (N493)? \nz.mem [870] : 
                            (N495)? \nz.mem [878] : 
                            (N497)? \nz.mem [886] : 
                            (N499)? \nz.mem [894] : 
                            (N501)? \nz.mem [902] : 
                            (N503)? \nz.mem [910] : 
                            (N505)? \nz.mem [918] : 
                            (N507)? \nz.mem [926] : 
                            (N509)? \nz.mem [934] : 
                            (N511)? \nz.mem [942] : 
                            (N513)? \nz.mem [950] : 
                            (N515)? \nz.mem [958] : 
                            (N517)? \nz.mem [966] : 
                            (N519)? \nz.mem [974] : 
                            (N521)? \nz.mem [982] : 
                            (N523)? \nz.mem [990] : 
                            (N525)? \nz.mem [998] : 
                            (N527)? \nz.mem [1006] : 
                            (N529)? \nz.mem [1014] : 
                            (N531)? \nz.mem [1022] : 
                            (N278)? \nz.mem [1030] : 
                            (N280)? \nz.mem [1038] : 
                            (N282)? \nz.mem [1046] : 
                            (N284)? \nz.mem [1054] : 
                            (N286)? \nz.mem [1062] : 
                            (N288)? \nz.mem [1070] : 
                            (N290)? \nz.mem [1078] : 
                            (N292)? \nz.mem [1086] : 
                            (N294)? \nz.mem [1094] : 
                            (N296)? \nz.mem [1102] : 
                            (N298)? \nz.mem [1110] : 
                            (N300)? \nz.mem [1118] : 
                            (N302)? \nz.mem [1126] : 
                            (N304)? \nz.mem [1134] : 
                            (N306)? \nz.mem [1142] : 
                            (N308)? \nz.mem [1150] : 
                            (N310)? \nz.mem [1158] : 
                            (N312)? \nz.mem [1166] : 
                            (N314)? \nz.mem [1174] : 
                            (N316)? \nz.mem [1182] : 
                            (N318)? \nz.mem [1190] : 
                            (N320)? \nz.mem [1198] : 
                            (N322)? \nz.mem [1206] : 
                            (N324)? \nz.mem [1214] : 
                            (N326)? \nz.mem [1222] : 
                            (N328)? \nz.mem [1230] : 
                            (N330)? \nz.mem [1238] : 
                            (N332)? \nz.mem [1246] : 
                            (N334)? \nz.mem [1254] : 
                            (N336)? \nz.mem [1262] : 
                            (N338)? \nz.mem [1270] : 
                            (N340)? \nz.mem [1278] : 
                            (N342)? \nz.mem [1286] : 
                            (N344)? \nz.mem [1294] : 
                            (N346)? \nz.mem [1302] : 
                            (N348)? \nz.mem [1310] : 
                            (N350)? \nz.mem [1318] : 
                            (N352)? \nz.mem [1326] : 
                            (N354)? \nz.mem [1334] : 
                            (N356)? \nz.mem [1342] : 
                            (N358)? \nz.mem [1350] : 
                            (N360)? \nz.mem [1358] : 
                            (N362)? \nz.mem [1366] : 
                            (N364)? \nz.mem [1374] : 
                            (N366)? \nz.mem [1382] : 
                            (N368)? \nz.mem [1390] : 
                            (N370)? \nz.mem [1398] : 
                            (N372)? \nz.mem [1406] : 
                            (N374)? \nz.mem [1414] : 
                            (N376)? \nz.mem [1422] : 
                            (N378)? \nz.mem [1430] : 
                            (N380)? \nz.mem [1438] : 
                            (N382)? \nz.mem [1446] : 
                            (N384)? \nz.mem [1454] : 
                            (N386)? \nz.mem [1462] : 
                            (N388)? \nz.mem [1470] : 
                            (N390)? \nz.mem [1478] : 
                            (N392)? \nz.mem [1486] : 
                            (N394)? \nz.mem [1494] : 
                            (N396)? \nz.mem [1502] : 
                            (N398)? \nz.mem [1510] : 
                            (N400)? \nz.mem [1518] : 
                            (N402)? \nz.mem [1526] : 
                            (N404)? \nz.mem [1534] : 
                            (N406)? \nz.mem [1542] : 
                            (N408)? \nz.mem [1550] : 
                            (N410)? \nz.mem [1558] : 
                            (N412)? \nz.mem [1566] : 
                            (N414)? \nz.mem [1574] : 
                            (N416)? \nz.mem [1582] : 
                            (N418)? \nz.mem [1590] : 
                            (N420)? \nz.mem [1598] : 
                            (N422)? \nz.mem [1606] : 
                            (N424)? \nz.mem [1614] : 
                            (N426)? \nz.mem [1622] : 
                            (N428)? \nz.mem [1630] : 
                            (N430)? \nz.mem [1638] : 
                            (N432)? \nz.mem [1646] : 
                            (N434)? \nz.mem [1654] : 
                            (N436)? \nz.mem [1662] : 
                            (N438)? \nz.mem [1670] : 
                            (N440)? \nz.mem [1678] : 
                            (N442)? \nz.mem [1686] : 
                            (N444)? \nz.mem [1694] : 
                            (N446)? \nz.mem [1702] : 
                            (N448)? \nz.mem [1710] : 
                            (N450)? \nz.mem [1718] : 
                            (N452)? \nz.mem [1726] : 
                            (N454)? \nz.mem [1734] : 
                            (N456)? \nz.mem [1742] : 
                            (N458)? \nz.mem [1750] : 
                            (N460)? \nz.mem [1758] : 
                            (N462)? \nz.mem [1766] : 
                            (N464)? \nz.mem [1774] : 
                            (N466)? \nz.mem [1782] : 
                            (N468)? \nz.mem [1790] : 
                            (N470)? \nz.mem [1798] : 
                            (N472)? \nz.mem [1806] : 
                            (N474)? \nz.mem [1814] : 
                            (N476)? \nz.mem [1822] : 
                            (N478)? \nz.mem [1830] : 
                            (N480)? \nz.mem [1838] : 
                            (N482)? \nz.mem [1846] : 
                            (N484)? \nz.mem [1854] : 
                            (N486)? \nz.mem [1862] : 
                            (N488)? \nz.mem [1870] : 
                            (N490)? \nz.mem [1878] : 
                            (N492)? \nz.mem [1886] : 
                            (N494)? \nz.mem [1894] : 
                            (N496)? \nz.mem [1902] : 
                            (N498)? \nz.mem [1910] : 
                            (N500)? \nz.mem [1918] : 
                            (N502)? \nz.mem [1926] : 
                            (N504)? \nz.mem [1934] : 
                            (N506)? \nz.mem [1942] : 
                            (N508)? \nz.mem [1950] : 
                            (N510)? \nz.mem [1958] : 
                            (N512)? \nz.mem [1966] : 
                            (N514)? \nz.mem [1974] : 
                            (N516)? \nz.mem [1982] : 
                            (N518)? \nz.mem [1990] : 
                            (N520)? \nz.mem [1998] : 
                            (N522)? \nz.mem [2006] : 
                            (N524)? \nz.mem [2014] : 
                            (N526)? \nz.mem [2022] : 
                            (N528)? \nz.mem [2030] : 
                            (N530)? \nz.mem [2038] : 
                            (N532)? \nz.mem [2046] : 1'b0;
  assign \nz.data_out [5] = (N277)? \nz.mem [5] : 
                            (N279)? \nz.mem [13] : 
                            (N281)? \nz.mem [21] : 
                            (N283)? \nz.mem [29] : 
                            (N285)? \nz.mem [37] : 
                            (N287)? \nz.mem [45] : 
                            (N289)? \nz.mem [53] : 
                            (N291)? \nz.mem [61] : 
                            (N293)? \nz.mem [69] : 
                            (N295)? \nz.mem [77] : 
                            (N297)? \nz.mem [85] : 
                            (N299)? \nz.mem [93] : 
                            (N301)? \nz.mem [101] : 
                            (N303)? \nz.mem [109] : 
                            (N305)? \nz.mem [117] : 
                            (N307)? \nz.mem [125] : 
                            (N309)? \nz.mem [133] : 
                            (N311)? \nz.mem [141] : 
                            (N313)? \nz.mem [149] : 
                            (N315)? \nz.mem [157] : 
                            (N317)? \nz.mem [165] : 
                            (N319)? \nz.mem [173] : 
                            (N321)? \nz.mem [181] : 
                            (N323)? \nz.mem [189] : 
                            (N325)? \nz.mem [197] : 
                            (N327)? \nz.mem [205] : 
                            (N329)? \nz.mem [213] : 
                            (N331)? \nz.mem [221] : 
                            (N333)? \nz.mem [229] : 
                            (N335)? \nz.mem [237] : 
                            (N337)? \nz.mem [245] : 
                            (N339)? \nz.mem [253] : 
                            (N341)? \nz.mem [261] : 
                            (N343)? \nz.mem [269] : 
                            (N345)? \nz.mem [277] : 
                            (N347)? \nz.mem [285] : 
                            (N349)? \nz.mem [293] : 
                            (N351)? \nz.mem [301] : 
                            (N353)? \nz.mem [309] : 
                            (N355)? \nz.mem [317] : 
                            (N357)? \nz.mem [325] : 
                            (N359)? \nz.mem [333] : 
                            (N361)? \nz.mem [341] : 
                            (N363)? \nz.mem [349] : 
                            (N365)? \nz.mem [357] : 
                            (N367)? \nz.mem [365] : 
                            (N369)? \nz.mem [373] : 
                            (N371)? \nz.mem [381] : 
                            (N373)? \nz.mem [389] : 
                            (N375)? \nz.mem [397] : 
                            (N377)? \nz.mem [405] : 
                            (N379)? \nz.mem [413] : 
                            (N381)? \nz.mem [421] : 
                            (N383)? \nz.mem [429] : 
                            (N385)? \nz.mem [437] : 
                            (N387)? \nz.mem [445] : 
                            (N389)? \nz.mem [453] : 
                            (N391)? \nz.mem [461] : 
                            (N393)? \nz.mem [469] : 
                            (N395)? \nz.mem [477] : 
                            (N397)? \nz.mem [485] : 
                            (N399)? \nz.mem [493] : 
                            (N401)? \nz.mem [501] : 
                            (N403)? \nz.mem [509] : 
                            (N405)? \nz.mem [517] : 
                            (N407)? \nz.mem [525] : 
                            (N409)? \nz.mem [533] : 
                            (N411)? \nz.mem [541] : 
                            (N413)? \nz.mem [549] : 
                            (N415)? \nz.mem [557] : 
                            (N417)? \nz.mem [565] : 
                            (N419)? \nz.mem [573] : 
                            (N421)? \nz.mem [581] : 
                            (N423)? \nz.mem [589] : 
                            (N425)? \nz.mem [597] : 
                            (N427)? \nz.mem [605] : 
                            (N429)? \nz.mem [613] : 
                            (N431)? \nz.mem [621] : 
                            (N433)? \nz.mem [629] : 
                            (N435)? \nz.mem [637] : 
                            (N437)? \nz.mem [645] : 
                            (N439)? \nz.mem [653] : 
                            (N441)? \nz.mem [661] : 
                            (N443)? \nz.mem [669] : 
                            (N445)? \nz.mem [677] : 
                            (N447)? \nz.mem [685] : 
                            (N449)? \nz.mem [693] : 
                            (N451)? \nz.mem [701] : 
                            (N453)? \nz.mem [709] : 
                            (N455)? \nz.mem [717] : 
                            (N457)? \nz.mem [725] : 
                            (N459)? \nz.mem [733] : 
                            (N461)? \nz.mem [741] : 
                            (N463)? \nz.mem [749] : 
                            (N465)? \nz.mem [757] : 
                            (N467)? \nz.mem [765] : 
                            (N469)? \nz.mem [773] : 
                            (N471)? \nz.mem [781] : 
                            (N473)? \nz.mem [789] : 
                            (N475)? \nz.mem [797] : 
                            (N477)? \nz.mem [805] : 
                            (N479)? \nz.mem [813] : 
                            (N481)? \nz.mem [821] : 
                            (N483)? \nz.mem [829] : 
                            (N485)? \nz.mem [837] : 
                            (N487)? \nz.mem [845] : 
                            (N489)? \nz.mem [853] : 
                            (N491)? \nz.mem [861] : 
                            (N493)? \nz.mem [869] : 
                            (N495)? \nz.mem [877] : 
                            (N497)? \nz.mem [885] : 
                            (N499)? \nz.mem [893] : 
                            (N501)? \nz.mem [901] : 
                            (N503)? \nz.mem [909] : 
                            (N505)? \nz.mem [917] : 
                            (N507)? \nz.mem [925] : 
                            (N509)? \nz.mem [933] : 
                            (N511)? \nz.mem [941] : 
                            (N513)? \nz.mem [949] : 
                            (N515)? \nz.mem [957] : 
                            (N517)? \nz.mem [965] : 
                            (N519)? \nz.mem [973] : 
                            (N521)? \nz.mem [981] : 
                            (N523)? \nz.mem [989] : 
                            (N525)? \nz.mem [997] : 
                            (N527)? \nz.mem [1005] : 
                            (N529)? \nz.mem [1013] : 
                            (N531)? \nz.mem [1021] : 
                            (N278)? \nz.mem [1029] : 
                            (N280)? \nz.mem [1037] : 
                            (N282)? \nz.mem [1045] : 
                            (N284)? \nz.mem [1053] : 
                            (N286)? \nz.mem [1061] : 
                            (N288)? \nz.mem [1069] : 
                            (N290)? \nz.mem [1077] : 
                            (N292)? \nz.mem [1085] : 
                            (N294)? \nz.mem [1093] : 
                            (N296)? \nz.mem [1101] : 
                            (N298)? \nz.mem [1109] : 
                            (N300)? \nz.mem [1117] : 
                            (N302)? \nz.mem [1125] : 
                            (N304)? \nz.mem [1133] : 
                            (N306)? \nz.mem [1141] : 
                            (N308)? \nz.mem [1149] : 
                            (N310)? \nz.mem [1157] : 
                            (N312)? \nz.mem [1165] : 
                            (N314)? \nz.mem [1173] : 
                            (N316)? \nz.mem [1181] : 
                            (N318)? \nz.mem [1189] : 
                            (N320)? \nz.mem [1197] : 
                            (N322)? \nz.mem [1205] : 
                            (N324)? \nz.mem [1213] : 
                            (N326)? \nz.mem [1221] : 
                            (N328)? \nz.mem [1229] : 
                            (N330)? \nz.mem [1237] : 
                            (N332)? \nz.mem [1245] : 
                            (N334)? \nz.mem [1253] : 
                            (N336)? \nz.mem [1261] : 
                            (N338)? \nz.mem [1269] : 
                            (N340)? \nz.mem [1277] : 
                            (N342)? \nz.mem [1285] : 
                            (N344)? \nz.mem [1293] : 
                            (N346)? \nz.mem [1301] : 
                            (N348)? \nz.mem [1309] : 
                            (N350)? \nz.mem [1317] : 
                            (N352)? \nz.mem [1325] : 
                            (N354)? \nz.mem [1333] : 
                            (N356)? \nz.mem [1341] : 
                            (N358)? \nz.mem [1349] : 
                            (N360)? \nz.mem [1357] : 
                            (N362)? \nz.mem [1365] : 
                            (N364)? \nz.mem [1373] : 
                            (N366)? \nz.mem [1381] : 
                            (N368)? \nz.mem [1389] : 
                            (N370)? \nz.mem [1397] : 
                            (N372)? \nz.mem [1405] : 
                            (N374)? \nz.mem [1413] : 
                            (N376)? \nz.mem [1421] : 
                            (N378)? \nz.mem [1429] : 
                            (N380)? \nz.mem [1437] : 
                            (N382)? \nz.mem [1445] : 
                            (N384)? \nz.mem [1453] : 
                            (N386)? \nz.mem [1461] : 
                            (N388)? \nz.mem [1469] : 
                            (N390)? \nz.mem [1477] : 
                            (N392)? \nz.mem [1485] : 
                            (N394)? \nz.mem [1493] : 
                            (N396)? \nz.mem [1501] : 
                            (N398)? \nz.mem [1509] : 
                            (N400)? \nz.mem [1517] : 
                            (N402)? \nz.mem [1525] : 
                            (N404)? \nz.mem [1533] : 
                            (N406)? \nz.mem [1541] : 
                            (N408)? \nz.mem [1549] : 
                            (N410)? \nz.mem [1557] : 
                            (N412)? \nz.mem [1565] : 
                            (N414)? \nz.mem [1573] : 
                            (N416)? \nz.mem [1581] : 
                            (N418)? \nz.mem [1589] : 
                            (N420)? \nz.mem [1597] : 
                            (N422)? \nz.mem [1605] : 
                            (N424)? \nz.mem [1613] : 
                            (N426)? \nz.mem [1621] : 
                            (N428)? \nz.mem [1629] : 
                            (N430)? \nz.mem [1637] : 
                            (N432)? \nz.mem [1645] : 
                            (N434)? \nz.mem [1653] : 
                            (N436)? \nz.mem [1661] : 
                            (N438)? \nz.mem [1669] : 
                            (N440)? \nz.mem [1677] : 
                            (N442)? \nz.mem [1685] : 
                            (N444)? \nz.mem [1693] : 
                            (N446)? \nz.mem [1701] : 
                            (N448)? \nz.mem [1709] : 
                            (N450)? \nz.mem [1717] : 
                            (N452)? \nz.mem [1725] : 
                            (N454)? \nz.mem [1733] : 
                            (N456)? \nz.mem [1741] : 
                            (N458)? \nz.mem [1749] : 
                            (N460)? \nz.mem [1757] : 
                            (N462)? \nz.mem [1765] : 
                            (N464)? \nz.mem [1773] : 
                            (N466)? \nz.mem [1781] : 
                            (N468)? \nz.mem [1789] : 
                            (N470)? \nz.mem [1797] : 
                            (N472)? \nz.mem [1805] : 
                            (N474)? \nz.mem [1813] : 
                            (N476)? \nz.mem [1821] : 
                            (N478)? \nz.mem [1829] : 
                            (N480)? \nz.mem [1837] : 
                            (N482)? \nz.mem [1845] : 
                            (N484)? \nz.mem [1853] : 
                            (N486)? \nz.mem [1861] : 
                            (N488)? \nz.mem [1869] : 
                            (N490)? \nz.mem [1877] : 
                            (N492)? \nz.mem [1885] : 
                            (N494)? \nz.mem [1893] : 
                            (N496)? \nz.mem [1901] : 
                            (N498)? \nz.mem [1909] : 
                            (N500)? \nz.mem [1917] : 
                            (N502)? \nz.mem [1925] : 
                            (N504)? \nz.mem [1933] : 
                            (N506)? \nz.mem [1941] : 
                            (N508)? \nz.mem [1949] : 
                            (N510)? \nz.mem [1957] : 
                            (N512)? \nz.mem [1965] : 
                            (N514)? \nz.mem [1973] : 
                            (N516)? \nz.mem [1981] : 
                            (N518)? \nz.mem [1989] : 
                            (N520)? \nz.mem [1997] : 
                            (N522)? \nz.mem [2005] : 
                            (N524)? \nz.mem [2013] : 
                            (N526)? \nz.mem [2021] : 
                            (N528)? \nz.mem [2029] : 
                            (N530)? \nz.mem [2037] : 
                            (N532)? \nz.mem [2045] : 1'b0;
  assign \nz.data_out [4] = (N277)? \nz.mem [4] : 
                            (N279)? \nz.mem [12] : 
                            (N281)? \nz.mem [20] : 
                            (N283)? \nz.mem [28] : 
                            (N285)? \nz.mem [36] : 
                            (N287)? \nz.mem [44] : 
                            (N289)? \nz.mem [52] : 
                            (N291)? \nz.mem [60] : 
                            (N293)? \nz.mem [68] : 
                            (N295)? \nz.mem [76] : 
                            (N297)? \nz.mem [84] : 
                            (N299)? \nz.mem [92] : 
                            (N301)? \nz.mem [100] : 
                            (N303)? \nz.mem [108] : 
                            (N305)? \nz.mem [116] : 
                            (N307)? \nz.mem [124] : 
                            (N309)? \nz.mem [132] : 
                            (N311)? \nz.mem [140] : 
                            (N313)? \nz.mem [148] : 
                            (N315)? \nz.mem [156] : 
                            (N317)? \nz.mem [164] : 
                            (N319)? \nz.mem [172] : 
                            (N321)? \nz.mem [180] : 
                            (N323)? \nz.mem [188] : 
                            (N325)? \nz.mem [196] : 
                            (N327)? \nz.mem [204] : 
                            (N329)? \nz.mem [212] : 
                            (N331)? \nz.mem [220] : 
                            (N333)? \nz.mem [228] : 
                            (N335)? \nz.mem [236] : 
                            (N337)? \nz.mem [244] : 
                            (N339)? \nz.mem [252] : 
                            (N341)? \nz.mem [260] : 
                            (N343)? \nz.mem [268] : 
                            (N345)? \nz.mem [276] : 
                            (N347)? \nz.mem [284] : 
                            (N349)? \nz.mem [292] : 
                            (N351)? \nz.mem [300] : 
                            (N353)? \nz.mem [308] : 
                            (N355)? \nz.mem [316] : 
                            (N357)? \nz.mem [324] : 
                            (N359)? \nz.mem [332] : 
                            (N361)? \nz.mem [340] : 
                            (N363)? \nz.mem [348] : 
                            (N365)? \nz.mem [356] : 
                            (N367)? \nz.mem [364] : 
                            (N369)? \nz.mem [372] : 
                            (N371)? \nz.mem [380] : 
                            (N373)? \nz.mem [388] : 
                            (N375)? \nz.mem [396] : 
                            (N377)? \nz.mem [404] : 
                            (N379)? \nz.mem [412] : 
                            (N381)? \nz.mem [420] : 
                            (N383)? \nz.mem [428] : 
                            (N385)? \nz.mem [436] : 
                            (N387)? \nz.mem [444] : 
                            (N389)? \nz.mem [452] : 
                            (N391)? \nz.mem [460] : 
                            (N393)? \nz.mem [468] : 
                            (N395)? \nz.mem [476] : 
                            (N397)? \nz.mem [484] : 
                            (N399)? \nz.mem [492] : 
                            (N401)? \nz.mem [500] : 
                            (N403)? \nz.mem [508] : 
                            (N405)? \nz.mem [516] : 
                            (N407)? \nz.mem [524] : 
                            (N409)? \nz.mem [532] : 
                            (N411)? \nz.mem [540] : 
                            (N413)? \nz.mem [548] : 
                            (N415)? \nz.mem [556] : 
                            (N417)? \nz.mem [564] : 
                            (N419)? \nz.mem [572] : 
                            (N421)? \nz.mem [580] : 
                            (N423)? \nz.mem [588] : 
                            (N425)? \nz.mem [596] : 
                            (N427)? \nz.mem [604] : 
                            (N429)? \nz.mem [612] : 
                            (N431)? \nz.mem [620] : 
                            (N433)? \nz.mem [628] : 
                            (N435)? \nz.mem [636] : 
                            (N437)? \nz.mem [644] : 
                            (N439)? \nz.mem [652] : 
                            (N441)? \nz.mem [660] : 
                            (N443)? \nz.mem [668] : 
                            (N445)? \nz.mem [676] : 
                            (N447)? \nz.mem [684] : 
                            (N449)? \nz.mem [692] : 
                            (N451)? \nz.mem [700] : 
                            (N453)? \nz.mem [708] : 
                            (N455)? \nz.mem [716] : 
                            (N457)? \nz.mem [724] : 
                            (N459)? \nz.mem [732] : 
                            (N461)? \nz.mem [740] : 
                            (N463)? \nz.mem [748] : 
                            (N465)? \nz.mem [756] : 
                            (N467)? \nz.mem [764] : 
                            (N469)? \nz.mem [772] : 
                            (N471)? \nz.mem [780] : 
                            (N473)? \nz.mem [788] : 
                            (N475)? \nz.mem [796] : 
                            (N477)? \nz.mem [804] : 
                            (N479)? \nz.mem [812] : 
                            (N481)? \nz.mem [820] : 
                            (N483)? \nz.mem [828] : 
                            (N485)? \nz.mem [836] : 
                            (N487)? \nz.mem [844] : 
                            (N489)? \nz.mem [852] : 
                            (N491)? \nz.mem [860] : 
                            (N493)? \nz.mem [868] : 
                            (N495)? \nz.mem [876] : 
                            (N497)? \nz.mem [884] : 
                            (N499)? \nz.mem [892] : 
                            (N501)? \nz.mem [900] : 
                            (N503)? \nz.mem [908] : 
                            (N505)? \nz.mem [916] : 
                            (N507)? \nz.mem [924] : 
                            (N509)? \nz.mem [932] : 
                            (N511)? \nz.mem [940] : 
                            (N513)? \nz.mem [948] : 
                            (N515)? \nz.mem [956] : 
                            (N517)? \nz.mem [964] : 
                            (N519)? \nz.mem [972] : 
                            (N521)? \nz.mem [980] : 
                            (N523)? \nz.mem [988] : 
                            (N525)? \nz.mem [996] : 
                            (N527)? \nz.mem [1004] : 
                            (N529)? \nz.mem [1012] : 
                            (N531)? \nz.mem [1020] : 
                            (N278)? \nz.mem [1028] : 
                            (N280)? \nz.mem [1036] : 
                            (N282)? \nz.mem [1044] : 
                            (N284)? \nz.mem [1052] : 
                            (N286)? \nz.mem [1060] : 
                            (N288)? \nz.mem [1068] : 
                            (N290)? \nz.mem [1076] : 
                            (N292)? \nz.mem [1084] : 
                            (N294)? \nz.mem [1092] : 
                            (N296)? \nz.mem [1100] : 
                            (N298)? \nz.mem [1108] : 
                            (N300)? \nz.mem [1116] : 
                            (N302)? \nz.mem [1124] : 
                            (N304)? \nz.mem [1132] : 
                            (N306)? \nz.mem [1140] : 
                            (N308)? \nz.mem [1148] : 
                            (N310)? \nz.mem [1156] : 
                            (N312)? \nz.mem [1164] : 
                            (N314)? \nz.mem [1172] : 
                            (N316)? \nz.mem [1180] : 
                            (N318)? \nz.mem [1188] : 
                            (N320)? \nz.mem [1196] : 
                            (N322)? \nz.mem [1204] : 
                            (N324)? \nz.mem [1212] : 
                            (N326)? \nz.mem [1220] : 
                            (N328)? \nz.mem [1228] : 
                            (N330)? \nz.mem [1236] : 
                            (N332)? \nz.mem [1244] : 
                            (N334)? \nz.mem [1252] : 
                            (N336)? \nz.mem [1260] : 
                            (N338)? \nz.mem [1268] : 
                            (N340)? \nz.mem [1276] : 
                            (N342)? \nz.mem [1284] : 
                            (N344)? \nz.mem [1292] : 
                            (N346)? \nz.mem [1300] : 
                            (N348)? \nz.mem [1308] : 
                            (N350)? \nz.mem [1316] : 
                            (N352)? \nz.mem [1324] : 
                            (N354)? \nz.mem [1332] : 
                            (N356)? \nz.mem [1340] : 
                            (N358)? \nz.mem [1348] : 
                            (N360)? \nz.mem [1356] : 
                            (N362)? \nz.mem [1364] : 
                            (N364)? \nz.mem [1372] : 
                            (N366)? \nz.mem [1380] : 
                            (N368)? \nz.mem [1388] : 
                            (N370)? \nz.mem [1396] : 
                            (N372)? \nz.mem [1404] : 
                            (N374)? \nz.mem [1412] : 
                            (N376)? \nz.mem [1420] : 
                            (N378)? \nz.mem [1428] : 
                            (N380)? \nz.mem [1436] : 
                            (N382)? \nz.mem [1444] : 
                            (N384)? \nz.mem [1452] : 
                            (N386)? \nz.mem [1460] : 
                            (N388)? \nz.mem [1468] : 
                            (N390)? \nz.mem [1476] : 
                            (N392)? \nz.mem [1484] : 
                            (N394)? \nz.mem [1492] : 
                            (N396)? \nz.mem [1500] : 
                            (N398)? \nz.mem [1508] : 
                            (N400)? \nz.mem [1516] : 
                            (N402)? \nz.mem [1524] : 
                            (N404)? \nz.mem [1532] : 
                            (N406)? \nz.mem [1540] : 
                            (N408)? \nz.mem [1548] : 
                            (N410)? \nz.mem [1556] : 
                            (N412)? \nz.mem [1564] : 
                            (N414)? \nz.mem [1572] : 
                            (N416)? \nz.mem [1580] : 
                            (N418)? \nz.mem [1588] : 
                            (N420)? \nz.mem [1596] : 
                            (N422)? \nz.mem [1604] : 
                            (N424)? \nz.mem [1612] : 
                            (N426)? \nz.mem [1620] : 
                            (N428)? \nz.mem [1628] : 
                            (N430)? \nz.mem [1636] : 
                            (N432)? \nz.mem [1644] : 
                            (N434)? \nz.mem [1652] : 
                            (N436)? \nz.mem [1660] : 
                            (N438)? \nz.mem [1668] : 
                            (N440)? \nz.mem [1676] : 
                            (N442)? \nz.mem [1684] : 
                            (N444)? \nz.mem [1692] : 
                            (N446)? \nz.mem [1700] : 
                            (N448)? \nz.mem [1708] : 
                            (N450)? \nz.mem [1716] : 
                            (N452)? \nz.mem [1724] : 
                            (N454)? \nz.mem [1732] : 
                            (N456)? \nz.mem [1740] : 
                            (N458)? \nz.mem [1748] : 
                            (N460)? \nz.mem [1756] : 
                            (N462)? \nz.mem [1764] : 
                            (N464)? \nz.mem [1772] : 
                            (N466)? \nz.mem [1780] : 
                            (N468)? \nz.mem [1788] : 
                            (N470)? \nz.mem [1796] : 
                            (N472)? \nz.mem [1804] : 
                            (N474)? \nz.mem [1812] : 
                            (N476)? \nz.mem [1820] : 
                            (N478)? \nz.mem [1828] : 
                            (N480)? \nz.mem [1836] : 
                            (N482)? \nz.mem [1844] : 
                            (N484)? \nz.mem [1852] : 
                            (N486)? \nz.mem [1860] : 
                            (N488)? \nz.mem [1868] : 
                            (N490)? \nz.mem [1876] : 
                            (N492)? \nz.mem [1884] : 
                            (N494)? \nz.mem [1892] : 
                            (N496)? \nz.mem [1900] : 
                            (N498)? \nz.mem [1908] : 
                            (N500)? \nz.mem [1916] : 
                            (N502)? \nz.mem [1924] : 
                            (N504)? \nz.mem [1932] : 
                            (N506)? \nz.mem [1940] : 
                            (N508)? \nz.mem [1948] : 
                            (N510)? \nz.mem [1956] : 
                            (N512)? \nz.mem [1964] : 
                            (N514)? \nz.mem [1972] : 
                            (N516)? \nz.mem [1980] : 
                            (N518)? \nz.mem [1988] : 
                            (N520)? \nz.mem [1996] : 
                            (N522)? \nz.mem [2004] : 
                            (N524)? \nz.mem [2012] : 
                            (N526)? \nz.mem [2020] : 
                            (N528)? \nz.mem [2028] : 
                            (N530)? \nz.mem [2036] : 
                            (N532)? \nz.mem [2044] : 1'b0;
  assign \nz.data_out [3] = (N277)? \nz.mem [3] : 
                            (N279)? \nz.mem [11] : 
                            (N281)? \nz.mem [19] : 
                            (N283)? \nz.mem [27] : 
                            (N285)? \nz.mem [35] : 
                            (N287)? \nz.mem [43] : 
                            (N289)? \nz.mem [51] : 
                            (N291)? \nz.mem [59] : 
                            (N293)? \nz.mem [67] : 
                            (N295)? \nz.mem [75] : 
                            (N297)? \nz.mem [83] : 
                            (N299)? \nz.mem [91] : 
                            (N301)? \nz.mem [99] : 
                            (N303)? \nz.mem [107] : 
                            (N305)? \nz.mem [115] : 
                            (N307)? \nz.mem [123] : 
                            (N309)? \nz.mem [131] : 
                            (N311)? \nz.mem [139] : 
                            (N313)? \nz.mem [147] : 
                            (N315)? \nz.mem [155] : 
                            (N317)? \nz.mem [163] : 
                            (N319)? \nz.mem [171] : 
                            (N321)? \nz.mem [179] : 
                            (N323)? \nz.mem [187] : 
                            (N325)? \nz.mem [195] : 
                            (N327)? \nz.mem [203] : 
                            (N329)? \nz.mem [211] : 
                            (N331)? \nz.mem [219] : 
                            (N333)? \nz.mem [227] : 
                            (N335)? \nz.mem [235] : 
                            (N337)? \nz.mem [243] : 
                            (N339)? \nz.mem [251] : 
                            (N341)? \nz.mem [259] : 
                            (N343)? \nz.mem [267] : 
                            (N345)? \nz.mem [275] : 
                            (N347)? \nz.mem [283] : 
                            (N349)? \nz.mem [291] : 
                            (N351)? \nz.mem [299] : 
                            (N353)? \nz.mem [307] : 
                            (N355)? \nz.mem [315] : 
                            (N357)? \nz.mem [323] : 
                            (N359)? \nz.mem [331] : 
                            (N361)? \nz.mem [339] : 
                            (N363)? \nz.mem [347] : 
                            (N365)? \nz.mem [355] : 
                            (N367)? \nz.mem [363] : 
                            (N369)? \nz.mem [371] : 
                            (N371)? \nz.mem [379] : 
                            (N373)? \nz.mem [387] : 
                            (N375)? \nz.mem [395] : 
                            (N377)? \nz.mem [403] : 
                            (N379)? \nz.mem [411] : 
                            (N381)? \nz.mem [419] : 
                            (N383)? \nz.mem [427] : 
                            (N385)? \nz.mem [435] : 
                            (N387)? \nz.mem [443] : 
                            (N389)? \nz.mem [451] : 
                            (N391)? \nz.mem [459] : 
                            (N393)? \nz.mem [467] : 
                            (N395)? \nz.mem [475] : 
                            (N397)? \nz.mem [483] : 
                            (N399)? \nz.mem [491] : 
                            (N401)? \nz.mem [499] : 
                            (N403)? \nz.mem [507] : 
                            (N405)? \nz.mem [515] : 
                            (N407)? \nz.mem [523] : 
                            (N409)? \nz.mem [531] : 
                            (N411)? \nz.mem [539] : 
                            (N413)? \nz.mem [547] : 
                            (N415)? \nz.mem [555] : 
                            (N417)? \nz.mem [563] : 
                            (N419)? \nz.mem [571] : 
                            (N421)? \nz.mem [579] : 
                            (N423)? \nz.mem [587] : 
                            (N425)? \nz.mem [595] : 
                            (N427)? \nz.mem [603] : 
                            (N429)? \nz.mem [611] : 
                            (N431)? \nz.mem [619] : 
                            (N433)? \nz.mem [627] : 
                            (N435)? \nz.mem [635] : 
                            (N437)? \nz.mem [643] : 
                            (N439)? \nz.mem [651] : 
                            (N441)? \nz.mem [659] : 
                            (N443)? \nz.mem [667] : 
                            (N445)? \nz.mem [675] : 
                            (N447)? \nz.mem [683] : 
                            (N449)? \nz.mem [691] : 
                            (N451)? \nz.mem [699] : 
                            (N453)? \nz.mem [707] : 
                            (N455)? \nz.mem [715] : 
                            (N457)? \nz.mem [723] : 
                            (N459)? \nz.mem [731] : 
                            (N461)? \nz.mem [739] : 
                            (N463)? \nz.mem [747] : 
                            (N465)? \nz.mem [755] : 
                            (N467)? \nz.mem [763] : 
                            (N469)? \nz.mem [771] : 
                            (N471)? \nz.mem [779] : 
                            (N473)? \nz.mem [787] : 
                            (N475)? \nz.mem [795] : 
                            (N477)? \nz.mem [803] : 
                            (N479)? \nz.mem [811] : 
                            (N481)? \nz.mem [819] : 
                            (N483)? \nz.mem [827] : 
                            (N485)? \nz.mem [835] : 
                            (N487)? \nz.mem [843] : 
                            (N489)? \nz.mem [851] : 
                            (N491)? \nz.mem [859] : 
                            (N493)? \nz.mem [867] : 
                            (N495)? \nz.mem [875] : 
                            (N497)? \nz.mem [883] : 
                            (N499)? \nz.mem [891] : 
                            (N501)? \nz.mem [899] : 
                            (N503)? \nz.mem [907] : 
                            (N505)? \nz.mem [915] : 
                            (N507)? \nz.mem [923] : 
                            (N509)? \nz.mem [931] : 
                            (N511)? \nz.mem [939] : 
                            (N513)? \nz.mem [947] : 
                            (N515)? \nz.mem [955] : 
                            (N517)? \nz.mem [963] : 
                            (N519)? \nz.mem [971] : 
                            (N521)? \nz.mem [979] : 
                            (N523)? \nz.mem [987] : 
                            (N525)? \nz.mem [995] : 
                            (N527)? \nz.mem [1003] : 
                            (N529)? \nz.mem [1011] : 
                            (N531)? \nz.mem [1019] : 
                            (N278)? \nz.mem [1027] : 
                            (N280)? \nz.mem [1035] : 
                            (N282)? \nz.mem [1043] : 
                            (N284)? \nz.mem [1051] : 
                            (N286)? \nz.mem [1059] : 
                            (N288)? \nz.mem [1067] : 
                            (N290)? \nz.mem [1075] : 
                            (N292)? \nz.mem [1083] : 
                            (N294)? \nz.mem [1091] : 
                            (N296)? \nz.mem [1099] : 
                            (N298)? \nz.mem [1107] : 
                            (N300)? \nz.mem [1115] : 
                            (N302)? \nz.mem [1123] : 
                            (N304)? \nz.mem [1131] : 
                            (N306)? \nz.mem [1139] : 
                            (N308)? \nz.mem [1147] : 
                            (N310)? \nz.mem [1155] : 
                            (N312)? \nz.mem [1163] : 
                            (N314)? \nz.mem [1171] : 
                            (N316)? \nz.mem [1179] : 
                            (N318)? \nz.mem [1187] : 
                            (N320)? \nz.mem [1195] : 
                            (N322)? \nz.mem [1203] : 
                            (N324)? \nz.mem [1211] : 
                            (N326)? \nz.mem [1219] : 
                            (N328)? \nz.mem [1227] : 
                            (N330)? \nz.mem [1235] : 
                            (N332)? \nz.mem [1243] : 
                            (N334)? \nz.mem [1251] : 
                            (N336)? \nz.mem [1259] : 
                            (N338)? \nz.mem [1267] : 
                            (N340)? \nz.mem [1275] : 
                            (N342)? \nz.mem [1283] : 
                            (N344)? \nz.mem [1291] : 
                            (N346)? \nz.mem [1299] : 
                            (N348)? \nz.mem [1307] : 
                            (N350)? \nz.mem [1315] : 
                            (N352)? \nz.mem [1323] : 
                            (N354)? \nz.mem [1331] : 
                            (N356)? \nz.mem [1339] : 
                            (N358)? \nz.mem [1347] : 
                            (N360)? \nz.mem [1355] : 
                            (N362)? \nz.mem [1363] : 
                            (N364)? \nz.mem [1371] : 
                            (N366)? \nz.mem [1379] : 
                            (N368)? \nz.mem [1387] : 
                            (N370)? \nz.mem [1395] : 
                            (N372)? \nz.mem [1403] : 
                            (N374)? \nz.mem [1411] : 
                            (N376)? \nz.mem [1419] : 
                            (N378)? \nz.mem [1427] : 
                            (N380)? \nz.mem [1435] : 
                            (N382)? \nz.mem [1443] : 
                            (N384)? \nz.mem [1451] : 
                            (N386)? \nz.mem [1459] : 
                            (N388)? \nz.mem [1467] : 
                            (N390)? \nz.mem [1475] : 
                            (N392)? \nz.mem [1483] : 
                            (N394)? \nz.mem [1491] : 
                            (N396)? \nz.mem [1499] : 
                            (N398)? \nz.mem [1507] : 
                            (N400)? \nz.mem [1515] : 
                            (N402)? \nz.mem [1523] : 
                            (N404)? \nz.mem [1531] : 
                            (N406)? \nz.mem [1539] : 
                            (N408)? \nz.mem [1547] : 
                            (N410)? \nz.mem [1555] : 
                            (N412)? \nz.mem [1563] : 
                            (N414)? \nz.mem [1571] : 
                            (N416)? \nz.mem [1579] : 
                            (N418)? \nz.mem [1587] : 
                            (N420)? \nz.mem [1595] : 
                            (N422)? \nz.mem [1603] : 
                            (N424)? \nz.mem [1611] : 
                            (N426)? \nz.mem [1619] : 
                            (N428)? \nz.mem [1627] : 
                            (N430)? \nz.mem [1635] : 
                            (N432)? \nz.mem [1643] : 
                            (N434)? \nz.mem [1651] : 
                            (N436)? \nz.mem [1659] : 
                            (N438)? \nz.mem [1667] : 
                            (N440)? \nz.mem [1675] : 
                            (N442)? \nz.mem [1683] : 
                            (N444)? \nz.mem [1691] : 
                            (N446)? \nz.mem [1699] : 
                            (N448)? \nz.mem [1707] : 
                            (N450)? \nz.mem [1715] : 
                            (N452)? \nz.mem [1723] : 
                            (N454)? \nz.mem [1731] : 
                            (N456)? \nz.mem [1739] : 
                            (N458)? \nz.mem [1747] : 
                            (N460)? \nz.mem [1755] : 
                            (N462)? \nz.mem [1763] : 
                            (N464)? \nz.mem [1771] : 
                            (N466)? \nz.mem [1779] : 
                            (N468)? \nz.mem [1787] : 
                            (N470)? \nz.mem [1795] : 
                            (N472)? \nz.mem [1803] : 
                            (N474)? \nz.mem [1811] : 
                            (N476)? \nz.mem [1819] : 
                            (N478)? \nz.mem [1827] : 
                            (N480)? \nz.mem [1835] : 
                            (N482)? \nz.mem [1843] : 
                            (N484)? \nz.mem [1851] : 
                            (N486)? \nz.mem [1859] : 
                            (N488)? \nz.mem [1867] : 
                            (N490)? \nz.mem [1875] : 
                            (N492)? \nz.mem [1883] : 
                            (N494)? \nz.mem [1891] : 
                            (N496)? \nz.mem [1899] : 
                            (N498)? \nz.mem [1907] : 
                            (N500)? \nz.mem [1915] : 
                            (N502)? \nz.mem [1923] : 
                            (N504)? \nz.mem [1931] : 
                            (N506)? \nz.mem [1939] : 
                            (N508)? \nz.mem [1947] : 
                            (N510)? \nz.mem [1955] : 
                            (N512)? \nz.mem [1963] : 
                            (N514)? \nz.mem [1971] : 
                            (N516)? \nz.mem [1979] : 
                            (N518)? \nz.mem [1987] : 
                            (N520)? \nz.mem [1995] : 
                            (N522)? \nz.mem [2003] : 
                            (N524)? \nz.mem [2011] : 
                            (N526)? \nz.mem [2019] : 
                            (N528)? \nz.mem [2027] : 
                            (N530)? \nz.mem [2035] : 
                            (N532)? \nz.mem [2043] : 1'b0;
  assign \nz.data_out [2] = (N277)? \nz.mem [2] : 
                            (N279)? \nz.mem [10] : 
                            (N281)? \nz.mem [18] : 
                            (N283)? \nz.mem [26] : 
                            (N285)? \nz.mem [34] : 
                            (N287)? \nz.mem [42] : 
                            (N289)? \nz.mem [50] : 
                            (N291)? \nz.mem [58] : 
                            (N293)? \nz.mem [66] : 
                            (N295)? \nz.mem [74] : 
                            (N297)? \nz.mem [82] : 
                            (N299)? \nz.mem [90] : 
                            (N301)? \nz.mem [98] : 
                            (N303)? \nz.mem [106] : 
                            (N305)? \nz.mem [114] : 
                            (N307)? \nz.mem [122] : 
                            (N309)? \nz.mem [130] : 
                            (N311)? \nz.mem [138] : 
                            (N313)? \nz.mem [146] : 
                            (N315)? \nz.mem [154] : 
                            (N317)? \nz.mem [162] : 
                            (N319)? \nz.mem [170] : 
                            (N321)? \nz.mem [178] : 
                            (N323)? \nz.mem [186] : 
                            (N325)? \nz.mem [194] : 
                            (N327)? \nz.mem [202] : 
                            (N329)? \nz.mem [210] : 
                            (N331)? \nz.mem [218] : 
                            (N333)? \nz.mem [226] : 
                            (N335)? \nz.mem [234] : 
                            (N337)? \nz.mem [242] : 
                            (N339)? \nz.mem [250] : 
                            (N341)? \nz.mem [258] : 
                            (N343)? \nz.mem [266] : 
                            (N345)? \nz.mem [274] : 
                            (N347)? \nz.mem [282] : 
                            (N349)? \nz.mem [290] : 
                            (N351)? \nz.mem [298] : 
                            (N353)? \nz.mem [306] : 
                            (N355)? \nz.mem [314] : 
                            (N357)? \nz.mem [322] : 
                            (N359)? \nz.mem [330] : 
                            (N361)? \nz.mem [338] : 
                            (N363)? \nz.mem [346] : 
                            (N365)? \nz.mem [354] : 
                            (N367)? \nz.mem [362] : 
                            (N369)? \nz.mem [370] : 
                            (N371)? \nz.mem [378] : 
                            (N373)? \nz.mem [386] : 
                            (N375)? \nz.mem [394] : 
                            (N377)? \nz.mem [402] : 
                            (N379)? \nz.mem [410] : 
                            (N381)? \nz.mem [418] : 
                            (N383)? \nz.mem [426] : 
                            (N385)? \nz.mem [434] : 
                            (N387)? \nz.mem [442] : 
                            (N389)? \nz.mem [450] : 
                            (N391)? \nz.mem [458] : 
                            (N393)? \nz.mem [466] : 
                            (N395)? \nz.mem [474] : 
                            (N397)? \nz.mem [482] : 
                            (N399)? \nz.mem [490] : 
                            (N401)? \nz.mem [498] : 
                            (N403)? \nz.mem [506] : 
                            (N405)? \nz.mem [514] : 
                            (N407)? \nz.mem [522] : 
                            (N409)? \nz.mem [530] : 
                            (N411)? \nz.mem [538] : 
                            (N413)? \nz.mem [546] : 
                            (N415)? \nz.mem [554] : 
                            (N417)? \nz.mem [562] : 
                            (N419)? \nz.mem [570] : 
                            (N421)? \nz.mem [578] : 
                            (N423)? \nz.mem [586] : 
                            (N425)? \nz.mem [594] : 
                            (N427)? \nz.mem [602] : 
                            (N429)? \nz.mem [610] : 
                            (N431)? \nz.mem [618] : 
                            (N433)? \nz.mem [626] : 
                            (N435)? \nz.mem [634] : 
                            (N437)? \nz.mem [642] : 
                            (N439)? \nz.mem [650] : 
                            (N441)? \nz.mem [658] : 
                            (N443)? \nz.mem [666] : 
                            (N445)? \nz.mem [674] : 
                            (N447)? \nz.mem [682] : 
                            (N449)? \nz.mem [690] : 
                            (N451)? \nz.mem [698] : 
                            (N453)? \nz.mem [706] : 
                            (N455)? \nz.mem [714] : 
                            (N457)? \nz.mem [722] : 
                            (N459)? \nz.mem [730] : 
                            (N461)? \nz.mem [738] : 
                            (N463)? \nz.mem [746] : 
                            (N465)? \nz.mem [754] : 
                            (N467)? \nz.mem [762] : 
                            (N469)? \nz.mem [770] : 
                            (N471)? \nz.mem [778] : 
                            (N473)? \nz.mem [786] : 
                            (N475)? \nz.mem [794] : 
                            (N477)? \nz.mem [802] : 
                            (N479)? \nz.mem [810] : 
                            (N481)? \nz.mem [818] : 
                            (N483)? \nz.mem [826] : 
                            (N485)? \nz.mem [834] : 
                            (N487)? \nz.mem [842] : 
                            (N489)? \nz.mem [850] : 
                            (N491)? \nz.mem [858] : 
                            (N493)? \nz.mem [866] : 
                            (N495)? \nz.mem [874] : 
                            (N497)? \nz.mem [882] : 
                            (N499)? \nz.mem [890] : 
                            (N501)? \nz.mem [898] : 
                            (N503)? \nz.mem [906] : 
                            (N505)? \nz.mem [914] : 
                            (N507)? \nz.mem [922] : 
                            (N509)? \nz.mem [930] : 
                            (N511)? \nz.mem [938] : 
                            (N513)? \nz.mem [946] : 
                            (N515)? \nz.mem [954] : 
                            (N517)? \nz.mem [962] : 
                            (N519)? \nz.mem [970] : 
                            (N521)? \nz.mem [978] : 
                            (N523)? \nz.mem [986] : 
                            (N525)? \nz.mem [994] : 
                            (N527)? \nz.mem [1002] : 
                            (N529)? \nz.mem [1010] : 
                            (N531)? \nz.mem [1018] : 
                            (N278)? \nz.mem [1026] : 
                            (N280)? \nz.mem [1034] : 
                            (N282)? \nz.mem [1042] : 
                            (N284)? \nz.mem [1050] : 
                            (N286)? \nz.mem [1058] : 
                            (N288)? \nz.mem [1066] : 
                            (N290)? \nz.mem [1074] : 
                            (N292)? \nz.mem [1082] : 
                            (N294)? \nz.mem [1090] : 
                            (N296)? \nz.mem [1098] : 
                            (N298)? \nz.mem [1106] : 
                            (N300)? \nz.mem [1114] : 
                            (N302)? \nz.mem [1122] : 
                            (N304)? \nz.mem [1130] : 
                            (N306)? \nz.mem [1138] : 
                            (N308)? \nz.mem [1146] : 
                            (N310)? \nz.mem [1154] : 
                            (N312)? \nz.mem [1162] : 
                            (N314)? \nz.mem [1170] : 
                            (N316)? \nz.mem [1178] : 
                            (N318)? \nz.mem [1186] : 
                            (N320)? \nz.mem [1194] : 
                            (N322)? \nz.mem [1202] : 
                            (N324)? \nz.mem [1210] : 
                            (N326)? \nz.mem [1218] : 
                            (N328)? \nz.mem [1226] : 
                            (N330)? \nz.mem [1234] : 
                            (N332)? \nz.mem [1242] : 
                            (N334)? \nz.mem [1250] : 
                            (N336)? \nz.mem [1258] : 
                            (N338)? \nz.mem [1266] : 
                            (N340)? \nz.mem [1274] : 
                            (N342)? \nz.mem [1282] : 
                            (N344)? \nz.mem [1290] : 
                            (N346)? \nz.mem [1298] : 
                            (N348)? \nz.mem [1306] : 
                            (N350)? \nz.mem [1314] : 
                            (N352)? \nz.mem [1322] : 
                            (N354)? \nz.mem [1330] : 
                            (N356)? \nz.mem [1338] : 
                            (N358)? \nz.mem [1346] : 
                            (N360)? \nz.mem [1354] : 
                            (N362)? \nz.mem [1362] : 
                            (N364)? \nz.mem [1370] : 
                            (N366)? \nz.mem [1378] : 
                            (N368)? \nz.mem [1386] : 
                            (N370)? \nz.mem [1394] : 
                            (N372)? \nz.mem [1402] : 
                            (N374)? \nz.mem [1410] : 
                            (N376)? \nz.mem [1418] : 
                            (N378)? \nz.mem [1426] : 
                            (N380)? \nz.mem [1434] : 
                            (N382)? \nz.mem [1442] : 
                            (N384)? \nz.mem [1450] : 
                            (N386)? \nz.mem [1458] : 
                            (N388)? \nz.mem [1466] : 
                            (N390)? \nz.mem [1474] : 
                            (N392)? \nz.mem [1482] : 
                            (N394)? \nz.mem [1490] : 
                            (N396)? \nz.mem [1498] : 
                            (N398)? \nz.mem [1506] : 
                            (N400)? \nz.mem [1514] : 
                            (N402)? \nz.mem [1522] : 
                            (N404)? \nz.mem [1530] : 
                            (N406)? \nz.mem [1538] : 
                            (N408)? \nz.mem [1546] : 
                            (N410)? \nz.mem [1554] : 
                            (N412)? \nz.mem [1562] : 
                            (N414)? \nz.mem [1570] : 
                            (N416)? \nz.mem [1578] : 
                            (N418)? \nz.mem [1586] : 
                            (N420)? \nz.mem [1594] : 
                            (N422)? \nz.mem [1602] : 
                            (N424)? \nz.mem [1610] : 
                            (N426)? \nz.mem [1618] : 
                            (N428)? \nz.mem [1626] : 
                            (N430)? \nz.mem [1634] : 
                            (N432)? \nz.mem [1642] : 
                            (N434)? \nz.mem [1650] : 
                            (N436)? \nz.mem [1658] : 
                            (N438)? \nz.mem [1666] : 
                            (N440)? \nz.mem [1674] : 
                            (N442)? \nz.mem [1682] : 
                            (N444)? \nz.mem [1690] : 
                            (N446)? \nz.mem [1698] : 
                            (N448)? \nz.mem [1706] : 
                            (N450)? \nz.mem [1714] : 
                            (N452)? \nz.mem [1722] : 
                            (N454)? \nz.mem [1730] : 
                            (N456)? \nz.mem [1738] : 
                            (N458)? \nz.mem [1746] : 
                            (N460)? \nz.mem [1754] : 
                            (N462)? \nz.mem [1762] : 
                            (N464)? \nz.mem [1770] : 
                            (N466)? \nz.mem [1778] : 
                            (N468)? \nz.mem [1786] : 
                            (N470)? \nz.mem [1794] : 
                            (N472)? \nz.mem [1802] : 
                            (N474)? \nz.mem [1810] : 
                            (N476)? \nz.mem [1818] : 
                            (N478)? \nz.mem [1826] : 
                            (N480)? \nz.mem [1834] : 
                            (N482)? \nz.mem [1842] : 
                            (N484)? \nz.mem [1850] : 
                            (N486)? \nz.mem [1858] : 
                            (N488)? \nz.mem [1866] : 
                            (N490)? \nz.mem [1874] : 
                            (N492)? \nz.mem [1882] : 
                            (N494)? \nz.mem [1890] : 
                            (N496)? \nz.mem [1898] : 
                            (N498)? \nz.mem [1906] : 
                            (N500)? \nz.mem [1914] : 
                            (N502)? \nz.mem [1922] : 
                            (N504)? \nz.mem [1930] : 
                            (N506)? \nz.mem [1938] : 
                            (N508)? \nz.mem [1946] : 
                            (N510)? \nz.mem [1954] : 
                            (N512)? \nz.mem [1962] : 
                            (N514)? \nz.mem [1970] : 
                            (N516)? \nz.mem [1978] : 
                            (N518)? \nz.mem [1986] : 
                            (N520)? \nz.mem [1994] : 
                            (N522)? \nz.mem [2002] : 
                            (N524)? \nz.mem [2010] : 
                            (N526)? \nz.mem [2018] : 
                            (N528)? \nz.mem [2026] : 
                            (N530)? \nz.mem [2034] : 
                            (N532)? \nz.mem [2042] : 1'b0;
  assign \nz.data_out [1] = (N277)? \nz.mem [1] : 
                            (N279)? \nz.mem [9] : 
                            (N281)? \nz.mem [17] : 
                            (N283)? \nz.mem [25] : 
                            (N285)? \nz.mem [33] : 
                            (N287)? \nz.mem [41] : 
                            (N289)? \nz.mem [49] : 
                            (N291)? \nz.mem [57] : 
                            (N293)? \nz.mem [65] : 
                            (N295)? \nz.mem [73] : 
                            (N297)? \nz.mem [81] : 
                            (N299)? \nz.mem [89] : 
                            (N301)? \nz.mem [97] : 
                            (N303)? \nz.mem [105] : 
                            (N305)? \nz.mem [113] : 
                            (N307)? \nz.mem [121] : 
                            (N309)? \nz.mem [129] : 
                            (N311)? \nz.mem [137] : 
                            (N313)? \nz.mem [145] : 
                            (N315)? \nz.mem [153] : 
                            (N317)? \nz.mem [161] : 
                            (N319)? \nz.mem [169] : 
                            (N321)? \nz.mem [177] : 
                            (N323)? \nz.mem [185] : 
                            (N325)? \nz.mem [193] : 
                            (N327)? \nz.mem [201] : 
                            (N329)? \nz.mem [209] : 
                            (N331)? \nz.mem [217] : 
                            (N333)? \nz.mem [225] : 
                            (N335)? \nz.mem [233] : 
                            (N337)? \nz.mem [241] : 
                            (N339)? \nz.mem [249] : 
                            (N341)? \nz.mem [257] : 
                            (N343)? \nz.mem [265] : 
                            (N345)? \nz.mem [273] : 
                            (N347)? \nz.mem [281] : 
                            (N349)? \nz.mem [289] : 
                            (N351)? \nz.mem [297] : 
                            (N353)? \nz.mem [305] : 
                            (N355)? \nz.mem [313] : 
                            (N357)? \nz.mem [321] : 
                            (N359)? \nz.mem [329] : 
                            (N361)? \nz.mem [337] : 
                            (N363)? \nz.mem [345] : 
                            (N365)? \nz.mem [353] : 
                            (N367)? \nz.mem [361] : 
                            (N369)? \nz.mem [369] : 
                            (N371)? \nz.mem [377] : 
                            (N373)? \nz.mem [385] : 
                            (N375)? \nz.mem [393] : 
                            (N377)? \nz.mem [401] : 
                            (N379)? \nz.mem [409] : 
                            (N381)? \nz.mem [417] : 
                            (N383)? \nz.mem [425] : 
                            (N385)? \nz.mem [433] : 
                            (N387)? \nz.mem [441] : 
                            (N389)? \nz.mem [449] : 
                            (N391)? \nz.mem [457] : 
                            (N393)? \nz.mem [465] : 
                            (N395)? \nz.mem [473] : 
                            (N397)? \nz.mem [481] : 
                            (N399)? \nz.mem [489] : 
                            (N401)? \nz.mem [497] : 
                            (N403)? \nz.mem [505] : 
                            (N405)? \nz.mem [513] : 
                            (N407)? \nz.mem [521] : 
                            (N409)? \nz.mem [529] : 
                            (N411)? \nz.mem [537] : 
                            (N413)? \nz.mem [545] : 
                            (N415)? \nz.mem [553] : 
                            (N417)? \nz.mem [561] : 
                            (N419)? \nz.mem [569] : 
                            (N421)? \nz.mem [577] : 
                            (N423)? \nz.mem [585] : 
                            (N425)? \nz.mem [593] : 
                            (N427)? \nz.mem [601] : 
                            (N429)? \nz.mem [609] : 
                            (N431)? \nz.mem [617] : 
                            (N433)? \nz.mem [625] : 
                            (N435)? \nz.mem [633] : 
                            (N437)? \nz.mem [641] : 
                            (N439)? \nz.mem [649] : 
                            (N441)? \nz.mem [657] : 
                            (N443)? \nz.mem [665] : 
                            (N445)? \nz.mem [673] : 
                            (N447)? \nz.mem [681] : 
                            (N449)? \nz.mem [689] : 
                            (N451)? \nz.mem [697] : 
                            (N453)? \nz.mem [705] : 
                            (N455)? \nz.mem [713] : 
                            (N457)? \nz.mem [721] : 
                            (N459)? \nz.mem [729] : 
                            (N461)? \nz.mem [737] : 
                            (N463)? \nz.mem [745] : 
                            (N465)? \nz.mem [753] : 
                            (N467)? \nz.mem [761] : 
                            (N469)? \nz.mem [769] : 
                            (N471)? \nz.mem [777] : 
                            (N473)? \nz.mem [785] : 
                            (N475)? \nz.mem [793] : 
                            (N477)? \nz.mem [801] : 
                            (N479)? \nz.mem [809] : 
                            (N481)? \nz.mem [817] : 
                            (N483)? \nz.mem [825] : 
                            (N485)? \nz.mem [833] : 
                            (N487)? \nz.mem [841] : 
                            (N489)? \nz.mem [849] : 
                            (N491)? \nz.mem [857] : 
                            (N493)? \nz.mem [865] : 
                            (N495)? \nz.mem [873] : 
                            (N497)? \nz.mem [881] : 
                            (N499)? \nz.mem [889] : 
                            (N501)? \nz.mem [897] : 
                            (N503)? \nz.mem [905] : 
                            (N505)? \nz.mem [913] : 
                            (N507)? \nz.mem [921] : 
                            (N509)? \nz.mem [929] : 
                            (N511)? \nz.mem [937] : 
                            (N513)? \nz.mem [945] : 
                            (N515)? \nz.mem [953] : 
                            (N517)? \nz.mem [961] : 
                            (N519)? \nz.mem [969] : 
                            (N521)? \nz.mem [977] : 
                            (N523)? \nz.mem [985] : 
                            (N525)? \nz.mem [993] : 
                            (N527)? \nz.mem [1001] : 
                            (N529)? \nz.mem [1009] : 
                            (N531)? \nz.mem [1017] : 
                            (N278)? \nz.mem [1025] : 
                            (N280)? \nz.mem [1033] : 
                            (N282)? \nz.mem [1041] : 
                            (N284)? \nz.mem [1049] : 
                            (N286)? \nz.mem [1057] : 
                            (N288)? \nz.mem [1065] : 
                            (N290)? \nz.mem [1073] : 
                            (N292)? \nz.mem [1081] : 
                            (N294)? \nz.mem [1089] : 
                            (N296)? \nz.mem [1097] : 
                            (N298)? \nz.mem [1105] : 
                            (N300)? \nz.mem [1113] : 
                            (N302)? \nz.mem [1121] : 
                            (N304)? \nz.mem [1129] : 
                            (N306)? \nz.mem [1137] : 
                            (N308)? \nz.mem [1145] : 
                            (N310)? \nz.mem [1153] : 
                            (N312)? \nz.mem [1161] : 
                            (N314)? \nz.mem [1169] : 
                            (N316)? \nz.mem [1177] : 
                            (N318)? \nz.mem [1185] : 
                            (N320)? \nz.mem [1193] : 
                            (N322)? \nz.mem [1201] : 
                            (N324)? \nz.mem [1209] : 
                            (N326)? \nz.mem [1217] : 
                            (N328)? \nz.mem [1225] : 
                            (N330)? \nz.mem [1233] : 
                            (N332)? \nz.mem [1241] : 
                            (N334)? \nz.mem [1249] : 
                            (N336)? \nz.mem [1257] : 
                            (N338)? \nz.mem [1265] : 
                            (N340)? \nz.mem [1273] : 
                            (N342)? \nz.mem [1281] : 
                            (N344)? \nz.mem [1289] : 
                            (N346)? \nz.mem [1297] : 
                            (N348)? \nz.mem [1305] : 
                            (N350)? \nz.mem [1313] : 
                            (N352)? \nz.mem [1321] : 
                            (N354)? \nz.mem [1329] : 
                            (N356)? \nz.mem [1337] : 
                            (N358)? \nz.mem [1345] : 
                            (N360)? \nz.mem [1353] : 
                            (N362)? \nz.mem [1361] : 
                            (N364)? \nz.mem [1369] : 
                            (N366)? \nz.mem [1377] : 
                            (N368)? \nz.mem [1385] : 
                            (N370)? \nz.mem [1393] : 
                            (N372)? \nz.mem [1401] : 
                            (N374)? \nz.mem [1409] : 
                            (N376)? \nz.mem [1417] : 
                            (N378)? \nz.mem [1425] : 
                            (N380)? \nz.mem [1433] : 
                            (N382)? \nz.mem [1441] : 
                            (N384)? \nz.mem [1449] : 
                            (N386)? \nz.mem [1457] : 
                            (N388)? \nz.mem [1465] : 
                            (N390)? \nz.mem [1473] : 
                            (N392)? \nz.mem [1481] : 
                            (N394)? \nz.mem [1489] : 
                            (N396)? \nz.mem [1497] : 
                            (N398)? \nz.mem [1505] : 
                            (N400)? \nz.mem [1513] : 
                            (N402)? \nz.mem [1521] : 
                            (N404)? \nz.mem [1529] : 
                            (N406)? \nz.mem [1537] : 
                            (N408)? \nz.mem [1545] : 
                            (N410)? \nz.mem [1553] : 
                            (N412)? \nz.mem [1561] : 
                            (N414)? \nz.mem [1569] : 
                            (N416)? \nz.mem [1577] : 
                            (N418)? \nz.mem [1585] : 
                            (N420)? \nz.mem [1593] : 
                            (N422)? \nz.mem [1601] : 
                            (N424)? \nz.mem [1609] : 
                            (N426)? \nz.mem [1617] : 
                            (N428)? \nz.mem [1625] : 
                            (N430)? \nz.mem [1633] : 
                            (N432)? \nz.mem [1641] : 
                            (N434)? \nz.mem [1649] : 
                            (N436)? \nz.mem [1657] : 
                            (N438)? \nz.mem [1665] : 
                            (N440)? \nz.mem [1673] : 
                            (N442)? \nz.mem [1681] : 
                            (N444)? \nz.mem [1689] : 
                            (N446)? \nz.mem [1697] : 
                            (N448)? \nz.mem [1705] : 
                            (N450)? \nz.mem [1713] : 
                            (N452)? \nz.mem [1721] : 
                            (N454)? \nz.mem [1729] : 
                            (N456)? \nz.mem [1737] : 
                            (N458)? \nz.mem [1745] : 
                            (N460)? \nz.mem [1753] : 
                            (N462)? \nz.mem [1761] : 
                            (N464)? \nz.mem [1769] : 
                            (N466)? \nz.mem [1777] : 
                            (N468)? \nz.mem [1785] : 
                            (N470)? \nz.mem [1793] : 
                            (N472)? \nz.mem [1801] : 
                            (N474)? \nz.mem [1809] : 
                            (N476)? \nz.mem [1817] : 
                            (N478)? \nz.mem [1825] : 
                            (N480)? \nz.mem [1833] : 
                            (N482)? \nz.mem [1841] : 
                            (N484)? \nz.mem [1849] : 
                            (N486)? \nz.mem [1857] : 
                            (N488)? \nz.mem [1865] : 
                            (N490)? \nz.mem [1873] : 
                            (N492)? \nz.mem [1881] : 
                            (N494)? \nz.mem [1889] : 
                            (N496)? \nz.mem [1897] : 
                            (N498)? \nz.mem [1905] : 
                            (N500)? \nz.mem [1913] : 
                            (N502)? \nz.mem [1921] : 
                            (N504)? \nz.mem [1929] : 
                            (N506)? \nz.mem [1937] : 
                            (N508)? \nz.mem [1945] : 
                            (N510)? \nz.mem [1953] : 
                            (N512)? \nz.mem [1961] : 
                            (N514)? \nz.mem [1969] : 
                            (N516)? \nz.mem [1977] : 
                            (N518)? \nz.mem [1985] : 
                            (N520)? \nz.mem [1993] : 
                            (N522)? \nz.mem [2001] : 
                            (N524)? \nz.mem [2009] : 
                            (N526)? \nz.mem [2017] : 
                            (N528)? \nz.mem [2025] : 
                            (N530)? \nz.mem [2033] : 
                            (N532)? \nz.mem [2041] : 1'b0;
  assign \nz.data_out [0] = (N277)? \nz.mem [0] : 
                            (N279)? \nz.mem [8] : 
                            (N281)? \nz.mem [16] : 
                            (N283)? \nz.mem [24] : 
                            (N285)? \nz.mem [32] : 
                            (N287)? \nz.mem [40] : 
                            (N289)? \nz.mem [48] : 
                            (N291)? \nz.mem [56] : 
                            (N293)? \nz.mem [64] : 
                            (N295)? \nz.mem [72] : 
                            (N297)? \nz.mem [80] : 
                            (N299)? \nz.mem [88] : 
                            (N301)? \nz.mem [96] : 
                            (N303)? \nz.mem [104] : 
                            (N305)? \nz.mem [112] : 
                            (N307)? \nz.mem [120] : 
                            (N309)? \nz.mem [128] : 
                            (N311)? \nz.mem [136] : 
                            (N313)? \nz.mem [144] : 
                            (N315)? \nz.mem [152] : 
                            (N317)? \nz.mem [160] : 
                            (N319)? \nz.mem [168] : 
                            (N321)? \nz.mem [176] : 
                            (N323)? \nz.mem [184] : 
                            (N325)? \nz.mem [192] : 
                            (N327)? \nz.mem [200] : 
                            (N329)? \nz.mem [208] : 
                            (N331)? \nz.mem [216] : 
                            (N333)? \nz.mem [224] : 
                            (N335)? \nz.mem [232] : 
                            (N337)? \nz.mem [240] : 
                            (N339)? \nz.mem [248] : 
                            (N341)? \nz.mem [256] : 
                            (N343)? \nz.mem [264] : 
                            (N345)? \nz.mem [272] : 
                            (N347)? \nz.mem [280] : 
                            (N349)? \nz.mem [288] : 
                            (N351)? \nz.mem [296] : 
                            (N353)? \nz.mem [304] : 
                            (N355)? \nz.mem [312] : 
                            (N357)? \nz.mem [320] : 
                            (N359)? \nz.mem [328] : 
                            (N361)? \nz.mem [336] : 
                            (N363)? \nz.mem [344] : 
                            (N365)? \nz.mem [352] : 
                            (N367)? \nz.mem [360] : 
                            (N369)? \nz.mem [368] : 
                            (N371)? \nz.mem [376] : 
                            (N373)? \nz.mem [384] : 
                            (N375)? \nz.mem [392] : 
                            (N377)? \nz.mem [400] : 
                            (N379)? \nz.mem [408] : 
                            (N381)? \nz.mem [416] : 
                            (N383)? \nz.mem [424] : 
                            (N385)? \nz.mem [432] : 
                            (N387)? \nz.mem [440] : 
                            (N389)? \nz.mem [448] : 
                            (N391)? \nz.mem [456] : 
                            (N393)? \nz.mem [464] : 
                            (N395)? \nz.mem [472] : 
                            (N397)? \nz.mem [480] : 
                            (N399)? \nz.mem [488] : 
                            (N401)? \nz.mem [496] : 
                            (N403)? \nz.mem [504] : 
                            (N405)? \nz.mem [512] : 
                            (N407)? \nz.mem [520] : 
                            (N409)? \nz.mem [528] : 
                            (N411)? \nz.mem [536] : 
                            (N413)? \nz.mem [544] : 
                            (N415)? \nz.mem [552] : 
                            (N417)? \nz.mem [560] : 
                            (N419)? \nz.mem [568] : 
                            (N421)? \nz.mem [576] : 
                            (N423)? \nz.mem [584] : 
                            (N425)? \nz.mem [592] : 
                            (N427)? \nz.mem [600] : 
                            (N429)? \nz.mem [608] : 
                            (N431)? \nz.mem [616] : 
                            (N433)? \nz.mem [624] : 
                            (N435)? \nz.mem [632] : 
                            (N437)? \nz.mem [640] : 
                            (N439)? \nz.mem [648] : 
                            (N441)? \nz.mem [656] : 
                            (N443)? \nz.mem [664] : 
                            (N445)? \nz.mem [672] : 
                            (N447)? \nz.mem [680] : 
                            (N449)? \nz.mem [688] : 
                            (N451)? \nz.mem [696] : 
                            (N453)? \nz.mem [704] : 
                            (N455)? \nz.mem [712] : 
                            (N457)? \nz.mem [720] : 
                            (N459)? \nz.mem [728] : 
                            (N461)? \nz.mem [736] : 
                            (N463)? \nz.mem [744] : 
                            (N465)? \nz.mem [752] : 
                            (N467)? \nz.mem [760] : 
                            (N469)? \nz.mem [768] : 
                            (N471)? \nz.mem [776] : 
                            (N473)? \nz.mem [784] : 
                            (N475)? \nz.mem [792] : 
                            (N477)? \nz.mem [800] : 
                            (N479)? \nz.mem [808] : 
                            (N481)? \nz.mem [816] : 
                            (N483)? \nz.mem [824] : 
                            (N485)? \nz.mem [832] : 
                            (N487)? \nz.mem [840] : 
                            (N489)? \nz.mem [848] : 
                            (N491)? \nz.mem [856] : 
                            (N493)? \nz.mem [864] : 
                            (N495)? \nz.mem [872] : 
                            (N497)? \nz.mem [880] : 
                            (N499)? \nz.mem [888] : 
                            (N501)? \nz.mem [896] : 
                            (N503)? \nz.mem [904] : 
                            (N505)? \nz.mem [912] : 
                            (N507)? \nz.mem [920] : 
                            (N509)? \nz.mem [928] : 
                            (N511)? \nz.mem [936] : 
                            (N513)? \nz.mem [944] : 
                            (N515)? \nz.mem [952] : 
                            (N517)? \nz.mem [960] : 
                            (N519)? \nz.mem [968] : 
                            (N521)? \nz.mem [976] : 
                            (N523)? \nz.mem [984] : 
                            (N525)? \nz.mem [992] : 
                            (N527)? \nz.mem [1000] : 
                            (N529)? \nz.mem [1008] : 
                            (N531)? \nz.mem [1016] : 
                            (N278)? \nz.mem [1024] : 
                            (N280)? \nz.mem [1032] : 
                            (N282)? \nz.mem [1040] : 
                            (N284)? \nz.mem [1048] : 
                            (N286)? \nz.mem [1056] : 
                            (N288)? \nz.mem [1064] : 
                            (N290)? \nz.mem [1072] : 
                            (N292)? \nz.mem [1080] : 
                            (N294)? \nz.mem [1088] : 
                            (N296)? \nz.mem [1096] : 
                            (N298)? \nz.mem [1104] : 
                            (N300)? \nz.mem [1112] : 
                            (N302)? \nz.mem [1120] : 
                            (N304)? \nz.mem [1128] : 
                            (N306)? \nz.mem [1136] : 
                            (N308)? \nz.mem [1144] : 
                            (N310)? \nz.mem [1152] : 
                            (N312)? \nz.mem [1160] : 
                            (N314)? \nz.mem [1168] : 
                            (N316)? \nz.mem [1176] : 
                            (N318)? \nz.mem [1184] : 
                            (N320)? \nz.mem [1192] : 
                            (N322)? \nz.mem [1200] : 
                            (N324)? \nz.mem [1208] : 
                            (N326)? \nz.mem [1216] : 
                            (N328)? \nz.mem [1224] : 
                            (N330)? \nz.mem [1232] : 
                            (N332)? \nz.mem [1240] : 
                            (N334)? \nz.mem [1248] : 
                            (N336)? \nz.mem [1256] : 
                            (N338)? \nz.mem [1264] : 
                            (N340)? \nz.mem [1272] : 
                            (N342)? \nz.mem [1280] : 
                            (N344)? \nz.mem [1288] : 
                            (N346)? \nz.mem [1296] : 
                            (N348)? \nz.mem [1304] : 
                            (N350)? \nz.mem [1312] : 
                            (N352)? \nz.mem [1320] : 
                            (N354)? \nz.mem [1328] : 
                            (N356)? \nz.mem [1336] : 
                            (N358)? \nz.mem [1344] : 
                            (N360)? \nz.mem [1352] : 
                            (N362)? \nz.mem [1360] : 
                            (N364)? \nz.mem [1368] : 
                            (N366)? \nz.mem [1376] : 
                            (N368)? \nz.mem [1384] : 
                            (N370)? \nz.mem [1392] : 
                            (N372)? \nz.mem [1400] : 
                            (N374)? \nz.mem [1408] : 
                            (N376)? \nz.mem [1416] : 
                            (N378)? \nz.mem [1424] : 
                            (N380)? \nz.mem [1432] : 
                            (N382)? \nz.mem [1440] : 
                            (N384)? \nz.mem [1448] : 
                            (N386)? \nz.mem [1456] : 
                            (N388)? \nz.mem [1464] : 
                            (N390)? \nz.mem [1472] : 
                            (N392)? \nz.mem [1480] : 
                            (N394)? \nz.mem [1488] : 
                            (N396)? \nz.mem [1496] : 
                            (N398)? \nz.mem [1504] : 
                            (N400)? \nz.mem [1512] : 
                            (N402)? \nz.mem [1520] : 
                            (N404)? \nz.mem [1528] : 
                            (N406)? \nz.mem [1536] : 
                            (N408)? \nz.mem [1544] : 
                            (N410)? \nz.mem [1552] : 
                            (N412)? \nz.mem [1560] : 
                            (N414)? \nz.mem [1568] : 
                            (N416)? \nz.mem [1576] : 
                            (N418)? \nz.mem [1584] : 
                            (N420)? \nz.mem [1592] : 
                            (N422)? \nz.mem [1600] : 
                            (N424)? \nz.mem [1608] : 
                            (N426)? \nz.mem [1616] : 
                            (N428)? \nz.mem [1624] : 
                            (N430)? \nz.mem [1632] : 
                            (N432)? \nz.mem [1640] : 
                            (N434)? \nz.mem [1648] : 
                            (N436)? \nz.mem [1656] : 
                            (N438)? \nz.mem [1664] : 
                            (N440)? \nz.mem [1672] : 
                            (N442)? \nz.mem [1680] : 
                            (N444)? \nz.mem [1688] : 
                            (N446)? \nz.mem [1696] : 
                            (N448)? \nz.mem [1704] : 
                            (N450)? \nz.mem [1712] : 
                            (N452)? \nz.mem [1720] : 
                            (N454)? \nz.mem [1728] : 
                            (N456)? \nz.mem [1736] : 
                            (N458)? \nz.mem [1744] : 
                            (N460)? \nz.mem [1752] : 
                            (N462)? \nz.mem [1760] : 
                            (N464)? \nz.mem [1768] : 
                            (N466)? \nz.mem [1776] : 
                            (N468)? \nz.mem [1784] : 
                            (N470)? \nz.mem [1792] : 
                            (N472)? \nz.mem [1800] : 
                            (N474)? \nz.mem [1808] : 
                            (N476)? \nz.mem [1816] : 
                            (N478)? \nz.mem [1824] : 
                            (N480)? \nz.mem [1832] : 
                            (N482)? \nz.mem [1840] : 
                            (N484)? \nz.mem [1848] : 
                            (N486)? \nz.mem [1856] : 
                            (N488)? \nz.mem [1864] : 
                            (N490)? \nz.mem [1872] : 
                            (N492)? \nz.mem [1880] : 
                            (N494)? \nz.mem [1888] : 
                            (N496)? \nz.mem [1896] : 
                            (N498)? \nz.mem [1904] : 
                            (N500)? \nz.mem [1912] : 
                            (N502)? \nz.mem [1920] : 
                            (N504)? \nz.mem [1928] : 
                            (N506)? \nz.mem [1936] : 
                            (N508)? \nz.mem [1944] : 
                            (N510)? \nz.mem [1952] : 
                            (N512)? \nz.mem [1960] : 
                            (N514)? \nz.mem [1968] : 
                            (N516)? \nz.mem [1976] : 
                            (N518)? \nz.mem [1984] : 
                            (N520)? \nz.mem [1992] : 
                            (N522)? \nz.mem [2000] : 
                            (N524)? \nz.mem [2008] : 
                            (N526)? \nz.mem [2016] : 
                            (N528)? \nz.mem [2024] : 
                            (N530)? \nz.mem [2032] : 
                            (N532)? \nz.mem [2040] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p8
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N1047 = addr_i[6] & addr_i[7];
  assign N1048 = N0 & addr_i[7];
  assign N0 = ~addr_i[6];
  assign N1049 = addr_i[6] & N1;
  assign N1 = ~addr_i[7];
  assign N1050 = N2 & N3;
  assign N2 = ~addr_i[6];
  assign N3 = ~addr_i[7];
  assign N1051 = addr_i[4] & addr_i[5];
  assign N1052 = N4 & addr_i[5];
  assign N4 = ~addr_i[4];
  assign N1053 = addr_i[4] & N5;
  assign N5 = ~addr_i[5];
  assign N1054 = N6 & N7;
  assign N6 = ~addr_i[4];
  assign N7 = ~addr_i[5];
  assign N1055 = N1047 & N1051;
  assign N1056 = N1047 & N1052;
  assign N1057 = N1047 & N1053;
  assign N1058 = N1047 & N1054;
  assign N1059 = N1048 & N1051;
  assign N1060 = N1048 & N1052;
  assign N1061 = N1048 & N1053;
  assign N1062 = N1048 & N1054;
  assign N1063 = N1049 & N1051;
  assign N1064 = N1049 & N1052;
  assign N1065 = N1049 & N1053;
  assign N1066 = N1049 & N1054;
  assign N1067 = N1050 & N1051;
  assign N1068 = N1050 & N1052;
  assign N1069 = N1050 & N1053;
  assign N1070 = N1050 & N1054;
  assign N1071 = addr_i[2] & addr_i[3];
  assign N1072 = N8 & addr_i[3];
  assign N8 = ~addr_i[2];
  assign N1073 = addr_i[2] & N9;
  assign N9 = ~addr_i[3];
  assign N1074 = N10 & N11;
  assign N10 = ~addr_i[2];
  assign N11 = ~addr_i[3];
  assign N1075 = addr_i[0] & addr_i[1];
  assign N1076 = N12 & addr_i[1];
  assign N12 = ~addr_i[0];
  assign N1077 = addr_i[0] & N13;
  assign N13 = ~addr_i[1];
  assign N1078 = N14 & N15;
  assign N14 = ~addr_i[0];
  assign N15 = ~addr_i[1];
  assign N1079 = N1071 & N1075;
  assign N1080 = N1071 & N1076;
  assign N1081 = N1071 & N1077;
  assign N1082 = N1071 & N1078;
  assign N1083 = N1072 & N1075;
  assign N1084 = N1072 & N1076;
  assign N1085 = N1072 & N1077;
  assign N1086 = N1072 & N1078;
  assign N1087 = N1073 & N1075;
  assign N1088 = N1073 & N1076;
  assign N1089 = N1073 & N1077;
  assign N1090 = N1073 & N1078;
  assign N1091 = N1074 & N1075;
  assign N1092 = N1074 & N1076;
  assign N1093 = N1074 & N1077;
  assign N1094 = N1074 & N1078;
  assign N790 = N1055 & N1079;
  assign N789 = N1055 & N1080;
  assign N788 = N1055 & N1081;
  assign N787 = N1055 & N1082;
  assign N786 = N1055 & N1083;
  assign N785 = N1055 & N1084;
  assign N784 = N1055 & N1085;
  assign N783 = N1055 & N1086;
  assign N782 = N1055 & N1087;
  assign N781 = N1055 & N1088;
  assign N780 = N1055 & N1089;
  assign N779 = N1055 & N1090;
  assign N778 = N1055 & N1091;
  assign N777 = N1055 & N1092;
  assign N776 = N1055 & N1093;
  assign N775 = N1055 & N1094;
  assign N774 = N1056 & N1079;
  assign N773 = N1056 & N1080;
  assign N772 = N1056 & N1081;
  assign N771 = N1056 & N1082;
  assign N770 = N1056 & N1083;
  assign N769 = N1056 & N1084;
  assign N768 = N1056 & N1085;
  assign N767 = N1056 & N1086;
  assign N766 = N1056 & N1087;
  assign N765 = N1056 & N1088;
  assign N764 = N1056 & N1089;
  assign N763 = N1056 & N1090;
  assign N762 = N1056 & N1091;
  assign N761 = N1056 & N1092;
  assign N760 = N1056 & N1093;
  assign N759 = N1056 & N1094;
  assign N758 = N1057 & N1079;
  assign N757 = N1057 & N1080;
  assign N756 = N1057 & N1081;
  assign N755 = N1057 & N1082;
  assign N754 = N1057 & N1083;
  assign N753 = N1057 & N1084;
  assign N752 = N1057 & N1085;
  assign N751 = N1057 & N1086;
  assign N750 = N1057 & N1087;
  assign N749 = N1057 & N1088;
  assign N748 = N1057 & N1089;
  assign N747 = N1057 & N1090;
  assign N746 = N1057 & N1091;
  assign N745 = N1057 & N1092;
  assign N744 = N1057 & N1093;
  assign N743 = N1057 & N1094;
  assign N742 = N1058 & N1079;
  assign N741 = N1058 & N1080;
  assign N740 = N1058 & N1081;
  assign N739 = N1058 & N1082;
  assign N738 = N1058 & N1083;
  assign N737 = N1058 & N1084;
  assign N736 = N1058 & N1085;
  assign N735 = N1058 & N1086;
  assign N734 = N1058 & N1087;
  assign N733 = N1058 & N1088;
  assign N732 = N1058 & N1089;
  assign N731 = N1058 & N1090;
  assign N730 = N1058 & N1091;
  assign N729 = N1058 & N1092;
  assign N728 = N1058 & N1093;
  assign N727 = N1058 & N1094;
  assign N726 = N1059 & N1079;
  assign N725 = N1059 & N1080;
  assign N724 = N1059 & N1081;
  assign N723 = N1059 & N1082;
  assign N722 = N1059 & N1083;
  assign N721 = N1059 & N1084;
  assign N720 = N1059 & N1085;
  assign N719 = N1059 & N1086;
  assign N718 = N1059 & N1087;
  assign N717 = N1059 & N1088;
  assign N716 = N1059 & N1089;
  assign N715 = N1059 & N1090;
  assign N714 = N1059 & N1091;
  assign N713 = N1059 & N1092;
  assign N712 = N1059 & N1093;
  assign N711 = N1059 & N1094;
  assign N710 = N1060 & N1079;
  assign N709 = N1060 & N1080;
  assign N708 = N1060 & N1081;
  assign N707 = N1060 & N1082;
  assign N706 = N1060 & N1083;
  assign N705 = N1060 & N1084;
  assign N704 = N1060 & N1085;
  assign N703 = N1060 & N1086;
  assign N702 = N1060 & N1087;
  assign N701 = N1060 & N1088;
  assign N700 = N1060 & N1089;
  assign N699 = N1060 & N1090;
  assign N698 = N1060 & N1091;
  assign N697 = N1060 & N1092;
  assign N696 = N1060 & N1093;
  assign N695 = N1060 & N1094;
  assign N694 = N1061 & N1079;
  assign N693 = N1061 & N1080;
  assign N692 = N1061 & N1081;
  assign N691 = N1061 & N1082;
  assign N690 = N1061 & N1083;
  assign N689 = N1061 & N1084;
  assign N688 = N1061 & N1085;
  assign N687 = N1061 & N1086;
  assign N686 = N1061 & N1087;
  assign N685 = N1061 & N1088;
  assign N684 = N1061 & N1089;
  assign N683 = N1061 & N1090;
  assign N682 = N1061 & N1091;
  assign N681 = N1061 & N1092;
  assign N680 = N1061 & N1093;
  assign N679 = N1061 & N1094;
  assign N678 = N1062 & N1079;
  assign N677 = N1062 & N1080;
  assign N676 = N1062 & N1081;
  assign N675 = N1062 & N1082;
  assign N674 = N1062 & N1083;
  assign N673 = N1062 & N1084;
  assign N672 = N1062 & N1085;
  assign N671 = N1062 & N1086;
  assign N670 = N1062 & N1087;
  assign N669 = N1062 & N1088;
  assign N668 = N1062 & N1089;
  assign N667 = N1062 & N1090;
  assign N666 = N1062 & N1091;
  assign N665 = N1062 & N1092;
  assign N664 = N1062 & N1093;
  assign N663 = N1062 & N1094;
  assign N662 = N1063 & N1079;
  assign N661 = N1063 & N1080;
  assign N660 = N1063 & N1081;
  assign N659 = N1063 & N1082;
  assign N658 = N1063 & N1083;
  assign N657 = N1063 & N1084;
  assign N656 = N1063 & N1085;
  assign N655 = N1063 & N1086;
  assign N654 = N1063 & N1087;
  assign N653 = N1063 & N1088;
  assign N652 = N1063 & N1089;
  assign N651 = N1063 & N1090;
  assign N650 = N1063 & N1091;
  assign N649 = N1063 & N1092;
  assign N648 = N1063 & N1093;
  assign N647 = N1063 & N1094;
  assign N646 = N1064 & N1079;
  assign N645 = N1064 & N1080;
  assign N644 = N1064 & N1081;
  assign N643 = N1064 & N1082;
  assign N642 = N1064 & N1083;
  assign N641 = N1064 & N1084;
  assign N640 = N1064 & N1085;
  assign N639 = N1064 & N1086;
  assign N638 = N1064 & N1087;
  assign N637 = N1064 & N1088;
  assign N636 = N1064 & N1089;
  assign N635 = N1064 & N1090;
  assign N634 = N1064 & N1091;
  assign N633 = N1064 & N1092;
  assign N632 = N1064 & N1093;
  assign N631 = N1064 & N1094;
  assign N630 = N1065 & N1079;
  assign N629 = N1065 & N1080;
  assign N628 = N1065 & N1081;
  assign N627 = N1065 & N1082;
  assign N626 = N1065 & N1083;
  assign N625 = N1065 & N1084;
  assign N624 = N1065 & N1085;
  assign N623 = N1065 & N1086;
  assign N622 = N1065 & N1087;
  assign N621 = N1065 & N1088;
  assign N620 = N1065 & N1089;
  assign N619 = N1065 & N1090;
  assign N618 = N1065 & N1091;
  assign N617 = N1065 & N1092;
  assign N616 = N1065 & N1093;
  assign N615 = N1065 & N1094;
  assign N614 = N1066 & N1079;
  assign N613 = N1066 & N1080;
  assign N612 = N1066 & N1081;
  assign N611 = N1066 & N1082;
  assign N610 = N1066 & N1083;
  assign N609 = N1066 & N1084;
  assign N608 = N1066 & N1085;
  assign N607 = N1066 & N1086;
  assign N606 = N1066 & N1087;
  assign N605 = N1066 & N1088;
  assign N604 = N1066 & N1089;
  assign N603 = N1066 & N1090;
  assign N602 = N1066 & N1091;
  assign N601 = N1066 & N1092;
  assign N600 = N1066 & N1093;
  assign N599 = N1066 & N1094;
  assign N598 = N1067 & N1079;
  assign N597 = N1067 & N1080;
  assign N596 = N1067 & N1081;
  assign N595 = N1067 & N1082;
  assign N594 = N1067 & N1083;
  assign N593 = N1067 & N1084;
  assign N592 = N1067 & N1085;
  assign N591 = N1067 & N1086;
  assign N590 = N1067 & N1087;
  assign N589 = N1067 & N1088;
  assign N588 = N1067 & N1089;
  assign N587 = N1067 & N1090;
  assign N586 = N1067 & N1091;
  assign N585 = N1067 & N1092;
  assign N584 = N1067 & N1093;
  assign N583 = N1067 & N1094;
  assign N582 = N1068 & N1079;
  assign N581 = N1068 & N1080;
  assign N580 = N1068 & N1081;
  assign N579 = N1068 & N1082;
  assign N578 = N1068 & N1083;
  assign N577 = N1068 & N1084;
  assign N576 = N1068 & N1085;
  assign N575 = N1068 & N1086;
  assign N574 = N1068 & N1087;
  assign N573 = N1068 & N1088;
  assign N572 = N1068 & N1089;
  assign N571 = N1068 & N1090;
  assign N570 = N1068 & N1091;
  assign N569 = N1068 & N1092;
  assign N568 = N1068 & N1093;
  assign N567 = N1068 & N1094;
  assign N566 = N1069 & N1079;
  assign N565 = N1069 & N1080;
  assign N564 = N1069 & N1081;
  assign N563 = N1069 & N1082;
  assign N562 = N1069 & N1083;
  assign N561 = N1069 & N1084;
  assign N560 = N1069 & N1085;
  assign N559 = N1069 & N1086;
  assign N558 = N1069 & N1087;
  assign N557 = N1069 & N1088;
  assign N556 = N1069 & N1089;
  assign N555 = N1069 & N1090;
  assign N554 = N1069 & N1091;
  assign N553 = N1069 & N1092;
  assign N552 = N1069 & N1093;
  assign N551 = N1069 & N1094;
  assign N550 = N1070 & N1079;
  assign N549 = N1070 & N1080;
  assign N548 = N1070 & N1081;
  assign N547 = N1070 & N1082;
  assign N546 = N1070 & N1083;
  assign N545 = N1070 & N1084;
  assign N544 = N1070 & N1085;
  assign N543 = N1070 & N1086;
  assign N542 = N1070 & N1087;
  assign N541 = N1070 & N1088;
  assign N540 = N1070 & N1089;
  assign N539 = N1070 & N1090;
  assign N538 = N1070 & N1091;
  assign N537 = N1070 & N1092;
  assign N536 = N1070 & N1093;
  assign N535 = N1070 & N1094;
  assign { N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791 } = (N16)? { N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N533;
  assign \nz.read_en  = v_i & N1095;
  assign N1095 = ~w_i;
  assign N17 = ~\nz.addr_r [0];
  assign N18 = ~\nz.addr_r [1];
  assign N19 = N17 & N18;
  assign N20 = N17 & \nz.addr_r [1];
  assign N21 = \nz.addr_r [0] & N18;
  assign N22 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N23 = ~\nz.addr_r [2];
  assign N24 = N19 & N23;
  assign N25 = N19 & \nz.addr_r [2];
  assign N26 = N21 & N23;
  assign N27 = N21 & \nz.addr_r [2];
  assign N28 = N20 & N23;
  assign N29 = N20 & \nz.addr_r [2];
  assign N30 = N22 & N23;
  assign N31 = N22 & \nz.addr_r [2];
  assign N32 = ~\nz.addr_r [3];
  assign N33 = N24 & N32;
  assign N34 = N24 & \nz.addr_r [3];
  assign N35 = N26 & N32;
  assign N36 = N26 & \nz.addr_r [3];
  assign N37 = N28 & N32;
  assign N38 = N28 & \nz.addr_r [3];
  assign N39 = N30 & N32;
  assign N40 = N30 & \nz.addr_r [3];
  assign N41 = N25 & N32;
  assign N42 = N25 & \nz.addr_r [3];
  assign N43 = N27 & N32;
  assign N44 = N27 & \nz.addr_r [3];
  assign N45 = N29 & N32;
  assign N46 = N29 & \nz.addr_r [3];
  assign N47 = N31 & N32;
  assign N48 = N31 & \nz.addr_r [3];
  assign N49 = ~\nz.addr_r [4];
  assign N50 = N33 & N49;
  assign N51 = N33 & \nz.addr_r [4];
  assign N52 = N35 & N49;
  assign N53 = N35 & \nz.addr_r [4];
  assign N54 = N37 & N49;
  assign N55 = N37 & \nz.addr_r [4];
  assign N56 = N39 & N49;
  assign N57 = N39 & \nz.addr_r [4];
  assign N58 = N41 & N49;
  assign N59 = N41 & \nz.addr_r [4];
  assign N60 = N43 & N49;
  assign N61 = N43 & \nz.addr_r [4];
  assign N62 = N45 & N49;
  assign N63 = N45 & \nz.addr_r [4];
  assign N64 = N47 & N49;
  assign N65 = N47 & \nz.addr_r [4];
  assign N66 = N34 & N49;
  assign N67 = N34 & \nz.addr_r [4];
  assign N68 = N36 & N49;
  assign N69 = N36 & \nz.addr_r [4];
  assign N70 = N38 & N49;
  assign N71 = N38 & \nz.addr_r [4];
  assign N72 = N40 & N49;
  assign N73 = N40 & \nz.addr_r [4];
  assign N74 = N42 & N49;
  assign N75 = N42 & \nz.addr_r [4];
  assign N76 = N44 & N49;
  assign N77 = N44 & \nz.addr_r [4];
  assign N78 = N46 & N49;
  assign N79 = N46 & \nz.addr_r [4];
  assign N80 = N48 & N49;
  assign N81 = N48 & \nz.addr_r [4];
  assign N82 = ~\nz.addr_r [5];
  assign N83 = N50 & N82;
  assign N84 = N50 & \nz.addr_r [5];
  assign N85 = N52 & N82;
  assign N86 = N52 & \nz.addr_r [5];
  assign N87 = N54 & N82;
  assign N88 = N54 & \nz.addr_r [5];
  assign N89 = N56 & N82;
  assign N90 = N56 & \nz.addr_r [5];
  assign N91 = N58 & N82;
  assign N92 = N58 & \nz.addr_r [5];
  assign N93 = N60 & N82;
  assign N94 = N60 & \nz.addr_r [5];
  assign N95 = N62 & N82;
  assign N96 = N62 & \nz.addr_r [5];
  assign N97 = N64 & N82;
  assign N98 = N64 & \nz.addr_r [5];
  assign N99 = N66 & N82;
  assign N100 = N66 & \nz.addr_r [5];
  assign N101 = N68 & N82;
  assign N102 = N68 & \nz.addr_r [5];
  assign N103 = N70 & N82;
  assign N104 = N70 & \nz.addr_r [5];
  assign N105 = N72 & N82;
  assign N106 = N72 & \nz.addr_r [5];
  assign N107 = N74 & N82;
  assign N108 = N74 & \nz.addr_r [5];
  assign N109 = N76 & N82;
  assign N110 = N76 & \nz.addr_r [5];
  assign N111 = N78 & N82;
  assign N112 = N78 & \nz.addr_r [5];
  assign N113 = N80 & N82;
  assign N114 = N80 & \nz.addr_r [5];
  assign N115 = N51 & N82;
  assign N116 = N51 & \nz.addr_r [5];
  assign N117 = N53 & N82;
  assign N118 = N53 & \nz.addr_r [5];
  assign N119 = N55 & N82;
  assign N120 = N55 & \nz.addr_r [5];
  assign N121 = N57 & N82;
  assign N122 = N57 & \nz.addr_r [5];
  assign N123 = N59 & N82;
  assign N124 = N59 & \nz.addr_r [5];
  assign N125 = N61 & N82;
  assign N126 = N61 & \nz.addr_r [5];
  assign N127 = N63 & N82;
  assign N128 = N63 & \nz.addr_r [5];
  assign N129 = N65 & N82;
  assign N130 = N65 & \nz.addr_r [5];
  assign N131 = N67 & N82;
  assign N132 = N67 & \nz.addr_r [5];
  assign N133 = N69 & N82;
  assign N134 = N69 & \nz.addr_r [5];
  assign N135 = N71 & N82;
  assign N136 = N71 & \nz.addr_r [5];
  assign N137 = N73 & N82;
  assign N138 = N73 & \nz.addr_r [5];
  assign N139 = N75 & N82;
  assign N140 = N75 & \nz.addr_r [5];
  assign N141 = N77 & N82;
  assign N142 = N77 & \nz.addr_r [5];
  assign N143 = N79 & N82;
  assign N144 = N79 & \nz.addr_r [5];
  assign N145 = N81 & N82;
  assign N146 = N81 & \nz.addr_r [5];
  assign N147 = ~\nz.addr_r [6];
  assign N148 = N83 & N147;
  assign N149 = N83 & \nz.addr_r [6];
  assign N150 = N85 & N147;
  assign N151 = N85 & \nz.addr_r [6];
  assign N152 = N87 & N147;
  assign N153 = N87 & \nz.addr_r [6];
  assign N154 = N89 & N147;
  assign N155 = N89 & \nz.addr_r [6];
  assign N156 = N91 & N147;
  assign N157 = N91 & \nz.addr_r [6];
  assign N158 = N93 & N147;
  assign N159 = N93 & \nz.addr_r [6];
  assign N160 = N95 & N147;
  assign N161 = N95 & \nz.addr_r [6];
  assign N162 = N97 & N147;
  assign N163 = N97 & \nz.addr_r [6];
  assign N164 = N99 & N147;
  assign N165 = N99 & \nz.addr_r [6];
  assign N166 = N101 & N147;
  assign N167 = N101 & \nz.addr_r [6];
  assign N168 = N103 & N147;
  assign N169 = N103 & \nz.addr_r [6];
  assign N170 = N105 & N147;
  assign N171 = N105 & \nz.addr_r [6];
  assign N172 = N107 & N147;
  assign N173 = N107 & \nz.addr_r [6];
  assign N174 = N109 & N147;
  assign N175 = N109 & \nz.addr_r [6];
  assign N176 = N111 & N147;
  assign N177 = N111 & \nz.addr_r [6];
  assign N178 = N113 & N147;
  assign N179 = N113 & \nz.addr_r [6];
  assign N180 = N115 & N147;
  assign N181 = N115 & \nz.addr_r [6];
  assign N182 = N117 & N147;
  assign N183 = N117 & \nz.addr_r [6];
  assign N184 = N119 & N147;
  assign N185 = N119 & \nz.addr_r [6];
  assign N186 = N121 & N147;
  assign N187 = N121 & \nz.addr_r [6];
  assign N188 = N123 & N147;
  assign N189 = N123 & \nz.addr_r [6];
  assign N190 = N125 & N147;
  assign N191 = N125 & \nz.addr_r [6];
  assign N192 = N127 & N147;
  assign N193 = N127 & \nz.addr_r [6];
  assign N194 = N129 & N147;
  assign N195 = N129 & \nz.addr_r [6];
  assign N196 = N131 & N147;
  assign N197 = N131 & \nz.addr_r [6];
  assign N198 = N133 & N147;
  assign N199 = N133 & \nz.addr_r [6];
  assign N200 = N135 & N147;
  assign N201 = N135 & \nz.addr_r [6];
  assign N202 = N137 & N147;
  assign N203 = N137 & \nz.addr_r [6];
  assign N204 = N139 & N147;
  assign N205 = N139 & \nz.addr_r [6];
  assign N206 = N141 & N147;
  assign N207 = N141 & \nz.addr_r [6];
  assign N208 = N143 & N147;
  assign N209 = N143 & \nz.addr_r [6];
  assign N210 = N145 & N147;
  assign N211 = N145 & \nz.addr_r [6];
  assign N212 = N84 & N147;
  assign N213 = N84 & \nz.addr_r [6];
  assign N214 = N86 & N147;
  assign N215 = N86 & \nz.addr_r [6];
  assign N216 = N88 & N147;
  assign N217 = N88 & \nz.addr_r [6];
  assign N218 = N90 & N147;
  assign N219 = N90 & \nz.addr_r [6];
  assign N220 = N92 & N147;
  assign N221 = N92 & \nz.addr_r [6];
  assign N222 = N94 & N147;
  assign N223 = N94 & \nz.addr_r [6];
  assign N224 = N96 & N147;
  assign N225 = N96 & \nz.addr_r [6];
  assign N226 = N98 & N147;
  assign N227 = N98 & \nz.addr_r [6];
  assign N228 = N100 & N147;
  assign N229 = N100 & \nz.addr_r [6];
  assign N230 = N102 & N147;
  assign N231 = N102 & \nz.addr_r [6];
  assign N232 = N104 & N147;
  assign N233 = N104 & \nz.addr_r [6];
  assign N234 = N106 & N147;
  assign N235 = N106 & \nz.addr_r [6];
  assign N236 = N108 & N147;
  assign N237 = N108 & \nz.addr_r [6];
  assign N238 = N110 & N147;
  assign N239 = N110 & \nz.addr_r [6];
  assign N240 = N112 & N147;
  assign N241 = N112 & \nz.addr_r [6];
  assign N242 = N114 & N147;
  assign N243 = N114 & \nz.addr_r [6];
  assign N244 = N116 & N147;
  assign N245 = N116 & \nz.addr_r [6];
  assign N246 = N118 & N147;
  assign N247 = N118 & \nz.addr_r [6];
  assign N248 = N120 & N147;
  assign N249 = N120 & \nz.addr_r [6];
  assign N250 = N122 & N147;
  assign N251 = N122 & \nz.addr_r [6];
  assign N252 = N124 & N147;
  assign N253 = N124 & \nz.addr_r [6];
  assign N254 = N126 & N147;
  assign N255 = N126 & \nz.addr_r [6];
  assign N256 = N128 & N147;
  assign N257 = N128 & \nz.addr_r [6];
  assign N258 = N130 & N147;
  assign N259 = N130 & \nz.addr_r [6];
  assign N260 = N132 & N147;
  assign N261 = N132 & \nz.addr_r [6];
  assign N262 = N134 & N147;
  assign N263 = N134 & \nz.addr_r [6];
  assign N264 = N136 & N147;
  assign N265 = N136 & \nz.addr_r [6];
  assign N266 = N138 & N147;
  assign N267 = N138 & \nz.addr_r [6];
  assign N268 = N140 & N147;
  assign N269 = N140 & \nz.addr_r [6];
  assign N270 = N142 & N147;
  assign N271 = N142 & \nz.addr_r [6];
  assign N272 = N144 & N147;
  assign N273 = N144 & \nz.addr_r [6];
  assign N274 = N146 & N147;
  assign N275 = N146 & \nz.addr_r [6];
  assign N276 = ~\nz.addr_r [7];
  assign N277 = N148 & N276;
  assign N278 = N148 & \nz.addr_r [7];
  assign N279 = N150 & N276;
  assign N280 = N150 & \nz.addr_r [7];
  assign N281 = N152 & N276;
  assign N282 = N152 & \nz.addr_r [7];
  assign N283 = N154 & N276;
  assign N284 = N154 & \nz.addr_r [7];
  assign N285 = N156 & N276;
  assign N286 = N156 & \nz.addr_r [7];
  assign N287 = N158 & N276;
  assign N288 = N158 & \nz.addr_r [7];
  assign N289 = N160 & N276;
  assign N290 = N160 & \nz.addr_r [7];
  assign N291 = N162 & N276;
  assign N292 = N162 & \nz.addr_r [7];
  assign N293 = N164 & N276;
  assign N294 = N164 & \nz.addr_r [7];
  assign N295 = N166 & N276;
  assign N296 = N166 & \nz.addr_r [7];
  assign N297 = N168 & N276;
  assign N298 = N168 & \nz.addr_r [7];
  assign N299 = N170 & N276;
  assign N300 = N170 & \nz.addr_r [7];
  assign N301 = N172 & N276;
  assign N302 = N172 & \nz.addr_r [7];
  assign N303 = N174 & N276;
  assign N304 = N174 & \nz.addr_r [7];
  assign N305 = N176 & N276;
  assign N306 = N176 & \nz.addr_r [7];
  assign N307 = N178 & N276;
  assign N308 = N178 & \nz.addr_r [7];
  assign N309 = N180 & N276;
  assign N310 = N180 & \nz.addr_r [7];
  assign N311 = N182 & N276;
  assign N312 = N182 & \nz.addr_r [7];
  assign N313 = N184 & N276;
  assign N314 = N184 & \nz.addr_r [7];
  assign N315 = N186 & N276;
  assign N316 = N186 & \nz.addr_r [7];
  assign N317 = N188 & N276;
  assign N318 = N188 & \nz.addr_r [7];
  assign N319 = N190 & N276;
  assign N320 = N190 & \nz.addr_r [7];
  assign N321 = N192 & N276;
  assign N322 = N192 & \nz.addr_r [7];
  assign N323 = N194 & N276;
  assign N324 = N194 & \nz.addr_r [7];
  assign N325 = N196 & N276;
  assign N326 = N196 & \nz.addr_r [7];
  assign N327 = N198 & N276;
  assign N328 = N198 & \nz.addr_r [7];
  assign N329 = N200 & N276;
  assign N330 = N200 & \nz.addr_r [7];
  assign N331 = N202 & N276;
  assign N332 = N202 & \nz.addr_r [7];
  assign N333 = N204 & N276;
  assign N334 = N204 & \nz.addr_r [7];
  assign N335 = N206 & N276;
  assign N336 = N206 & \nz.addr_r [7];
  assign N337 = N208 & N276;
  assign N338 = N208 & \nz.addr_r [7];
  assign N339 = N210 & N276;
  assign N340 = N210 & \nz.addr_r [7];
  assign N341 = N212 & N276;
  assign N342 = N212 & \nz.addr_r [7];
  assign N343 = N214 & N276;
  assign N344 = N214 & \nz.addr_r [7];
  assign N345 = N216 & N276;
  assign N346 = N216 & \nz.addr_r [7];
  assign N347 = N218 & N276;
  assign N348 = N218 & \nz.addr_r [7];
  assign N349 = N220 & N276;
  assign N350 = N220 & \nz.addr_r [7];
  assign N351 = N222 & N276;
  assign N352 = N222 & \nz.addr_r [7];
  assign N353 = N224 & N276;
  assign N354 = N224 & \nz.addr_r [7];
  assign N355 = N226 & N276;
  assign N356 = N226 & \nz.addr_r [7];
  assign N357 = N228 & N276;
  assign N358 = N228 & \nz.addr_r [7];
  assign N359 = N230 & N276;
  assign N360 = N230 & \nz.addr_r [7];
  assign N361 = N232 & N276;
  assign N362 = N232 & \nz.addr_r [7];
  assign N363 = N234 & N276;
  assign N364 = N234 & \nz.addr_r [7];
  assign N365 = N236 & N276;
  assign N366 = N236 & \nz.addr_r [7];
  assign N367 = N238 & N276;
  assign N368 = N238 & \nz.addr_r [7];
  assign N369 = N240 & N276;
  assign N370 = N240 & \nz.addr_r [7];
  assign N371 = N242 & N276;
  assign N372 = N242 & \nz.addr_r [7];
  assign N373 = N244 & N276;
  assign N374 = N244 & \nz.addr_r [7];
  assign N375 = N246 & N276;
  assign N376 = N246 & \nz.addr_r [7];
  assign N377 = N248 & N276;
  assign N378 = N248 & \nz.addr_r [7];
  assign N379 = N250 & N276;
  assign N380 = N250 & \nz.addr_r [7];
  assign N381 = N252 & N276;
  assign N382 = N252 & \nz.addr_r [7];
  assign N383 = N254 & N276;
  assign N384 = N254 & \nz.addr_r [7];
  assign N385 = N256 & N276;
  assign N386 = N256 & \nz.addr_r [7];
  assign N387 = N258 & N276;
  assign N388 = N258 & \nz.addr_r [7];
  assign N389 = N260 & N276;
  assign N390 = N260 & \nz.addr_r [7];
  assign N391 = N262 & N276;
  assign N392 = N262 & \nz.addr_r [7];
  assign N393 = N264 & N276;
  assign N394 = N264 & \nz.addr_r [7];
  assign N395 = N266 & N276;
  assign N396 = N266 & \nz.addr_r [7];
  assign N397 = N268 & N276;
  assign N398 = N268 & \nz.addr_r [7];
  assign N399 = N270 & N276;
  assign N400 = N270 & \nz.addr_r [7];
  assign N401 = N272 & N276;
  assign N402 = N272 & \nz.addr_r [7];
  assign N403 = N274 & N276;
  assign N404 = N274 & \nz.addr_r [7];
  assign N405 = N149 & N276;
  assign N406 = N149 & \nz.addr_r [7];
  assign N407 = N151 & N276;
  assign N408 = N151 & \nz.addr_r [7];
  assign N409 = N153 & N276;
  assign N410 = N153 & \nz.addr_r [7];
  assign N411 = N155 & N276;
  assign N412 = N155 & \nz.addr_r [7];
  assign N413 = N157 & N276;
  assign N414 = N157 & \nz.addr_r [7];
  assign N415 = N159 & N276;
  assign N416 = N159 & \nz.addr_r [7];
  assign N417 = N161 & N276;
  assign N418 = N161 & \nz.addr_r [7];
  assign N419 = N163 & N276;
  assign N420 = N163 & \nz.addr_r [7];
  assign N421 = N165 & N276;
  assign N422 = N165 & \nz.addr_r [7];
  assign N423 = N167 & N276;
  assign N424 = N167 & \nz.addr_r [7];
  assign N425 = N169 & N276;
  assign N426 = N169 & \nz.addr_r [7];
  assign N427 = N171 & N276;
  assign N428 = N171 & \nz.addr_r [7];
  assign N429 = N173 & N276;
  assign N430 = N173 & \nz.addr_r [7];
  assign N431 = N175 & N276;
  assign N432 = N175 & \nz.addr_r [7];
  assign N433 = N177 & N276;
  assign N434 = N177 & \nz.addr_r [7];
  assign N435 = N179 & N276;
  assign N436 = N179 & \nz.addr_r [7];
  assign N437 = N181 & N276;
  assign N438 = N181 & \nz.addr_r [7];
  assign N439 = N183 & N276;
  assign N440 = N183 & \nz.addr_r [7];
  assign N441 = N185 & N276;
  assign N442 = N185 & \nz.addr_r [7];
  assign N443 = N187 & N276;
  assign N444 = N187 & \nz.addr_r [7];
  assign N445 = N189 & N276;
  assign N446 = N189 & \nz.addr_r [7];
  assign N447 = N191 & N276;
  assign N448 = N191 & \nz.addr_r [7];
  assign N449 = N193 & N276;
  assign N450 = N193 & \nz.addr_r [7];
  assign N451 = N195 & N276;
  assign N452 = N195 & \nz.addr_r [7];
  assign N453 = N197 & N276;
  assign N454 = N197 & \nz.addr_r [7];
  assign N455 = N199 & N276;
  assign N456 = N199 & \nz.addr_r [7];
  assign N457 = N201 & N276;
  assign N458 = N201 & \nz.addr_r [7];
  assign N459 = N203 & N276;
  assign N460 = N203 & \nz.addr_r [7];
  assign N461 = N205 & N276;
  assign N462 = N205 & \nz.addr_r [7];
  assign N463 = N207 & N276;
  assign N464 = N207 & \nz.addr_r [7];
  assign N465 = N209 & N276;
  assign N466 = N209 & \nz.addr_r [7];
  assign N467 = N211 & N276;
  assign N468 = N211 & \nz.addr_r [7];
  assign N469 = N213 & N276;
  assign N470 = N213 & \nz.addr_r [7];
  assign N471 = N215 & N276;
  assign N472 = N215 & \nz.addr_r [7];
  assign N473 = N217 & N276;
  assign N474 = N217 & \nz.addr_r [7];
  assign N475 = N219 & N276;
  assign N476 = N219 & \nz.addr_r [7];
  assign N477 = N221 & N276;
  assign N478 = N221 & \nz.addr_r [7];
  assign N479 = N223 & N276;
  assign N480 = N223 & \nz.addr_r [7];
  assign N481 = N225 & N276;
  assign N482 = N225 & \nz.addr_r [7];
  assign N483 = N227 & N276;
  assign N484 = N227 & \nz.addr_r [7];
  assign N485 = N229 & N276;
  assign N486 = N229 & \nz.addr_r [7];
  assign N487 = N231 & N276;
  assign N488 = N231 & \nz.addr_r [7];
  assign N489 = N233 & N276;
  assign N490 = N233 & \nz.addr_r [7];
  assign N491 = N235 & N276;
  assign N492 = N235 & \nz.addr_r [7];
  assign N493 = N237 & N276;
  assign N494 = N237 & \nz.addr_r [7];
  assign N495 = N239 & N276;
  assign N496 = N239 & \nz.addr_r [7];
  assign N497 = N241 & N276;
  assign N498 = N241 & \nz.addr_r [7];
  assign N499 = N243 & N276;
  assign N500 = N243 & \nz.addr_r [7];
  assign N501 = N245 & N276;
  assign N502 = N245 & \nz.addr_r [7];
  assign N503 = N247 & N276;
  assign N504 = N247 & \nz.addr_r [7];
  assign N505 = N249 & N276;
  assign N506 = N249 & \nz.addr_r [7];
  assign N507 = N251 & N276;
  assign N508 = N251 & \nz.addr_r [7];
  assign N509 = N253 & N276;
  assign N510 = N253 & \nz.addr_r [7];
  assign N511 = N255 & N276;
  assign N512 = N255 & \nz.addr_r [7];
  assign N513 = N257 & N276;
  assign N514 = N257 & \nz.addr_r [7];
  assign N515 = N259 & N276;
  assign N516 = N259 & \nz.addr_r [7];
  assign N517 = N261 & N276;
  assign N518 = N261 & \nz.addr_r [7];
  assign N519 = N263 & N276;
  assign N520 = N263 & \nz.addr_r [7];
  assign N521 = N265 & N276;
  assign N522 = N265 & \nz.addr_r [7];
  assign N523 = N267 & N276;
  assign N524 = N267 & \nz.addr_r [7];
  assign N525 = N269 & N276;
  assign N526 = N269 & \nz.addr_r [7];
  assign N527 = N271 & N276;
  assign N528 = N271 & \nz.addr_r [7];
  assign N529 = N273 & N276;
  assign N530 = N273 & \nz.addr_r [7];
  assign N531 = N275 & N276;
  assign N532 = N275 & \nz.addr_r [7];
  assign N533 = v_i & w_i;
  assign N534 = ~N533;

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_7_sv2v_reg  <= addr_i[7];
      \nz.addr_r_6_sv2v_reg  <= addr_i[6];
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N1046) begin
      \nz.mem_2047_sv2v_reg  <= data_i[7];
      \nz.mem_2046_sv2v_reg  <= data_i[6];
      \nz.mem_2045_sv2v_reg  <= data_i[5];
      \nz.mem_2044_sv2v_reg  <= data_i[4];
      \nz.mem_2043_sv2v_reg  <= data_i[3];
      \nz.mem_2042_sv2v_reg  <= data_i[2];
      \nz.mem_2041_sv2v_reg  <= data_i[1];
      \nz.mem_2040_sv2v_reg  <= data_i[0];
    end 
    if(N1045) begin
      \nz.mem_2039_sv2v_reg  <= data_i[7];
      \nz.mem_2038_sv2v_reg  <= data_i[6];
      \nz.mem_2037_sv2v_reg  <= data_i[5];
      \nz.mem_2036_sv2v_reg  <= data_i[4];
      \nz.mem_2035_sv2v_reg  <= data_i[3];
      \nz.mem_2034_sv2v_reg  <= data_i[2];
      \nz.mem_2033_sv2v_reg  <= data_i[1];
      \nz.mem_2032_sv2v_reg  <= data_i[0];
    end 
    if(N1044) begin
      \nz.mem_2031_sv2v_reg  <= data_i[7];
      \nz.mem_2030_sv2v_reg  <= data_i[6];
      \nz.mem_2029_sv2v_reg  <= data_i[5];
      \nz.mem_2028_sv2v_reg  <= data_i[4];
      \nz.mem_2027_sv2v_reg  <= data_i[3];
      \nz.mem_2026_sv2v_reg  <= data_i[2];
      \nz.mem_2025_sv2v_reg  <= data_i[1];
      \nz.mem_2024_sv2v_reg  <= data_i[0];
    end 
    if(N1043) begin
      \nz.mem_2023_sv2v_reg  <= data_i[7];
      \nz.mem_2022_sv2v_reg  <= data_i[6];
      \nz.mem_2021_sv2v_reg  <= data_i[5];
      \nz.mem_2020_sv2v_reg  <= data_i[4];
      \nz.mem_2019_sv2v_reg  <= data_i[3];
      \nz.mem_2018_sv2v_reg  <= data_i[2];
      \nz.mem_2017_sv2v_reg  <= data_i[1];
      \nz.mem_2016_sv2v_reg  <= data_i[0];
    end 
    if(N1042) begin
      \nz.mem_2015_sv2v_reg  <= data_i[7];
      \nz.mem_2014_sv2v_reg  <= data_i[6];
      \nz.mem_2013_sv2v_reg  <= data_i[5];
      \nz.mem_2012_sv2v_reg  <= data_i[4];
      \nz.mem_2011_sv2v_reg  <= data_i[3];
      \nz.mem_2010_sv2v_reg  <= data_i[2];
      \nz.mem_2009_sv2v_reg  <= data_i[1];
      \nz.mem_2008_sv2v_reg  <= data_i[0];
    end 
    if(N1041) begin
      \nz.mem_2007_sv2v_reg  <= data_i[7];
      \nz.mem_2006_sv2v_reg  <= data_i[6];
      \nz.mem_2005_sv2v_reg  <= data_i[5];
      \nz.mem_2004_sv2v_reg  <= data_i[4];
      \nz.mem_2003_sv2v_reg  <= data_i[3];
      \nz.mem_2002_sv2v_reg  <= data_i[2];
      \nz.mem_2001_sv2v_reg  <= data_i[1];
      \nz.mem_2000_sv2v_reg  <= data_i[0];
    end 
    if(N1040) begin
      \nz.mem_1999_sv2v_reg  <= data_i[7];
      \nz.mem_1998_sv2v_reg  <= data_i[6];
      \nz.mem_1997_sv2v_reg  <= data_i[5];
      \nz.mem_1996_sv2v_reg  <= data_i[4];
      \nz.mem_1995_sv2v_reg  <= data_i[3];
      \nz.mem_1994_sv2v_reg  <= data_i[2];
      \nz.mem_1993_sv2v_reg  <= data_i[1];
      \nz.mem_1992_sv2v_reg  <= data_i[0];
    end 
    if(N1039) begin
      \nz.mem_1991_sv2v_reg  <= data_i[7];
      \nz.mem_1990_sv2v_reg  <= data_i[6];
      \nz.mem_1989_sv2v_reg  <= data_i[5];
      \nz.mem_1988_sv2v_reg  <= data_i[4];
      \nz.mem_1987_sv2v_reg  <= data_i[3];
      \nz.mem_1986_sv2v_reg  <= data_i[2];
      \nz.mem_1985_sv2v_reg  <= data_i[1];
      \nz.mem_1984_sv2v_reg  <= data_i[0];
    end 
    if(N1038) begin
      \nz.mem_1983_sv2v_reg  <= data_i[7];
      \nz.mem_1982_sv2v_reg  <= data_i[6];
      \nz.mem_1981_sv2v_reg  <= data_i[5];
      \nz.mem_1980_sv2v_reg  <= data_i[4];
      \nz.mem_1979_sv2v_reg  <= data_i[3];
      \nz.mem_1978_sv2v_reg  <= data_i[2];
      \nz.mem_1977_sv2v_reg  <= data_i[1];
      \nz.mem_1976_sv2v_reg  <= data_i[0];
    end 
    if(N1037) begin
      \nz.mem_1975_sv2v_reg  <= data_i[7];
      \nz.mem_1974_sv2v_reg  <= data_i[6];
      \nz.mem_1973_sv2v_reg  <= data_i[5];
      \nz.mem_1972_sv2v_reg  <= data_i[4];
      \nz.mem_1971_sv2v_reg  <= data_i[3];
      \nz.mem_1970_sv2v_reg  <= data_i[2];
      \nz.mem_1969_sv2v_reg  <= data_i[1];
      \nz.mem_1968_sv2v_reg  <= data_i[0];
    end 
    if(N1036) begin
      \nz.mem_1967_sv2v_reg  <= data_i[7];
      \nz.mem_1966_sv2v_reg  <= data_i[6];
      \nz.mem_1965_sv2v_reg  <= data_i[5];
      \nz.mem_1964_sv2v_reg  <= data_i[4];
      \nz.mem_1963_sv2v_reg  <= data_i[3];
      \nz.mem_1962_sv2v_reg  <= data_i[2];
      \nz.mem_1961_sv2v_reg  <= data_i[1];
      \nz.mem_1960_sv2v_reg  <= data_i[0];
    end 
    if(N1035) begin
      \nz.mem_1959_sv2v_reg  <= data_i[7];
      \nz.mem_1958_sv2v_reg  <= data_i[6];
      \nz.mem_1957_sv2v_reg  <= data_i[5];
      \nz.mem_1956_sv2v_reg  <= data_i[4];
      \nz.mem_1955_sv2v_reg  <= data_i[3];
      \nz.mem_1954_sv2v_reg  <= data_i[2];
      \nz.mem_1953_sv2v_reg  <= data_i[1];
      \nz.mem_1952_sv2v_reg  <= data_i[0];
    end 
    if(N1034) begin
      \nz.mem_1951_sv2v_reg  <= data_i[7];
      \nz.mem_1950_sv2v_reg  <= data_i[6];
      \nz.mem_1949_sv2v_reg  <= data_i[5];
      \nz.mem_1948_sv2v_reg  <= data_i[4];
      \nz.mem_1947_sv2v_reg  <= data_i[3];
      \nz.mem_1946_sv2v_reg  <= data_i[2];
      \nz.mem_1945_sv2v_reg  <= data_i[1];
      \nz.mem_1944_sv2v_reg  <= data_i[0];
    end 
    if(N1033) begin
      \nz.mem_1943_sv2v_reg  <= data_i[7];
      \nz.mem_1942_sv2v_reg  <= data_i[6];
      \nz.mem_1941_sv2v_reg  <= data_i[5];
      \nz.mem_1940_sv2v_reg  <= data_i[4];
      \nz.mem_1939_sv2v_reg  <= data_i[3];
      \nz.mem_1938_sv2v_reg  <= data_i[2];
      \nz.mem_1937_sv2v_reg  <= data_i[1];
      \nz.mem_1936_sv2v_reg  <= data_i[0];
    end 
    if(N1032) begin
      \nz.mem_1935_sv2v_reg  <= data_i[7];
      \nz.mem_1934_sv2v_reg  <= data_i[6];
      \nz.mem_1933_sv2v_reg  <= data_i[5];
      \nz.mem_1932_sv2v_reg  <= data_i[4];
      \nz.mem_1931_sv2v_reg  <= data_i[3];
      \nz.mem_1930_sv2v_reg  <= data_i[2];
      \nz.mem_1929_sv2v_reg  <= data_i[1];
      \nz.mem_1928_sv2v_reg  <= data_i[0];
    end 
    if(N1031) begin
      \nz.mem_1927_sv2v_reg  <= data_i[7];
      \nz.mem_1926_sv2v_reg  <= data_i[6];
      \nz.mem_1925_sv2v_reg  <= data_i[5];
      \nz.mem_1924_sv2v_reg  <= data_i[4];
      \nz.mem_1923_sv2v_reg  <= data_i[3];
      \nz.mem_1922_sv2v_reg  <= data_i[2];
      \nz.mem_1921_sv2v_reg  <= data_i[1];
      \nz.mem_1920_sv2v_reg  <= data_i[0];
    end 
    if(N1030) begin
      \nz.mem_1919_sv2v_reg  <= data_i[7];
      \nz.mem_1918_sv2v_reg  <= data_i[6];
      \nz.mem_1917_sv2v_reg  <= data_i[5];
      \nz.mem_1916_sv2v_reg  <= data_i[4];
      \nz.mem_1915_sv2v_reg  <= data_i[3];
      \nz.mem_1914_sv2v_reg  <= data_i[2];
      \nz.mem_1913_sv2v_reg  <= data_i[1];
      \nz.mem_1912_sv2v_reg  <= data_i[0];
    end 
    if(N1029) begin
      \nz.mem_1911_sv2v_reg  <= data_i[7];
      \nz.mem_1910_sv2v_reg  <= data_i[6];
      \nz.mem_1909_sv2v_reg  <= data_i[5];
      \nz.mem_1908_sv2v_reg  <= data_i[4];
      \nz.mem_1907_sv2v_reg  <= data_i[3];
      \nz.mem_1906_sv2v_reg  <= data_i[2];
      \nz.mem_1905_sv2v_reg  <= data_i[1];
      \nz.mem_1904_sv2v_reg  <= data_i[0];
    end 
    if(N1028) begin
      \nz.mem_1903_sv2v_reg  <= data_i[7];
      \nz.mem_1902_sv2v_reg  <= data_i[6];
      \nz.mem_1901_sv2v_reg  <= data_i[5];
      \nz.mem_1900_sv2v_reg  <= data_i[4];
      \nz.mem_1899_sv2v_reg  <= data_i[3];
      \nz.mem_1898_sv2v_reg  <= data_i[2];
      \nz.mem_1897_sv2v_reg  <= data_i[1];
      \nz.mem_1896_sv2v_reg  <= data_i[0];
    end 
    if(N1027) begin
      \nz.mem_1895_sv2v_reg  <= data_i[7];
      \nz.mem_1894_sv2v_reg  <= data_i[6];
      \nz.mem_1893_sv2v_reg  <= data_i[5];
      \nz.mem_1892_sv2v_reg  <= data_i[4];
      \nz.mem_1891_sv2v_reg  <= data_i[3];
      \nz.mem_1890_sv2v_reg  <= data_i[2];
      \nz.mem_1889_sv2v_reg  <= data_i[1];
      \nz.mem_1888_sv2v_reg  <= data_i[0];
    end 
    if(N1026) begin
      \nz.mem_1887_sv2v_reg  <= data_i[7];
      \nz.mem_1886_sv2v_reg  <= data_i[6];
      \nz.mem_1885_sv2v_reg  <= data_i[5];
      \nz.mem_1884_sv2v_reg  <= data_i[4];
      \nz.mem_1883_sv2v_reg  <= data_i[3];
      \nz.mem_1882_sv2v_reg  <= data_i[2];
      \nz.mem_1881_sv2v_reg  <= data_i[1];
      \nz.mem_1880_sv2v_reg  <= data_i[0];
    end 
    if(N1025) begin
      \nz.mem_1879_sv2v_reg  <= data_i[7];
      \nz.mem_1878_sv2v_reg  <= data_i[6];
      \nz.mem_1877_sv2v_reg  <= data_i[5];
      \nz.mem_1876_sv2v_reg  <= data_i[4];
      \nz.mem_1875_sv2v_reg  <= data_i[3];
      \nz.mem_1874_sv2v_reg  <= data_i[2];
      \nz.mem_1873_sv2v_reg  <= data_i[1];
      \nz.mem_1872_sv2v_reg  <= data_i[0];
    end 
    if(N1024) begin
      \nz.mem_1871_sv2v_reg  <= data_i[7];
      \nz.mem_1870_sv2v_reg  <= data_i[6];
      \nz.mem_1869_sv2v_reg  <= data_i[5];
      \nz.mem_1868_sv2v_reg  <= data_i[4];
      \nz.mem_1867_sv2v_reg  <= data_i[3];
      \nz.mem_1866_sv2v_reg  <= data_i[2];
      \nz.mem_1865_sv2v_reg  <= data_i[1];
      \nz.mem_1864_sv2v_reg  <= data_i[0];
    end 
    if(N1023) begin
      \nz.mem_1863_sv2v_reg  <= data_i[7];
      \nz.mem_1862_sv2v_reg  <= data_i[6];
      \nz.mem_1861_sv2v_reg  <= data_i[5];
      \nz.mem_1860_sv2v_reg  <= data_i[4];
      \nz.mem_1859_sv2v_reg  <= data_i[3];
      \nz.mem_1858_sv2v_reg  <= data_i[2];
      \nz.mem_1857_sv2v_reg  <= data_i[1];
      \nz.mem_1856_sv2v_reg  <= data_i[0];
    end 
    if(N1022) begin
      \nz.mem_1855_sv2v_reg  <= data_i[7];
      \nz.mem_1854_sv2v_reg  <= data_i[6];
      \nz.mem_1853_sv2v_reg  <= data_i[5];
      \nz.mem_1852_sv2v_reg  <= data_i[4];
      \nz.mem_1851_sv2v_reg  <= data_i[3];
      \nz.mem_1850_sv2v_reg  <= data_i[2];
      \nz.mem_1849_sv2v_reg  <= data_i[1];
      \nz.mem_1848_sv2v_reg  <= data_i[0];
    end 
    if(N1021) begin
      \nz.mem_1847_sv2v_reg  <= data_i[7];
      \nz.mem_1846_sv2v_reg  <= data_i[6];
      \nz.mem_1845_sv2v_reg  <= data_i[5];
      \nz.mem_1844_sv2v_reg  <= data_i[4];
      \nz.mem_1843_sv2v_reg  <= data_i[3];
      \nz.mem_1842_sv2v_reg  <= data_i[2];
      \nz.mem_1841_sv2v_reg  <= data_i[1];
      \nz.mem_1840_sv2v_reg  <= data_i[0];
    end 
    if(N1020) begin
      \nz.mem_1839_sv2v_reg  <= data_i[7];
      \nz.mem_1838_sv2v_reg  <= data_i[6];
      \nz.mem_1837_sv2v_reg  <= data_i[5];
      \nz.mem_1836_sv2v_reg  <= data_i[4];
      \nz.mem_1835_sv2v_reg  <= data_i[3];
      \nz.mem_1834_sv2v_reg  <= data_i[2];
      \nz.mem_1833_sv2v_reg  <= data_i[1];
      \nz.mem_1832_sv2v_reg  <= data_i[0];
    end 
    if(N1019) begin
      \nz.mem_1831_sv2v_reg  <= data_i[7];
      \nz.mem_1830_sv2v_reg  <= data_i[6];
      \nz.mem_1829_sv2v_reg  <= data_i[5];
      \nz.mem_1828_sv2v_reg  <= data_i[4];
      \nz.mem_1827_sv2v_reg  <= data_i[3];
      \nz.mem_1826_sv2v_reg  <= data_i[2];
      \nz.mem_1825_sv2v_reg  <= data_i[1];
      \nz.mem_1824_sv2v_reg  <= data_i[0];
    end 
    if(N1018) begin
      \nz.mem_1823_sv2v_reg  <= data_i[7];
      \nz.mem_1822_sv2v_reg  <= data_i[6];
      \nz.mem_1821_sv2v_reg  <= data_i[5];
      \nz.mem_1820_sv2v_reg  <= data_i[4];
      \nz.mem_1819_sv2v_reg  <= data_i[3];
      \nz.mem_1818_sv2v_reg  <= data_i[2];
      \nz.mem_1817_sv2v_reg  <= data_i[1];
      \nz.mem_1816_sv2v_reg  <= data_i[0];
    end 
    if(N1017) begin
      \nz.mem_1815_sv2v_reg  <= data_i[7];
      \nz.mem_1814_sv2v_reg  <= data_i[6];
      \nz.mem_1813_sv2v_reg  <= data_i[5];
      \nz.mem_1812_sv2v_reg  <= data_i[4];
      \nz.mem_1811_sv2v_reg  <= data_i[3];
      \nz.mem_1810_sv2v_reg  <= data_i[2];
      \nz.mem_1809_sv2v_reg  <= data_i[1];
      \nz.mem_1808_sv2v_reg  <= data_i[0];
    end 
    if(N1016) begin
      \nz.mem_1807_sv2v_reg  <= data_i[7];
      \nz.mem_1806_sv2v_reg  <= data_i[6];
      \nz.mem_1805_sv2v_reg  <= data_i[5];
      \nz.mem_1804_sv2v_reg  <= data_i[4];
      \nz.mem_1803_sv2v_reg  <= data_i[3];
      \nz.mem_1802_sv2v_reg  <= data_i[2];
      \nz.mem_1801_sv2v_reg  <= data_i[1];
      \nz.mem_1800_sv2v_reg  <= data_i[0];
    end 
    if(N1015) begin
      \nz.mem_1799_sv2v_reg  <= data_i[7];
      \nz.mem_1798_sv2v_reg  <= data_i[6];
      \nz.mem_1797_sv2v_reg  <= data_i[5];
      \nz.mem_1796_sv2v_reg  <= data_i[4];
      \nz.mem_1795_sv2v_reg  <= data_i[3];
      \nz.mem_1794_sv2v_reg  <= data_i[2];
      \nz.mem_1793_sv2v_reg  <= data_i[1];
      \nz.mem_1792_sv2v_reg  <= data_i[0];
    end 
    if(N1014) begin
      \nz.mem_1791_sv2v_reg  <= data_i[7];
      \nz.mem_1790_sv2v_reg  <= data_i[6];
      \nz.mem_1789_sv2v_reg  <= data_i[5];
      \nz.mem_1788_sv2v_reg  <= data_i[4];
      \nz.mem_1787_sv2v_reg  <= data_i[3];
      \nz.mem_1786_sv2v_reg  <= data_i[2];
      \nz.mem_1785_sv2v_reg  <= data_i[1];
      \nz.mem_1784_sv2v_reg  <= data_i[0];
    end 
    if(N1013) begin
      \nz.mem_1783_sv2v_reg  <= data_i[7];
      \nz.mem_1782_sv2v_reg  <= data_i[6];
      \nz.mem_1781_sv2v_reg  <= data_i[5];
      \nz.mem_1780_sv2v_reg  <= data_i[4];
      \nz.mem_1779_sv2v_reg  <= data_i[3];
      \nz.mem_1778_sv2v_reg  <= data_i[2];
      \nz.mem_1777_sv2v_reg  <= data_i[1];
      \nz.mem_1776_sv2v_reg  <= data_i[0];
    end 
    if(N1012) begin
      \nz.mem_1775_sv2v_reg  <= data_i[7];
      \nz.mem_1774_sv2v_reg  <= data_i[6];
      \nz.mem_1773_sv2v_reg  <= data_i[5];
      \nz.mem_1772_sv2v_reg  <= data_i[4];
      \nz.mem_1771_sv2v_reg  <= data_i[3];
      \nz.mem_1770_sv2v_reg  <= data_i[2];
      \nz.mem_1769_sv2v_reg  <= data_i[1];
      \nz.mem_1768_sv2v_reg  <= data_i[0];
    end 
    if(N1011) begin
      \nz.mem_1767_sv2v_reg  <= data_i[7];
      \nz.mem_1766_sv2v_reg  <= data_i[6];
      \nz.mem_1765_sv2v_reg  <= data_i[5];
      \nz.mem_1764_sv2v_reg  <= data_i[4];
      \nz.mem_1763_sv2v_reg  <= data_i[3];
      \nz.mem_1762_sv2v_reg  <= data_i[2];
      \nz.mem_1761_sv2v_reg  <= data_i[1];
      \nz.mem_1760_sv2v_reg  <= data_i[0];
    end 
    if(N1010) begin
      \nz.mem_1759_sv2v_reg  <= data_i[7];
      \nz.mem_1758_sv2v_reg  <= data_i[6];
      \nz.mem_1757_sv2v_reg  <= data_i[5];
      \nz.mem_1756_sv2v_reg  <= data_i[4];
      \nz.mem_1755_sv2v_reg  <= data_i[3];
      \nz.mem_1754_sv2v_reg  <= data_i[2];
      \nz.mem_1753_sv2v_reg  <= data_i[1];
      \nz.mem_1752_sv2v_reg  <= data_i[0];
    end 
    if(N1009) begin
      \nz.mem_1751_sv2v_reg  <= data_i[7];
      \nz.mem_1750_sv2v_reg  <= data_i[6];
      \nz.mem_1749_sv2v_reg  <= data_i[5];
      \nz.mem_1748_sv2v_reg  <= data_i[4];
      \nz.mem_1747_sv2v_reg  <= data_i[3];
      \nz.mem_1746_sv2v_reg  <= data_i[2];
      \nz.mem_1745_sv2v_reg  <= data_i[1];
      \nz.mem_1744_sv2v_reg  <= data_i[0];
    end 
    if(N1008) begin
      \nz.mem_1743_sv2v_reg  <= data_i[7];
      \nz.mem_1742_sv2v_reg  <= data_i[6];
      \nz.mem_1741_sv2v_reg  <= data_i[5];
      \nz.mem_1740_sv2v_reg  <= data_i[4];
      \nz.mem_1739_sv2v_reg  <= data_i[3];
      \nz.mem_1738_sv2v_reg  <= data_i[2];
      \nz.mem_1737_sv2v_reg  <= data_i[1];
      \nz.mem_1736_sv2v_reg  <= data_i[0];
    end 
    if(N1007) begin
      \nz.mem_1735_sv2v_reg  <= data_i[7];
      \nz.mem_1734_sv2v_reg  <= data_i[6];
      \nz.mem_1733_sv2v_reg  <= data_i[5];
      \nz.mem_1732_sv2v_reg  <= data_i[4];
      \nz.mem_1731_sv2v_reg  <= data_i[3];
      \nz.mem_1730_sv2v_reg  <= data_i[2];
      \nz.mem_1729_sv2v_reg  <= data_i[1];
      \nz.mem_1728_sv2v_reg  <= data_i[0];
    end 
    if(N1006) begin
      \nz.mem_1727_sv2v_reg  <= data_i[7];
      \nz.mem_1726_sv2v_reg  <= data_i[6];
      \nz.mem_1725_sv2v_reg  <= data_i[5];
      \nz.mem_1724_sv2v_reg  <= data_i[4];
      \nz.mem_1723_sv2v_reg  <= data_i[3];
      \nz.mem_1722_sv2v_reg  <= data_i[2];
      \nz.mem_1721_sv2v_reg  <= data_i[1];
      \nz.mem_1720_sv2v_reg  <= data_i[0];
    end 
    if(N1005) begin
      \nz.mem_1719_sv2v_reg  <= data_i[7];
      \nz.mem_1718_sv2v_reg  <= data_i[6];
      \nz.mem_1717_sv2v_reg  <= data_i[5];
      \nz.mem_1716_sv2v_reg  <= data_i[4];
      \nz.mem_1715_sv2v_reg  <= data_i[3];
      \nz.mem_1714_sv2v_reg  <= data_i[2];
      \nz.mem_1713_sv2v_reg  <= data_i[1];
      \nz.mem_1712_sv2v_reg  <= data_i[0];
    end 
    if(N1004) begin
      \nz.mem_1711_sv2v_reg  <= data_i[7];
      \nz.mem_1710_sv2v_reg  <= data_i[6];
      \nz.mem_1709_sv2v_reg  <= data_i[5];
      \nz.mem_1708_sv2v_reg  <= data_i[4];
      \nz.mem_1707_sv2v_reg  <= data_i[3];
      \nz.mem_1706_sv2v_reg  <= data_i[2];
      \nz.mem_1705_sv2v_reg  <= data_i[1];
      \nz.mem_1704_sv2v_reg  <= data_i[0];
    end 
    if(N1003) begin
      \nz.mem_1703_sv2v_reg  <= data_i[7];
      \nz.mem_1702_sv2v_reg  <= data_i[6];
      \nz.mem_1701_sv2v_reg  <= data_i[5];
      \nz.mem_1700_sv2v_reg  <= data_i[4];
      \nz.mem_1699_sv2v_reg  <= data_i[3];
      \nz.mem_1698_sv2v_reg  <= data_i[2];
      \nz.mem_1697_sv2v_reg  <= data_i[1];
      \nz.mem_1696_sv2v_reg  <= data_i[0];
    end 
    if(N1002) begin
      \nz.mem_1695_sv2v_reg  <= data_i[7];
      \nz.mem_1694_sv2v_reg  <= data_i[6];
      \nz.mem_1693_sv2v_reg  <= data_i[5];
      \nz.mem_1692_sv2v_reg  <= data_i[4];
      \nz.mem_1691_sv2v_reg  <= data_i[3];
      \nz.mem_1690_sv2v_reg  <= data_i[2];
      \nz.mem_1689_sv2v_reg  <= data_i[1];
      \nz.mem_1688_sv2v_reg  <= data_i[0];
    end 
    if(N1001) begin
      \nz.mem_1687_sv2v_reg  <= data_i[7];
      \nz.mem_1686_sv2v_reg  <= data_i[6];
      \nz.mem_1685_sv2v_reg  <= data_i[5];
      \nz.mem_1684_sv2v_reg  <= data_i[4];
      \nz.mem_1683_sv2v_reg  <= data_i[3];
      \nz.mem_1682_sv2v_reg  <= data_i[2];
      \nz.mem_1681_sv2v_reg  <= data_i[1];
      \nz.mem_1680_sv2v_reg  <= data_i[0];
    end 
    if(N1000) begin
      \nz.mem_1679_sv2v_reg  <= data_i[7];
      \nz.mem_1678_sv2v_reg  <= data_i[6];
      \nz.mem_1677_sv2v_reg  <= data_i[5];
      \nz.mem_1676_sv2v_reg  <= data_i[4];
      \nz.mem_1675_sv2v_reg  <= data_i[3];
      \nz.mem_1674_sv2v_reg  <= data_i[2];
      \nz.mem_1673_sv2v_reg  <= data_i[1];
      \nz.mem_1672_sv2v_reg  <= data_i[0];
    end 
    if(N999) begin
      \nz.mem_1671_sv2v_reg  <= data_i[7];
      \nz.mem_1670_sv2v_reg  <= data_i[6];
      \nz.mem_1669_sv2v_reg  <= data_i[5];
      \nz.mem_1668_sv2v_reg  <= data_i[4];
      \nz.mem_1667_sv2v_reg  <= data_i[3];
      \nz.mem_1666_sv2v_reg  <= data_i[2];
      \nz.mem_1665_sv2v_reg  <= data_i[1];
      \nz.mem_1664_sv2v_reg  <= data_i[0];
    end 
    if(N998) begin
      \nz.mem_1663_sv2v_reg  <= data_i[7];
      \nz.mem_1662_sv2v_reg  <= data_i[6];
      \nz.mem_1661_sv2v_reg  <= data_i[5];
      \nz.mem_1660_sv2v_reg  <= data_i[4];
      \nz.mem_1659_sv2v_reg  <= data_i[3];
      \nz.mem_1658_sv2v_reg  <= data_i[2];
      \nz.mem_1657_sv2v_reg  <= data_i[1];
      \nz.mem_1656_sv2v_reg  <= data_i[0];
    end 
    if(N997) begin
      \nz.mem_1655_sv2v_reg  <= data_i[7];
      \nz.mem_1654_sv2v_reg  <= data_i[6];
      \nz.mem_1653_sv2v_reg  <= data_i[5];
      \nz.mem_1652_sv2v_reg  <= data_i[4];
      \nz.mem_1651_sv2v_reg  <= data_i[3];
      \nz.mem_1650_sv2v_reg  <= data_i[2];
      \nz.mem_1649_sv2v_reg  <= data_i[1];
      \nz.mem_1648_sv2v_reg  <= data_i[0];
    end 
    if(N996) begin
      \nz.mem_1647_sv2v_reg  <= data_i[7];
      \nz.mem_1646_sv2v_reg  <= data_i[6];
      \nz.mem_1645_sv2v_reg  <= data_i[5];
      \nz.mem_1644_sv2v_reg  <= data_i[4];
      \nz.mem_1643_sv2v_reg  <= data_i[3];
      \nz.mem_1642_sv2v_reg  <= data_i[2];
      \nz.mem_1641_sv2v_reg  <= data_i[1];
      \nz.mem_1640_sv2v_reg  <= data_i[0];
    end 
    if(N995) begin
      \nz.mem_1639_sv2v_reg  <= data_i[7];
      \nz.mem_1638_sv2v_reg  <= data_i[6];
      \nz.mem_1637_sv2v_reg  <= data_i[5];
      \nz.mem_1636_sv2v_reg  <= data_i[4];
      \nz.mem_1635_sv2v_reg  <= data_i[3];
      \nz.mem_1634_sv2v_reg  <= data_i[2];
      \nz.mem_1633_sv2v_reg  <= data_i[1];
      \nz.mem_1632_sv2v_reg  <= data_i[0];
    end 
    if(N994) begin
      \nz.mem_1631_sv2v_reg  <= data_i[7];
      \nz.mem_1630_sv2v_reg  <= data_i[6];
      \nz.mem_1629_sv2v_reg  <= data_i[5];
      \nz.mem_1628_sv2v_reg  <= data_i[4];
      \nz.mem_1627_sv2v_reg  <= data_i[3];
      \nz.mem_1626_sv2v_reg  <= data_i[2];
      \nz.mem_1625_sv2v_reg  <= data_i[1];
      \nz.mem_1624_sv2v_reg  <= data_i[0];
    end 
    if(N993) begin
      \nz.mem_1623_sv2v_reg  <= data_i[7];
      \nz.mem_1622_sv2v_reg  <= data_i[6];
      \nz.mem_1621_sv2v_reg  <= data_i[5];
      \nz.mem_1620_sv2v_reg  <= data_i[4];
      \nz.mem_1619_sv2v_reg  <= data_i[3];
      \nz.mem_1618_sv2v_reg  <= data_i[2];
      \nz.mem_1617_sv2v_reg  <= data_i[1];
      \nz.mem_1616_sv2v_reg  <= data_i[0];
    end 
    if(N992) begin
      \nz.mem_1615_sv2v_reg  <= data_i[7];
      \nz.mem_1614_sv2v_reg  <= data_i[6];
      \nz.mem_1613_sv2v_reg  <= data_i[5];
      \nz.mem_1612_sv2v_reg  <= data_i[4];
      \nz.mem_1611_sv2v_reg  <= data_i[3];
      \nz.mem_1610_sv2v_reg  <= data_i[2];
      \nz.mem_1609_sv2v_reg  <= data_i[1];
      \nz.mem_1608_sv2v_reg  <= data_i[0];
    end 
    if(N991) begin
      \nz.mem_1607_sv2v_reg  <= data_i[7];
      \nz.mem_1606_sv2v_reg  <= data_i[6];
      \nz.mem_1605_sv2v_reg  <= data_i[5];
      \nz.mem_1604_sv2v_reg  <= data_i[4];
      \nz.mem_1603_sv2v_reg  <= data_i[3];
      \nz.mem_1602_sv2v_reg  <= data_i[2];
      \nz.mem_1601_sv2v_reg  <= data_i[1];
      \nz.mem_1600_sv2v_reg  <= data_i[0];
    end 
    if(N990) begin
      \nz.mem_1599_sv2v_reg  <= data_i[7];
      \nz.mem_1598_sv2v_reg  <= data_i[6];
      \nz.mem_1597_sv2v_reg  <= data_i[5];
      \nz.mem_1596_sv2v_reg  <= data_i[4];
      \nz.mem_1595_sv2v_reg  <= data_i[3];
      \nz.mem_1594_sv2v_reg  <= data_i[2];
      \nz.mem_1593_sv2v_reg  <= data_i[1];
      \nz.mem_1592_sv2v_reg  <= data_i[0];
    end 
    if(N989) begin
      \nz.mem_1591_sv2v_reg  <= data_i[7];
      \nz.mem_1590_sv2v_reg  <= data_i[6];
      \nz.mem_1589_sv2v_reg  <= data_i[5];
      \nz.mem_1588_sv2v_reg  <= data_i[4];
      \nz.mem_1587_sv2v_reg  <= data_i[3];
      \nz.mem_1586_sv2v_reg  <= data_i[2];
      \nz.mem_1585_sv2v_reg  <= data_i[1];
      \nz.mem_1584_sv2v_reg  <= data_i[0];
    end 
    if(N988) begin
      \nz.mem_1583_sv2v_reg  <= data_i[7];
      \nz.mem_1582_sv2v_reg  <= data_i[6];
      \nz.mem_1581_sv2v_reg  <= data_i[5];
      \nz.mem_1580_sv2v_reg  <= data_i[4];
      \nz.mem_1579_sv2v_reg  <= data_i[3];
      \nz.mem_1578_sv2v_reg  <= data_i[2];
      \nz.mem_1577_sv2v_reg  <= data_i[1];
      \nz.mem_1576_sv2v_reg  <= data_i[0];
    end 
    if(N987) begin
      \nz.mem_1575_sv2v_reg  <= data_i[7];
      \nz.mem_1574_sv2v_reg  <= data_i[6];
      \nz.mem_1573_sv2v_reg  <= data_i[5];
      \nz.mem_1572_sv2v_reg  <= data_i[4];
      \nz.mem_1571_sv2v_reg  <= data_i[3];
      \nz.mem_1570_sv2v_reg  <= data_i[2];
      \nz.mem_1569_sv2v_reg  <= data_i[1];
      \nz.mem_1568_sv2v_reg  <= data_i[0];
    end 
    if(N986) begin
      \nz.mem_1567_sv2v_reg  <= data_i[7];
      \nz.mem_1566_sv2v_reg  <= data_i[6];
      \nz.mem_1565_sv2v_reg  <= data_i[5];
      \nz.mem_1564_sv2v_reg  <= data_i[4];
      \nz.mem_1563_sv2v_reg  <= data_i[3];
      \nz.mem_1562_sv2v_reg  <= data_i[2];
      \nz.mem_1561_sv2v_reg  <= data_i[1];
      \nz.mem_1560_sv2v_reg  <= data_i[0];
    end 
    if(N985) begin
      \nz.mem_1559_sv2v_reg  <= data_i[7];
      \nz.mem_1558_sv2v_reg  <= data_i[6];
      \nz.mem_1557_sv2v_reg  <= data_i[5];
      \nz.mem_1556_sv2v_reg  <= data_i[4];
      \nz.mem_1555_sv2v_reg  <= data_i[3];
      \nz.mem_1554_sv2v_reg  <= data_i[2];
      \nz.mem_1553_sv2v_reg  <= data_i[1];
      \nz.mem_1552_sv2v_reg  <= data_i[0];
    end 
    if(N984) begin
      \nz.mem_1551_sv2v_reg  <= data_i[7];
      \nz.mem_1550_sv2v_reg  <= data_i[6];
      \nz.mem_1549_sv2v_reg  <= data_i[5];
      \nz.mem_1548_sv2v_reg  <= data_i[4];
      \nz.mem_1547_sv2v_reg  <= data_i[3];
      \nz.mem_1546_sv2v_reg  <= data_i[2];
      \nz.mem_1545_sv2v_reg  <= data_i[1];
      \nz.mem_1544_sv2v_reg  <= data_i[0];
    end 
    if(N983) begin
      \nz.mem_1543_sv2v_reg  <= data_i[7];
      \nz.mem_1542_sv2v_reg  <= data_i[6];
      \nz.mem_1541_sv2v_reg  <= data_i[5];
      \nz.mem_1540_sv2v_reg  <= data_i[4];
      \nz.mem_1539_sv2v_reg  <= data_i[3];
      \nz.mem_1538_sv2v_reg  <= data_i[2];
      \nz.mem_1537_sv2v_reg  <= data_i[1];
      \nz.mem_1536_sv2v_reg  <= data_i[0];
    end 
    if(N982) begin
      \nz.mem_1535_sv2v_reg  <= data_i[7];
      \nz.mem_1534_sv2v_reg  <= data_i[6];
      \nz.mem_1533_sv2v_reg  <= data_i[5];
      \nz.mem_1532_sv2v_reg  <= data_i[4];
      \nz.mem_1531_sv2v_reg  <= data_i[3];
      \nz.mem_1530_sv2v_reg  <= data_i[2];
      \nz.mem_1529_sv2v_reg  <= data_i[1];
      \nz.mem_1528_sv2v_reg  <= data_i[0];
    end 
    if(N981) begin
      \nz.mem_1527_sv2v_reg  <= data_i[7];
      \nz.mem_1526_sv2v_reg  <= data_i[6];
      \nz.mem_1525_sv2v_reg  <= data_i[5];
      \nz.mem_1524_sv2v_reg  <= data_i[4];
      \nz.mem_1523_sv2v_reg  <= data_i[3];
      \nz.mem_1522_sv2v_reg  <= data_i[2];
      \nz.mem_1521_sv2v_reg  <= data_i[1];
      \nz.mem_1520_sv2v_reg  <= data_i[0];
    end 
    if(N980) begin
      \nz.mem_1519_sv2v_reg  <= data_i[7];
      \nz.mem_1518_sv2v_reg  <= data_i[6];
      \nz.mem_1517_sv2v_reg  <= data_i[5];
      \nz.mem_1516_sv2v_reg  <= data_i[4];
      \nz.mem_1515_sv2v_reg  <= data_i[3];
      \nz.mem_1514_sv2v_reg  <= data_i[2];
      \nz.mem_1513_sv2v_reg  <= data_i[1];
      \nz.mem_1512_sv2v_reg  <= data_i[0];
    end 
    if(N979) begin
      \nz.mem_1511_sv2v_reg  <= data_i[7];
      \nz.mem_1510_sv2v_reg  <= data_i[6];
      \nz.mem_1509_sv2v_reg  <= data_i[5];
      \nz.mem_1508_sv2v_reg  <= data_i[4];
      \nz.mem_1507_sv2v_reg  <= data_i[3];
      \nz.mem_1506_sv2v_reg  <= data_i[2];
      \nz.mem_1505_sv2v_reg  <= data_i[1];
      \nz.mem_1504_sv2v_reg  <= data_i[0];
    end 
    if(N978) begin
      \nz.mem_1503_sv2v_reg  <= data_i[7];
      \nz.mem_1502_sv2v_reg  <= data_i[6];
      \nz.mem_1501_sv2v_reg  <= data_i[5];
      \nz.mem_1500_sv2v_reg  <= data_i[4];
      \nz.mem_1499_sv2v_reg  <= data_i[3];
      \nz.mem_1498_sv2v_reg  <= data_i[2];
      \nz.mem_1497_sv2v_reg  <= data_i[1];
      \nz.mem_1496_sv2v_reg  <= data_i[0];
    end 
    if(N977) begin
      \nz.mem_1495_sv2v_reg  <= data_i[7];
      \nz.mem_1494_sv2v_reg  <= data_i[6];
      \nz.mem_1493_sv2v_reg  <= data_i[5];
      \nz.mem_1492_sv2v_reg  <= data_i[4];
      \nz.mem_1491_sv2v_reg  <= data_i[3];
      \nz.mem_1490_sv2v_reg  <= data_i[2];
      \nz.mem_1489_sv2v_reg  <= data_i[1];
      \nz.mem_1488_sv2v_reg  <= data_i[0];
    end 
    if(N976) begin
      \nz.mem_1487_sv2v_reg  <= data_i[7];
      \nz.mem_1486_sv2v_reg  <= data_i[6];
      \nz.mem_1485_sv2v_reg  <= data_i[5];
      \nz.mem_1484_sv2v_reg  <= data_i[4];
      \nz.mem_1483_sv2v_reg  <= data_i[3];
      \nz.mem_1482_sv2v_reg  <= data_i[2];
      \nz.mem_1481_sv2v_reg  <= data_i[1];
      \nz.mem_1480_sv2v_reg  <= data_i[0];
    end 
    if(N975) begin
      \nz.mem_1479_sv2v_reg  <= data_i[7];
      \nz.mem_1478_sv2v_reg  <= data_i[6];
      \nz.mem_1477_sv2v_reg  <= data_i[5];
      \nz.mem_1476_sv2v_reg  <= data_i[4];
      \nz.mem_1475_sv2v_reg  <= data_i[3];
      \nz.mem_1474_sv2v_reg  <= data_i[2];
      \nz.mem_1473_sv2v_reg  <= data_i[1];
      \nz.mem_1472_sv2v_reg  <= data_i[0];
    end 
    if(N974) begin
      \nz.mem_1471_sv2v_reg  <= data_i[7];
      \nz.mem_1470_sv2v_reg  <= data_i[6];
      \nz.mem_1469_sv2v_reg  <= data_i[5];
      \nz.mem_1468_sv2v_reg  <= data_i[4];
      \nz.mem_1467_sv2v_reg  <= data_i[3];
      \nz.mem_1466_sv2v_reg  <= data_i[2];
      \nz.mem_1465_sv2v_reg  <= data_i[1];
      \nz.mem_1464_sv2v_reg  <= data_i[0];
    end 
    if(N973) begin
      \nz.mem_1463_sv2v_reg  <= data_i[7];
      \nz.mem_1462_sv2v_reg  <= data_i[6];
      \nz.mem_1461_sv2v_reg  <= data_i[5];
      \nz.mem_1460_sv2v_reg  <= data_i[4];
      \nz.mem_1459_sv2v_reg  <= data_i[3];
      \nz.mem_1458_sv2v_reg  <= data_i[2];
      \nz.mem_1457_sv2v_reg  <= data_i[1];
      \nz.mem_1456_sv2v_reg  <= data_i[0];
    end 
    if(N972) begin
      \nz.mem_1455_sv2v_reg  <= data_i[7];
      \nz.mem_1454_sv2v_reg  <= data_i[6];
      \nz.mem_1453_sv2v_reg  <= data_i[5];
      \nz.mem_1452_sv2v_reg  <= data_i[4];
      \nz.mem_1451_sv2v_reg  <= data_i[3];
      \nz.mem_1450_sv2v_reg  <= data_i[2];
      \nz.mem_1449_sv2v_reg  <= data_i[1];
      \nz.mem_1448_sv2v_reg  <= data_i[0];
    end 
    if(N971) begin
      \nz.mem_1447_sv2v_reg  <= data_i[7];
      \nz.mem_1446_sv2v_reg  <= data_i[6];
      \nz.mem_1445_sv2v_reg  <= data_i[5];
      \nz.mem_1444_sv2v_reg  <= data_i[4];
      \nz.mem_1443_sv2v_reg  <= data_i[3];
      \nz.mem_1442_sv2v_reg  <= data_i[2];
      \nz.mem_1441_sv2v_reg  <= data_i[1];
      \nz.mem_1440_sv2v_reg  <= data_i[0];
    end 
    if(N970) begin
      \nz.mem_1439_sv2v_reg  <= data_i[7];
      \nz.mem_1438_sv2v_reg  <= data_i[6];
      \nz.mem_1437_sv2v_reg  <= data_i[5];
      \nz.mem_1436_sv2v_reg  <= data_i[4];
      \nz.mem_1435_sv2v_reg  <= data_i[3];
      \nz.mem_1434_sv2v_reg  <= data_i[2];
      \nz.mem_1433_sv2v_reg  <= data_i[1];
      \nz.mem_1432_sv2v_reg  <= data_i[0];
    end 
    if(N969) begin
      \nz.mem_1431_sv2v_reg  <= data_i[7];
      \nz.mem_1430_sv2v_reg  <= data_i[6];
      \nz.mem_1429_sv2v_reg  <= data_i[5];
      \nz.mem_1428_sv2v_reg  <= data_i[4];
      \nz.mem_1427_sv2v_reg  <= data_i[3];
      \nz.mem_1426_sv2v_reg  <= data_i[2];
      \nz.mem_1425_sv2v_reg  <= data_i[1];
      \nz.mem_1424_sv2v_reg  <= data_i[0];
    end 
    if(N968) begin
      \nz.mem_1423_sv2v_reg  <= data_i[7];
      \nz.mem_1422_sv2v_reg  <= data_i[6];
      \nz.mem_1421_sv2v_reg  <= data_i[5];
      \nz.mem_1420_sv2v_reg  <= data_i[4];
      \nz.mem_1419_sv2v_reg  <= data_i[3];
      \nz.mem_1418_sv2v_reg  <= data_i[2];
      \nz.mem_1417_sv2v_reg  <= data_i[1];
      \nz.mem_1416_sv2v_reg  <= data_i[0];
    end 
    if(N967) begin
      \nz.mem_1415_sv2v_reg  <= data_i[7];
      \nz.mem_1414_sv2v_reg  <= data_i[6];
      \nz.mem_1413_sv2v_reg  <= data_i[5];
      \nz.mem_1412_sv2v_reg  <= data_i[4];
      \nz.mem_1411_sv2v_reg  <= data_i[3];
      \nz.mem_1410_sv2v_reg  <= data_i[2];
      \nz.mem_1409_sv2v_reg  <= data_i[1];
      \nz.mem_1408_sv2v_reg  <= data_i[0];
    end 
    if(N966) begin
      \nz.mem_1407_sv2v_reg  <= data_i[7];
      \nz.mem_1406_sv2v_reg  <= data_i[6];
      \nz.mem_1405_sv2v_reg  <= data_i[5];
      \nz.mem_1404_sv2v_reg  <= data_i[4];
      \nz.mem_1403_sv2v_reg  <= data_i[3];
      \nz.mem_1402_sv2v_reg  <= data_i[2];
      \nz.mem_1401_sv2v_reg  <= data_i[1];
      \nz.mem_1400_sv2v_reg  <= data_i[0];
    end 
    if(N965) begin
      \nz.mem_1399_sv2v_reg  <= data_i[7];
      \nz.mem_1398_sv2v_reg  <= data_i[6];
      \nz.mem_1397_sv2v_reg  <= data_i[5];
      \nz.mem_1396_sv2v_reg  <= data_i[4];
      \nz.mem_1395_sv2v_reg  <= data_i[3];
      \nz.mem_1394_sv2v_reg  <= data_i[2];
      \nz.mem_1393_sv2v_reg  <= data_i[1];
      \nz.mem_1392_sv2v_reg  <= data_i[0];
    end 
    if(N964) begin
      \nz.mem_1391_sv2v_reg  <= data_i[7];
      \nz.mem_1390_sv2v_reg  <= data_i[6];
      \nz.mem_1389_sv2v_reg  <= data_i[5];
      \nz.mem_1388_sv2v_reg  <= data_i[4];
      \nz.mem_1387_sv2v_reg  <= data_i[3];
      \nz.mem_1386_sv2v_reg  <= data_i[2];
      \nz.mem_1385_sv2v_reg  <= data_i[1];
      \nz.mem_1384_sv2v_reg  <= data_i[0];
    end 
    if(N963) begin
      \nz.mem_1383_sv2v_reg  <= data_i[7];
      \nz.mem_1382_sv2v_reg  <= data_i[6];
      \nz.mem_1381_sv2v_reg  <= data_i[5];
      \nz.mem_1380_sv2v_reg  <= data_i[4];
      \nz.mem_1379_sv2v_reg  <= data_i[3];
      \nz.mem_1378_sv2v_reg  <= data_i[2];
      \nz.mem_1377_sv2v_reg  <= data_i[1];
      \nz.mem_1376_sv2v_reg  <= data_i[0];
    end 
    if(N962) begin
      \nz.mem_1375_sv2v_reg  <= data_i[7];
      \nz.mem_1374_sv2v_reg  <= data_i[6];
      \nz.mem_1373_sv2v_reg  <= data_i[5];
      \nz.mem_1372_sv2v_reg  <= data_i[4];
      \nz.mem_1371_sv2v_reg  <= data_i[3];
      \nz.mem_1370_sv2v_reg  <= data_i[2];
      \nz.mem_1369_sv2v_reg  <= data_i[1];
      \nz.mem_1368_sv2v_reg  <= data_i[0];
    end 
    if(N961) begin
      \nz.mem_1367_sv2v_reg  <= data_i[7];
      \nz.mem_1366_sv2v_reg  <= data_i[6];
      \nz.mem_1365_sv2v_reg  <= data_i[5];
      \nz.mem_1364_sv2v_reg  <= data_i[4];
      \nz.mem_1363_sv2v_reg  <= data_i[3];
      \nz.mem_1362_sv2v_reg  <= data_i[2];
      \nz.mem_1361_sv2v_reg  <= data_i[1];
      \nz.mem_1360_sv2v_reg  <= data_i[0];
    end 
    if(N960) begin
      \nz.mem_1359_sv2v_reg  <= data_i[7];
      \nz.mem_1358_sv2v_reg  <= data_i[6];
      \nz.mem_1357_sv2v_reg  <= data_i[5];
      \nz.mem_1356_sv2v_reg  <= data_i[4];
      \nz.mem_1355_sv2v_reg  <= data_i[3];
      \nz.mem_1354_sv2v_reg  <= data_i[2];
      \nz.mem_1353_sv2v_reg  <= data_i[1];
      \nz.mem_1352_sv2v_reg  <= data_i[0];
    end 
    if(N959) begin
      \nz.mem_1351_sv2v_reg  <= data_i[7];
      \nz.mem_1350_sv2v_reg  <= data_i[6];
      \nz.mem_1349_sv2v_reg  <= data_i[5];
      \nz.mem_1348_sv2v_reg  <= data_i[4];
      \nz.mem_1347_sv2v_reg  <= data_i[3];
      \nz.mem_1346_sv2v_reg  <= data_i[2];
      \nz.mem_1345_sv2v_reg  <= data_i[1];
      \nz.mem_1344_sv2v_reg  <= data_i[0];
    end 
    if(N958) begin
      \nz.mem_1343_sv2v_reg  <= data_i[7];
      \nz.mem_1342_sv2v_reg  <= data_i[6];
      \nz.mem_1341_sv2v_reg  <= data_i[5];
      \nz.mem_1340_sv2v_reg  <= data_i[4];
      \nz.mem_1339_sv2v_reg  <= data_i[3];
      \nz.mem_1338_sv2v_reg  <= data_i[2];
      \nz.mem_1337_sv2v_reg  <= data_i[1];
      \nz.mem_1336_sv2v_reg  <= data_i[0];
    end 
    if(N957) begin
      \nz.mem_1335_sv2v_reg  <= data_i[7];
      \nz.mem_1334_sv2v_reg  <= data_i[6];
      \nz.mem_1333_sv2v_reg  <= data_i[5];
      \nz.mem_1332_sv2v_reg  <= data_i[4];
      \nz.mem_1331_sv2v_reg  <= data_i[3];
      \nz.mem_1330_sv2v_reg  <= data_i[2];
      \nz.mem_1329_sv2v_reg  <= data_i[1];
      \nz.mem_1328_sv2v_reg  <= data_i[0];
    end 
    if(N956) begin
      \nz.mem_1327_sv2v_reg  <= data_i[7];
      \nz.mem_1326_sv2v_reg  <= data_i[6];
      \nz.mem_1325_sv2v_reg  <= data_i[5];
      \nz.mem_1324_sv2v_reg  <= data_i[4];
      \nz.mem_1323_sv2v_reg  <= data_i[3];
      \nz.mem_1322_sv2v_reg  <= data_i[2];
      \nz.mem_1321_sv2v_reg  <= data_i[1];
      \nz.mem_1320_sv2v_reg  <= data_i[0];
    end 
    if(N955) begin
      \nz.mem_1319_sv2v_reg  <= data_i[7];
      \nz.mem_1318_sv2v_reg  <= data_i[6];
      \nz.mem_1317_sv2v_reg  <= data_i[5];
      \nz.mem_1316_sv2v_reg  <= data_i[4];
      \nz.mem_1315_sv2v_reg  <= data_i[3];
      \nz.mem_1314_sv2v_reg  <= data_i[2];
      \nz.mem_1313_sv2v_reg  <= data_i[1];
      \nz.mem_1312_sv2v_reg  <= data_i[0];
    end 
    if(N954) begin
      \nz.mem_1311_sv2v_reg  <= data_i[7];
      \nz.mem_1310_sv2v_reg  <= data_i[6];
      \nz.mem_1309_sv2v_reg  <= data_i[5];
      \nz.mem_1308_sv2v_reg  <= data_i[4];
      \nz.mem_1307_sv2v_reg  <= data_i[3];
      \nz.mem_1306_sv2v_reg  <= data_i[2];
      \nz.mem_1305_sv2v_reg  <= data_i[1];
      \nz.mem_1304_sv2v_reg  <= data_i[0];
    end 
    if(N953) begin
      \nz.mem_1303_sv2v_reg  <= data_i[7];
      \nz.mem_1302_sv2v_reg  <= data_i[6];
      \nz.mem_1301_sv2v_reg  <= data_i[5];
      \nz.mem_1300_sv2v_reg  <= data_i[4];
      \nz.mem_1299_sv2v_reg  <= data_i[3];
      \nz.mem_1298_sv2v_reg  <= data_i[2];
      \nz.mem_1297_sv2v_reg  <= data_i[1];
      \nz.mem_1296_sv2v_reg  <= data_i[0];
    end 
    if(N952) begin
      \nz.mem_1295_sv2v_reg  <= data_i[7];
      \nz.mem_1294_sv2v_reg  <= data_i[6];
      \nz.mem_1293_sv2v_reg  <= data_i[5];
      \nz.mem_1292_sv2v_reg  <= data_i[4];
      \nz.mem_1291_sv2v_reg  <= data_i[3];
      \nz.mem_1290_sv2v_reg  <= data_i[2];
      \nz.mem_1289_sv2v_reg  <= data_i[1];
      \nz.mem_1288_sv2v_reg  <= data_i[0];
    end 
    if(N951) begin
      \nz.mem_1287_sv2v_reg  <= data_i[7];
      \nz.mem_1286_sv2v_reg  <= data_i[6];
      \nz.mem_1285_sv2v_reg  <= data_i[5];
      \nz.mem_1284_sv2v_reg  <= data_i[4];
      \nz.mem_1283_sv2v_reg  <= data_i[3];
      \nz.mem_1282_sv2v_reg  <= data_i[2];
      \nz.mem_1281_sv2v_reg  <= data_i[1];
      \nz.mem_1280_sv2v_reg  <= data_i[0];
    end 
    if(N950) begin
      \nz.mem_1279_sv2v_reg  <= data_i[7];
      \nz.mem_1278_sv2v_reg  <= data_i[6];
      \nz.mem_1277_sv2v_reg  <= data_i[5];
      \nz.mem_1276_sv2v_reg  <= data_i[4];
      \nz.mem_1275_sv2v_reg  <= data_i[3];
      \nz.mem_1274_sv2v_reg  <= data_i[2];
      \nz.mem_1273_sv2v_reg  <= data_i[1];
      \nz.mem_1272_sv2v_reg  <= data_i[0];
    end 
    if(N949) begin
      \nz.mem_1271_sv2v_reg  <= data_i[7];
      \nz.mem_1270_sv2v_reg  <= data_i[6];
      \nz.mem_1269_sv2v_reg  <= data_i[5];
      \nz.mem_1268_sv2v_reg  <= data_i[4];
      \nz.mem_1267_sv2v_reg  <= data_i[3];
      \nz.mem_1266_sv2v_reg  <= data_i[2];
      \nz.mem_1265_sv2v_reg  <= data_i[1];
      \nz.mem_1264_sv2v_reg  <= data_i[0];
    end 
    if(N948) begin
      \nz.mem_1263_sv2v_reg  <= data_i[7];
      \nz.mem_1262_sv2v_reg  <= data_i[6];
      \nz.mem_1261_sv2v_reg  <= data_i[5];
      \nz.mem_1260_sv2v_reg  <= data_i[4];
      \nz.mem_1259_sv2v_reg  <= data_i[3];
      \nz.mem_1258_sv2v_reg  <= data_i[2];
      \nz.mem_1257_sv2v_reg  <= data_i[1];
      \nz.mem_1256_sv2v_reg  <= data_i[0];
    end 
    if(N947) begin
      \nz.mem_1255_sv2v_reg  <= data_i[7];
      \nz.mem_1254_sv2v_reg  <= data_i[6];
      \nz.mem_1253_sv2v_reg  <= data_i[5];
      \nz.mem_1252_sv2v_reg  <= data_i[4];
      \nz.mem_1251_sv2v_reg  <= data_i[3];
      \nz.mem_1250_sv2v_reg  <= data_i[2];
      \nz.mem_1249_sv2v_reg  <= data_i[1];
      \nz.mem_1248_sv2v_reg  <= data_i[0];
    end 
    if(N946) begin
      \nz.mem_1247_sv2v_reg  <= data_i[7];
      \nz.mem_1246_sv2v_reg  <= data_i[6];
      \nz.mem_1245_sv2v_reg  <= data_i[5];
      \nz.mem_1244_sv2v_reg  <= data_i[4];
      \nz.mem_1243_sv2v_reg  <= data_i[3];
      \nz.mem_1242_sv2v_reg  <= data_i[2];
      \nz.mem_1241_sv2v_reg  <= data_i[1];
      \nz.mem_1240_sv2v_reg  <= data_i[0];
    end 
    if(N945) begin
      \nz.mem_1239_sv2v_reg  <= data_i[7];
      \nz.mem_1238_sv2v_reg  <= data_i[6];
      \nz.mem_1237_sv2v_reg  <= data_i[5];
      \nz.mem_1236_sv2v_reg  <= data_i[4];
      \nz.mem_1235_sv2v_reg  <= data_i[3];
      \nz.mem_1234_sv2v_reg  <= data_i[2];
      \nz.mem_1233_sv2v_reg  <= data_i[1];
      \nz.mem_1232_sv2v_reg  <= data_i[0];
    end 
    if(N944) begin
      \nz.mem_1231_sv2v_reg  <= data_i[7];
      \nz.mem_1230_sv2v_reg  <= data_i[6];
      \nz.mem_1229_sv2v_reg  <= data_i[5];
      \nz.mem_1228_sv2v_reg  <= data_i[4];
      \nz.mem_1227_sv2v_reg  <= data_i[3];
      \nz.mem_1226_sv2v_reg  <= data_i[2];
      \nz.mem_1225_sv2v_reg  <= data_i[1];
      \nz.mem_1224_sv2v_reg  <= data_i[0];
    end 
    if(N943) begin
      \nz.mem_1223_sv2v_reg  <= data_i[7];
      \nz.mem_1222_sv2v_reg  <= data_i[6];
      \nz.mem_1221_sv2v_reg  <= data_i[5];
      \nz.mem_1220_sv2v_reg  <= data_i[4];
      \nz.mem_1219_sv2v_reg  <= data_i[3];
      \nz.mem_1218_sv2v_reg  <= data_i[2];
      \nz.mem_1217_sv2v_reg  <= data_i[1];
      \nz.mem_1216_sv2v_reg  <= data_i[0];
    end 
    if(N942) begin
      \nz.mem_1215_sv2v_reg  <= data_i[7];
      \nz.mem_1214_sv2v_reg  <= data_i[6];
      \nz.mem_1213_sv2v_reg  <= data_i[5];
      \nz.mem_1212_sv2v_reg  <= data_i[4];
      \nz.mem_1211_sv2v_reg  <= data_i[3];
      \nz.mem_1210_sv2v_reg  <= data_i[2];
      \nz.mem_1209_sv2v_reg  <= data_i[1];
      \nz.mem_1208_sv2v_reg  <= data_i[0];
    end 
    if(N941) begin
      \nz.mem_1207_sv2v_reg  <= data_i[7];
      \nz.mem_1206_sv2v_reg  <= data_i[6];
      \nz.mem_1205_sv2v_reg  <= data_i[5];
      \nz.mem_1204_sv2v_reg  <= data_i[4];
      \nz.mem_1203_sv2v_reg  <= data_i[3];
      \nz.mem_1202_sv2v_reg  <= data_i[2];
      \nz.mem_1201_sv2v_reg  <= data_i[1];
      \nz.mem_1200_sv2v_reg  <= data_i[0];
    end 
    if(N940) begin
      \nz.mem_1199_sv2v_reg  <= data_i[7];
      \nz.mem_1198_sv2v_reg  <= data_i[6];
      \nz.mem_1197_sv2v_reg  <= data_i[5];
      \nz.mem_1196_sv2v_reg  <= data_i[4];
      \nz.mem_1195_sv2v_reg  <= data_i[3];
      \nz.mem_1194_sv2v_reg  <= data_i[2];
      \nz.mem_1193_sv2v_reg  <= data_i[1];
      \nz.mem_1192_sv2v_reg  <= data_i[0];
    end 
    if(N939) begin
      \nz.mem_1191_sv2v_reg  <= data_i[7];
      \nz.mem_1190_sv2v_reg  <= data_i[6];
      \nz.mem_1189_sv2v_reg  <= data_i[5];
      \nz.mem_1188_sv2v_reg  <= data_i[4];
      \nz.mem_1187_sv2v_reg  <= data_i[3];
      \nz.mem_1186_sv2v_reg  <= data_i[2];
      \nz.mem_1185_sv2v_reg  <= data_i[1];
      \nz.mem_1184_sv2v_reg  <= data_i[0];
    end 
    if(N938) begin
      \nz.mem_1183_sv2v_reg  <= data_i[7];
      \nz.mem_1182_sv2v_reg  <= data_i[6];
      \nz.mem_1181_sv2v_reg  <= data_i[5];
      \nz.mem_1180_sv2v_reg  <= data_i[4];
      \nz.mem_1179_sv2v_reg  <= data_i[3];
      \nz.mem_1178_sv2v_reg  <= data_i[2];
      \nz.mem_1177_sv2v_reg  <= data_i[1];
      \nz.mem_1176_sv2v_reg  <= data_i[0];
    end 
    if(N937) begin
      \nz.mem_1175_sv2v_reg  <= data_i[7];
      \nz.mem_1174_sv2v_reg  <= data_i[6];
      \nz.mem_1173_sv2v_reg  <= data_i[5];
      \nz.mem_1172_sv2v_reg  <= data_i[4];
      \nz.mem_1171_sv2v_reg  <= data_i[3];
      \nz.mem_1170_sv2v_reg  <= data_i[2];
      \nz.mem_1169_sv2v_reg  <= data_i[1];
      \nz.mem_1168_sv2v_reg  <= data_i[0];
    end 
    if(N936) begin
      \nz.mem_1167_sv2v_reg  <= data_i[7];
      \nz.mem_1166_sv2v_reg  <= data_i[6];
      \nz.mem_1165_sv2v_reg  <= data_i[5];
      \nz.mem_1164_sv2v_reg  <= data_i[4];
      \nz.mem_1163_sv2v_reg  <= data_i[3];
      \nz.mem_1162_sv2v_reg  <= data_i[2];
      \nz.mem_1161_sv2v_reg  <= data_i[1];
      \nz.mem_1160_sv2v_reg  <= data_i[0];
    end 
    if(N935) begin
      \nz.mem_1159_sv2v_reg  <= data_i[7];
      \nz.mem_1158_sv2v_reg  <= data_i[6];
      \nz.mem_1157_sv2v_reg  <= data_i[5];
      \nz.mem_1156_sv2v_reg  <= data_i[4];
      \nz.mem_1155_sv2v_reg  <= data_i[3];
      \nz.mem_1154_sv2v_reg  <= data_i[2];
      \nz.mem_1153_sv2v_reg  <= data_i[1];
      \nz.mem_1152_sv2v_reg  <= data_i[0];
    end 
    if(N934) begin
      \nz.mem_1151_sv2v_reg  <= data_i[7];
      \nz.mem_1150_sv2v_reg  <= data_i[6];
      \nz.mem_1149_sv2v_reg  <= data_i[5];
      \nz.mem_1148_sv2v_reg  <= data_i[4];
      \nz.mem_1147_sv2v_reg  <= data_i[3];
      \nz.mem_1146_sv2v_reg  <= data_i[2];
      \nz.mem_1145_sv2v_reg  <= data_i[1];
      \nz.mem_1144_sv2v_reg  <= data_i[0];
    end 
    if(N933) begin
      \nz.mem_1143_sv2v_reg  <= data_i[7];
      \nz.mem_1142_sv2v_reg  <= data_i[6];
      \nz.mem_1141_sv2v_reg  <= data_i[5];
      \nz.mem_1140_sv2v_reg  <= data_i[4];
      \nz.mem_1139_sv2v_reg  <= data_i[3];
      \nz.mem_1138_sv2v_reg  <= data_i[2];
      \nz.mem_1137_sv2v_reg  <= data_i[1];
      \nz.mem_1136_sv2v_reg  <= data_i[0];
    end 
    if(N932) begin
      \nz.mem_1135_sv2v_reg  <= data_i[7];
      \nz.mem_1134_sv2v_reg  <= data_i[6];
      \nz.mem_1133_sv2v_reg  <= data_i[5];
      \nz.mem_1132_sv2v_reg  <= data_i[4];
      \nz.mem_1131_sv2v_reg  <= data_i[3];
      \nz.mem_1130_sv2v_reg  <= data_i[2];
      \nz.mem_1129_sv2v_reg  <= data_i[1];
      \nz.mem_1128_sv2v_reg  <= data_i[0];
    end 
    if(N931) begin
      \nz.mem_1127_sv2v_reg  <= data_i[7];
      \nz.mem_1126_sv2v_reg  <= data_i[6];
      \nz.mem_1125_sv2v_reg  <= data_i[5];
      \nz.mem_1124_sv2v_reg  <= data_i[4];
      \nz.mem_1123_sv2v_reg  <= data_i[3];
      \nz.mem_1122_sv2v_reg  <= data_i[2];
      \nz.mem_1121_sv2v_reg  <= data_i[1];
      \nz.mem_1120_sv2v_reg  <= data_i[0];
    end 
    if(N930) begin
      \nz.mem_1119_sv2v_reg  <= data_i[7];
      \nz.mem_1118_sv2v_reg  <= data_i[6];
      \nz.mem_1117_sv2v_reg  <= data_i[5];
      \nz.mem_1116_sv2v_reg  <= data_i[4];
      \nz.mem_1115_sv2v_reg  <= data_i[3];
      \nz.mem_1114_sv2v_reg  <= data_i[2];
      \nz.mem_1113_sv2v_reg  <= data_i[1];
      \nz.mem_1112_sv2v_reg  <= data_i[0];
    end 
    if(N929) begin
      \nz.mem_1111_sv2v_reg  <= data_i[7];
      \nz.mem_1110_sv2v_reg  <= data_i[6];
      \nz.mem_1109_sv2v_reg  <= data_i[5];
      \nz.mem_1108_sv2v_reg  <= data_i[4];
      \nz.mem_1107_sv2v_reg  <= data_i[3];
      \nz.mem_1106_sv2v_reg  <= data_i[2];
      \nz.mem_1105_sv2v_reg  <= data_i[1];
      \nz.mem_1104_sv2v_reg  <= data_i[0];
    end 
    if(N928) begin
      \nz.mem_1103_sv2v_reg  <= data_i[7];
      \nz.mem_1102_sv2v_reg  <= data_i[6];
      \nz.mem_1101_sv2v_reg  <= data_i[5];
      \nz.mem_1100_sv2v_reg  <= data_i[4];
      \nz.mem_1099_sv2v_reg  <= data_i[3];
      \nz.mem_1098_sv2v_reg  <= data_i[2];
      \nz.mem_1097_sv2v_reg  <= data_i[1];
      \nz.mem_1096_sv2v_reg  <= data_i[0];
    end 
    if(N927) begin
      \nz.mem_1095_sv2v_reg  <= data_i[7];
      \nz.mem_1094_sv2v_reg  <= data_i[6];
      \nz.mem_1093_sv2v_reg  <= data_i[5];
      \nz.mem_1092_sv2v_reg  <= data_i[4];
      \nz.mem_1091_sv2v_reg  <= data_i[3];
      \nz.mem_1090_sv2v_reg  <= data_i[2];
      \nz.mem_1089_sv2v_reg  <= data_i[1];
      \nz.mem_1088_sv2v_reg  <= data_i[0];
    end 
    if(N926) begin
      \nz.mem_1087_sv2v_reg  <= data_i[7];
      \nz.mem_1086_sv2v_reg  <= data_i[6];
      \nz.mem_1085_sv2v_reg  <= data_i[5];
      \nz.mem_1084_sv2v_reg  <= data_i[4];
      \nz.mem_1083_sv2v_reg  <= data_i[3];
      \nz.mem_1082_sv2v_reg  <= data_i[2];
      \nz.mem_1081_sv2v_reg  <= data_i[1];
      \nz.mem_1080_sv2v_reg  <= data_i[0];
    end 
    if(N925) begin
      \nz.mem_1079_sv2v_reg  <= data_i[7];
      \nz.mem_1078_sv2v_reg  <= data_i[6];
      \nz.mem_1077_sv2v_reg  <= data_i[5];
      \nz.mem_1076_sv2v_reg  <= data_i[4];
      \nz.mem_1075_sv2v_reg  <= data_i[3];
      \nz.mem_1074_sv2v_reg  <= data_i[2];
      \nz.mem_1073_sv2v_reg  <= data_i[1];
      \nz.mem_1072_sv2v_reg  <= data_i[0];
    end 
    if(N924) begin
      \nz.mem_1071_sv2v_reg  <= data_i[7];
      \nz.mem_1070_sv2v_reg  <= data_i[6];
      \nz.mem_1069_sv2v_reg  <= data_i[5];
      \nz.mem_1068_sv2v_reg  <= data_i[4];
      \nz.mem_1067_sv2v_reg  <= data_i[3];
      \nz.mem_1066_sv2v_reg  <= data_i[2];
      \nz.mem_1065_sv2v_reg  <= data_i[1];
      \nz.mem_1064_sv2v_reg  <= data_i[0];
    end 
    if(N923) begin
      \nz.mem_1063_sv2v_reg  <= data_i[7];
      \nz.mem_1062_sv2v_reg  <= data_i[6];
      \nz.mem_1061_sv2v_reg  <= data_i[5];
      \nz.mem_1060_sv2v_reg  <= data_i[4];
      \nz.mem_1059_sv2v_reg  <= data_i[3];
      \nz.mem_1058_sv2v_reg  <= data_i[2];
      \nz.mem_1057_sv2v_reg  <= data_i[1];
      \nz.mem_1056_sv2v_reg  <= data_i[0];
    end 
    if(N922) begin
      \nz.mem_1055_sv2v_reg  <= data_i[7];
      \nz.mem_1054_sv2v_reg  <= data_i[6];
      \nz.mem_1053_sv2v_reg  <= data_i[5];
      \nz.mem_1052_sv2v_reg  <= data_i[4];
      \nz.mem_1051_sv2v_reg  <= data_i[3];
      \nz.mem_1050_sv2v_reg  <= data_i[2];
      \nz.mem_1049_sv2v_reg  <= data_i[1];
      \nz.mem_1048_sv2v_reg  <= data_i[0];
    end 
    if(N921) begin
      \nz.mem_1047_sv2v_reg  <= data_i[7];
      \nz.mem_1046_sv2v_reg  <= data_i[6];
      \nz.mem_1045_sv2v_reg  <= data_i[5];
      \nz.mem_1044_sv2v_reg  <= data_i[4];
      \nz.mem_1043_sv2v_reg  <= data_i[3];
      \nz.mem_1042_sv2v_reg  <= data_i[2];
      \nz.mem_1041_sv2v_reg  <= data_i[1];
      \nz.mem_1040_sv2v_reg  <= data_i[0];
    end 
    if(N920) begin
      \nz.mem_1039_sv2v_reg  <= data_i[7];
      \nz.mem_1038_sv2v_reg  <= data_i[6];
      \nz.mem_1037_sv2v_reg  <= data_i[5];
      \nz.mem_1036_sv2v_reg  <= data_i[4];
      \nz.mem_1035_sv2v_reg  <= data_i[3];
      \nz.mem_1034_sv2v_reg  <= data_i[2];
      \nz.mem_1033_sv2v_reg  <= data_i[1];
      \nz.mem_1032_sv2v_reg  <= data_i[0];
    end 
    if(N919) begin
      \nz.mem_1031_sv2v_reg  <= data_i[7];
      \nz.mem_1030_sv2v_reg  <= data_i[6];
      \nz.mem_1029_sv2v_reg  <= data_i[5];
      \nz.mem_1028_sv2v_reg  <= data_i[4];
      \nz.mem_1027_sv2v_reg  <= data_i[3];
      \nz.mem_1026_sv2v_reg  <= data_i[2];
      \nz.mem_1025_sv2v_reg  <= data_i[1];
      \nz.mem_1024_sv2v_reg  <= data_i[0];
    end 
    if(N918) begin
      \nz.mem_1023_sv2v_reg  <= data_i[7];
      \nz.mem_1022_sv2v_reg  <= data_i[6];
      \nz.mem_1021_sv2v_reg  <= data_i[5];
      \nz.mem_1020_sv2v_reg  <= data_i[4];
      \nz.mem_1019_sv2v_reg  <= data_i[3];
      \nz.mem_1018_sv2v_reg  <= data_i[2];
      \nz.mem_1017_sv2v_reg  <= data_i[1];
      \nz.mem_1016_sv2v_reg  <= data_i[0];
    end 
    if(N917) begin
      \nz.mem_1015_sv2v_reg  <= data_i[7];
      \nz.mem_1014_sv2v_reg  <= data_i[6];
      \nz.mem_1013_sv2v_reg  <= data_i[5];
      \nz.mem_1012_sv2v_reg  <= data_i[4];
      \nz.mem_1011_sv2v_reg  <= data_i[3];
      \nz.mem_1010_sv2v_reg  <= data_i[2];
      \nz.mem_1009_sv2v_reg  <= data_i[1];
      \nz.mem_1008_sv2v_reg  <= data_i[0];
    end 
    if(N916) begin
      \nz.mem_1007_sv2v_reg  <= data_i[7];
      \nz.mem_1006_sv2v_reg  <= data_i[6];
      \nz.mem_1005_sv2v_reg  <= data_i[5];
      \nz.mem_1004_sv2v_reg  <= data_i[4];
      \nz.mem_1003_sv2v_reg  <= data_i[3];
      \nz.mem_1002_sv2v_reg  <= data_i[2];
      \nz.mem_1001_sv2v_reg  <= data_i[1];
      \nz.mem_1000_sv2v_reg  <= data_i[0];
    end 
    if(N915) begin
      \nz.mem_999_sv2v_reg  <= data_i[7];
      \nz.mem_998_sv2v_reg  <= data_i[6];
      \nz.mem_997_sv2v_reg  <= data_i[5];
      \nz.mem_996_sv2v_reg  <= data_i[4];
      \nz.mem_995_sv2v_reg  <= data_i[3];
      \nz.mem_994_sv2v_reg  <= data_i[2];
      \nz.mem_993_sv2v_reg  <= data_i[1];
      \nz.mem_992_sv2v_reg  <= data_i[0];
    end 
    if(N914) begin
      \nz.mem_991_sv2v_reg  <= data_i[7];
      \nz.mem_990_sv2v_reg  <= data_i[6];
      \nz.mem_989_sv2v_reg  <= data_i[5];
      \nz.mem_988_sv2v_reg  <= data_i[4];
      \nz.mem_987_sv2v_reg  <= data_i[3];
      \nz.mem_986_sv2v_reg  <= data_i[2];
      \nz.mem_985_sv2v_reg  <= data_i[1];
      \nz.mem_984_sv2v_reg  <= data_i[0];
    end 
    if(N913) begin
      \nz.mem_983_sv2v_reg  <= data_i[7];
      \nz.mem_982_sv2v_reg  <= data_i[6];
      \nz.mem_981_sv2v_reg  <= data_i[5];
      \nz.mem_980_sv2v_reg  <= data_i[4];
      \nz.mem_979_sv2v_reg  <= data_i[3];
      \nz.mem_978_sv2v_reg  <= data_i[2];
      \nz.mem_977_sv2v_reg  <= data_i[1];
      \nz.mem_976_sv2v_reg  <= data_i[0];
    end 
    if(N912) begin
      \nz.mem_975_sv2v_reg  <= data_i[7];
      \nz.mem_974_sv2v_reg  <= data_i[6];
      \nz.mem_973_sv2v_reg  <= data_i[5];
      \nz.mem_972_sv2v_reg  <= data_i[4];
      \nz.mem_971_sv2v_reg  <= data_i[3];
      \nz.mem_970_sv2v_reg  <= data_i[2];
      \nz.mem_969_sv2v_reg  <= data_i[1];
      \nz.mem_968_sv2v_reg  <= data_i[0];
    end 
    if(N911) begin
      \nz.mem_967_sv2v_reg  <= data_i[7];
      \nz.mem_966_sv2v_reg  <= data_i[6];
      \nz.mem_965_sv2v_reg  <= data_i[5];
      \nz.mem_964_sv2v_reg  <= data_i[4];
      \nz.mem_963_sv2v_reg  <= data_i[3];
      \nz.mem_962_sv2v_reg  <= data_i[2];
      \nz.mem_961_sv2v_reg  <= data_i[1];
      \nz.mem_960_sv2v_reg  <= data_i[0];
    end 
    if(N910) begin
      \nz.mem_959_sv2v_reg  <= data_i[7];
      \nz.mem_958_sv2v_reg  <= data_i[6];
      \nz.mem_957_sv2v_reg  <= data_i[5];
      \nz.mem_956_sv2v_reg  <= data_i[4];
      \nz.mem_955_sv2v_reg  <= data_i[3];
      \nz.mem_954_sv2v_reg  <= data_i[2];
      \nz.mem_953_sv2v_reg  <= data_i[1];
      \nz.mem_952_sv2v_reg  <= data_i[0];
    end 
    if(N909) begin
      \nz.mem_951_sv2v_reg  <= data_i[7];
      \nz.mem_950_sv2v_reg  <= data_i[6];
      \nz.mem_949_sv2v_reg  <= data_i[5];
      \nz.mem_948_sv2v_reg  <= data_i[4];
      \nz.mem_947_sv2v_reg  <= data_i[3];
      \nz.mem_946_sv2v_reg  <= data_i[2];
      \nz.mem_945_sv2v_reg  <= data_i[1];
      \nz.mem_944_sv2v_reg  <= data_i[0];
    end 
    if(N908) begin
      \nz.mem_943_sv2v_reg  <= data_i[7];
      \nz.mem_942_sv2v_reg  <= data_i[6];
      \nz.mem_941_sv2v_reg  <= data_i[5];
      \nz.mem_940_sv2v_reg  <= data_i[4];
      \nz.mem_939_sv2v_reg  <= data_i[3];
      \nz.mem_938_sv2v_reg  <= data_i[2];
      \nz.mem_937_sv2v_reg  <= data_i[1];
      \nz.mem_936_sv2v_reg  <= data_i[0];
    end 
    if(N907) begin
      \nz.mem_935_sv2v_reg  <= data_i[7];
      \nz.mem_934_sv2v_reg  <= data_i[6];
      \nz.mem_933_sv2v_reg  <= data_i[5];
      \nz.mem_932_sv2v_reg  <= data_i[4];
      \nz.mem_931_sv2v_reg  <= data_i[3];
      \nz.mem_930_sv2v_reg  <= data_i[2];
      \nz.mem_929_sv2v_reg  <= data_i[1];
      \nz.mem_928_sv2v_reg  <= data_i[0];
    end 
    if(N906) begin
      \nz.mem_927_sv2v_reg  <= data_i[7];
      \nz.mem_926_sv2v_reg  <= data_i[6];
      \nz.mem_925_sv2v_reg  <= data_i[5];
      \nz.mem_924_sv2v_reg  <= data_i[4];
      \nz.mem_923_sv2v_reg  <= data_i[3];
      \nz.mem_922_sv2v_reg  <= data_i[2];
      \nz.mem_921_sv2v_reg  <= data_i[1];
      \nz.mem_920_sv2v_reg  <= data_i[0];
    end 
    if(N905) begin
      \nz.mem_919_sv2v_reg  <= data_i[7];
      \nz.mem_918_sv2v_reg  <= data_i[6];
      \nz.mem_917_sv2v_reg  <= data_i[5];
      \nz.mem_916_sv2v_reg  <= data_i[4];
      \nz.mem_915_sv2v_reg  <= data_i[3];
      \nz.mem_914_sv2v_reg  <= data_i[2];
      \nz.mem_913_sv2v_reg  <= data_i[1];
      \nz.mem_912_sv2v_reg  <= data_i[0];
    end 
    if(N904) begin
      \nz.mem_911_sv2v_reg  <= data_i[7];
      \nz.mem_910_sv2v_reg  <= data_i[6];
      \nz.mem_909_sv2v_reg  <= data_i[5];
      \nz.mem_908_sv2v_reg  <= data_i[4];
      \nz.mem_907_sv2v_reg  <= data_i[3];
      \nz.mem_906_sv2v_reg  <= data_i[2];
      \nz.mem_905_sv2v_reg  <= data_i[1];
      \nz.mem_904_sv2v_reg  <= data_i[0];
    end 
    if(N903) begin
      \nz.mem_903_sv2v_reg  <= data_i[7];
      \nz.mem_902_sv2v_reg  <= data_i[6];
      \nz.mem_901_sv2v_reg  <= data_i[5];
      \nz.mem_900_sv2v_reg  <= data_i[4];
      \nz.mem_899_sv2v_reg  <= data_i[3];
      \nz.mem_898_sv2v_reg  <= data_i[2];
      \nz.mem_897_sv2v_reg  <= data_i[1];
      \nz.mem_896_sv2v_reg  <= data_i[0];
    end 
    if(N902) begin
      \nz.mem_895_sv2v_reg  <= data_i[7];
      \nz.mem_894_sv2v_reg  <= data_i[6];
      \nz.mem_893_sv2v_reg  <= data_i[5];
      \nz.mem_892_sv2v_reg  <= data_i[4];
      \nz.mem_891_sv2v_reg  <= data_i[3];
      \nz.mem_890_sv2v_reg  <= data_i[2];
      \nz.mem_889_sv2v_reg  <= data_i[1];
      \nz.mem_888_sv2v_reg  <= data_i[0];
    end 
    if(N901) begin
      \nz.mem_887_sv2v_reg  <= data_i[7];
      \nz.mem_886_sv2v_reg  <= data_i[6];
      \nz.mem_885_sv2v_reg  <= data_i[5];
      \nz.mem_884_sv2v_reg  <= data_i[4];
      \nz.mem_883_sv2v_reg  <= data_i[3];
      \nz.mem_882_sv2v_reg  <= data_i[2];
      \nz.mem_881_sv2v_reg  <= data_i[1];
      \nz.mem_880_sv2v_reg  <= data_i[0];
    end 
    if(N900) begin
      \nz.mem_879_sv2v_reg  <= data_i[7];
      \nz.mem_878_sv2v_reg  <= data_i[6];
      \nz.mem_877_sv2v_reg  <= data_i[5];
      \nz.mem_876_sv2v_reg  <= data_i[4];
      \nz.mem_875_sv2v_reg  <= data_i[3];
      \nz.mem_874_sv2v_reg  <= data_i[2];
      \nz.mem_873_sv2v_reg  <= data_i[1];
      \nz.mem_872_sv2v_reg  <= data_i[0];
    end 
    if(N899) begin
      \nz.mem_871_sv2v_reg  <= data_i[7];
      \nz.mem_870_sv2v_reg  <= data_i[6];
      \nz.mem_869_sv2v_reg  <= data_i[5];
      \nz.mem_868_sv2v_reg  <= data_i[4];
      \nz.mem_867_sv2v_reg  <= data_i[3];
      \nz.mem_866_sv2v_reg  <= data_i[2];
      \nz.mem_865_sv2v_reg  <= data_i[1];
      \nz.mem_864_sv2v_reg  <= data_i[0];
    end 
    if(N898) begin
      \nz.mem_863_sv2v_reg  <= data_i[7];
      \nz.mem_862_sv2v_reg  <= data_i[6];
      \nz.mem_861_sv2v_reg  <= data_i[5];
      \nz.mem_860_sv2v_reg  <= data_i[4];
      \nz.mem_859_sv2v_reg  <= data_i[3];
      \nz.mem_858_sv2v_reg  <= data_i[2];
      \nz.mem_857_sv2v_reg  <= data_i[1];
      \nz.mem_856_sv2v_reg  <= data_i[0];
    end 
    if(N897) begin
      \nz.mem_855_sv2v_reg  <= data_i[7];
      \nz.mem_854_sv2v_reg  <= data_i[6];
      \nz.mem_853_sv2v_reg  <= data_i[5];
      \nz.mem_852_sv2v_reg  <= data_i[4];
      \nz.mem_851_sv2v_reg  <= data_i[3];
      \nz.mem_850_sv2v_reg  <= data_i[2];
      \nz.mem_849_sv2v_reg  <= data_i[1];
      \nz.mem_848_sv2v_reg  <= data_i[0];
    end 
    if(N896) begin
      \nz.mem_847_sv2v_reg  <= data_i[7];
      \nz.mem_846_sv2v_reg  <= data_i[6];
      \nz.mem_845_sv2v_reg  <= data_i[5];
      \nz.mem_844_sv2v_reg  <= data_i[4];
      \nz.mem_843_sv2v_reg  <= data_i[3];
      \nz.mem_842_sv2v_reg  <= data_i[2];
      \nz.mem_841_sv2v_reg  <= data_i[1];
      \nz.mem_840_sv2v_reg  <= data_i[0];
    end 
    if(N895) begin
      \nz.mem_839_sv2v_reg  <= data_i[7];
      \nz.mem_838_sv2v_reg  <= data_i[6];
      \nz.mem_837_sv2v_reg  <= data_i[5];
      \nz.mem_836_sv2v_reg  <= data_i[4];
      \nz.mem_835_sv2v_reg  <= data_i[3];
      \nz.mem_834_sv2v_reg  <= data_i[2];
      \nz.mem_833_sv2v_reg  <= data_i[1];
      \nz.mem_832_sv2v_reg  <= data_i[0];
    end 
    if(N894) begin
      \nz.mem_831_sv2v_reg  <= data_i[7];
      \nz.mem_830_sv2v_reg  <= data_i[6];
      \nz.mem_829_sv2v_reg  <= data_i[5];
      \nz.mem_828_sv2v_reg  <= data_i[4];
      \nz.mem_827_sv2v_reg  <= data_i[3];
      \nz.mem_826_sv2v_reg  <= data_i[2];
      \nz.mem_825_sv2v_reg  <= data_i[1];
      \nz.mem_824_sv2v_reg  <= data_i[0];
    end 
    if(N893) begin
      \nz.mem_823_sv2v_reg  <= data_i[7];
      \nz.mem_822_sv2v_reg  <= data_i[6];
      \nz.mem_821_sv2v_reg  <= data_i[5];
      \nz.mem_820_sv2v_reg  <= data_i[4];
      \nz.mem_819_sv2v_reg  <= data_i[3];
      \nz.mem_818_sv2v_reg  <= data_i[2];
      \nz.mem_817_sv2v_reg  <= data_i[1];
      \nz.mem_816_sv2v_reg  <= data_i[0];
    end 
    if(N892) begin
      \nz.mem_815_sv2v_reg  <= data_i[7];
      \nz.mem_814_sv2v_reg  <= data_i[6];
      \nz.mem_813_sv2v_reg  <= data_i[5];
      \nz.mem_812_sv2v_reg  <= data_i[4];
      \nz.mem_811_sv2v_reg  <= data_i[3];
      \nz.mem_810_sv2v_reg  <= data_i[2];
      \nz.mem_809_sv2v_reg  <= data_i[1];
      \nz.mem_808_sv2v_reg  <= data_i[0];
    end 
    if(N891) begin
      \nz.mem_807_sv2v_reg  <= data_i[7];
      \nz.mem_806_sv2v_reg  <= data_i[6];
      \nz.mem_805_sv2v_reg  <= data_i[5];
      \nz.mem_804_sv2v_reg  <= data_i[4];
      \nz.mem_803_sv2v_reg  <= data_i[3];
      \nz.mem_802_sv2v_reg  <= data_i[2];
      \nz.mem_801_sv2v_reg  <= data_i[1];
      \nz.mem_800_sv2v_reg  <= data_i[0];
    end 
    if(N890) begin
      \nz.mem_799_sv2v_reg  <= data_i[7];
      \nz.mem_798_sv2v_reg  <= data_i[6];
      \nz.mem_797_sv2v_reg  <= data_i[5];
      \nz.mem_796_sv2v_reg  <= data_i[4];
      \nz.mem_795_sv2v_reg  <= data_i[3];
      \nz.mem_794_sv2v_reg  <= data_i[2];
      \nz.mem_793_sv2v_reg  <= data_i[1];
      \nz.mem_792_sv2v_reg  <= data_i[0];
    end 
    if(N889) begin
      \nz.mem_791_sv2v_reg  <= data_i[7];
      \nz.mem_790_sv2v_reg  <= data_i[6];
      \nz.mem_789_sv2v_reg  <= data_i[5];
      \nz.mem_788_sv2v_reg  <= data_i[4];
      \nz.mem_787_sv2v_reg  <= data_i[3];
      \nz.mem_786_sv2v_reg  <= data_i[2];
      \nz.mem_785_sv2v_reg  <= data_i[1];
      \nz.mem_784_sv2v_reg  <= data_i[0];
    end 
    if(N888) begin
      \nz.mem_783_sv2v_reg  <= data_i[7];
      \nz.mem_782_sv2v_reg  <= data_i[6];
      \nz.mem_781_sv2v_reg  <= data_i[5];
      \nz.mem_780_sv2v_reg  <= data_i[4];
      \nz.mem_779_sv2v_reg  <= data_i[3];
      \nz.mem_778_sv2v_reg  <= data_i[2];
      \nz.mem_777_sv2v_reg  <= data_i[1];
      \nz.mem_776_sv2v_reg  <= data_i[0];
    end 
    if(N887) begin
      \nz.mem_775_sv2v_reg  <= data_i[7];
      \nz.mem_774_sv2v_reg  <= data_i[6];
      \nz.mem_773_sv2v_reg  <= data_i[5];
      \nz.mem_772_sv2v_reg  <= data_i[4];
      \nz.mem_771_sv2v_reg  <= data_i[3];
      \nz.mem_770_sv2v_reg  <= data_i[2];
      \nz.mem_769_sv2v_reg  <= data_i[1];
      \nz.mem_768_sv2v_reg  <= data_i[0];
    end 
    if(N886) begin
      \nz.mem_767_sv2v_reg  <= data_i[7];
      \nz.mem_766_sv2v_reg  <= data_i[6];
      \nz.mem_765_sv2v_reg  <= data_i[5];
      \nz.mem_764_sv2v_reg  <= data_i[4];
      \nz.mem_763_sv2v_reg  <= data_i[3];
      \nz.mem_762_sv2v_reg  <= data_i[2];
      \nz.mem_761_sv2v_reg  <= data_i[1];
      \nz.mem_760_sv2v_reg  <= data_i[0];
    end 
    if(N885) begin
      \nz.mem_759_sv2v_reg  <= data_i[7];
      \nz.mem_758_sv2v_reg  <= data_i[6];
      \nz.mem_757_sv2v_reg  <= data_i[5];
      \nz.mem_756_sv2v_reg  <= data_i[4];
      \nz.mem_755_sv2v_reg  <= data_i[3];
      \nz.mem_754_sv2v_reg  <= data_i[2];
      \nz.mem_753_sv2v_reg  <= data_i[1];
      \nz.mem_752_sv2v_reg  <= data_i[0];
    end 
    if(N884) begin
      \nz.mem_751_sv2v_reg  <= data_i[7];
      \nz.mem_750_sv2v_reg  <= data_i[6];
      \nz.mem_749_sv2v_reg  <= data_i[5];
      \nz.mem_748_sv2v_reg  <= data_i[4];
      \nz.mem_747_sv2v_reg  <= data_i[3];
      \nz.mem_746_sv2v_reg  <= data_i[2];
      \nz.mem_745_sv2v_reg  <= data_i[1];
      \nz.mem_744_sv2v_reg  <= data_i[0];
    end 
    if(N883) begin
      \nz.mem_743_sv2v_reg  <= data_i[7];
      \nz.mem_742_sv2v_reg  <= data_i[6];
      \nz.mem_741_sv2v_reg  <= data_i[5];
      \nz.mem_740_sv2v_reg  <= data_i[4];
      \nz.mem_739_sv2v_reg  <= data_i[3];
      \nz.mem_738_sv2v_reg  <= data_i[2];
      \nz.mem_737_sv2v_reg  <= data_i[1];
      \nz.mem_736_sv2v_reg  <= data_i[0];
    end 
    if(N882) begin
      \nz.mem_735_sv2v_reg  <= data_i[7];
      \nz.mem_734_sv2v_reg  <= data_i[6];
      \nz.mem_733_sv2v_reg  <= data_i[5];
      \nz.mem_732_sv2v_reg  <= data_i[4];
      \nz.mem_731_sv2v_reg  <= data_i[3];
      \nz.mem_730_sv2v_reg  <= data_i[2];
      \nz.mem_729_sv2v_reg  <= data_i[1];
      \nz.mem_728_sv2v_reg  <= data_i[0];
    end 
    if(N881) begin
      \nz.mem_727_sv2v_reg  <= data_i[7];
      \nz.mem_726_sv2v_reg  <= data_i[6];
      \nz.mem_725_sv2v_reg  <= data_i[5];
      \nz.mem_724_sv2v_reg  <= data_i[4];
      \nz.mem_723_sv2v_reg  <= data_i[3];
      \nz.mem_722_sv2v_reg  <= data_i[2];
      \nz.mem_721_sv2v_reg  <= data_i[1];
      \nz.mem_720_sv2v_reg  <= data_i[0];
    end 
    if(N880) begin
      \nz.mem_719_sv2v_reg  <= data_i[7];
      \nz.mem_718_sv2v_reg  <= data_i[6];
      \nz.mem_717_sv2v_reg  <= data_i[5];
      \nz.mem_716_sv2v_reg  <= data_i[4];
      \nz.mem_715_sv2v_reg  <= data_i[3];
      \nz.mem_714_sv2v_reg  <= data_i[2];
      \nz.mem_713_sv2v_reg  <= data_i[1];
      \nz.mem_712_sv2v_reg  <= data_i[0];
    end 
    if(N879) begin
      \nz.mem_711_sv2v_reg  <= data_i[7];
      \nz.mem_710_sv2v_reg  <= data_i[6];
      \nz.mem_709_sv2v_reg  <= data_i[5];
      \nz.mem_708_sv2v_reg  <= data_i[4];
      \nz.mem_707_sv2v_reg  <= data_i[3];
      \nz.mem_706_sv2v_reg  <= data_i[2];
      \nz.mem_705_sv2v_reg  <= data_i[1];
      \nz.mem_704_sv2v_reg  <= data_i[0];
    end 
    if(N878) begin
      \nz.mem_703_sv2v_reg  <= data_i[7];
      \nz.mem_702_sv2v_reg  <= data_i[6];
      \nz.mem_701_sv2v_reg  <= data_i[5];
      \nz.mem_700_sv2v_reg  <= data_i[4];
      \nz.mem_699_sv2v_reg  <= data_i[3];
      \nz.mem_698_sv2v_reg  <= data_i[2];
      \nz.mem_697_sv2v_reg  <= data_i[1];
      \nz.mem_696_sv2v_reg  <= data_i[0];
    end 
    if(N877) begin
      \nz.mem_695_sv2v_reg  <= data_i[7];
      \nz.mem_694_sv2v_reg  <= data_i[6];
      \nz.mem_693_sv2v_reg  <= data_i[5];
      \nz.mem_692_sv2v_reg  <= data_i[4];
      \nz.mem_691_sv2v_reg  <= data_i[3];
      \nz.mem_690_sv2v_reg  <= data_i[2];
      \nz.mem_689_sv2v_reg  <= data_i[1];
      \nz.mem_688_sv2v_reg  <= data_i[0];
    end 
    if(N876) begin
      \nz.mem_687_sv2v_reg  <= data_i[7];
      \nz.mem_686_sv2v_reg  <= data_i[6];
      \nz.mem_685_sv2v_reg  <= data_i[5];
      \nz.mem_684_sv2v_reg  <= data_i[4];
      \nz.mem_683_sv2v_reg  <= data_i[3];
      \nz.mem_682_sv2v_reg  <= data_i[2];
      \nz.mem_681_sv2v_reg  <= data_i[1];
      \nz.mem_680_sv2v_reg  <= data_i[0];
    end 
    if(N875) begin
      \nz.mem_679_sv2v_reg  <= data_i[7];
      \nz.mem_678_sv2v_reg  <= data_i[6];
      \nz.mem_677_sv2v_reg  <= data_i[5];
      \nz.mem_676_sv2v_reg  <= data_i[4];
      \nz.mem_675_sv2v_reg  <= data_i[3];
      \nz.mem_674_sv2v_reg  <= data_i[2];
      \nz.mem_673_sv2v_reg  <= data_i[1];
      \nz.mem_672_sv2v_reg  <= data_i[0];
    end 
    if(N874) begin
      \nz.mem_671_sv2v_reg  <= data_i[7];
      \nz.mem_670_sv2v_reg  <= data_i[6];
      \nz.mem_669_sv2v_reg  <= data_i[5];
      \nz.mem_668_sv2v_reg  <= data_i[4];
      \nz.mem_667_sv2v_reg  <= data_i[3];
      \nz.mem_666_sv2v_reg  <= data_i[2];
      \nz.mem_665_sv2v_reg  <= data_i[1];
      \nz.mem_664_sv2v_reg  <= data_i[0];
    end 
    if(N873) begin
      \nz.mem_663_sv2v_reg  <= data_i[7];
      \nz.mem_662_sv2v_reg  <= data_i[6];
      \nz.mem_661_sv2v_reg  <= data_i[5];
      \nz.mem_660_sv2v_reg  <= data_i[4];
      \nz.mem_659_sv2v_reg  <= data_i[3];
      \nz.mem_658_sv2v_reg  <= data_i[2];
      \nz.mem_657_sv2v_reg  <= data_i[1];
      \nz.mem_656_sv2v_reg  <= data_i[0];
    end 
    if(N872) begin
      \nz.mem_655_sv2v_reg  <= data_i[7];
      \nz.mem_654_sv2v_reg  <= data_i[6];
      \nz.mem_653_sv2v_reg  <= data_i[5];
      \nz.mem_652_sv2v_reg  <= data_i[4];
      \nz.mem_651_sv2v_reg  <= data_i[3];
      \nz.mem_650_sv2v_reg  <= data_i[2];
      \nz.mem_649_sv2v_reg  <= data_i[1];
      \nz.mem_648_sv2v_reg  <= data_i[0];
    end 
    if(N871) begin
      \nz.mem_647_sv2v_reg  <= data_i[7];
      \nz.mem_646_sv2v_reg  <= data_i[6];
      \nz.mem_645_sv2v_reg  <= data_i[5];
      \nz.mem_644_sv2v_reg  <= data_i[4];
      \nz.mem_643_sv2v_reg  <= data_i[3];
      \nz.mem_642_sv2v_reg  <= data_i[2];
      \nz.mem_641_sv2v_reg  <= data_i[1];
      \nz.mem_640_sv2v_reg  <= data_i[0];
    end 
    if(N870) begin
      \nz.mem_639_sv2v_reg  <= data_i[7];
      \nz.mem_638_sv2v_reg  <= data_i[6];
      \nz.mem_637_sv2v_reg  <= data_i[5];
      \nz.mem_636_sv2v_reg  <= data_i[4];
      \nz.mem_635_sv2v_reg  <= data_i[3];
      \nz.mem_634_sv2v_reg  <= data_i[2];
      \nz.mem_633_sv2v_reg  <= data_i[1];
      \nz.mem_632_sv2v_reg  <= data_i[0];
    end 
    if(N869) begin
      \nz.mem_631_sv2v_reg  <= data_i[7];
      \nz.mem_630_sv2v_reg  <= data_i[6];
      \nz.mem_629_sv2v_reg  <= data_i[5];
      \nz.mem_628_sv2v_reg  <= data_i[4];
      \nz.mem_627_sv2v_reg  <= data_i[3];
      \nz.mem_626_sv2v_reg  <= data_i[2];
      \nz.mem_625_sv2v_reg  <= data_i[1];
      \nz.mem_624_sv2v_reg  <= data_i[0];
    end 
    if(N868) begin
      \nz.mem_623_sv2v_reg  <= data_i[7];
      \nz.mem_622_sv2v_reg  <= data_i[6];
      \nz.mem_621_sv2v_reg  <= data_i[5];
      \nz.mem_620_sv2v_reg  <= data_i[4];
      \nz.mem_619_sv2v_reg  <= data_i[3];
      \nz.mem_618_sv2v_reg  <= data_i[2];
      \nz.mem_617_sv2v_reg  <= data_i[1];
      \nz.mem_616_sv2v_reg  <= data_i[0];
    end 
    if(N867) begin
      \nz.mem_615_sv2v_reg  <= data_i[7];
      \nz.mem_614_sv2v_reg  <= data_i[6];
      \nz.mem_613_sv2v_reg  <= data_i[5];
      \nz.mem_612_sv2v_reg  <= data_i[4];
      \nz.mem_611_sv2v_reg  <= data_i[3];
      \nz.mem_610_sv2v_reg  <= data_i[2];
      \nz.mem_609_sv2v_reg  <= data_i[1];
      \nz.mem_608_sv2v_reg  <= data_i[0];
    end 
    if(N866) begin
      \nz.mem_607_sv2v_reg  <= data_i[7];
      \nz.mem_606_sv2v_reg  <= data_i[6];
      \nz.mem_605_sv2v_reg  <= data_i[5];
      \nz.mem_604_sv2v_reg  <= data_i[4];
      \nz.mem_603_sv2v_reg  <= data_i[3];
      \nz.mem_602_sv2v_reg  <= data_i[2];
      \nz.mem_601_sv2v_reg  <= data_i[1];
      \nz.mem_600_sv2v_reg  <= data_i[0];
    end 
    if(N865) begin
      \nz.mem_599_sv2v_reg  <= data_i[7];
      \nz.mem_598_sv2v_reg  <= data_i[6];
      \nz.mem_597_sv2v_reg  <= data_i[5];
      \nz.mem_596_sv2v_reg  <= data_i[4];
      \nz.mem_595_sv2v_reg  <= data_i[3];
      \nz.mem_594_sv2v_reg  <= data_i[2];
      \nz.mem_593_sv2v_reg  <= data_i[1];
      \nz.mem_592_sv2v_reg  <= data_i[0];
    end 
    if(N864) begin
      \nz.mem_591_sv2v_reg  <= data_i[7];
      \nz.mem_590_sv2v_reg  <= data_i[6];
      \nz.mem_589_sv2v_reg  <= data_i[5];
      \nz.mem_588_sv2v_reg  <= data_i[4];
      \nz.mem_587_sv2v_reg  <= data_i[3];
      \nz.mem_586_sv2v_reg  <= data_i[2];
      \nz.mem_585_sv2v_reg  <= data_i[1];
      \nz.mem_584_sv2v_reg  <= data_i[0];
    end 
    if(N863) begin
      \nz.mem_583_sv2v_reg  <= data_i[7];
      \nz.mem_582_sv2v_reg  <= data_i[6];
      \nz.mem_581_sv2v_reg  <= data_i[5];
      \nz.mem_580_sv2v_reg  <= data_i[4];
      \nz.mem_579_sv2v_reg  <= data_i[3];
      \nz.mem_578_sv2v_reg  <= data_i[2];
      \nz.mem_577_sv2v_reg  <= data_i[1];
      \nz.mem_576_sv2v_reg  <= data_i[0];
    end 
    if(N862) begin
      \nz.mem_575_sv2v_reg  <= data_i[7];
      \nz.mem_574_sv2v_reg  <= data_i[6];
      \nz.mem_573_sv2v_reg  <= data_i[5];
      \nz.mem_572_sv2v_reg  <= data_i[4];
      \nz.mem_571_sv2v_reg  <= data_i[3];
      \nz.mem_570_sv2v_reg  <= data_i[2];
      \nz.mem_569_sv2v_reg  <= data_i[1];
      \nz.mem_568_sv2v_reg  <= data_i[0];
    end 
    if(N861) begin
      \nz.mem_567_sv2v_reg  <= data_i[7];
      \nz.mem_566_sv2v_reg  <= data_i[6];
      \nz.mem_565_sv2v_reg  <= data_i[5];
      \nz.mem_564_sv2v_reg  <= data_i[4];
      \nz.mem_563_sv2v_reg  <= data_i[3];
      \nz.mem_562_sv2v_reg  <= data_i[2];
      \nz.mem_561_sv2v_reg  <= data_i[1];
      \nz.mem_560_sv2v_reg  <= data_i[0];
    end 
    if(N860) begin
      \nz.mem_559_sv2v_reg  <= data_i[7];
      \nz.mem_558_sv2v_reg  <= data_i[6];
      \nz.mem_557_sv2v_reg  <= data_i[5];
      \nz.mem_556_sv2v_reg  <= data_i[4];
      \nz.mem_555_sv2v_reg  <= data_i[3];
      \nz.mem_554_sv2v_reg  <= data_i[2];
      \nz.mem_553_sv2v_reg  <= data_i[1];
      \nz.mem_552_sv2v_reg  <= data_i[0];
    end 
    if(N859) begin
      \nz.mem_551_sv2v_reg  <= data_i[7];
      \nz.mem_550_sv2v_reg  <= data_i[6];
      \nz.mem_549_sv2v_reg  <= data_i[5];
      \nz.mem_548_sv2v_reg  <= data_i[4];
      \nz.mem_547_sv2v_reg  <= data_i[3];
      \nz.mem_546_sv2v_reg  <= data_i[2];
      \nz.mem_545_sv2v_reg  <= data_i[1];
      \nz.mem_544_sv2v_reg  <= data_i[0];
    end 
    if(N858) begin
      \nz.mem_543_sv2v_reg  <= data_i[7];
      \nz.mem_542_sv2v_reg  <= data_i[6];
      \nz.mem_541_sv2v_reg  <= data_i[5];
      \nz.mem_540_sv2v_reg  <= data_i[4];
      \nz.mem_539_sv2v_reg  <= data_i[3];
      \nz.mem_538_sv2v_reg  <= data_i[2];
      \nz.mem_537_sv2v_reg  <= data_i[1];
      \nz.mem_536_sv2v_reg  <= data_i[0];
    end 
    if(N857) begin
      \nz.mem_535_sv2v_reg  <= data_i[7];
      \nz.mem_534_sv2v_reg  <= data_i[6];
      \nz.mem_533_sv2v_reg  <= data_i[5];
      \nz.mem_532_sv2v_reg  <= data_i[4];
      \nz.mem_531_sv2v_reg  <= data_i[3];
      \nz.mem_530_sv2v_reg  <= data_i[2];
      \nz.mem_529_sv2v_reg  <= data_i[1];
      \nz.mem_528_sv2v_reg  <= data_i[0];
    end 
    if(N856) begin
      \nz.mem_527_sv2v_reg  <= data_i[7];
      \nz.mem_526_sv2v_reg  <= data_i[6];
      \nz.mem_525_sv2v_reg  <= data_i[5];
      \nz.mem_524_sv2v_reg  <= data_i[4];
      \nz.mem_523_sv2v_reg  <= data_i[3];
      \nz.mem_522_sv2v_reg  <= data_i[2];
      \nz.mem_521_sv2v_reg  <= data_i[1];
      \nz.mem_520_sv2v_reg  <= data_i[0];
    end 
    if(N855) begin
      \nz.mem_519_sv2v_reg  <= data_i[7];
      \nz.mem_518_sv2v_reg  <= data_i[6];
      \nz.mem_517_sv2v_reg  <= data_i[5];
      \nz.mem_516_sv2v_reg  <= data_i[4];
      \nz.mem_515_sv2v_reg  <= data_i[3];
      \nz.mem_514_sv2v_reg  <= data_i[2];
      \nz.mem_513_sv2v_reg  <= data_i[1];
      \nz.mem_512_sv2v_reg  <= data_i[0];
    end 
    if(N854) begin
      \nz.mem_511_sv2v_reg  <= data_i[7];
      \nz.mem_510_sv2v_reg  <= data_i[6];
      \nz.mem_509_sv2v_reg  <= data_i[5];
      \nz.mem_508_sv2v_reg  <= data_i[4];
      \nz.mem_507_sv2v_reg  <= data_i[3];
      \nz.mem_506_sv2v_reg  <= data_i[2];
      \nz.mem_505_sv2v_reg  <= data_i[1];
      \nz.mem_504_sv2v_reg  <= data_i[0];
    end 
    if(N853) begin
      \nz.mem_503_sv2v_reg  <= data_i[7];
      \nz.mem_502_sv2v_reg  <= data_i[6];
      \nz.mem_501_sv2v_reg  <= data_i[5];
      \nz.mem_500_sv2v_reg  <= data_i[4];
      \nz.mem_499_sv2v_reg  <= data_i[3];
      \nz.mem_498_sv2v_reg  <= data_i[2];
      \nz.mem_497_sv2v_reg  <= data_i[1];
      \nz.mem_496_sv2v_reg  <= data_i[0];
    end 
    if(N852) begin
      \nz.mem_495_sv2v_reg  <= data_i[7];
      \nz.mem_494_sv2v_reg  <= data_i[6];
      \nz.mem_493_sv2v_reg  <= data_i[5];
      \nz.mem_492_sv2v_reg  <= data_i[4];
      \nz.mem_491_sv2v_reg  <= data_i[3];
      \nz.mem_490_sv2v_reg  <= data_i[2];
      \nz.mem_489_sv2v_reg  <= data_i[1];
      \nz.mem_488_sv2v_reg  <= data_i[0];
    end 
    if(N851) begin
      \nz.mem_487_sv2v_reg  <= data_i[7];
      \nz.mem_486_sv2v_reg  <= data_i[6];
      \nz.mem_485_sv2v_reg  <= data_i[5];
      \nz.mem_484_sv2v_reg  <= data_i[4];
      \nz.mem_483_sv2v_reg  <= data_i[3];
      \nz.mem_482_sv2v_reg  <= data_i[2];
      \nz.mem_481_sv2v_reg  <= data_i[1];
      \nz.mem_480_sv2v_reg  <= data_i[0];
    end 
    if(N850) begin
      \nz.mem_479_sv2v_reg  <= data_i[7];
      \nz.mem_478_sv2v_reg  <= data_i[6];
      \nz.mem_477_sv2v_reg  <= data_i[5];
      \nz.mem_476_sv2v_reg  <= data_i[4];
      \nz.mem_475_sv2v_reg  <= data_i[3];
      \nz.mem_474_sv2v_reg  <= data_i[2];
      \nz.mem_473_sv2v_reg  <= data_i[1];
      \nz.mem_472_sv2v_reg  <= data_i[0];
    end 
    if(N849) begin
      \nz.mem_471_sv2v_reg  <= data_i[7];
      \nz.mem_470_sv2v_reg  <= data_i[6];
      \nz.mem_469_sv2v_reg  <= data_i[5];
      \nz.mem_468_sv2v_reg  <= data_i[4];
      \nz.mem_467_sv2v_reg  <= data_i[3];
      \nz.mem_466_sv2v_reg  <= data_i[2];
      \nz.mem_465_sv2v_reg  <= data_i[1];
      \nz.mem_464_sv2v_reg  <= data_i[0];
    end 
    if(N848) begin
      \nz.mem_463_sv2v_reg  <= data_i[7];
      \nz.mem_462_sv2v_reg  <= data_i[6];
      \nz.mem_461_sv2v_reg  <= data_i[5];
      \nz.mem_460_sv2v_reg  <= data_i[4];
      \nz.mem_459_sv2v_reg  <= data_i[3];
      \nz.mem_458_sv2v_reg  <= data_i[2];
      \nz.mem_457_sv2v_reg  <= data_i[1];
      \nz.mem_456_sv2v_reg  <= data_i[0];
    end 
    if(N847) begin
      \nz.mem_455_sv2v_reg  <= data_i[7];
      \nz.mem_454_sv2v_reg  <= data_i[6];
      \nz.mem_453_sv2v_reg  <= data_i[5];
      \nz.mem_452_sv2v_reg  <= data_i[4];
      \nz.mem_451_sv2v_reg  <= data_i[3];
      \nz.mem_450_sv2v_reg  <= data_i[2];
      \nz.mem_449_sv2v_reg  <= data_i[1];
      \nz.mem_448_sv2v_reg  <= data_i[0];
    end 
    if(N846) begin
      \nz.mem_447_sv2v_reg  <= data_i[7];
      \nz.mem_446_sv2v_reg  <= data_i[6];
      \nz.mem_445_sv2v_reg  <= data_i[5];
      \nz.mem_444_sv2v_reg  <= data_i[4];
      \nz.mem_443_sv2v_reg  <= data_i[3];
      \nz.mem_442_sv2v_reg  <= data_i[2];
      \nz.mem_441_sv2v_reg  <= data_i[1];
      \nz.mem_440_sv2v_reg  <= data_i[0];
    end 
    if(N845) begin
      \nz.mem_439_sv2v_reg  <= data_i[7];
      \nz.mem_438_sv2v_reg  <= data_i[6];
      \nz.mem_437_sv2v_reg  <= data_i[5];
      \nz.mem_436_sv2v_reg  <= data_i[4];
      \nz.mem_435_sv2v_reg  <= data_i[3];
      \nz.mem_434_sv2v_reg  <= data_i[2];
      \nz.mem_433_sv2v_reg  <= data_i[1];
      \nz.mem_432_sv2v_reg  <= data_i[0];
    end 
    if(N844) begin
      \nz.mem_431_sv2v_reg  <= data_i[7];
      \nz.mem_430_sv2v_reg  <= data_i[6];
      \nz.mem_429_sv2v_reg  <= data_i[5];
      \nz.mem_428_sv2v_reg  <= data_i[4];
      \nz.mem_427_sv2v_reg  <= data_i[3];
      \nz.mem_426_sv2v_reg  <= data_i[2];
      \nz.mem_425_sv2v_reg  <= data_i[1];
      \nz.mem_424_sv2v_reg  <= data_i[0];
    end 
    if(N843) begin
      \nz.mem_423_sv2v_reg  <= data_i[7];
      \nz.mem_422_sv2v_reg  <= data_i[6];
      \nz.mem_421_sv2v_reg  <= data_i[5];
      \nz.mem_420_sv2v_reg  <= data_i[4];
      \nz.mem_419_sv2v_reg  <= data_i[3];
      \nz.mem_418_sv2v_reg  <= data_i[2];
      \nz.mem_417_sv2v_reg  <= data_i[1];
      \nz.mem_416_sv2v_reg  <= data_i[0];
    end 
    if(N842) begin
      \nz.mem_415_sv2v_reg  <= data_i[7];
      \nz.mem_414_sv2v_reg  <= data_i[6];
      \nz.mem_413_sv2v_reg  <= data_i[5];
      \nz.mem_412_sv2v_reg  <= data_i[4];
      \nz.mem_411_sv2v_reg  <= data_i[3];
      \nz.mem_410_sv2v_reg  <= data_i[2];
      \nz.mem_409_sv2v_reg  <= data_i[1];
      \nz.mem_408_sv2v_reg  <= data_i[0];
    end 
    if(N841) begin
      \nz.mem_407_sv2v_reg  <= data_i[7];
      \nz.mem_406_sv2v_reg  <= data_i[6];
      \nz.mem_405_sv2v_reg  <= data_i[5];
      \nz.mem_404_sv2v_reg  <= data_i[4];
      \nz.mem_403_sv2v_reg  <= data_i[3];
      \nz.mem_402_sv2v_reg  <= data_i[2];
      \nz.mem_401_sv2v_reg  <= data_i[1];
      \nz.mem_400_sv2v_reg  <= data_i[0];
    end 
    if(N840) begin
      \nz.mem_399_sv2v_reg  <= data_i[7];
      \nz.mem_398_sv2v_reg  <= data_i[6];
      \nz.mem_397_sv2v_reg  <= data_i[5];
      \nz.mem_396_sv2v_reg  <= data_i[4];
      \nz.mem_395_sv2v_reg  <= data_i[3];
      \nz.mem_394_sv2v_reg  <= data_i[2];
      \nz.mem_393_sv2v_reg  <= data_i[1];
      \nz.mem_392_sv2v_reg  <= data_i[0];
    end 
    if(N839) begin
      \nz.mem_391_sv2v_reg  <= data_i[7];
      \nz.mem_390_sv2v_reg  <= data_i[6];
      \nz.mem_389_sv2v_reg  <= data_i[5];
      \nz.mem_388_sv2v_reg  <= data_i[4];
      \nz.mem_387_sv2v_reg  <= data_i[3];
      \nz.mem_386_sv2v_reg  <= data_i[2];
      \nz.mem_385_sv2v_reg  <= data_i[1];
      \nz.mem_384_sv2v_reg  <= data_i[0];
    end 
    if(N838) begin
      \nz.mem_383_sv2v_reg  <= data_i[7];
      \nz.mem_382_sv2v_reg  <= data_i[6];
      \nz.mem_381_sv2v_reg  <= data_i[5];
      \nz.mem_380_sv2v_reg  <= data_i[4];
      \nz.mem_379_sv2v_reg  <= data_i[3];
      \nz.mem_378_sv2v_reg  <= data_i[2];
      \nz.mem_377_sv2v_reg  <= data_i[1];
      \nz.mem_376_sv2v_reg  <= data_i[0];
    end 
    if(N837) begin
      \nz.mem_375_sv2v_reg  <= data_i[7];
      \nz.mem_374_sv2v_reg  <= data_i[6];
      \nz.mem_373_sv2v_reg  <= data_i[5];
      \nz.mem_372_sv2v_reg  <= data_i[4];
      \nz.mem_371_sv2v_reg  <= data_i[3];
      \nz.mem_370_sv2v_reg  <= data_i[2];
      \nz.mem_369_sv2v_reg  <= data_i[1];
      \nz.mem_368_sv2v_reg  <= data_i[0];
    end 
    if(N836) begin
      \nz.mem_367_sv2v_reg  <= data_i[7];
      \nz.mem_366_sv2v_reg  <= data_i[6];
      \nz.mem_365_sv2v_reg  <= data_i[5];
      \nz.mem_364_sv2v_reg  <= data_i[4];
      \nz.mem_363_sv2v_reg  <= data_i[3];
      \nz.mem_362_sv2v_reg  <= data_i[2];
      \nz.mem_361_sv2v_reg  <= data_i[1];
      \nz.mem_360_sv2v_reg  <= data_i[0];
    end 
    if(N835) begin
      \nz.mem_359_sv2v_reg  <= data_i[7];
      \nz.mem_358_sv2v_reg  <= data_i[6];
      \nz.mem_357_sv2v_reg  <= data_i[5];
      \nz.mem_356_sv2v_reg  <= data_i[4];
      \nz.mem_355_sv2v_reg  <= data_i[3];
      \nz.mem_354_sv2v_reg  <= data_i[2];
      \nz.mem_353_sv2v_reg  <= data_i[1];
      \nz.mem_352_sv2v_reg  <= data_i[0];
    end 
    if(N834) begin
      \nz.mem_351_sv2v_reg  <= data_i[7];
      \nz.mem_350_sv2v_reg  <= data_i[6];
      \nz.mem_349_sv2v_reg  <= data_i[5];
      \nz.mem_348_sv2v_reg  <= data_i[4];
      \nz.mem_347_sv2v_reg  <= data_i[3];
      \nz.mem_346_sv2v_reg  <= data_i[2];
      \nz.mem_345_sv2v_reg  <= data_i[1];
      \nz.mem_344_sv2v_reg  <= data_i[0];
    end 
    if(N833) begin
      \nz.mem_343_sv2v_reg  <= data_i[7];
      \nz.mem_342_sv2v_reg  <= data_i[6];
      \nz.mem_341_sv2v_reg  <= data_i[5];
      \nz.mem_340_sv2v_reg  <= data_i[4];
      \nz.mem_339_sv2v_reg  <= data_i[3];
      \nz.mem_338_sv2v_reg  <= data_i[2];
      \nz.mem_337_sv2v_reg  <= data_i[1];
      \nz.mem_336_sv2v_reg  <= data_i[0];
    end 
    if(N832) begin
      \nz.mem_335_sv2v_reg  <= data_i[7];
      \nz.mem_334_sv2v_reg  <= data_i[6];
      \nz.mem_333_sv2v_reg  <= data_i[5];
      \nz.mem_332_sv2v_reg  <= data_i[4];
      \nz.mem_331_sv2v_reg  <= data_i[3];
      \nz.mem_330_sv2v_reg  <= data_i[2];
      \nz.mem_329_sv2v_reg  <= data_i[1];
      \nz.mem_328_sv2v_reg  <= data_i[0];
    end 
    if(N831) begin
      \nz.mem_327_sv2v_reg  <= data_i[7];
      \nz.mem_326_sv2v_reg  <= data_i[6];
      \nz.mem_325_sv2v_reg  <= data_i[5];
      \nz.mem_324_sv2v_reg  <= data_i[4];
      \nz.mem_323_sv2v_reg  <= data_i[3];
      \nz.mem_322_sv2v_reg  <= data_i[2];
      \nz.mem_321_sv2v_reg  <= data_i[1];
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N830) begin
      \nz.mem_319_sv2v_reg  <= data_i[7];
      \nz.mem_318_sv2v_reg  <= data_i[6];
      \nz.mem_317_sv2v_reg  <= data_i[5];
      \nz.mem_316_sv2v_reg  <= data_i[4];
      \nz.mem_315_sv2v_reg  <= data_i[3];
      \nz.mem_314_sv2v_reg  <= data_i[2];
      \nz.mem_313_sv2v_reg  <= data_i[1];
      \nz.mem_312_sv2v_reg  <= data_i[0];
    end 
    if(N829) begin
      \nz.mem_311_sv2v_reg  <= data_i[7];
      \nz.mem_310_sv2v_reg  <= data_i[6];
      \nz.mem_309_sv2v_reg  <= data_i[5];
      \nz.mem_308_sv2v_reg  <= data_i[4];
      \nz.mem_307_sv2v_reg  <= data_i[3];
      \nz.mem_306_sv2v_reg  <= data_i[2];
      \nz.mem_305_sv2v_reg  <= data_i[1];
      \nz.mem_304_sv2v_reg  <= data_i[0];
    end 
    if(N828) begin
      \nz.mem_303_sv2v_reg  <= data_i[7];
      \nz.mem_302_sv2v_reg  <= data_i[6];
      \nz.mem_301_sv2v_reg  <= data_i[5];
      \nz.mem_300_sv2v_reg  <= data_i[4];
      \nz.mem_299_sv2v_reg  <= data_i[3];
      \nz.mem_298_sv2v_reg  <= data_i[2];
      \nz.mem_297_sv2v_reg  <= data_i[1];
      \nz.mem_296_sv2v_reg  <= data_i[0];
    end 
    if(N827) begin
      \nz.mem_295_sv2v_reg  <= data_i[7];
      \nz.mem_294_sv2v_reg  <= data_i[6];
      \nz.mem_293_sv2v_reg  <= data_i[5];
      \nz.mem_292_sv2v_reg  <= data_i[4];
      \nz.mem_291_sv2v_reg  <= data_i[3];
      \nz.mem_290_sv2v_reg  <= data_i[2];
      \nz.mem_289_sv2v_reg  <= data_i[1];
      \nz.mem_288_sv2v_reg  <= data_i[0];
    end 
    if(N826) begin
      \nz.mem_287_sv2v_reg  <= data_i[7];
      \nz.mem_286_sv2v_reg  <= data_i[6];
      \nz.mem_285_sv2v_reg  <= data_i[5];
      \nz.mem_284_sv2v_reg  <= data_i[4];
      \nz.mem_283_sv2v_reg  <= data_i[3];
      \nz.mem_282_sv2v_reg  <= data_i[2];
      \nz.mem_281_sv2v_reg  <= data_i[1];
      \nz.mem_280_sv2v_reg  <= data_i[0];
    end 
    if(N825) begin
      \nz.mem_279_sv2v_reg  <= data_i[7];
      \nz.mem_278_sv2v_reg  <= data_i[6];
      \nz.mem_277_sv2v_reg  <= data_i[5];
      \nz.mem_276_sv2v_reg  <= data_i[4];
      \nz.mem_275_sv2v_reg  <= data_i[3];
      \nz.mem_274_sv2v_reg  <= data_i[2];
      \nz.mem_273_sv2v_reg  <= data_i[1];
      \nz.mem_272_sv2v_reg  <= data_i[0];
    end 
    if(N824) begin
      \nz.mem_271_sv2v_reg  <= data_i[7];
      \nz.mem_270_sv2v_reg  <= data_i[6];
      \nz.mem_269_sv2v_reg  <= data_i[5];
      \nz.mem_268_sv2v_reg  <= data_i[4];
      \nz.mem_267_sv2v_reg  <= data_i[3];
      \nz.mem_266_sv2v_reg  <= data_i[2];
      \nz.mem_265_sv2v_reg  <= data_i[1];
      \nz.mem_264_sv2v_reg  <= data_i[0];
    end 
    if(N823) begin
      \nz.mem_263_sv2v_reg  <= data_i[7];
      \nz.mem_262_sv2v_reg  <= data_i[6];
      \nz.mem_261_sv2v_reg  <= data_i[5];
      \nz.mem_260_sv2v_reg  <= data_i[4];
      \nz.mem_259_sv2v_reg  <= data_i[3];
      \nz.mem_258_sv2v_reg  <= data_i[2];
      \nz.mem_257_sv2v_reg  <= data_i[1];
      \nz.mem_256_sv2v_reg  <= data_i[0];
    end 
    if(N822) begin
      \nz.mem_255_sv2v_reg  <= data_i[7];
      \nz.mem_254_sv2v_reg  <= data_i[6];
      \nz.mem_253_sv2v_reg  <= data_i[5];
      \nz.mem_252_sv2v_reg  <= data_i[4];
      \nz.mem_251_sv2v_reg  <= data_i[3];
      \nz.mem_250_sv2v_reg  <= data_i[2];
      \nz.mem_249_sv2v_reg  <= data_i[1];
      \nz.mem_248_sv2v_reg  <= data_i[0];
    end 
    if(N821) begin
      \nz.mem_247_sv2v_reg  <= data_i[7];
      \nz.mem_246_sv2v_reg  <= data_i[6];
      \nz.mem_245_sv2v_reg  <= data_i[5];
      \nz.mem_244_sv2v_reg  <= data_i[4];
      \nz.mem_243_sv2v_reg  <= data_i[3];
      \nz.mem_242_sv2v_reg  <= data_i[2];
      \nz.mem_241_sv2v_reg  <= data_i[1];
      \nz.mem_240_sv2v_reg  <= data_i[0];
    end 
    if(N820) begin
      \nz.mem_239_sv2v_reg  <= data_i[7];
      \nz.mem_238_sv2v_reg  <= data_i[6];
      \nz.mem_237_sv2v_reg  <= data_i[5];
      \nz.mem_236_sv2v_reg  <= data_i[4];
      \nz.mem_235_sv2v_reg  <= data_i[3];
      \nz.mem_234_sv2v_reg  <= data_i[2];
      \nz.mem_233_sv2v_reg  <= data_i[1];
      \nz.mem_232_sv2v_reg  <= data_i[0];
    end 
    if(N819) begin
      \nz.mem_231_sv2v_reg  <= data_i[7];
      \nz.mem_230_sv2v_reg  <= data_i[6];
      \nz.mem_229_sv2v_reg  <= data_i[5];
      \nz.mem_228_sv2v_reg  <= data_i[4];
      \nz.mem_227_sv2v_reg  <= data_i[3];
      \nz.mem_226_sv2v_reg  <= data_i[2];
      \nz.mem_225_sv2v_reg  <= data_i[1];
      \nz.mem_224_sv2v_reg  <= data_i[0];
    end 
    if(N818) begin
      \nz.mem_223_sv2v_reg  <= data_i[7];
      \nz.mem_222_sv2v_reg  <= data_i[6];
      \nz.mem_221_sv2v_reg  <= data_i[5];
      \nz.mem_220_sv2v_reg  <= data_i[4];
      \nz.mem_219_sv2v_reg  <= data_i[3];
      \nz.mem_218_sv2v_reg  <= data_i[2];
      \nz.mem_217_sv2v_reg  <= data_i[1];
      \nz.mem_216_sv2v_reg  <= data_i[0];
    end 
    if(N817) begin
      \nz.mem_215_sv2v_reg  <= data_i[7];
      \nz.mem_214_sv2v_reg  <= data_i[6];
      \nz.mem_213_sv2v_reg  <= data_i[5];
      \nz.mem_212_sv2v_reg  <= data_i[4];
      \nz.mem_211_sv2v_reg  <= data_i[3];
      \nz.mem_210_sv2v_reg  <= data_i[2];
      \nz.mem_209_sv2v_reg  <= data_i[1];
      \nz.mem_208_sv2v_reg  <= data_i[0];
    end 
    if(N816) begin
      \nz.mem_207_sv2v_reg  <= data_i[7];
      \nz.mem_206_sv2v_reg  <= data_i[6];
      \nz.mem_205_sv2v_reg  <= data_i[5];
      \nz.mem_204_sv2v_reg  <= data_i[4];
      \nz.mem_203_sv2v_reg  <= data_i[3];
      \nz.mem_202_sv2v_reg  <= data_i[2];
      \nz.mem_201_sv2v_reg  <= data_i[1];
      \nz.mem_200_sv2v_reg  <= data_i[0];
    end 
    if(N815) begin
      \nz.mem_199_sv2v_reg  <= data_i[7];
      \nz.mem_198_sv2v_reg  <= data_i[6];
      \nz.mem_197_sv2v_reg  <= data_i[5];
      \nz.mem_196_sv2v_reg  <= data_i[4];
      \nz.mem_195_sv2v_reg  <= data_i[3];
      \nz.mem_194_sv2v_reg  <= data_i[2];
      \nz.mem_193_sv2v_reg  <= data_i[1];
      \nz.mem_192_sv2v_reg  <= data_i[0];
    end 
    if(N814) begin
      \nz.mem_191_sv2v_reg  <= data_i[7];
      \nz.mem_190_sv2v_reg  <= data_i[6];
      \nz.mem_189_sv2v_reg  <= data_i[5];
      \nz.mem_188_sv2v_reg  <= data_i[4];
      \nz.mem_187_sv2v_reg  <= data_i[3];
      \nz.mem_186_sv2v_reg  <= data_i[2];
      \nz.mem_185_sv2v_reg  <= data_i[1];
      \nz.mem_184_sv2v_reg  <= data_i[0];
    end 
    if(N813) begin
      \nz.mem_183_sv2v_reg  <= data_i[7];
      \nz.mem_182_sv2v_reg  <= data_i[6];
      \nz.mem_181_sv2v_reg  <= data_i[5];
      \nz.mem_180_sv2v_reg  <= data_i[4];
      \nz.mem_179_sv2v_reg  <= data_i[3];
      \nz.mem_178_sv2v_reg  <= data_i[2];
      \nz.mem_177_sv2v_reg  <= data_i[1];
      \nz.mem_176_sv2v_reg  <= data_i[0];
    end 
    if(N812) begin
      \nz.mem_175_sv2v_reg  <= data_i[7];
      \nz.mem_174_sv2v_reg  <= data_i[6];
      \nz.mem_173_sv2v_reg  <= data_i[5];
      \nz.mem_172_sv2v_reg  <= data_i[4];
      \nz.mem_171_sv2v_reg  <= data_i[3];
      \nz.mem_170_sv2v_reg  <= data_i[2];
      \nz.mem_169_sv2v_reg  <= data_i[1];
      \nz.mem_168_sv2v_reg  <= data_i[0];
    end 
    if(N811) begin
      \nz.mem_167_sv2v_reg  <= data_i[7];
      \nz.mem_166_sv2v_reg  <= data_i[6];
      \nz.mem_165_sv2v_reg  <= data_i[5];
      \nz.mem_164_sv2v_reg  <= data_i[4];
      \nz.mem_163_sv2v_reg  <= data_i[3];
      \nz.mem_162_sv2v_reg  <= data_i[2];
      \nz.mem_161_sv2v_reg  <= data_i[1];
      \nz.mem_160_sv2v_reg  <= data_i[0];
    end 
    if(N810) begin
      \nz.mem_159_sv2v_reg  <= data_i[7];
      \nz.mem_158_sv2v_reg  <= data_i[6];
      \nz.mem_157_sv2v_reg  <= data_i[5];
      \nz.mem_156_sv2v_reg  <= data_i[4];
      \nz.mem_155_sv2v_reg  <= data_i[3];
      \nz.mem_154_sv2v_reg  <= data_i[2];
      \nz.mem_153_sv2v_reg  <= data_i[1];
      \nz.mem_152_sv2v_reg  <= data_i[0];
    end 
    if(N809) begin
      \nz.mem_151_sv2v_reg  <= data_i[7];
      \nz.mem_150_sv2v_reg  <= data_i[6];
      \nz.mem_149_sv2v_reg  <= data_i[5];
      \nz.mem_148_sv2v_reg  <= data_i[4];
      \nz.mem_147_sv2v_reg  <= data_i[3];
      \nz.mem_146_sv2v_reg  <= data_i[2];
      \nz.mem_145_sv2v_reg  <= data_i[1];
      \nz.mem_144_sv2v_reg  <= data_i[0];
    end 
    if(N808) begin
      \nz.mem_143_sv2v_reg  <= data_i[7];
      \nz.mem_142_sv2v_reg  <= data_i[6];
      \nz.mem_141_sv2v_reg  <= data_i[5];
      \nz.mem_140_sv2v_reg  <= data_i[4];
      \nz.mem_139_sv2v_reg  <= data_i[3];
      \nz.mem_138_sv2v_reg  <= data_i[2];
      \nz.mem_137_sv2v_reg  <= data_i[1];
      \nz.mem_136_sv2v_reg  <= data_i[0];
    end 
    if(N807) begin
      \nz.mem_135_sv2v_reg  <= data_i[7];
      \nz.mem_134_sv2v_reg  <= data_i[6];
      \nz.mem_133_sv2v_reg  <= data_i[5];
      \nz.mem_132_sv2v_reg  <= data_i[4];
      \nz.mem_131_sv2v_reg  <= data_i[3];
      \nz.mem_130_sv2v_reg  <= data_i[2];
      \nz.mem_129_sv2v_reg  <= data_i[1];
      \nz.mem_128_sv2v_reg  <= data_i[0];
    end 
    if(N806) begin
      \nz.mem_127_sv2v_reg  <= data_i[7];
      \nz.mem_126_sv2v_reg  <= data_i[6];
      \nz.mem_125_sv2v_reg  <= data_i[5];
      \nz.mem_124_sv2v_reg  <= data_i[4];
      \nz.mem_123_sv2v_reg  <= data_i[3];
      \nz.mem_122_sv2v_reg  <= data_i[2];
      \nz.mem_121_sv2v_reg  <= data_i[1];
      \nz.mem_120_sv2v_reg  <= data_i[0];
    end 
    if(N805) begin
      \nz.mem_119_sv2v_reg  <= data_i[7];
      \nz.mem_118_sv2v_reg  <= data_i[6];
      \nz.mem_117_sv2v_reg  <= data_i[5];
      \nz.mem_116_sv2v_reg  <= data_i[4];
      \nz.mem_115_sv2v_reg  <= data_i[3];
      \nz.mem_114_sv2v_reg  <= data_i[2];
      \nz.mem_113_sv2v_reg  <= data_i[1];
      \nz.mem_112_sv2v_reg  <= data_i[0];
    end 
    if(N804) begin
      \nz.mem_111_sv2v_reg  <= data_i[7];
      \nz.mem_110_sv2v_reg  <= data_i[6];
      \nz.mem_109_sv2v_reg  <= data_i[5];
      \nz.mem_108_sv2v_reg  <= data_i[4];
      \nz.mem_107_sv2v_reg  <= data_i[3];
      \nz.mem_106_sv2v_reg  <= data_i[2];
      \nz.mem_105_sv2v_reg  <= data_i[1];
      \nz.mem_104_sv2v_reg  <= data_i[0];
    end 
    if(N803) begin
      \nz.mem_103_sv2v_reg  <= data_i[7];
      \nz.mem_102_sv2v_reg  <= data_i[6];
      \nz.mem_101_sv2v_reg  <= data_i[5];
      \nz.mem_100_sv2v_reg  <= data_i[4];
      \nz.mem_99_sv2v_reg  <= data_i[3];
      \nz.mem_98_sv2v_reg  <= data_i[2];
      \nz.mem_97_sv2v_reg  <= data_i[1];
      \nz.mem_96_sv2v_reg  <= data_i[0];
    end 
    if(N802) begin
      \nz.mem_95_sv2v_reg  <= data_i[7];
      \nz.mem_94_sv2v_reg  <= data_i[6];
      \nz.mem_93_sv2v_reg  <= data_i[5];
      \nz.mem_92_sv2v_reg  <= data_i[4];
      \nz.mem_91_sv2v_reg  <= data_i[3];
      \nz.mem_90_sv2v_reg  <= data_i[2];
      \nz.mem_89_sv2v_reg  <= data_i[1];
      \nz.mem_88_sv2v_reg  <= data_i[0];
    end 
    if(N801) begin
      \nz.mem_87_sv2v_reg  <= data_i[7];
      \nz.mem_86_sv2v_reg  <= data_i[6];
      \nz.mem_85_sv2v_reg  <= data_i[5];
      \nz.mem_84_sv2v_reg  <= data_i[4];
      \nz.mem_83_sv2v_reg  <= data_i[3];
      \nz.mem_82_sv2v_reg  <= data_i[2];
      \nz.mem_81_sv2v_reg  <= data_i[1];
      \nz.mem_80_sv2v_reg  <= data_i[0];
    end 
    if(N800) begin
      \nz.mem_79_sv2v_reg  <= data_i[7];
      \nz.mem_78_sv2v_reg  <= data_i[6];
      \nz.mem_77_sv2v_reg  <= data_i[5];
      \nz.mem_76_sv2v_reg  <= data_i[4];
      \nz.mem_75_sv2v_reg  <= data_i[3];
      \nz.mem_74_sv2v_reg  <= data_i[2];
      \nz.mem_73_sv2v_reg  <= data_i[1];
      \nz.mem_72_sv2v_reg  <= data_i[0];
    end 
    if(N799) begin
      \nz.mem_71_sv2v_reg  <= data_i[7];
      \nz.mem_70_sv2v_reg  <= data_i[6];
      \nz.mem_69_sv2v_reg  <= data_i[5];
      \nz.mem_68_sv2v_reg  <= data_i[4];
      \nz.mem_67_sv2v_reg  <= data_i[3];
      \nz.mem_66_sv2v_reg  <= data_i[2];
      \nz.mem_65_sv2v_reg  <= data_i[1];
      \nz.mem_64_sv2v_reg  <= data_i[0];
    end 
    if(N798) begin
      \nz.mem_63_sv2v_reg  <= data_i[7];
      \nz.mem_62_sv2v_reg  <= data_i[6];
      \nz.mem_61_sv2v_reg  <= data_i[5];
      \nz.mem_60_sv2v_reg  <= data_i[4];
      \nz.mem_59_sv2v_reg  <= data_i[3];
      \nz.mem_58_sv2v_reg  <= data_i[2];
      \nz.mem_57_sv2v_reg  <= data_i[1];
      \nz.mem_56_sv2v_reg  <= data_i[0];
    end 
    if(N797) begin
      \nz.mem_55_sv2v_reg  <= data_i[7];
      \nz.mem_54_sv2v_reg  <= data_i[6];
      \nz.mem_53_sv2v_reg  <= data_i[5];
      \nz.mem_52_sv2v_reg  <= data_i[4];
      \nz.mem_51_sv2v_reg  <= data_i[3];
      \nz.mem_50_sv2v_reg  <= data_i[2];
      \nz.mem_49_sv2v_reg  <= data_i[1];
      \nz.mem_48_sv2v_reg  <= data_i[0];
    end 
    if(N796) begin
      \nz.mem_47_sv2v_reg  <= data_i[7];
      \nz.mem_46_sv2v_reg  <= data_i[6];
      \nz.mem_45_sv2v_reg  <= data_i[5];
      \nz.mem_44_sv2v_reg  <= data_i[4];
      \nz.mem_43_sv2v_reg  <= data_i[3];
      \nz.mem_42_sv2v_reg  <= data_i[2];
      \nz.mem_41_sv2v_reg  <= data_i[1];
      \nz.mem_40_sv2v_reg  <= data_i[0];
    end 
    if(N795) begin
      \nz.mem_39_sv2v_reg  <= data_i[7];
      \nz.mem_38_sv2v_reg  <= data_i[6];
      \nz.mem_37_sv2v_reg  <= data_i[5];
      \nz.mem_36_sv2v_reg  <= data_i[4];
      \nz.mem_35_sv2v_reg  <= data_i[3];
      \nz.mem_34_sv2v_reg  <= data_i[2];
      \nz.mem_33_sv2v_reg  <= data_i[1];
      \nz.mem_32_sv2v_reg  <= data_i[0];
    end 
    if(N794) begin
      \nz.mem_31_sv2v_reg  <= data_i[7];
      \nz.mem_30_sv2v_reg  <= data_i[6];
      \nz.mem_29_sv2v_reg  <= data_i[5];
      \nz.mem_28_sv2v_reg  <= data_i[4];
      \nz.mem_27_sv2v_reg  <= data_i[3];
      \nz.mem_26_sv2v_reg  <= data_i[2];
      \nz.mem_25_sv2v_reg  <= data_i[1];
      \nz.mem_24_sv2v_reg  <= data_i[0];
    end 
    if(N793) begin
      \nz.mem_23_sv2v_reg  <= data_i[7];
      \nz.mem_22_sv2v_reg  <= data_i[6];
      \nz.mem_21_sv2v_reg  <= data_i[5];
      \nz.mem_20_sv2v_reg  <= data_i[4];
      \nz.mem_19_sv2v_reg  <= data_i[3];
      \nz.mem_18_sv2v_reg  <= data_i[2];
      \nz.mem_17_sv2v_reg  <= data_i[1];
      \nz.mem_16_sv2v_reg  <= data_i[0];
    end 
    if(N792) begin
      \nz.mem_15_sv2v_reg  <= data_i[7];
      \nz.mem_14_sv2v_reg  <= data_i[6];
      \nz.mem_13_sv2v_reg  <= data_i[5];
      \nz.mem_12_sv2v_reg  <= data_i[4];
      \nz.mem_11_sv2v_reg  <= data_i[3];
      \nz.mem_10_sv2v_reg  <= data_i[2];
      \nz.mem_9_sv2v_reg  <= data_i[1];
      \nz.mem_8_sv2v_reg  <= data_i[0];
    end 
    if(N791) begin
      \nz.mem_7_sv2v_reg  <= data_i[7];
      \nz.mem_6_sv2v_reg  <= data_i[6];
      \nz.mem_5_sv2v_reg  <= data_i[5];
      \nz.mem_4_sv2v_reg  <= data_i[4];
      \nz.mem_3_sv2v_reg  <= data_i[3];
      \nz.mem_2_sv2v_reg  <= data_i[2];
      \nz.mem_1_sv2v_reg  <= data_i[1];
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [7:0] data_o;

  bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1_verbose_p0
  synth
  (
    .clk_i(clk_i),
    .v_i(v_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p128
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [127:0] data_i;
  input [15:0] write_mask_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [127:0] data_o;
  wire N0,N1,_0_net__0_,_1_net_,N2,N3,_2_net__0_,_3_net_,N4,_4_net__0_,_5_net_,N5,
  _6_net__0_,_7_net_,N6,_8_net__0_,_9_net_,N7,_10_net__0_,_11_net_,N8,_12_net__0_,
  _13_net_,N9,_14_net__0_,_15_net_,N10,_16_net__0_,_17_net_,N11,_18_net__0_,_19_net_,
  N12,_20_net__0_,_21_net_,N13,_22_net__0_,_23_net_,N14,_24_net__0_,_25_net_,N15,
  _26_net__0_,_27_net_,N16,_28_net__0_,_29_net_,N17,_30_net__0_,_31_net_,N18;

  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_0_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[7:0]),
    .addr_i(addr_i),
    .v_i(_0_net__0_),
    .w_i(_1_net_),
    .data_o(data_o[7:0])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_1_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[15:8]),
    .addr_i(addr_i),
    .v_i(_2_net__0_),
    .w_i(_3_net_),
    .data_o(data_o[15:8])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_2_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[23:16]),
    .addr_i(addr_i),
    .v_i(_4_net__0_),
    .w_i(_5_net_),
    .data_o(data_o[23:16])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_3_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[31:24]),
    .addr_i(addr_i),
    .v_i(_6_net__0_),
    .w_i(_7_net_),
    .data_o(data_o[31:24])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_4_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[39:32]),
    .addr_i(addr_i),
    .v_i(_8_net__0_),
    .w_i(_9_net_),
    .data_o(data_o[39:32])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_5_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[47:40]),
    .addr_i(addr_i),
    .v_i(_10_net__0_),
    .w_i(_11_net_),
    .data_o(data_o[47:40])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_6_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[55:48]),
    .addr_i(addr_i),
    .v_i(_12_net__0_),
    .w_i(_13_net_),
    .data_o(data_o[55:48])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_7_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[63:56]),
    .addr_i(addr_i),
    .v_i(_14_net__0_),
    .w_i(_15_net_),
    .data_o(data_o[63:56])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_8_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[71:64]),
    .addr_i(addr_i),
    .v_i(_16_net__0_),
    .w_i(_17_net_),
    .data_o(data_o[71:64])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_9_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[79:72]),
    .addr_i(addr_i),
    .v_i(_18_net__0_),
    .w_i(_19_net_),
    .data_o(data_o[79:72])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_10_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[87:80]),
    .addr_i(addr_i),
    .v_i(_20_net__0_),
    .w_i(_21_net_),
    .data_o(data_o[87:80])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_11_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[95:88]),
    .addr_i(addr_i),
    .v_i(_22_net__0_),
    .w_i(_23_net_),
    .data_o(data_o[95:88])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_12_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[103:96]),
    .addr_i(addr_i),
    .v_i(_24_net__0_),
    .w_i(_25_net_),
    .data_o(data_o[103:96])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_13_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[111:104]),
    .addr_i(addr_i),
    .v_i(_26_net__0_),
    .w_i(_27_net_),
    .data_o(data_o[111:104])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_14_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[119:112]),
    .addr_i(addr_i),
    .v_i(_28_net__0_),
    .w_i(_29_net_),
    .data_o(data_o[119:112])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_15_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[127:120]),
    .addr_i(addr_i),
    .v_i(_30_net__0_),
    .w_i(_31_net_),
    .data_o(data_o[127:120])
  );

  assign N3 = (N0)? write_mask_i[0] : 
              (N1)? 1'b1 : 1'b0;
  assign N0 = w_i;
  assign N1 = N2;
  assign N4 = (N0)? write_mask_i[1] : 
              (N1)? 1'b1 : 1'b0;
  assign N5 = (N0)? write_mask_i[2] : 
              (N1)? 1'b1 : 1'b0;
  assign N6 = (N0)? write_mask_i[3] : 
              (N1)? 1'b1 : 1'b0;
  assign N7 = (N0)? write_mask_i[4] : 
              (N1)? 1'b1 : 1'b0;
  assign N8 = (N0)? write_mask_i[5] : 
              (N1)? 1'b1 : 1'b0;
  assign N9 = (N0)? write_mask_i[6] : 
              (N1)? 1'b1 : 1'b0;
  assign N10 = (N0)? write_mask_i[7] : 
               (N1)? 1'b1 : 1'b0;
  assign N11 = (N0)? write_mask_i[8] : 
               (N1)? 1'b1 : 1'b0;
  assign N12 = (N0)? write_mask_i[9] : 
               (N1)? 1'b1 : 1'b0;
  assign N13 = (N0)? write_mask_i[10] : 
               (N1)? 1'b1 : 1'b0;
  assign N14 = (N0)? write_mask_i[11] : 
               (N1)? 1'b1 : 1'b0;
  assign N15 = (N0)? write_mask_i[12] : 
               (N1)? 1'b1 : 1'b0;
  assign N16 = (N0)? write_mask_i[13] : 
               (N1)? 1'b1 : 1'b0;
  assign N17 = (N0)? write_mask_i[14] : 
               (N1)? 1'b1 : 1'b0;
  assign N18 = (N0)? write_mask_i[15] : 
               (N1)? 1'b1 : 1'b0;
  assign _1_net_ = w_i & write_mask_i[0];
  assign N2 = ~w_i;
  assign _0_net__0_ = v_i & N3;
  assign _3_net_ = w_i & write_mask_i[1];
  assign _2_net__0_ = v_i & N4;
  assign _5_net_ = w_i & write_mask_i[2];
  assign _4_net__0_ = v_i & N5;
  assign _7_net_ = w_i & write_mask_i[3];
  assign _6_net__0_ = v_i & N6;
  assign _9_net_ = w_i & write_mask_i[4];
  assign _8_net__0_ = v_i & N7;
  assign _11_net_ = w_i & write_mask_i[5];
  assign _10_net__0_ = v_i & N8;
  assign _13_net_ = w_i & write_mask_i[6];
  assign _12_net__0_ = v_i & N9;
  assign _15_net_ = w_i & write_mask_i[7];
  assign _14_net__0_ = v_i & N10;
  assign _17_net_ = w_i & write_mask_i[8];
  assign _16_net__0_ = v_i & N11;
  assign _19_net_ = w_i & write_mask_i[9];
  assign _18_net__0_ = v_i & N12;
  assign _21_net_ = w_i & write_mask_i[10];
  assign _20_net__0_ = v_i & N13;
  assign _23_net_ = w_i & write_mask_i[11];
  assign _22_net__0_ = v_i & N14;
  assign _25_net_ = w_i & write_mask_i[12];
  assign _24_net__0_ = v_i & N15;
  assign _27_net_ = w_i & write_mask_i[13];
  assign _26_net__0_ = v_i & N16;
  assign _29_net_ = w_i & write_mask_i[14];
  assign _28_net__0_ = v_i & N17;
  assign _31_net_ = w_i & write_mask_i[15];
  assign _30_net__0_ = v_i & N18;

endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p128_latch_last_read_p1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [127:0] data_i;
  input [15:0] write_mask_i;
  output [127:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [127:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p128
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_en_width_p16_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [15:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input en_i;
  wire [15:0] data_o;
  reg data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,
  data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,
  data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p16
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [15:0] data_i;
  output [15:0] data_o;
  input clk_i;
  input en_i;
  wire [15:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p16_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p16_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [15:0] data_i;
  input [5:0] addr_i;
  input [15:0] w_mask_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [15:0] data_o,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,\nz.read_en ,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,\nz.llr.read_en_r ,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,
  N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,
  N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,
  N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,
  N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,
  N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,
  N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,
  N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
  N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,
  N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,
  N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
  N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,
  N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,
  N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
  N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,
  N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,
  N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
  N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,
  N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,
  N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
  N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,
  N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,
  N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
  N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,
  N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,
  N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
  N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,
  N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,
  N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
  N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,
  N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,
  N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
  N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,
  N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,
  N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
  N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,
  N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,
  N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
  N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,
  N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,
  N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
  N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,
  N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,
  N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
  N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,
  N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,
  N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
  N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,
  N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,
  N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
  N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,
  N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,
  N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
  N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,
  N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,
  N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
  N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,
  N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,
  N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
  N2419,N2420,N2421;
  wire [5:0] \nz.addr_r ;
  wire [1023:0] \nz.mem ;
  reg \nz.addr_r_5_sv2v_reg ,\nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,
  \nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,
  \nz.mem_1023_sv2v_reg ,\nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,
  \nz.mem_1016_sv2v_reg ,\nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,
  \nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,
  \nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,
  \nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,
  \nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,
  \nz.mem_984_sv2v_reg ,\nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,
  \nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,
  \nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,
  \nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,
  \nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,
  \nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,
  \nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,
  \nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,
  \nz.mem_944_sv2v_reg ,\nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,
  \nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,
  \nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,
  \nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,
  \nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,
  \nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,
  \nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,
  \nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,
  \nz.mem_904_sv2v_reg ,\nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,
  \nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,
  \nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,
  \nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,
  \nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,
  \nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,
  \nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,
  \nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,
  \nz.mem_864_sv2v_reg ,\nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,
  \nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,
  \nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,
  \nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,
  \nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,
  \nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,
  \nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,
  \nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,
  \nz.mem_824_sv2v_reg ,\nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,
  \nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,
  \nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,
  \nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,
  \nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,
  \nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,
  \nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,
  \nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,
  \nz.mem_784_sv2v_reg ,\nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,
  \nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,
  \nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,
  \nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,
  \nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,
  \nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,
  \nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,
  \nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,
  \nz.mem_744_sv2v_reg ,\nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,
  \nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,
  \nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,
  \nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,
  \nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,
  \nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,
  \nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,
  \nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,
  \nz.mem_704_sv2v_reg ,\nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,
  \nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,
  \nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,
  \nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,
  \nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,
  \nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,
  \nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,
  \nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,
  \nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,
  \nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,
  \nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,
  \nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,
  \nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,
  \nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,
  \nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,
  \nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,
  \nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,
  \nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,
  \nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,
  \nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,
  \nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,
  \nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,
  \nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,
  \nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,
  \nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,
  \nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,
  \nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,
  \nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,
  \nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,
  \nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,
  \nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,
  \nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,
  \nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,
  \nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,
  \nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,
  \nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,
  \nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,
  \nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,
  \nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,
  \nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,
  \nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,
  \nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,
  \nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,
  \nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,
  \nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,
  \nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,
  \nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,
  \nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,
  \nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,
  \nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,
  \nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,
  \nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,
  \nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,
  \nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,
  \nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,
  \nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,
  \nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,
  \nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,
  \nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,
  \nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,
  \nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,
  \nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,
  \nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,
  \nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,
  \nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,
  \nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,
  \nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,
  \nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,
  \nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,
  \nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,
  \nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,
  \nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,
  \nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,
  \nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,
  \nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,
  \nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,
  \nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,
  \nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,
  \nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,
  \nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,
  \nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,
  \nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,
  \nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,
  \nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,
  \nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,
  \nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,
  \nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,
  \nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,
  \nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,
  \nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,
  \nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,
  \nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [15] = (N91)? \nz.mem [15] : 
                             (N93)? \nz.mem [31] : 
                             (N95)? \nz.mem [47] : 
                             (N97)? \nz.mem [63] : 
                             (N99)? \nz.mem [79] : 
                             (N101)? \nz.mem [95] : 
                             (N103)? \nz.mem [111] : 
                             (N105)? \nz.mem [127] : 
                             (N107)? \nz.mem [143] : 
                             (N109)? \nz.mem [159] : 
                             (N111)? \nz.mem [175] : 
                             (N113)? \nz.mem [191] : 
                             (N115)? \nz.mem [207] : 
                             (N117)? \nz.mem [223] : 
                             (N119)? \nz.mem [239] : 
                             (N121)? \nz.mem [255] : 
                             (N123)? \nz.mem [271] : 
                             (N125)? \nz.mem [287] : 
                             (N127)? \nz.mem [303] : 
                             (N129)? \nz.mem [319] : 
                             (N131)? \nz.mem [335] : 
                             (N133)? \nz.mem [351] : 
                             (N135)? \nz.mem [367] : 
                             (N137)? \nz.mem [383] : 
                             (N139)? \nz.mem [399] : 
                             (N141)? \nz.mem [415] : 
                             (N143)? \nz.mem [431] : 
                             (N145)? \nz.mem [447] : 
                             (N147)? \nz.mem [463] : 
                             (N149)? \nz.mem [479] : 
                             (N151)? \nz.mem [495] : 
                             (N153)? \nz.mem [511] : 
                             (N92)? \nz.mem [527] : 
                             (N94)? \nz.mem [543] : 
                             (N96)? \nz.mem [559] : 
                             (N98)? \nz.mem [575] : 
                             (N100)? \nz.mem [591] : 
                             (N102)? \nz.mem [607] : 
                             (N104)? \nz.mem [623] : 
                             (N106)? \nz.mem [639] : 
                             (N108)? \nz.mem [655] : 
                             (N110)? \nz.mem [671] : 
                             (N112)? \nz.mem [687] : 
                             (N114)? \nz.mem [703] : 
                             (N116)? \nz.mem [719] : 
                             (N118)? \nz.mem [735] : 
                             (N120)? \nz.mem [751] : 
                             (N122)? \nz.mem [767] : 
                             (N124)? \nz.mem [783] : 
                             (N126)? \nz.mem [799] : 
                             (N128)? \nz.mem [815] : 
                             (N130)? \nz.mem [831] : 
                             (N132)? \nz.mem [847] : 
                             (N134)? \nz.mem [863] : 
                             (N136)? \nz.mem [879] : 
                             (N138)? \nz.mem [895] : 
                             (N140)? \nz.mem [911] : 
                             (N142)? \nz.mem [927] : 
                             (N144)? \nz.mem [943] : 
                             (N146)? \nz.mem [959] : 
                             (N148)? \nz.mem [975] : 
                             (N150)? \nz.mem [991] : 
                             (N152)? \nz.mem [1007] : 
                             (N154)? \nz.mem [1023] : 1'b0;
  assign \nz.data_out [14] = (N91)? \nz.mem [14] : 
                             (N93)? \nz.mem [30] : 
                             (N95)? \nz.mem [46] : 
                             (N97)? \nz.mem [62] : 
                             (N99)? \nz.mem [78] : 
                             (N101)? \nz.mem [94] : 
                             (N103)? \nz.mem [110] : 
                             (N105)? \nz.mem [126] : 
                             (N107)? \nz.mem [142] : 
                             (N109)? \nz.mem [158] : 
                             (N111)? \nz.mem [174] : 
                             (N113)? \nz.mem [190] : 
                             (N115)? \nz.mem [206] : 
                             (N117)? \nz.mem [222] : 
                             (N119)? \nz.mem [238] : 
                             (N121)? \nz.mem [254] : 
                             (N123)? \nz.mem [270] : 
                             (N125)? \nz.mem [286] : 
                             (N127)? \nz.mem [302] : 
                             (N129)? \nz.mem [318] : 
                             (N131)? \nz.mem [334] : 
                             (N133)? \nz.mem [350] : 
                             (N135)? \nz.mem [366] : 
                             (N137)? \nz.mem [382] : 
                             (N139)? \nz.mem [398] : 
                             (N141)? \nz.mem [414] : 
                             (N143)? \nz.mem [430] : 
                             (N145)? \nz.mem [446] : 
                             (N147)? \nz.mem [462] : 
                             (N149)? \nz.mem [478] : 
                             (N151)? \nz.mem [494] : 
                             (N153)? \nz.mem [510] : 
                             (N92)? \nz.mem [526] : 
                             (N94)? \nz.mem [542] : 
                             (N96)? \nz.mem [558] : 
                             (N98)? \nz.mem [574] : 
                             (N100)? \nz.mem [590] : 
                             (N102)? \nz.mem [606] : 
                             (N104)? \nz.mem [622] : 
                             (N106)? \nz.mem [638] : 
                             (N108)? \nz.mem [654] : 
                             (N110)? \nz.mem [670] : 
                             (N112)? \nz.mem [686] : 
                             (N114)? \nz.mem [702] : 
                             (N116)? \nz.mem [718] : 
                             (N118)? \nz.mem [734] : 
                             (N120)? \nz.mem [750] : 
                             (N122)? \nz.mem [766] : 
                             (N124)? \nz.mem [782] : 
                             (N126)? \nz.mem [798] : 
                             (N128)? \nz.mem [814] : 
                             (N130)? \nz.mem [830] : 
                             (N132)? \nz.mem [846] : 
                             (N134)? \nz.mem [862] : 
                             (N136)? \nz.mem [878] : 
                             (N138)? \nz.mem [894] : 
                             (N140)? \nz.mem [910] : 
                             (N142)? \nz.mem [926] : 
                             (N144)? \nz.mem [942] : 
                             (N146)? \nz.mem [958] : 
                             (N148)? \nz.mem [974] : 
                             (N150)? \nz.mem [990] : 
                             (N152)? \nz.mem [1006] : 
                             (N154)? \nz.mem [1022] : 1'b0;
  assign \nz.data_out [13] = (N91)? \nz.mem [13] : 
                             (N93)? \nz.mem [29] : 
                             (N95)? \nz.mem [45] : 
                             (N97)? \nz.mem [61] : 
                             (N99)? \nz.mem [77] : 
                             (N101)? \nz.mem [93] : 
                             (N103)? \nz.mem [109] : 
                             (N105)? \nz.mem [125] : 
                             (N107)? \nz.mem [141] : 
                             (N109)? \nz.mem [157] : 
                             (N111)? \nz.mem [173] : 
                             (N113)? \nz.mem [189] : 
                             (N115)? \nz.mem [205] : 
                             (N117)? \nz.mem [221] : 
                             (N119)? \nz.mem [237] : 
                             (N121)? \nz.mem [253] : 
                             (N123)? \nz.mem [269] : 
                             (N125)? \nz.mem [285] : 
                             (N127)? \nz.mem [301] : 
                             (N129)? \nz.mem [317] : 
                             (N131)? \nz.mem [333] : 
                             (N133)? \nz.mem [349] : 
                             (N135)? \nz.mem [365] : 
                             (N137)? \nz.mem [381] : 
                             (N139)? \nz.mem [397] : 
                             (N141)? \nz.mem [413] : 
                             (N143)? \nz.mem [429] : 
                             (N145)? \nz.mem [445] : 
                             (N147)? \nz.mem [461] : 
                             (N149)? \nz.mem [477] : 
                             (N151)? \nz.mem [493] : 
                             (N153)? \nz.mem [509] : 
                             (N92)? \nz.mem [525] : 
                             (N94)? \nz.mem [541] : 
                             (N96)? \nz.mem [557] : 
                             (N98)? \nz.mem [573] : 
                             (N100)? \nz.mem [589] : 
                             (N102)? \nz.mem [605] : 
                             (N104)? \nz.mem [621] : 
                             (N106)? \nz.mem [637] : 
                             (N108)? \nz.mem [653] : 
                             (N110)? \nz.mem [669] : 
                             (N112)? \nz.mem [685] : 
                             (N114)? \nz.mem [701] : 
                             (N116)? \nz.mem [717] : 
                             (N118)? \nz.mem [733] : 
                             (N120)? \nz.mem [749] : 
                             (N122)? \nz.mem [765] : 
                             (N124)? \nz.mem [781] : 
                             (N126)? \nz.mem [797] : 
                             (N128)? \nz.mem [813] : 
                             (N130)? \nz.mem [829] : 
                             (N132)? \nz.mem [845] : 
                             (N134)? \nz.mem [861] : 
                             (N136)? \nz.mem [877] : 
                             (N138)? \nz.mem [893] : 
                             (N140)? \nz.mem [909] : 
                             (N142)? \nz.mem [925] : 
                             (N144)? \nz.mem [941] : 
                             (N146)? \nz.mem [957] : 
                             (N148)? \nz.mem [973] : 
                             (N150)? \nz.mem [989] : 
                             (N152)? \nz.mem [1005] : 
                             (N154)? \nz.mem [1021] : 1'b0;
  assign \nz.data_out [12] = (N91)? \nz.mem [12] : 
                             (N93)? \nz.mem [28] : 
                             (N95)? \nz.mem [44] : 
                             (N97)? \nz.mem [60] : 
                             (N99)? \nz.mem [76] : 
                             (N101)? \nz.mem [92] : 
                             (N103)? \nz.mem [108] : 
                             (N105)? \nz.mem [124] : 
                             (N107)? \nz.mem [140] : 
                             (N109)? \nz.mem [156] : 
                             (N111)? \nz.mem [172] : 
                             (N113)? \nz.mem [188] : 
                             (N115)? \nz.mem [204] : 
                             (N117)? \nz.mem [220] : 
                             (N119)? \nz.mem [236] : 
                             (N121)? \nz.mem [252] : 
                             (N123)? \nz.mem [268] : 
                             (N125)? \nz.mem [284] : 
                             (N127)? \nz.mem [300] : 
                             (N129)? \nz.mem [316] : 
                             (N131)? \nz.mem [332] : 
                             (N133)? \nz.mem [348] : 
                             (N135)? \nz.mem [364] : 
                             (N137)? \nz.mem [380] : 
                             (N139)? \nz.mem [396] : 
                             (N141)? \nz.mem [412] : 
                             (N143)? \nz.mem [428] : 
                             (N145)? \nz.mem [444] : 
                             (N147)? \nz.mem [460] : 
                             (N149)? \nz.mem [476] : 
                             (N151)? \nz.mem [492] : 
                             (N153)? \nz.mem [508] : 
                             (N92)? \nz.mem [524] : 
                             (N94)? \nz.mem [540] : 
                             (N96)? \nz.mem [556] : 
                             (N98)? \nz.mem [572] : 
                             (N100)? \nz.mem [588] : 
                             (N102)? \nz.mem [604] : 
                             (N104)? \nz.mem [620] : 
                             (N106)? \nz.mem [636] : 
                             (N108)? \nz.mem [652] : 
                             (N110)? \nz.mem [668] : 
                             (N112)? \nz.mem [684] : 
                             (N114)? \nz.mem [700] : 
                             (N116)? \nz.mem [716] : 
                             (N118)? \nz.mem [732] : 
                             (N120)? \nz.mem [748] : 
                             (N122)? \nz.mem [764] : 
                             (N124)? \nz.mem [780] : 
                             (N126)? \nz.mem [796] : 
                             (N128)? \nz.mem [812] : 
                             (N130)? \nz.mem [828] : 
                             (N132)? \nz.mem [844] : 
                             (N134)? \nz.mem [860] : 
                             (N136)? \nz.mem [876] : 
                             (N138)? \nz.mem [892] : 
                             (N140)? \nz.mem [908] : 
                             (N142)? \nz.mem [924] : 
                             (N144)? \nz.mem [940] : 
                             (N146)? \nz.mem [956] : 
                             (N148)? \nz.mem [972] : 
                             (N150)? \nz.mem [988] : 
                             (N152)? \nz.mem [1004] : 
                             (N154)? \nz.mem [1020] : 1'b0;
  assign \nz.data_out [11] = (N91)? \nz.mem [11] : 
                             (N93)? \nz.mem [27] : 
                             (N95)? \nz.mem [43] : 
                             (N97)? \nz.mem [59] : 
                             (N99)? \nz.mem [75] : 
                             (N101)? \nz.mem [91] : 
                             (N103)? \nz.mem [107] : 
                             (N105)? \nz.mem [123] : 
                             (N107)? \nz.mem [139] : 
                             (N109)? \nz.mem [155] : 
                             (N111)? \nz.mem [171] : 
                             (N113)? \nz.mem [187] : 
                             (N115)? \nz.mem [203] : 
                             (N117)? \nz.mem [219] : 
                             (N119)? \nz.mem [235] : 
                             (N121)? \nz.mem [251] : 
                             (N123)? \nz.mem [267] : 
                             (N125)? \nz.mem [283] : 
                             (N127)? \nz.mem [299] : 
                             (N129)? \nz.mem [315] : 
                             (N131)? \nz.mem [331] : 
                             (N133)? \nz.mem [347] : 
                             (N135)? \nz.mem [363] : 
                             (N137)? \nz.mem [379] : 
                             (N139)? \nz.mem [395] : 
                             (N141)? \nz.mem [411] : 
                             (N143)? \nz.mem [427] : 
                             (N145)? \nz.mem [443] : 
                             (N147)? \nz.mem [459] : 
                             (N149)? \nz.mem [475] : 
                             (N151)? \nz.mem [491] : 
                             (N153)? \nz.mem [507] : 
                             (N92)? \nz.mem [523] : 
                             (N94)? \nz.mem [539] : 
                             (N96)? \nz.mem [555] : 
                             (N98)? \nz.mem [571] : 
                             (N100)? \nz.mem [587] : 
                             (N102)? \nz.mem [603] : 
                             (N104)? \nz.mem [619] : 
                             (N106)? \nz.mem [635] : 
                             (N108)? \nz.mem [651] : 
                             (N110)? \nz.mem [667] : 
                             (N112)? \nz.mem [683] : 
                             (N114)? \nz.mem [699] : 
                             (N116)? \nz.mem [715] : 
                             (N118)? \nz.mem [731] : 
                             (N120)? \nz.mem [747] : 
                             (N122)? \nz.mem [763] : 
                             (N124)? \nz.mem [779] : 
                             (N126)? \nz.mem [795] : 
                             (N128)? \nz.mem [811] : 
                             (N130)? \nz.mem [827] : 
                             (N132)? \nz.mem [843] : 
                             (N134)? \nz.mem [859] : 
                             (N136)? \nz.mem [875] : 
                             (N138)? \nz.mem [891] : 
                             (N140)? \nz.mem [907] : 
                             (N142)? \nz.mem [923] : 
                             (N144)? \nz.mem [939] : 
                             (N146)? \nz.mem [955] : 
                             (N148)? \nz.mem [971] : 
                             (N150)? \nz.mem [987] : 
                             (N152)? \nz.mem [1003] : 
                             (N154)? \nz.mem [1019] : 1'b0;
  assign \nz.data_out [10] = (N91)? \nz.mem [10] : 
                             (N93)? \nz.mem [26] : 
                             (N95)? \nz.mem [42] : 
                             (N97)? \nz.mem [58] : 
                             (N99)? \nz.mem [74] : 
                             (N101)? \nz.mem [90] : 
                             (N103)? \nz.mem [106] : 
                             (N105)? \nz.mem [122] : 
                             (N107)? \nz.mem [138] : 
                             (N109)? \nz.mem [154] : 
                             (N111)? \nz.mem [170] : 
                             (N113)? \nz.mem [186] : 
                             (N115)? \nz.mem [202] : 
                             (N117)? \nz.mem [218] : 
                             (N119)? \nz.mem [234] : 
                             (N121)? \nz.mem [250] : 
                             (N123)? \nz.mem [266] : 
                             (N125)? \nz.mem [282] : 
                             (N127)? \nz.mem [298] : 
                             (N129)? \nz.mem [314] : 
                             (N131)? \nz.mem [330] : 
                             (N133)? \nz.mem [346] : 
                             (N135)? \nz.mem [362] : 
                             (N137)? \nz.mem [378] : 
                             (N139)? \nz.mem [394] : 
                             (N141)? \nz.mem [410] : 
                             (N143)? \nz.mem [426] : 
                             (N145)? \nz.mem [442] : 
                             (N147)? \nz.mem [458] : 
                             (N149)? \nz.mem [474] : 
                             (N151)? \nz.mem [490] : 
                             (N153)? \nz.mem [506] : 
                             (N92)? \nz.mem [522] : 
                             (N94)? \nz.mem [538] : 
                             (N96)? \nz.mem [554] : 
                             (N98)? \nz.mem [570] : 
                             (N100)? \nz.mem [586] : 
                             (N102)? \nz.mem [602] : 
                             (N104)? \nz.mem [618] : 
                             (N106)? \nz.mem [634] : 
                             (N108)? \nz.mem [650] : 
                             (N110)? \nz.mem [666] : 
                             (N112)? \nz.mem [682] : 
                             (N114)? \nz.mem [698] : 
                             (N116)? \nz.mem [714] : 
                             (N118)? \nz.mem [730] : 
                             (N120)? \nz.mem [746] : 
                             (N122)? \nz.mem [762] : 
                             (N124)? \nz.mem [778] : 
                             (N126)? \nz.mem [794] : 
                             (N128)? \nz.mem [810] : 
                             (N130)? \nz.mem [826] : 
                             (N132)? \nz.mem [842] : 
                             (N134)? \nz.mem [858] : 
                             (N136)? \nz.mem [874] : 
                             (N138)? \nz.mem [890] : 
                             (N140)? \nz.mem [906] : 
                             (N142)? \nz.mem [922] : 
                             (N144)? \nz.mem [938] : 
                             (N146)? \nz.mem [954] : 
                             (N148)? \nz.mem [970] : 
                             (N150)? \nz.mem [986] : 
                             (N152)? \nz.mem [1002] : 
                             (N154)? \nz.mem [1018] : 1'b0;
  assign \nz.data_out [9] = (N91)? \nz.mem [9] : 
                            (N93)? \nz.mem [25] : 
                            (N95)? \nz.mem [41] : 
                            (N97)? \nz.mem [57] : 
                            (N99)? \nz.mem [73] : 
                            (N101)? \nz.mem [89] : 
                            (N103)? \nz.mem [105] : 
                            (N105)? \nz.mem [121] : 
                            (N107)? \nz.mem [137] : 
                            (N109)? \nz.mem [153] : 
                            (N111)? \nz.mem [169] : 
                            (N113)? \nz.mem [185] : 
                            (N115)? \nz.mem [201] : 
                            (N117)? \nz.mem [217] : 
                            (N119)? \nz.mem [233] : 
                            (N121)? \nz.mem [249] : 
                            (N123)? \nz.mem [265] : 
                            (N125)? \nz.mem [281] : 
                            (N127)? \nz.mem [297] : 
                            (N129)? \nz.mem [313] : 
                            (N131)? \nz.mem [329] : 
                            (N133)? \nz.mem [345] : 
                            (N135)? \nz.mem [361] : 
                            (N137)? \nz.mem [377] : 
                            (N139)? \nz.mem [393] : 
                            (N141)? \nz.mem [409] : 
                            (N143)? \nz.mem [425] : 
                            (N145)? \nz.mem [441] : 
                            (N147)? \nz.mem [457] : 
                            (N149)? \nz.mem [473] : 
                            (N151)? \nz.mem [489] : 
                            (N153)? \nz.mem [505] : 
                            (N92)? \nz.mem [521] : 
                            (N94)? \nz.mem [537] : 
                            (N96)? \nz.mem [553] : 
                            (N98)? \nz.mem [569] : 
                            (N100)? \nz.mem [585] : 
                            (N102)? \nz.mem [601] : 
                            (N104)? \nz.mem [617] : 
                            (N106)? \nz.mem [633] : 
                            (N108)? \nz.mem [649] : 
                            (N110)? \nz.mem [665] : 
                            (N112)? \nz.mem [681] : 
                            (N114)? \nz.mem [697] : 
                            (N116)? \nz.mem [713] : 
                            (N118)? \nz.mem [729] : 
                            (N120)? \nz.mem [745] : 
                            (N122)? \nz.mem [761] : 
                            (N124)? \nz.mem [777] : 
                            (N126)? \nz.mem [793] : 
                            (N128)? \nz.mem [809] : 
                            (N130)? \nz.mem [825] : 
                            (N132)? \nz.mem [841] : 
                            (N134)? \nz.mem [857] : 
                            (N136)? \nz.mem [873] : 
                            (N138)? \nz.mem [889] : 
                            (N140)? \nz.mem [905] : 
                            (N142)? \nz.mem [921] : 
                            (N144)? \nz.mem [937] : 
                            (N146)? \nz.mem [953] : 
                            (N148)? \nz.mem [969] : 
                            (N150)? \nz.mem [985] : 
                            (N152)? \nz.mem [1001] : 
                            (N154)? \nz.mem [1017] : 1'b0;
  assign \nz.data_out [8] = (N91)? \nz.mem [8] : 
                            (N93)? \nz.mem [24] : 
                            (N95)? \nz.mem [40] : 
                            (N97)? \nz.mem [56] : 
                            (N99)? \nz.mem [72] : 
                            (N101)? \nz.mem [88] : 
                            (N103)? \nz.mem [104] : 
                            (N105)? \nz.mem [120] : 
                            (N107)? \nz.mem [136] : 
                            (N109)? \nz.mem [152] : 
                            (N111)? \nz.mem [168] : 
                            (N113)? \nz.mem [184] : 
                            (N115)? \nz.mem [200] : 
                            (N117)? \nz.mem [216] : 
                            (N119)? \nz.mem [232] : 
                            (N121)? \nz.mem [248] : 
                            (N123)? \nz.mem [264] : 
                            (N125)? \nz.mem [280] : 
                            (N127)? \nz.mem [296] : 
                            (N129)? \nz.mem [312] : 
                            (N131)? \nz.mem [328] : 
                            (N133)? \nz.mem [344] : 
                            (N135)? \nz.mem [360] : 
                            (N137)? \nz.mem [376] : 
                            (N139)? \nz.mem [392] : 
                            (N141)? \nz.mem [408] : 
                            (N143)? \nz.mem [424] : 
                            (N145)? \nz.mem [440] : 
                            (N147)? \nz.mem [456] : 
                            (N149)? \nz.mem [472] : 
                            (N151)? \nz.mem [488] : 
                            (N153)? \nz.mem [504] : 
                            (N92)? \nz.mem [520] : 
                            (N94)? \nz.mem [536] : 
                            (N96)? \nz.mem [552] : 
                            (N98)? \nz.mem [568] : 
                            (N100)? \nz.mem [584] : 
                            (N102)? \nz.mem [600] : 
                            (N104)? \nz.mem [616] : 
                            (N106)? \nz.mem [632] : 
                            (N108)? \nz.mem [648] : 
                            (N110)? \nz.mem [664] : 
                            (N112)? \nz.mem [680] : 
                            (N114)? \nz.mem [696] : 
                            (N116)? \nz.mem [712] : 
                            (N118)? \nz.mem [728] : 
                            (N120)? \nz.mem [744] : 
                            (N122)? \nz.mem [760] : 
                            (N124)? \nz.mem [776] : 
                            (N126)? \nz.mem [792] : 
                            (N128)? \nz.mem [808] : 
                            (N130)? \nz.mem [824] : 
                            (N132)? \nz.mem [840] : 
                            (N134)? \nz.mem [856] : 
                            (N136)? \nz.mem [872] : 
                            (N138)? \nz.mem [888] : 
                            (N140)? \nz.mem [904] : 
                            (N142)? \nz.mem [920] : 
                            (N144)? \nz.mem [936] : 
                            (N146)? \nz.mem [952] : 
                            (N148)? \nz.mem [968] : 
                            (N150)? \nz.mem [984] : 
                            (N152)? \nz.mem [1000] : 
                            (N154)? \nz.mem [1016] : 1'b0;
  assign \nz.data_out [7] = (N91)? \nz.mem [7] : 
                            (N93)? \nz.mem [23] : 
                            (N95)? \nz.mem [39] : 
                            (N97)? \nz.mem [55] : 
                            (N99)? \nz.mem [71] : 
                            (N101)? \nz.mem [87] : 
                            (N103)? \nz.mem [103] : 
                            (N105)? \nz.mem [119] : 
                            (N107)? \nz.mem [135] : 
                            (N109)? \nz.mem [151] : 
                            (N111)? \nz.mem [167] : 
                            (N113)? \nz.mem [183] : 
                            (N115)? \nz.mem [199] : 
                            (N117)? \nz.mem [215] : 
                            (N119)? \nz.mem [231] : 
                            (N121)? \nz.mem [247] : 
                            (N123)? \nz.mem [263] : 
                            (N125)? \nz.mem [279] : 
                            (N127)? \nz.mem [295] : 
                            (N129)? \nz.mem [311] : 
                            (N131)? \nz.mem [327] : 
                            (N133)? \nz.mem [343] : 
                            (N135)? \nz.mem [359] : 
                            (N137)? \nz.mem [375] : 
                            (N139)? \nz.mem [391] : 
                            (N141)? \nz.mem [407] : 
                            (N143)? \nz.mem [423] : 
                            (N145)? \nz.mem [439] : 
                            (N147)? \nz.mem [455] : 
                            (N149)? \nz.mem [471] : 
                            (N151)? \nz.mem [487] : 
                            (N153)? \nz.mem [503] : 
                            (N92)? \nz.mem [519] : 
                            (N94)? \nz.mem [535] : 
                            (N96)? \nz.mem [551] : 
                            (N98)? \nz.mem [567] : 
                            (N100)? \nz.mem [583] : 
                            (N102)? \nz.mem [599] : 
                            (N104)? \nz.mem [615] : 
                            (N106)? \nz.mem [631] : 
                            (N108)? \nz.mem [647] : 
                            (N110)? \nz.mem [663] : 
                            (N112)? \nz.mem [679] : 
                            (N114)? \nz.mem [695] : 
                            (N116)? \nz.mem [711] : 
                            (N118)? \nz.mem [727] : 
                            (N120)? \nz.mem [743] : 
                            (N122)? \nz.mem [759] : 
                            (N124)? \nz.mem [775] : 
                            (N126)? \nz.mem [791] : 
                            (N128)? \nz.mem [807] : 
                            (N130)? \nz.mem [823] : 
                            (N132)? \nz.mem [839] : 
                            (N134)? \nz.mem [855] : 
                            (N136)? \nz.mem [871] : 
                            (N138)? \nz.mem [887] : 
                            (N140)? \nz.mem [903] : 
                            (N142)? \nz.mem [919] : 
                            (N144)? \nz.mem [935] : 
                            (N146)? \nz.mem [951] : 
                            (N148)? \nz.mem [967] : 
                            (N150)? \nz.mem [983] : 
                            (N152)? \nz.mem [999] : 
                            (N154)? \nz.mem [1015] : 1'b0;
  assign \nz.data_out [6] = (N91)? \nz.mem [6] : 
                            (N93)? \nz.mem [22] : 
                            (N95)? \nz.mem [38] : 
                            (N97)? \nz.mem [54] : 
                            (N99)? \nz.mem [70] : 
                            (N101)? \nz.mem [86] : 
                            (N103)? \nz.mem [102] : 
                            (N105)? \nz.mem [118] : 
                            (N107)? \nz.mem [134] : 
                            (N109)? \nz.mem [150] : 
                            (N111)? \nz.mem [166] : 
                            (N113)? \nz.mem [182] : 
                            (N115)? \nz.mem [198] : 
                            (N117)? \nz.mem [214] : 
                            (N119)? \nz.mem [230] : 
                            (N121)? \nz.mem [246] : 
                            (N123)? \nz.mem [262] : 
                            (N125)? \nz.mem [278] : 
                            (N127)? \nz.mem [294] : 
                            (N129)? \nz.mem [310] : 
                            (N131)? \nz.mem [326] : 
                            (N133)? \nz.mem [342] : 
                            (N135)? \nz.mem [358] : 
                            (N137)? \nz.mem [374] : 
                            (N139)? \nz.mem [390] : 
                            (N141)? \nz.mem [406] : 
                            (N143)? \nz.mem [422] : 
                            (N145)? \nz.mem [438] : 
                            (N147)? \nz.mem [454] : 
                            (N149)? \nz.mem [470] : 
                            (N151)? \nz.mem [486] : 
                            (N153)? \nz.mem [502] : 
                            (N92)? \nz.mem [518] : 
                            (N94)? \nz.mem [534] : 
                            (N96)? \nz.mem [550] : 
                            (N98)? \nz.mem [566] : 
                            (N100)? \nz.mem [582] : 
                            (N102)? \nz.mem [598] : 
                            (N104)? \nz.mem [614] : 
                            (N106)? \nz.mem [630] : 
                            (N108)? \nz.mem [646] : 
                            (N110)? \nz.mem [662] : 
                            (N112)? \nz.mem [678] : 
                            (N114)? \nz.mem [694] : 
                            (N116)? \nz.mem [710] : 
                            (N118)? \nz.mem [726] : 
                            (N120)? \nz.mem [742] : 
                            (N122)? \nz.mem [758] : 
                            (N124)? \nz.mem [774] : 
                            (N126)? \nz.mem [790] : 
                            (N128)? \nz.mem [806] : 
                            (N130)? \nz.mem [822] : 
                            (N132)? \nz.mem [838] : 
                            (N134)? \nz.mem [854] : 
                            (N136)? \nz.mem [870] : 
                            (N138)? \nz.mem [886] : 
                            (N140)? \nz.mem [902] : 
                            (N142)? \nz.mem [918] : 
                            (N144)? \nz.mem [934] : 
                            (N146)? \nz.mem [950] : 
                            (N148)? \nz.mem [966] : 
                            (N150)? \nz.mem [982] : 
                            (N152)? \nz.mem [998] : 
                            (N154)? \nz.mem [1014] : 1'b0;
  assign \nz.data_out [5] = (N91)? \nz.mem [5] : 
                            (N93)? \nz.mem [21] : 
                            (N95)? \nz.mem [37] : 
                            (N97)? \nz.mem [53] : 
                            (N99)? \nz.mem [69] : 
                            (N101)? \nz.mem [85] : 
                            (N103)? \nz.mem [101] : 
                            (N105)? \nz.mem [117] : 
                            (N107)? \nz.mem [133] : 
                            (N109)? \nz.mem [149] : 
                            (N111)? \nz.mem [165] : 
                            (N113)? \nz.mem [181] : 
                            (N115)? \nz.mem [197] : 
                            (N117)? \nz.mem [213] : 
                            (N119)? \nz.mem [229] : 
                            (N121)? \nz.mem [245] : 
                            (N123)? \nz.mem [261] : 
                            (N125)? \nz.mem [277] : 
                            (N127)? \nz.mem [293] : 
                            (N129)? \nz.mem [309] : 
                            (N131)? \nz.mem [325] : 
                            (N133)? \nz.mem [341] : 
                            (N135)? \nz.mem [357] : 
                            (N137)? \nz.mem [373] : 
                            (N139)? \nz.mem [389] : 
                            (N141)? \nz.mem [405] : 
                            (N143)? \nz.mem [421] : 
                            (N145)? \nz.mem [437] : 
                            (N147)? \nz.mem [453] : 
                            (N149)? \nz.mem [469] : 
                            (N151)? \nz.mem [485] : 
                            (N153)? \nz.mem [501] : 
                            (N92)? \nz.mem [517] : 
                            (N94)? \nz.mem [533] : 
                            (N96)? \nz.mem [549] : 
                            (N98)? \nz.mem [565] : 
                            (N100)? \nz.mem [581] : 
                            (N102)? \nz.mem [597] : 
                            (N104)? \nz.mem [613] : 
                            (N106)? \nz.mem [629] : 
                            (N108)? \nz.mem [645] : 
                            (N110)? \nz.mem [661] : 
                            (N112)? \nz.mem [677] : 
                            (N114)? \nz.mem [693] : 
                            (N116)? \nz.mem [709] : 
                            (N118)? \nz.mem [725] : 
                            (N120)? \nz.mem [741] : 
                            (N122)? \nz.mem [757] : 
                            (N124)? \nz.mem [773] : 
                            (N126)? \nz.mem [789] : 
                            (N128)? \nz.mem [805] : 
                            (N130)? \nz.mem [821] : 
                            (N132)? \nz.mem [837] : 
                            (N134)? \nz.mem [853] : 
                            (N136)? \nz.mem [869] : 
                            (N138)? \nz.mem [885] : 
                            (N140)? \nz.mem [901] : 
                            (N142)? \nz.mem [917] : 
                            (N144)? \nz.mem [933] : 
                            (N146)? \nz.mem [949] : 
                            (N148)? \nz.mem [965] : 
                            (N150)? \nz.mem [981] : 
                            (N152)? \nz.mem [997] : 
                            (N154)? \nz.mem [1013] : 1'b0;
  assign \nz.data_out [4] = (N91)? \nz.mem [4] : 
                            (N93)? \nz.mem [20] : 
                            (N95)? \nz.mem [36] : 
                            (N97)? \nz.mem [52] : 
                            (N99)? \nz.mem [68] : 
                            (N101)? \nz.mem [84] : 
                            (N103)? \nz.mem [100] : 
                            (N105)? \nz.mem [116] : 
                            (N107)? \nz.mem [132] : 
                            (N109)? \nz.mem [148] : 
                            (N111)? \nz.mem [164] : 
                            (N113)? \nz.mem [180] : 
                            (N115)? \nz.mem [196] : 
                            (N117)? \nz.mem [212] : 
                            (N119)? \nz.mem [228] : 
                            (N121)? \nz.mem [244] : 
                            (N123)? \nz.mem [260] : 
                            (N125)? \nz.mem [276] : 
                            (N127)? \nz.mem [292] : 
                            (N129)? \nz.mem [308] : 
                            (N131)? \nz.mem [324] : 
                            (N133)? \nz.mem [340] : 
                            (N135)? \nz.mem [356] : 
                            (N137)? \nz.mem [372] : 
                            (N139)? \nz.mem [388] : 
                            (N141)? \nz.mem [404] : 
                            (N143)? \nz.mem [420] : 
                            (N145)? \nz.mem [436] : 
                            (N147)? \nz.mem [452] : 
                            (N149)? \nz.mem [468] : 
                            (N151)? \nz.mem [484] : 
                            (N153)? \nz.mem [500] : 
                            (N92)? \nz.mem [516] : 
                            (N94)? \nz.mem [532] : 
                            (N96)? \nz.mem [548] : 
                            (N98)? \nz.mem [564] : 
                            (N100)? \nz.mem [580] : 
                            (N102)? \nz.mem [596] : 
                            (N104)? \nz.mem [612] : 
                            (N106)? \nz.mem [628] : 
                            (N108)? \nz.mem [644] : 
                            (N110)? \nz.mem [660] : 
                            (N112)? \nz.mem [676] : 
                            (N114)? \nz.mem [692] : 
                            (N116)? \nz.mem [708] : 
                            (N118)? \nz.mem [724] : 
                            (N120)? \nz.mem [740] : 
                            (N122)? \nz.mem [756] : 
                            (N124)? \nz.mem [772] : 
                            (N126)? \nz.mem [788] : 
                            (N128)? \nz.mem [804] : 
                            (N130)? \nz.mem [820] : 
                            (N132)? \nz.mem [836] : 
                            (N134)? \nz.mem [852] : 
                            (N136)? \nz.mem [868] : 
                            (N138)? \nz.mem [884] : 
                            (N140)? \nz.mem [900] : 
                            (N142)? \nz.mem [916] : 
                            (N144)? \nz.mem [932] : 
                            (N146)? \nz.mem [948] : 
                            (N148)? \nz.mem [964] : 
                            (N150)? \nz.mem [980] : 
                            (N152)? \nz.mem [996] : 
                            (N154)? \nz.mem [1012] : 1'b0;
  assign \nz.data_out [3] = (N91)? \nz.mem [3] : 
                            (N93)? \nz.mem [19] : 
                            (N95)? \nz.mem [35] : 
                            (N97)? \nz.mem [51] : 
                            (N99)? \nz.mem [67] : 
                            (N101)? \nz.mem [83] : 
                            (N103)? \nz.mem [99] : 
                            (N105)? \nz.mem [115] : 
                            (N107)? \nz.mem [131] : 
                            (N109)? \nz.mem [147] : 
                            (N111)? \nz.mem [163] : 
                            (N113)? \nz.mem [179] : 
                            (N115)? \nz.mem [195] : 
                            (N117)? \nz.mem [211] : 
                            (N119)? \nz.mem [227] : 
                            (N121)? \nz.mem [243] : 
                            (N123)? \nz.mem [259] : 
                            (N125)? \nz.mem [275] : 
                            (N127)? \nz.mem [291] : 
                            (N129)? \nz.mem [307] : 
                            (N131)? \nz.mem [323] : 
                            (N133)? \nz.mem [339] : 
                            (N135)? \nz.mem [355] : 
                            (N137)? \nz.mem [371] : 
                            (N139)? \nz.mem [387] : 
                            (N141)? \nz.mem [403] : 
                            (N143)? \nz.mem [419] : 
                            (N145)? \nz.mem [435] : 
                            (N147)? \nz.mem [451] : 
                            (N149)? \nz.mem [467] : 
                            (N151)? \nz.mem [483] : 
                            (N153)? \nz.mem [499] : 
                            (N92)? \nz.mem [515] : 
                            (N94)? \nz.mem [531] : 
                            (N96)? \nz.mem [547] : 
                            (N98)? \nz.mem [563] : 
                            (N100)? \nz.mem [579] : 
                            (N102)? \nz.mem [595] : 
                            (N104)? \nz.mem [611] : 
                            (N106)? \nz.mem [627] : 
                            (N108)? \nz.mem [643] : 
                            (N110)? \nz.mem [659] : 
                            (N112)? \nz.mem [675] : 
                            (N114)? \nz.mem [691] : 
                            (N116)? \nz.mem [707] : 
                            (N118)? \nz.mem [723] : 
                            (N120)? \nz.mem [739] : 
                            (N122)? \nz.mem [755] : 
                            (N124)? \nz.mem [771] : 
                            (N126)? \nz.mem [787] : 
                            (N128)? \nz.mem [803] : 
                            (N130)? \nz.mem [819] : 
                            (N132)? \nz.mem [835] : 
                            (N134)? \nz.mem [851] : 
                            (N136)? \nz.mem [867] : 
                            (N138)? \nz.mem [883] : 
                            (N140)? \nz.mem [899] : 
                            (N142)? \nz.mem [915] : 
                            (N144)? \nz.mem [931] : 
                            (N146)? \nz.mem [947] : 
                            (N148)? \nz.mem [963] : 
                            (N150)? \nz.mem [979] : 
                            (N152)? \nz.mem [995] : 
                            (N154)? \nz.mem [1011] : 1'b0;
  assign \nz.data_out [2] = (N91)? \nz.mem [2] : 
                            (N93)? \nz.mem [18] : 
                            (N95)? \nz.mem [34] : 
                            (N97)? \nz.mem [50] : 
                            (N99)? \nz.mem [66] : 
                            (N101)? \nz.mem [82] : 
                            (N103)? \nz.mem [98] : 
                            (N105)? \nz.mem [114] : 
                            (N107)? \nz.mem [130] : 
                            (N109)? \nz.mem [146] : 
                            (N111)? \nz.mem [162] : 
                            (N113)? \nz.mem [178] : 
                            (N115)? \nz.mem [194] : 
                            (N117)? \nz.mem [210] : 
                            (N119)? \nz.mem [226] : 
                            (N121)? \nz.mem [242] : 
                            (N123)? \nz.mem [258] : 
                            (N125)? \nz.mem [274] : 
                            (N127)? \nz.mem [290] : 
                            (N129)? \nz.mem [306] : 
                            (N131)? \nz.mem [322] : 
                            (N133)? \nz.mem [338] : 
                            (N135)? \nz.mem [354] : 
                            (N137)? \nz.mem [370] : 
                            (N139)? \nz.mem [386] : 
                            (N141)? \nz.mem [402] : 
                            (N143)? \nz.mem [418] : 
                            (N145)? \nz.mem [434] : 
                            (N147)? \nz.mem [450] : 
                            (N149)? \nz.mem [466] : 
                            (N151)? \nz.mem [482] : 
                            (N153)? \nz.mem [498] : 
                            (N92)? \nz.mem [514] : 
                            (N94)? \nz.mem [530] : 
                            (N96)? \nz.mem [546] : 
                            (N98)? \nz.mem [562] : 
                            (N100)? \nz.mem [578] : 
                            (N102)? \nz.mem [594] : 
                            (N104)? \nz.mem [610] : 
                            (N106)? \nz.mem [626] : 
                            (N108)? \nz.mem [642] : 
                            (N110)? \nz.mem [658] : 
                            (N112)? \nz.mem [674] : 
                            (N114)? \nz.mem [690] : 
                            (N116)? \nz.mem [706] : 
                            (N118)? \nz.mem [722] : 
                            (N120)? \nz.mem [738] : 
                            (N122)? \nz.mem [754] : 
                            (N124)? \nz.mem [770] : 
                            (N126)? \nz.mem [786] : 
                            (N128)? \nz.mem [802] : 
                            (N130)? \nz.mem [818] : 
                            (N132)? \nz.mem [834] : 
                            (N134)? \nz.mem [850] : 
                            (N136)? \nz.mem [866] : 
                            (N138)? \nz.mem [882] : 
                            (N140)? \nz.mem [898] : 
                            (N142)? \nz.mem [914] : 
                            (N144)? \nz.mem [930] : 
                            (N146)? \nz.mem [946] : 
                            (N148)? \nz.mem [962] : 
                            (N150)? \nz.mem [978] : 
                            (N152)? \nz.mem [994] : 
                            (N154)? \nz.mem [1010] : 1'b0;
  assign \nz.data_out [1] = (N91)? \nz.mem [1] : 
                            (N93)? \nz.mem [17] : 
                            (N95)? \nz.mem [33] : 
                            (N97)? \nz.mem [49] : 
                            (N99)? \nz.mem [65] : 
                            (N101)? \nz.mem [81] : 
                            (N103)? \nz.mem [97] : 
                            (N105)? \nz.mem [113] : 
                            (N107)? \nz.mem [129] : 
                            (N109)? \nz.mem [145] : 
                            (N111)? \nz.mem [161] : 
                            (N113)? \nz.mem [177] : 
                            (N115)? \nz.mem [193] : 
                            (N117)? \nz.mem [209] : 
                            (N119)? \nz.mem [225] : 
                            (N121)? \nz.mem [241] : 
                            (N123)? \nz.mem [257] : 
                            (N125)? \nz.mem [273] : 
                            (N127)? \nz.mem [289] : 
                            (N129)? \nz.mem [305] : 
                            (N131)? \nz.mem [321] : 
                            (N133)? \nz.mem [337] : 
                            (N135)? \nz.mem [353] : 
                            (N137)? \nz.mem [369] : 
                            (N139)? \nz.mem [385] : 
                            (N141)? \nz.mem [401] : 
                            (N143)? \nz.mem [417] : 
                            (N145)? \nz.mem [433] : 
                            (N147)? \nz.mem [449] : 
                            (N149)? \nz.mem [465] : 
                            (N151)? \nz.mem [481] : 
                            (N153)? \nz.mem [497] : 
                            (N92)? \nz.mem [513] : 
                            (N94)? \nz.mem [529] : 
                            (N96)? \nz.mem [545] : 
                            (N98)? \nz.mem [561] : 
                            (N100)? \nz.mem [577] : 
                            (N102)? \nz.mem [593] : 
                            (N104)? \nz.mem [609] : 
                            (N106)? \nz.mem [625] : 
                            (N108)? \nz.mem [641] : 
                            (N110)? \nz.mem [657] : 
                            (N112)? \nz.mem [673] : 
                            (N114)? \nz.mem [689] : 
                            (N116)? \nz.mem [705] : 
                            (N118)? \nz.mem [721] : 
                            (N120)? \nz.mem [737] : 
                            (N122)? \nz.mem [753] : 
                            (N124)? \nz.mem [769] : 
                            (N126)? \nz.mem [785] : 
                            (N128)? \nz.mem [801] : 
                            (N130)? \nz.mem [817] : 
                            (N132)? \nz.mem [833] : 
                            (N134)? \nz.mem [849] : 
                            (N136)? \nz.mem [865] : 
                            (N138)? \nz.mem [881] : 
                            (N140)? \nz.mem [897] : 
                            (N142)? \nz.mem [913] : 
                            (N144)? \nz.mem [929] : 
                            (N146)? \nz.mem [945] : 
                            (N148)? \nz.mem [961] : 
                            (N150)? \nz.mem [977] : 
                            (N152)? \nz.mem [993] : 
                            (N154)? \nz.mem [1009] : 1'b0;
  assign \nz.data_out [0] = (N91)? \nz.mem [0] : 
                            (N93)? \nz.mem [16] : 
                            (N95)? \nz.mem [32] : 
                            (N97)? \nz.mem [48] : 
                            (N99)? \nz.mem [64] : 
                            (N101)? \nz.mem [80] : 
                            (N103)? \nz.mem [96] : 
                            (N105)? \nz.mem [112] : 
                            (N107)? \nz.mem [128] : 
                            (N109)? \nz.mem [144] : 
                            (N111)? \nz.mem [160] : 
                            (N113)? \nz.mem [176] : 
                            (N115)? \nz.mem [192] : 
                            (N117)? \nz.mem [208] : 
                            (N119)? \nz.mem [224] : 
                            (N121)? \nz.mem [240] : 
                            (N123)? \nz.mem [256] : 
                            (N125)? \nz.mem [272] : 
                            (N127)? \nz.mem [288] : 
                            (N129)? \nz.mem [304] : 
                            (N131)? \nz.mem [320] : 
                            (N133)? \nz.mem [336] : 
                            (N135)? \nz.mem [352] : 
                            (N137)? \nz.mem [368] : 
                            (N139)? \nz.mem [384] : 
                            (N141)? \nz.mem [400] : 
                            (N143)? \nz.mem [416] : 
                            (N145)? \nz.mem [432] : 
                            (N147)? \nz.mem [448] : 
                            (N149)? \nz.mem [464] : 
                            (N151)? \nz.mem [480] : 
                            (N153)? \nz.mem [496] : 
                            (N92)? \nz.mem [512] : 
                            (N94)? \nz.mem [528] : 
                            (N96)? \nz.mem [544] : 
                            (N98)? \nz.mem [560] : 
                            (N100)? \nz.mem [576] : 
                            (N102)? \nz.mem [592] : 
                            (N104)? \nz.mem [608] : 
                            (N106)? \nz.mem [624] : 
                            (N108)? \nz.mem [640] : 
                            (N110)? \nz.mem [656] : 
                            (N112)? \nz.mem [672] : 
                            (N114)? \nz.mem [688] : 
                            (N116)? \nz.mem [704] : 
                            (N118)? \nz.mem [720] : 
                            (N120)? \nz.mem [736] : 
                            (N122)? \nz.mem [752] : 
                            (N124)? \nz.mem [768] : 
                            (N126)? \nz.mem [784] : 
                            (N128)? \nz.mem [800] : 
                            (N130)? \nz.mem [816] : 
                            (N132)? \nz.mem [832] : 
                            (N134)? \nz.mem [848] : 
                            (N136)? \nz.mem [864] : 
                            (N138)? \nz.mem [880] : 
                            (N140)? \nz.mem [896] : 
                            (N142)? \nz.mem [912] : 
                            (N144)? \nz.mem [928] : 
                            (N146)? \nz.mem [944] : 
                            (N148)? \nz.mem [960] : 
                            (N150)? \nz.mem [976] : 
                            (N152)? \nz.mem [992] : 
                            (N154)? \nz.mem [1008] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p16
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N2379 = addr_i[5] & N2396;
  assign N2380 = addr_i[5] & N2397;
  assign N2381 = addr_i[5] & N2398;
  assign N2382 = addr_i[2] & N2409;
  assign N2383 = addr_i[2] & N2410;
  assign N2384 = addr_i[2] & N2411;
  assign N391 = N2379 & N2382;
  assign N390 = N2379 & N2383;
  assign N389 = N2379 & N2384;
  assign N388 = N2379 & N2416;
  assign N387 = N2379 & N2417;
  assign N386 = N2379 & N2418;
  assign N385 = N2379 & N2419;
  assign N384 = N2379 & N2420;
  assign N383 = N2380 & N2382;
  assign N382 = N2380 & N2383;
  assign N381 = N2380 & N2384;
  assign N380 = N2380 & N2416;
  assign N379 = N2380 & N2417;
  assign N378 = N2380 & N2418;
  assign N377 = N2380 & N2419;
  assign N376 = N2380 & N2420;
  assign N375 = N2381 & N2382;
  assign N374 = N2381 & N2383;
  assign N373 = N2381 & N2384;
  assign N372 = N2381 & N2416;
  assign N371 = N2381 & N2417;
  assign N370 = N2381 & N2418;
  assign N369 = N2381 & N2419;
  assign N368 = N2381 & N2420;
  assign N367 = N2403 & N2382;
  assign N366 = N2403 & N2383;
  assign N365 = N2403 & N2384;
  assign N364 = N2404 & N2382;
  assign N363 = N2404 & N2383;
  assign N362 = N2404 & N2384;
  assign N361 = N2405 & N2382;
  assign N360 = N2405 & N2383;
  assign N359 = N2405 & N2384;
  assign N358 = N2406 & N2382;
  assign N357 = N2406 & N2383;
  assign N356 = N2406 & N2384;
  assign N355 = N2407 & N2382;
  assign N354 = N2407 & N2383;
  assign N353 = N2407 & N2384;
  assign N2385 = addr_i[5] & N2399;
  assign N2386 = N2395 & N2396;
  assign N2387 = N2395 & N2397;
  assign N2388 = N2395 & N2398;
  assign N2389 = N2395 & N2399;
  assign N2390 = addr_i[2] & N2412;
  assign N2391 = N2408 & N2409;
  assign N2392 = N2408 & N2410;
  assign N2393 = N2408 & N2411;
  assign N2394 = N2408 & N2412;
  assign N1161 = N2400 & N2390;
  assign N1160 = N2400 & N2391;
  assign N1159 = N2400 & N2392;
  assign N1158 = N2400 & N2393;
  assign N1157 = N2400 & N2394;
  assign N1156 = N2401 & N2390;
  assign N1155 = N2401 & N2391;
  assign N1154 = N2401 & N2392;
  assign N1153 = N2401 & N2393;
  assign N1152 = N2401 & N2394;
  assign N1151 = N2402 & N2390;
  assign N1150 = N2402 & N2391;
  assign N1149 = N2402 & N2392;
  assign N1148 = N2402 & N2393;
  assign N1147 = N2402 & N2394;
  assign N1146 = N2385 & N2413;
  assign N1145 = N2385 & N2414;
  assign N1144 = N2385 & N2415;
  assign N1143 = N2385 & N2390;
  assign N1142 = N2385 & N2391;
  assign N1141 = N2385 & N2392;
  assign N1140 = N2385 & N2393;
  assign N1139 = N2385 & N2394;
  assign N1138 = N2386 & N2413;
  assign N1137 = N2386 & N2414;
  assign N1136 = N2386 & N2415;
  assign N1135 = N2386 & N2390;
  assign N1134 = N2386 & N2391;
  assign N1133 = N2386 & N2392;
  assign N1132 = N2386 & N2393;
  assign N1131 = N2386 & N2394;
  assign N1130 = N2387 & N2413;
  assign N1129 = N2387 & N2414;
  assign N1128 = N2387 & N2415;
  assign N1127 = N2387 & N2390;
  assign N1126 = N2387 & N2391;
  assign N1125 = N2387 & N2392;
  assign N1124 = N2387 & N2393;
  assign N1123 = N2387 & N2394;
  assign N1122 = N2388 & N2413;
  assign N1121 = N2388 & N2414;
  assign N1120 = N2388 & N2415;
  assign N1119 = N2388 & N2390;
  assign N1118 = N2388 & N2391;
  assign N1117 = N2388 & N2392;
  assign N1116 = N2388 & N2393;
  assign N1115 = N2388 & N2394;
  assign N1114 = N2389 & N2413;
  assign N1113 = N2389 & N2414;
  assign N1112 = N2389 & N2415;
  assign N1111 = N2389 & N2390;
  assign N1110 = N2389 & N2391;
  assign N1109 = N2389 & N2392;
  assign N1108 = N2389 & N2393;
  assign N1107 = N2389 & N2394;
  assign N2395 = ~addr_i[5];
  assign N2396 = addr_i[3] & addr_i[4];
  assign N2397 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N2398 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N2399 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N2400 = addr_i[5] & N2396;
  assign N2401 = addr_i[5] & N2397;
  assign N2402 = addr_i[5] & N2398;
  assign N2403 = addr_i[5] & N2399;
  assign N2404 = N2395 & N2396;
  assign N2405 = N2395 & N2397;
  assign N2406 = N2395 & N2398;
  assign N2407 = N2395 & N2399;
  assign N2408 = ~addr_i[2];
  assign N2409 = addr_i[0] & addr_i[1];
  assign N2410 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N2411 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N2412 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N2413 = addr_i[2] & N2409;
  assign N2414 = addr_i[2] & N2410;
  assign N2415 = addr_i[2] & N2411;
  assign N2416 = addr_i[2] & N2412;
  assign N2417 = N2408 & N2409;
  assign N2418 = N2408 & N2410;
  assign N2419 = N2408 & N2411;
  assign N2420 = N2408 & N2412;
  assign N1290 = N2400 & N2413;
  assign N1289 = N2400 & N2414;
  assign N1288 = N2400 & N2415;
  assign N1287 = N2400 & N2416;
  assign N1286 = N2400 & N2417;
  assign N1285 = N2400 & N2418;
  assign N1284 = N2400 & N2419;
  assign N1283 = N2400 & N2420;
  assign N1282 = N2401 & N2413;
  assign N1281 = N2401 & N2414;
  assign N1280 = N2401 & N2415;
  assign N1279 = N2401 & N2416;
  assign N1278 = N2401 & N2417;
  assign N1277 = N2401 & N2418;
  assign N1276 = N2401 & N2419;
  assign N1275 = N2401 & N2420;
  assign N1274 = N2402 & N2413;
  assign N1273 = N2402 & N2414;
  assign N1272 = N2402 & N2415;
  assign N1271 = N2402 & N2416;
  assign N1270 = N2402 & N2417;
  assign N1269 = N2402 & N2418;
  assign N1268 = N2402 & N2419;
  assign N1267 = N2402 & N2420;
  assign N1266 = N2403 & N2413;
  assign N1265 = N2403 & N2414;
  assign N1264 = N2403 & N2415;
  assign N1263 = N2403 & N2416;
  assign N1262 = N2403 & N2417;
  assign N1261 = N2403 & N2418;
  assign N1260 = N2403 & N2419;
  assign N1259 = N2403 & N2420;
  assign N1258 = N2404 & N2413;
  assign N1257 = N2404 & N2414;
  assign N1256 = N2404 & N2415;
  assign N1255 = N2404 & N2416;
  assign N1254 = N2404 & N2417;
  assign N1253 = N2404 & N2418;
  assign N1252 = N2404 & N2419;
  assign N1251 = N2404 & N2420;
  assign N1250 = N2405 & N2413;
  assign N1249 = N2405 & N2414;
  assign N1248 = N2405 & N2415;
  assign N1247 = N2405 & N2416;
  assign N1246 = N2405 & N2417;
  assign N1245 = N2405 & N2418;
  assign N1244 = N2405 & N2419;
  assign N1243 = N2405 & N2420;
  assign N1242 = N2406 & N2413;
  assign N1241 = N2406 & N2414;
  assign N1240 = N2406 & N2415;
  assign N1239 = N2406 & N2416;
  assign N1238 = N2406 & N2417;
  assign N1237 = N2406 & N2418;
  assign N1236 = N2406 & N2419;
  assign N1235 = N2406 & N2420;
  assign N1234 = N2407 & N2413;
  assign N1233 = N2407 & N2414;
  assign N1232 = N2407 & N2415;
  assign N1231 = N2407 & N2416;
  assign N1230 = N2407 & N2417;
  assign N1229 = N2407 & N2418;
  assign N1228 = N2407 & N2419;
  assign N1227 = N2407 & N2420;
  assign { N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158 } = (N8)? { N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N1263, N1262, N1261, N1260, N1259, N364, N363, N362, N1255, N1254, N1253, N1252, N1251, N361, N360, N359, N1247, N1246, N1245, N1244, N1243, N358, N357, N356, N1239, N1238, N1237, N1236, N1235, N355, N354, N353, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N157)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223 } = (N9)? { N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N1263, N1262, N1261, N1260, N1259, N364, N363, N362, N1255, N1254, N1253, N1252, N1251, N361, N360, N359, N1247, N1246, N1245, N1244, N1243, N358, N357, N356, N1239, N1238, N1237, N1236, N1235, N355, N354, N353, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N222)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288 } = (N10)? { N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N1263, N1262, N1261, N1260, N1259, N364, N363, N362, N1255, N1254, N1253, N1252, N1251, N361, N360, N359, N1247, N1246, N1245, N1244, N1243, N358, N357, N356, N1239, N1238, N1237, N1236, N1235, N355, N354, N353, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N287)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392 } = (N11)? { N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N1263, N1262, N1261, N1260, N1259, N364, N363, N362, N1255, N1254, N1253, N1252, N1251, N361, N360, N359, N1247, N1246, N1245, N1244, N1243, N358, N357, N356, N1239, N1238, N1237, N1236, N1235, N355, N354, N353, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N352)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457 } = (N12)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N456)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522 } = (N13)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N521)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587 } = (N14)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N586)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652 } = (N15)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N651)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = w_mask_i[7];
  assign { N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717 } = (N16)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N716)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[8];
  assign { N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782 } = (N17)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N781)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[9];
  assign { N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847 } = (N18)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N846)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[10];
  assign { N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912 } = (N19)? { N1290, N1289, N1288, N1161, N1160, N1159, N1158, N1157, N1282, N1281, N1280, N1156, N1155, N1154, N1153, N1152, N1274, N1273, N1272, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N911)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[11];
  assign { N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977 } = (N20)? { N1290, N1289, N1288, N1161, N1160, N1159, N1158, N1157, N1282, N1281, N1280, N1156, N1155, N1154, N1153, N1152, N1274, N1273, N1272, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                       (N976)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[12];
  assign { N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042 } = (N21)? { N1290, N1289, N1288, N1161, N1160, N1159, N1158, N1157, N1282, N1281, N1280, N1156, N1155, N1154, N1153, N1152, N1274, N1273, N1272, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1041)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[13];
  assign { N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162 } = (N22)? { N1290, N1289, N1288, N1161, N1160, N1159, N1158, N1157, N1282, N1281, N1280, N1156, N1155, N1154, N1153, N1152, N1274, N1273, N1272, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1106)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[14];
  assign { N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291 } = (N23)? { N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1226)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = w_mask_i[15];
  assign { N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355 } = (N24)? { N1354, N1225, N1105, N1040, N975, N910, N845, N780, N715, N650, N585, N520, N455, N351, N286, N221, N1353, N1224, N1104, N1039, N974, N909, N844, N779, N714, N649, N584, N519, N454, N350, N285, N220, N1352, N1223, N1103, N1038, N973, N908, N843, N778, N713, N648, N583, N518, N453, N349, N284, N219, N1351, N1222, N1102, N1037, N972, N907, N842, N777, N712, N647, N582, N517, N452, N348, N283, N218, N1350, N1221, N1101, N1036, N971, N906, N841, N776, N711, N646, N581, N516, N451, N347, N282, N217, N1349, N1220, N1100, N1035, N970, N905, N840, N775, N710, N645, N580, N515, N450, N346, N281, N216, N1348, N1219, N1099, N1034, N969, N904, N839, N774, N709, N644, N579, N514, N449, N345, N280, N215, N1347, N1218, N1098, N1033, N968, N903, N838, N773, N708, N643, N578, N513, N448, N344, N279, N214, N1346, N1217, N1097, N1032, N967, N902, N837, N772, N707, N642, N577, N512, N447, N343, N278, N213, N1345, N1216, N1096, N1031, N966, N901, N836, N771, N706, N641, N576, N511, N446, N342, N277, N212, N1344, N1215, N1095, N1030, N965, N900, N835, N770, N705, N640, N575, N510, N445, N341, N276, N211, N1343, N1214, N1094, N1029, N964, N899, N834, N769, N704, N639, N574, N509, N444, N340, N275, N210, N1342, N1213, N1093, N1028, N963, N898, N833, N768, N703, N638, N573, N508, N443, N339, N274, N209, N1341, N1212, N1092, N1027, N962, N897, N832, N767, N702, N637, N572, N507, N442, N338, N273, N208, N1340, N1211, N1091, N1026, N961, N896, N831, N766, N701, N636, N571, N506, N441, N337, N272, N207, N1339, N1210, N1090, N1025, N960, N895, N830, N765, N700, N635, N570, N505, N440, N336, N271, N206, N1338, N1209, N1089, N1024, N959, N894, N829, N764, N699, N634, N569, N504, N439, N335, N270, N205, N1337, N1208, N1088, N1023, N958, N893, N828, N763, N698, N633, N568, N503, N438, N334, N269, N204, N1336, N1207, N1087, N1022, N957, N892, N827, N762, N697, N632, N567, N502, N437, N333, N268, N203, N1335, N1206, N1086, N1021, N956, N891, N826, N761, N696, N631, N566, N501, N436, N332, N267, N202, N1334, N1205, N1085, N1020, N955, N890, N825, N760, N695, N630, N565, N500, N435, N331, N266, N201, N1333, N1204, N1084, N1019, N954, N889, N824, N759, N694, N629, N564, N499, N434, N330, N265, N200, N1332, N1203, N1083, N1018, N953, N888, N823, N758, N693, N628, N563, N498, N433, N329, N264, N199, N1331, N1202, N1082, N1017, N952, N887, N822, N757, N692, N627, N562, N497, N432, N328, N263, N198, N1330, N1201, N1081, N1016, N951, N886, N821, N756, N691, N626, N561, N496, N431, N327, N262, N197, N1329, N1200, N1080, N1015, N950, N885, N820, N755, N690, N625, N560, N495, N430, N326, N261, N196, N1328, N1199, N1079, N1014, N949, N884, N819, N754, N689, N624, N559, N494, N429, N325, N260, N195, N1327, N1198, N1078, N1013, N948, N883, N818, N753, N688, N623, N558, N493, N428, N324, N259, N194, N1326, N1197, N1077, N1012, N947, N882, N817, N752, N687, N622, N557, N492, N427, N323, N258, N193, N1325, N1196, N1076, N1011, N946, N881, N816, N751, N686, N621, N556, N491, N426, N322, N257, N192, N1324, N1195, N1075, N1010, N945, N880, N815, N750, N685, N620, N555, N490, N425, N321, N256, N191, N1323, N1194, N1074, N1009, N944, N879, N814, N749, N684, N619, N554, N489, N424, N320, N255, N190, N1322, N1193, N1073, N1008, N943, N878, N813, N748, N683, N618, N553, N488, N423, N319, N254, N189, N1321, N1192, N1072, N1007, N942, N877, N812, N747, N682, N617, N552, N487, N422, N318, N253, N188, N1320, N1191, N1071, N1006, N941, N876, N811, N746, N681, N616, N551, N486, N421, N317, N252, N187, N1319, N1190, N1070, N1005, N940, N875, N810, N745, N680, N615, N550, N485, N420, N316, N251, N186, N1318, N1189, N1069, N1004, N939, N874, N809, N744, N679, N614, N549, N484, N419, N315, N250, N185, N1317, N1188, N1068, N1003, N938, N873, N808, N743, N678, N613, N548, N483, N418, N314, N249, N184, N1316, N1187, N1067, N1002, N937, N872, N807, N742, N677, N612, N547, N482, N417, N313, N248, N183, N1315, N1186, N1066, N1001, N936, N871, N806, N741, N676, N611, N546, N481, N416, N312, N247, N182, N1314, N1185, N1065, N1000, N935, N870, N805, N740, N675, N610, N545, N480, N415, N311, N246, N181, N1313, N1184, N1064, N999, N934, N869, N804, N739, N674, N609, N544, N479, N414, N310, N245, N180, N1312, N1183, N1063, N998, N933, N868, N803, N738, N673, N608, N543, N478, N413, N309, N244, N179, N1311, N1182, N1062, N997, N932, N867, N802, N737, N672, N607, N542, N477, N412, N308, N243, N178, N1310, N1181, N1061, N996, N931, N866, N801, N736, N671, N606, N541, N476, N411, N307, N242, N177, N1309, N1180, N1060, N995, N930, N865, N800, N735, N670, N605, N540, N475, N410, N306, N241, N176, N1308, N1179, N1059, N994, N929, N864, N799, N734, N669, N604, N539, N474, N409, N305, N240, N175, N1307, N1178, N1058, N993, N928, N863, N798, N733, N668, N603, N538, N473, N408, N304, N239, N174, N1306, N1177, N1057, N992, N927, N862, N797, N732, N667, N602, N537, N472, N407, N303, N238, N173, N1305, N1176, N1056, N991, N926, N861, N796, N731, N666, N601, N536, N471, N406, N302, N237, N172, N1304, N1175, N1055, N990, N925, N860, N795, N730, N665, N600, N535, N470, N405, N301, N236, N171, N1303, N1174, N1054, N989, N924, N859, N794, N729, N664, N599, N534, N469, N404, N300, N235, N170, N1302, N1173, N1053, N988, N923, N858, N793, N728, N663, N598, N533, N468, N403, N299, N234, N169, N1301, N1172, N1052, N987, N922, N857, N792, N727, N662, N597, N532, N467, N402, N298, N233, N168, N1300, N1171, N1051, N986, N921, N856, N791, N726, N661, N596, N531, N466, N401, N297, N232, N167, N1299, N1170, N1050, N985, N920, N855, N790, N725, N660, N595, N530, N465, N400, N296, N231, N166, N1298, N1169, N1049, N984, N919, N854, N789, N724, N659, N594, N529, N464, N399, N295, N230, N165, N1297, N1168, N1048, N983, N918, N853, N788, N723, N658, N593, N528, N463, N398, N294, N229, N164, N1296, N1167, N1047, N982, N917, N852, N787, N722, N657, N592, N527, N462, N397, N293, N228, N163, N1295, N1166, N1046, N981, N916, N851, N786, N721, N656, N591, N526, N461, N396, N292, N227, N162, N1294, N1165, N1045, N980, N915, N850, N785, N720, N655, N590, N525, N460, N395, N291, N226, N161, N1293, N1164, N1044, N979, N914, N849, N784, N719, N654, N589, N524, N459, N394, N290, N225, N160, N1292, N1163, N1043, N978, N913, N848, N783, N718, N653, N588, N523, N458, N393, N289, N224, N159, N1291, N1162, N1042, N977, N912, N847, N782, N717, N652, N587, N522, N457, N392, N288, N223, N158 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N156)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N24 = N155;
  assign \nz.read_en  = v_i & N2421;
  assign N2421 = ~w_i;
  assign N25 = ~\nz.addr_r [0];
  assign N26 = ~\nz.addr_r [1];
  assign N27 = N25 & N26;
  assign N28 = N25 & \nz.addr_r [1];
  assign N29 = \nz.addr_r [0] & N26;
  assign N30 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N31 = ~\nz.addr_r [2];
  assign N32 = N27 & N31;
  assign N33 = N27 & \nz.addr_r [2];
  assign N34 = N29 & N31;
  assign N35 = N29 & \nz.addr_r [2];
  assign N36 = N28 & N31;
  assign N37 = N28 & \nz.addr_r [2];
  assign N38 = N30 & N31;
  assign N39 = N30 & \nz.addr_r [2];
  assign N40 = ~\nz.addr_r [3];
  assign N41 = N32 & N40;
  assign N42 = N32 & \nz.addr_r [3];
  assign N43 = N34 & N40;
  assign N44 = N34 & \nz.addr_r [3];
  assign N45 = N36 & N40;
  assign N46 = N36 & \nz.addr_r [3];
  assign N47 = N38 & N40;
  assign N48 = N38 & \nz.addr_r [3];
  assign N49 = N33 & N40;
  assign N50 = N33 & \nz.addr_r [3];
  assign N51 = N35 & N40;
  assign N52 = N35 & \nz.addr_r [3];
  assign N53 = N37 & N40;
  assign N54 = N37 & \nz.addr_r [3];
  assign N55 = N39 & N40;
  assign N56 = N39 & \nz.addr_r [3];
  assign N57 = ~\nz.addr_r [4];
  assign N58 = N41 & N57;
  assign N59 = N41 & \nz.addr_r [4];
  assign N60 = N43 & N57;
  assign N61 = N43 & \nz.addr_r [4];
  assign N62 = N45 & N57;
  assign N63 = N45 & \nz.addr_r [4];
  assign N64 = N47 & N57;
  assign N65 = N47 & \nz.addr_r [4];
  assign N66 = N49 & N57;
  assign N67 = N49 & \nz.addr_r [4];
  assign N68 = N51 & N57;
  assign N69 = N51 & \nz.addr_r [4];
  assign N70 = N53 & N57;
  assign N71 = N53 & \nz.addr_r [4];
  assign N72 = N55 & N57;
  assign N73 = N55 & \nz.addr_r [4];
  assign N74 = N42 & N57;
  assign N75 = N42 & \nz.addr_r [4];
  assign N76 = N44 & N57;
  assign N77 = N44 & \nz.addr_r [4];
  assign N78 = N46 & N57;
  assign N79 = N46 & \nz.addr_r [4];
  assign N80 = N48 & N57;
  assign N81 = N48 & \nz.addr_r [4];
  assign N82 = N50 & N57;
  assign N83 = N50 & \nz.addr_r [4];
  assign N84 = N52 & N57;
  assign N85 = N52 & \nz.addr_r [4];
  assign N86 = N54 & N57;
  assign N87 = N54 & \nz.addr_r [4];
  assign N88 = N56 & N57;
  assign N89 = N56 & \nz.addr_r [4];
  assign N90 = ~\nz.addr_r [5];
  assign N91 = N58 & N90;
  assign N92 = N58 & \nz.addr_r [5];
  assign N93 = N60 & N90;
  assign N94 = N60 & \nz.addr_r [5];
  assign N95 = N62 & N90;
  assign N96 = N62 & \nz.addr_r [5];
  assign N97 = N64 & N90;
  assign N98 = N64 & \nz.addr_r [5];
  assign N99 = N66 & N90;
  assign N100 = N66 & \nz.addr_r [5];
  assign N101 = N68 & N90;
  assign N102 = N68 & \nz.addr_r [5];
  assign N103 = N70 & N90;
  assign N104 = N70 & \nz.addr_r [5];
  assign N105 = N72 & N90;
  assign N106 = N72 & \nz.addr_r [5];
  assign N107 = N74 & N90;
  assign N108 = N74 & \nz.addr_r [5];
  assign N109 = N76 & N90;
  assign N110 = N76 & \nz.addr_r [5];
  assign N111 = N78 & N90;
  assign N112 = N78 & \nz.addr_r [5];
  assign N113 = N80 & N90;
  assign N114 = N80 & \nz.addr_r [5];
  assign N115 = N82 & N90;
  assign N116 = N82 & \nz.addr_r [5];
  assign N117 = N84 & N90;
  assign N118 = N84 & \nz.addr_r [5];
  assign N119 = N86 & N90;
  assign N120 = N86 & \nz.addr_r [5];
  assign N121 = N88 & N90;
  assign N122 = N88 & \nz.addr_r [5];
  assign N123 = N59 & N90;
  assign N124 = N59 & \nz.addr_r [5];
  assign N125 = N61 & N90;
  assign N126 = N61 & \nz.addr_r [5];
  assign N127 = N63 & N90;
  assign N128 = N63 & \nz.addr_r [5];
  assign N129 = N65 & N90;
  assign N130 = N65 & \nz.addr_r [5];
  assign N131 = N67 & N90;
  assign N132 = N67 & \nz.addr_r [5];
  assign N133 = N69 & N90;
  assign N134 = N69 & \nz.addr_r [5];
  assign N135 = N71 & N90;
  assign N136 = N71 & \nz.addr_r [5];
  assign N137 = N73 & N90;
  assign N138 = N73 & \nz.addr_r [5];
  assign N139 = N75 & N90;
  assign N140 = N75 & \nz.addr_r [5];
  assign N141 = N77 & N90;
  assign N142 = N77 & \nz.addr_r [5];
  assign N143 = N79 & N90;
  assign N144 = N79 & \nz.addr_r [5];
  assign N145 = N81 & N90;
  assign N146 = N81 & \nz.addr_r [5];
  assign N147 = N83 & N90;
  assign N148 = N83 & \nz.addr_r [5];
  assign N149 = N85 & N90;
  assign N150 = N85 & \nz.addr_r [5];
  assign N151 = N87 & N90;
  assign N152 = N87 & \nz.addr_r [5];
  assign N153 = N89 & N90;
  assign N154 = N89 & \nz.addr_r [5];
  assign N155 = v_i & w_i;
  assign N156 = ~N155;
  assign N157 = ~w_mask_i[0];
  assign N222 = ~w_mask_i[1];
  assign N287 = ~w_mask_i[2];
  assign N352 = ~w_mask_i[3];
  assign N456 = ~w_mask_i[4];
  assign N521 = ~w_mask_i[5];
  assign N586 = ~w_mask_i[6];
  assign N651 = ~w_mask_i[7];
  assign N716 = ~w_mask_i[8];
  assign N781 = ~w_mask_i[9];
  assign N846 = ~w_mask_i[10];
  assign N911 = ~w_mask_i[11];
  assign N976 = ~w_mask_i[12];
  assign N1041 = ~w_mask_i[13];
  assign N1106 = ~w_mask_i[14];
  assign N1226 = ~w_mask_i[15];

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N2378) begin
      \nz.mem_1023_sv2v_reg  <= data_i[15];
    end 
    if(N2377) begin
      \nz.mem_1022_sv2v_reg  <= data_i[14];
    end 
    if(N2376) begin
      \nz.mem_1021_sv2v_reg  <= data_i[13];
    end 
    if(N2375) begin
      \nz.mem_1020_sv2v_reg  <= data_i[12];
    end 
    if(N2374) begin
      \nz.mem_1019_sv2v_reg  <= data_i[11];
    end 
    if(N2373) begin
      \nz.mem_1018_sv2v_reg  <= data_i[10];
    end 
    if(N2372) begin
      \nz.mem_1017_sv2v_reg  <= data_i[9];
    end 
    if(N2371) begin
      \nz.mem_1016_sv2v_reg  <= data_i[8];
    end 
    if(N2370) begin
      \nz.mem_1015_sv2v_reg  <= data_i[7];
    end 
    if(N2369) begin
      \nz.mem_1014_sv2v_reg  <= data_i[6];
    end 
    if(N2368) begin
      \nz.mem_1013_sv2v_reg  <= data_i[5];
    end 
    if(N2367) begin
      \nz.mem_1012_sv2v_reg  <= data_i[4];
    end 
    if(N2366) begin
      \nz.mem_1011_sv2v_reg  <= data_i[3];
    end 
    if(N2365) begin
      \nz.mem_1010_sv2v_reg  <= data_i[2];
    end 
    if(N2364) begin
      \nz.mem_1009_sv2v_reg  <= data_i[1];
    end 
    if(N2363) begin
      \nz.mem_1008_sv2v_reg  <= data_i[0];
    end 
    if(N2362) begin
      \nz.mem_1007_sv2v_reg  <= data_i[15];
    end 
    if(N2361) begin
      \nz.mem_1006_sv2v_reg  <= data_i[14];
    end 
    if(N2360) begin
      \nz.mem_1005_sv2v_reg  <= data_i[13];
    end 
    if(N2359) begin
      \nz.mem_1004_sv2v_reg  <= data_i[12];
    end 
    if(N2358) begin
      \nz.mem_1003_sv2v_reg  <= data_i[11];
    end 
    if(N2357) begin
      \nz.mem_1002_sv2v_reg  <= data_i[10];
    end 
    if(N2356) begin
      \nz.mem_1001_sv2v_reg  <= data_i[9];
    end 
    if(N2355) begin
      \nz.mem_1000_sv2v_reg  <= data_i[8];
    end 
    if(N2354) begin
      \nz.mem_999_sv2v_reg  <= data_i[7];
    end 
    if(N2353) begin
      \nz.mem_998_sv2v_reg  <= data_i[6];
    end 
    if(N2352) begin
      \nz.mem_997_sv2v_reg  <= data_i[5];
    end 
    if(N2351) begin
      \nz.mem_996_sv2v_reg  <= data_i[4];
    end 
    if(N2350) begin
      \nz.mem_995_sv2v_reg  <= data_i[3];
    end 
    if(N2349) begin
      \nz.mem_994_sv2v_reg  <= data_i[2];
    end 
    if(N2348) begin
      \nz.mem_993_sv2v_reg  <= data_i[1];
    end 
    if(N2347) begin
      \nz.mem_992_sv2v_reg  <= data_i[0];
    end 
    if(N2346) begin
      \nz.mem_991_sv2v_reg  <= data_i[15];
    end 
    if(N2345) begin
      \nz.mem_990_sv2v_reg  <= data_i[14];
    end 
    if(N2344) begin
      \nz.mem_989_sv2v_reg  <= data_i[13];
    end 
    if(N2343) begin
      \nz.mem_988_sv2v_reg  <= data_i[12];
    end 
    if(N2342) begin
      \nz.mem_987_sv2v_reg  <= data_i[11];
    end 
    if(N2341) begin
      \nz.mem_986_sv2v_reg  <= data_i[10];
    end 
    if(N2340) begin
      \nz.mem_985_sv2v_reg  <= data_i[9];
    end 
    if(N2339) begin
      \nz.mem_984_sv2v_reg  <= data_i[8];
    end 
    if(N2338) begin
      \nz.mem_983_sv2v_reg  <= data_i[7];
    end 
    if(N2337) begin
      \nz.mem_982_sv2v_reg  <= data_i[6];
    end 
    if(N2336) begin
      \nz.mem_981_sv2v_reg  <= data_i[5];
    end 
    if(N2335) begin
      \nz.mem_980_sv2v_reg  <= data_i[4];
    end 
    if(N2334) begin
      \nz.mem_979_sv2v_reg  <= data_i[3];
    end 
    if(N2333) begin
      \nz.mem_978_sv2v_reg  <= data_i[2];
    end 
    if(N2332) begin
      \nz.mem_977_sv2v_reg  <= data_i[1];
    end 
    if(N2331) begin
      \nz.mem_976_sv2v_reg  <= data_i[0];
    end 
    if(N2330) begin
      \nz.mem_975_sv2v_reg  <= data_i[15];
    end 
    if(N2329) begin
      \nz.mem_974_sv2v_reg  <= data_i[14];
    end 
    if(N2328) begin
      \nz.mem_973_sv2v_reg  <= data_i[13];
    end 
    if(N2327) begin
      \nz.mem_972_sv2v_reg  <= data_i[12];
    end 
    if(N2326) begin
      \nz.mem_971_sv2v_reg  <= data_i[11];
    end 
    if(N2325) begin
      \nz.mem_970_sv2v_reg  <= data_i[10];
    end 
    if(N2324) begin
      \nz.mem_969_sv2v_reg  <= data_i[9];
    end 
    if(N2323) begin
      \nz.mem_968_sv2v_reg  <= data_i[8];
    end 
    if(N2322) begin
      \nz.mem_967_sv2v_reg  <= data_i[7];
    end 
    if(N2321) begin
      \nz.mem_966_sv2v_reg  <= data_i[6];
    end 
    if(N2320) begin
      \nz.mem_965_sv2v_reg  <= data_i[5];
    end 
    if(N2319) begin
      \nz.mem_964_sv2v_reg  <= data_i[4];
    end 
    if(N2318) begin
      \nz.mem_963_sv2v_reg  <= data_i[3];
    end 
    if(N2317) begin
      \nz.mem_962_sv2v_reg  <= data_i[2];
    end 
    if(N2316) begin
      \nz.mem_961_sv2v_reg  <= data_i[1];
    end 
    if(N2315) begin
      \nz.mem_960_sv2v_reg  <= data_i[0];
    end 
    if(N2314) begin
      \nz.mem_959_sv2v_reg  <= data_i[15];
    end 
    if(N2313) begin
      \nz.mem_958_sv2v_reg  <= data_i[14];
    end 
    if(N2312) begin
      \nz.mem_957_sv2v_reg  <= data_i[13];
    end 
    if(N2311) begin
      \nz.mem_956_sv2v_reg  <= data_i[12];
    end 
    if(N2310) begin
      \nz.mem_955_sv2v_reg  <= data_i[11];
    end 
    if(N2309) begin
      \nz.mem_954_sv2v_reg  <= data_i[10];
    end 
    if(N2308) begin
      \nz.mem_953_sv2v_reg  <= data_i[9];
    end 
    if(N2307) begin
      \nz.mem_952_sv2v_reg  <= data_i[8];
    end 
    if(N2306) begin
      \nz.mem_951_sv2v_reg  <= data_i[7];
    end 
    if(N2305) begin
      \nz.mem_950_sv2v_reg  <= data_i[6];
    end 
    if(N2304) begin
      \nz.mem_949_sv2v_reg  <= data_i[5];
    end 
    if(N2303) begin
      \nz.mem_948_sv2v_reg  <= data_i[4];
    end 
    if(N2302) begin
      \nz.mem_947_sv2v_reg  <= data_i[3];
    end 
    if(N2301) begin
      \nz.mem_946_sv2v_reg  <= data_i[2];
    end 
    if(N2300) begin
      \nz.mem_945_sv2v_reg  <= data_i[1];
    end 
    if(N2299) begin
      \nz.mem_944_sv2v_reg  <= data_i[0];
    end 
    if(N2298) begin
      \nz.mem_943_sv2v_reg  <= data_i[15];
    end 
    if(N2297) begin
      \nz.mem_942_sv2v_reg  <= data_i[14];
    end 
    if(N2296) begin
      \nz.mem_941_sv2v_reg  <= data_i[13];
    end 
    if(N2295) begin
      \nz.mem_940_sv2v_reg  <= data_i[12];
    end 
    if(N2294) begin
      \nz.mem_939_sv2v_reg  <= data_i[11];
    end 
    if(N2293) begin
      \nz.mem_938_sv2v_reg  <= data_i[10];
    end 
    if(N2292) begin
      \nz.mem_937_sv2v_reg  <= data_i[9];
    end 
    if(N2291) begin
      \nz.mem_936_sv2v_reg  <= data_i[8];
    end 
    if(N2290) begin
      \nz.mem_935_sv2v_reg  <= data_i[7];
    end 
    if(N2289) begin
      \nz.mem_934_sv2v_reg  <= data_i[6];
    end 
    if(N2288) begin
      \nz.mem_933_sv2v_reg  <= data_i[5];
    end 
    if(N2287) begin
      \nz.mem_932_sv2v_reg  <= data_i[4];
    end 
    if(N2286) begin
      \nz.mem_931_sv2v_reg  <= data_i[3];
    end 
    if(N2285) begin
      \nz.mem_930_sv2v_reg  <= data_i[2];
    end 
    if(N2284) begin
      \nz.mem_929_sv2v_reg  <= data_i[1];
    end 
    if(N2283) begin
      \nz.mem_928_sv2v_reg  <= data_i[0];
    end 
    if(N2282) begin
      \nz.mem_927_sv2v_reg  <= data_i[15];
    end 
    if(N2281) begin
      \nz.mem_926_sv2v_reg  <= data_i[14];
    end 
    if(N2280) begin
      \nz.mem_925_sv2v_reg  <= data_i[13];
    end 
    if(N2279) begin
      \nz.mem_924_sv2v_reg  <= data_i[12];
    end 
    if(N2278) begin
      \nz.mem_923_sv2v_reg  <= data_i[11];
    end 
    if(N2277) begin
      \nz.mem_922_sv2v_reg  <= data_i[10];
    end 
    if(N2276) begin
      \nz.mem_921_sv2v_reg  <= data_i[9];
    end 
    if(N2275) begin
      \nz.mem_920_sv2v_reg  <= data_i[8];
    end 
    if(N2274) begin
      \nz.mem_919_sv2v_reg  <= data_i[7];
    end 
    if(N2273) begin
      \nz.mem_918_sv2v_reg  <= data_i[6];
    end 
    if(N2272) begin
      \nz.mem_917_sv2v_reg  <= data_i[5];
    end 
    if(N2271) begin
      \nz.mem_916_sv2v_reg  <= data_i[4];
    end 
    if(N2270) begin
      \nz.mem_915_sv2v_reg  <= data_i[3];
    end 
    if(N2269) begin
      \nz.mem_914_sv2v_reg  <= data_i[2];
    end 
    if(N2268) begin
      \nz.mem_913_sv2v_reg  <= data_i[1];
    end 
    if(N2267) begin
      \nz.mem_912_sv2v_reg  <= data_i[0];
    end 
    if(N2266) begin
      \nz.mem_911_sv2v_reg  <= data_i[15];
    end 
    if(N2265) begin
      \nz.mem_910_sv2v_reg  <= data_i[14];
    end 
    if(N2264) begin
      \nz.mem_909_sv2v_reg  <= data_i[13];
    end 
    if(N2263) begin
      \nz.mem_908_sv2v_reg  <= data_i[12];
    end 
    if(N2262) begin
      \nz.mem_907_sv2v_reg  <= data_i[11];
    end 
    if(N2261) begin
      \nz.mem_906_sv2v_reg  <= data_i[10];
    end 
    if(N2260) begin
      \nz.mem_905_sv2v_reg  <= data_i[9];
    end 
    if(N2259) begin
      \nz.mem_904_sv2v_reg  <= data_i[8];
    end 
    if(N2258) begin
      \nz.mem_903_sv2v_reg  <= data_i[7];
    end 
    if(N2257) begin
      \nz.mem_902_sv2v_reg  <= data_i[6];
    end 
    if(N2256) begin
      \nz.mem_901_sv2v_reg  <= data_i[5];
    end 
    if(N2255) begin
      \nz.mem_900_sv2v_reg  <= data_i[4];
    end 
    if(N2254) begin
      \nz.mem_899_sv2v_reg  <= data_i[3];
    end 
    if(N2253) begin
      \nz.mem_898_sv2v_reg  <= data_i[2];
    end 
    if(N2252) begin
      \nz.mem_897_sv2v_reg  <= data_i[1];
    end 
    if(N2251) begin
      \nz.mem_896_sv2v_reg  <= data_i[0];
    end 
    if(N2250) begin
      \nz.mem_895_sv2v_reg  <= data_i[15];
    end 
    if(N2249) begin
      \nz.mem_894_sv2v_reg  <= data_i[14];
    end 
    if(N2248) begin
      \nz.mem_893_sv2v_reg  <= data_i[13];
    end 
    if(N2247) begin
      \nz.mem_892_sv2v_reg  <= data_i[12];
    end 
    if(N2246) begin
      \nz.mem_891_sv2v_reg  <= data_i[11];
    end 
    if(N2245) begin
      \nz.mem_890_sv2v_reg  <= data_i[10];
    end 
    if(N2244) begin
      \nz.mem_889_sv2v_reg  <= data_i[9];
    end 
    if(N2243) begin
      \nz.mem_888_sv2v_reg  <= data_i[8];
    end 
    if(N2242) begin
      \nz.mem_887_sv2v_reg  <= data_i[7];
    end 
    if(N2241) begin
      \nz.mem_886_sv2v_reg  <= data_i[6];
    end 
    if(N2240) begin
      \nz.mem_885_sv2v_reg  <= data_i[5];
    end 
    if(N2239) begin
      \nz.mem_884_sv2v_reg  <= data_i[4];
    end 
    if(N2238) begin
      \nz.mem_883_sv2v_reg  <= data_i[3];
    end 
    if(N2237) begin
      \nz.mem_882_sv2v_reg  <= data_i[2];
    end 
    if(N2236) begin
      \nz.mem_881_sv2v_reg  <= data_i[1];
    end 
    if(N2235) begin
      \nz.mem_880_sv2v_reg  <= data_i[0];
    end 
    if(N2234) begin
      \nz.mem_879_sv2v_reg  <= data_i[15];
    end 
    if(N2233) begin
      \nz.mem_878_sv2v_reg  <= data_i[14];
    end 
    if(N2232) begin
      \nz.mem_877_sv2v_reg  <= data_i[13];
    end 
    if(N2231) begin
      \nz.mem_876_sv2v_reg  <= data_i[12];
    end 
    if(N2230) begin
      \nz.mem_875_sv2v_reg  <= data_i[11];
    end 
    if(N2229) begin
      \nz.mem_874_sv2v_reg  <= data_i[10];
    end 
    if(N2228) begin
      \nz.mem_873_sv2v_reg  <= data_i[9];
    end 
    if(N2227) begin
      \nz.mem_872_sv2v_reg  <= data_i[8];
    end 
    if(N2226) begin
      \nz.mem_871_sv2v_reg  <= data_i[7];
    end 
    if(N2225) begin
      \nz.mem_870_sv2v_reg  <= data_i[6];
    end 
    if(N2224) begin
      \nz.mem_869_sv2v_reg  <= data_i[5];
    end 
    if(N2223) begin
      \nz.mem_868_sv2v_reg  <= data_i[4];
    end 
    if(N2222) begin
      \nz.mem_867_sv2v_reg  <= data_i[3];
    end 
    if(N2221) begin
      \nz.mem_866_sv2v_reg  <= data_i[2];
    end 
    if(N2220) begin
      \nz.mem_865_sv2v_reg  <= data_i[1];
    end 
    if(N2219) begin
      \nz.mem_864_sv2v_reg  <= data_i[0];
    end 
    if(N2218) begin
      \nz.mem_863_sv2v_reg  <= data_i[15];
    end 
    if(N2217) begin
      \nz.mem_862_sv2v_reg  <= data_i[14];
    end 
    if(N2216) begin
      \nz.mem_861_sv2v_reg  <= data_i[13];
    end 
    if(N2215) begin
      \nz.mem_860_sv2v_reg  <= data_i[12];
    end 
    if(N2214) begin
      \nz.mem_859_sv2v_reg  <= data_i[11];
    end 
    if(N2213) begin
      \nz.mem_858_sv2v_reg  <= data_i[10];
    end 
    if(N2212) begin
      \nz.mem_857_sv2v_reg  <= data_i[9];
    end 
    if(N2211) begin
      \nz.mem_856_sv2v_reg  <= data_i[8];
    end 
    if(N2210) begin
      \nz.mem_855_sv2v_reg  <= data_i[7];
    end 
    if(N2209) begin
      \nz.mem_854_sv2v_reg  <= data_i[6];
    end 
    if(N2208) begin
      \nz.mem_853_sv2v_reg  <= data_i[5];
    end 
    if(N2207) begin
      \nz.mem_852_sv2v_reg  <= data_i[4];
    end 
    if(N2206) begin
      \nz.mem_851_sv2v_reg  <= data_i[3];
    end 
    if(N2205) begin
      \nz.mem_850_sv2v_reg  <= data_i[2];
    end 
    if(N2204) begin
      \nz.mem_849_sv2v_reg  <= data_i[1];
    end 
    if(N2203) begin
      \nz.mem_848_sv2v_reg  <= data_i[0];
    end 
    if(N2202) begin
      \nz.mem_847_sv2v_reg  <= data_i[15];
    end 
    if(N2201) begin
      \nz.mem_846_sv2v_reg  <= data_i[14];
    end 
    if(N2200) begin
      \nz.mem_845_sv2v_reg  <= data_i[13];
    end 
    if(N2199) begin
      \nz.mem_844_sv2v_reg  <= data_i[12];
    end 
    if(N2198) begin
      \nz.mem_843_sv2v_reg  <= data_i[11];
    end 
    if(N2197) begin
      \nz.mem_842_sv2v_reg  <= data_i[10];
    end 
    if(N2196) begin
      \nz.mem_841_sv2v_reg  <= data_i[9];
    end 
    if(N2195) begin
      \nz.mem_840_sv2v_reg  <= data_i[8];
    end 
    if(N2194) begin
      \nz.mem_839_sv2v_reg  <= data_i[7];
    end 
    if(N2193) begin
      \nz.mem_838_sv2v_reg  <= data_i[6];
    end 
    if(N2192) begin
      \nz.mem_837_sv2v_reg  <= data_i[5];
    end 
    if(N2191) begin
      \nz.mem_836_sv2v_reg  <= data_i[4];
    end 
    if(N2190) begin
      \nz.mem_835_sv2v_reg  <= data_i[3];
    end 
    if(N2189) begin
      \nz.mem_834_sv2v_reg  <= data_i[2];
    end 
    if(N2188) begin
      \nz.mem_833_sv2v_reg  <= data_i[1];
    end 
    if(N2187) begin
      \nz.mem_832_sv2v_reg  <= data_i[0];
    end 
    if(N2186) begin
      \nz.mem_831_sv2v_reg  <= data_i[15];
    end 
    if(N2185) begin
      \nz.mem_830_sv2v_reg  <= data_i[14];
    end 
    if(N2184) begin
      \nz.mem_829_sv2v_reg  <= data_i[13];
    end 
    if(N2183) begin
      \nz.mem_828_sv2v_reg  <= data_i[12];
    end 
    if(N2182) begin
      \nz.mem_827_sv2v_reg  <= data_i[11];
    end 
    if(N2181) begin
      \nz.mem_826_sv2v_reg  <= data_i[10];
    end 
    if(N2180) begin
      \nz.mem_825_sv2v_reg  <= data_i[9];
    end 
    if(N2179) begin
      \nz.mem_824_sv2v_reg  <= data_i[8];
    end 
    if(N2178) begin
      \nz.mem_823_sv2v_reg  <= data_i[7];
    end 
    if(N2177) begin
      \nz.mem_822_sv2v_reg  <= data_i[6];
    end 
    if(N2176) begin
      \nz.mem_821_sv2v_reg  <= data_i[5];
    end 
    if(N2175) begin
      \nz.mem_820_sv2v_reg  <= data_i[4];
    end 
    if(N2174) begin
      \nz.mem_819_sv2v_reg  <= data_i[3];
    end 
    if(N2173) begin
      \nz.mem_818_sv2v_reg  <= data_i[2];
    end 
    if(N2172) begin
      \nz.mem_817_sv2v_reg  <= data_i[1];
    end 
    if(N2171) begin
      \nz.mem_816_sv2v_reg  <= data_i[0];
    end 
    if(N2170) begin
      \nz.mem_815_sv2v_reg  <= data_i[15];
    end 
    if(N2169) begin
      \nz.mem_814_sv2v_reg  <= data_i[14];
    end 
    if(N2168) begin
      \nz.mem_813_sv2v_reg  <= data_i[13];
    end 
    if(N2167) begin
      \nz.mem_812_sv2v_reg  <= data_i[12];
    end 
    if(N2166) begin
      \nz.mem_811_sv2v_reg  <= data_i[11];
    end 
    if(N2165) begin
      \nz.mem_810_sv2v_reg  <= data_i[10];
    end 
    if(N2164) begin
      \nz.mem_809_sv2v_reg  <= data_i[9];
    end 
    if(N2163) begin
      \nz.mem_808_sv2v_reg  <= data_i[8];
    end 
    if(N2162) begin
      \nz.mem_807_sv2v_reg  <= data_i[7];
    end 
    if(N2161) begin
      \nz.mem_806_sv2v_reg  <= data_i[6];
    end 
    if(N2160) begin
      \nz.mem_805_sv2v_reg  <= data_i[5];
    end 
    if(N2159) begin
      \nz.mem_804_sv2v_reg  <= data_i[4];
    end 
    if(N2158) begin
      \nz.mem_803_sv2v_reg  <= data_i[3];
    end 
    if(N2157) begin
      \nz.mem_802_sv2v_reg  <= data_i[2];
    end 
    if(N2156) begin
      \nz.mem_801_sv2v_reg  <= data_i[1];
    end 
    if(N2155) begin
      \nz.mem_800_sv2v_reg  <= data_i[0];
    end 
    if(N2154) begin
      \nz.mem_799_sv2v_reg  <= data_i[15];
    end 
    if(N2153) begin
      \nz.mem_798_sv2v_reg  <= data_i[14];
    end 
    if(N2152) begin
      \nz.mem_797_sv2v_reg  <= data_i[13];
    end 
    if(N2151) begin
      \nz.mem_796_sv2v_reg  <= data_i[12];
    end 
    if(N2150) begin
      \nz.mem_795_sv2v_reg  <= data_i[11];
    end 
    if(N2149) begin
      \nz.mem_794_sv2v_reg  <= data_i[10];
    end 
    if(N2148) begin
      \nz.mem_793_sv2v_reg  <= data_i[9];
    end 
    if(N2147) begin
      \nz.mem_792_sv2v_reg  <= data_i[8];
    end 
    if(N2146) begin
      \nz.mem_791_sv2v_reg  <= data_i[7];
    end 
    if(N2145) begin
      \nz.mem_790_sv2v_reg  <= data_i[6];
    end 
    if(N2144) begin
      \nz.mem_789_sv2v_reg  <= data_i[5];
    end 
    if(N2143) begin
      \nz.mem_788_sv2v_reg  <= data_i[4];
    end 
    if(N2142) begin
      \nz.mem_787_sv2v_reg  <= data_i[3];
    end 
    if(N2141) begin
      \nz.mem_786_sv2v_reg  <= data_i[2];
    end 
    if(N2140) begin
      \nz.mem_785_sv2v_reg  <= data_i[1];
    end 
    if(N2139) begin
      \nz.mem_784_sv2v_reg  <= data_i[0];
    end 
    if(N2138) begin
      \nz.mem_783_sv2v_reg  <= data_i[15];
    end 
    if(N2137) begin
      \nz.mem_782_sv2v_reg  <= data_i[14];
    end 
    if(N2136) begin
      \nz.mem_781_sv2v_reg  <= data_i[13];
    end 
    if(N2135) begin
      \nz.mem_780_sv2v_reg  <= data_i[12];
    end 
    if(N2134) begin
      \nz.mem_779_sv2v_reg  <= data_i[11];
    end 
    if(N2133) begin
      \nz.mem_778_sv2v_reg  <= data_i[10];
    end 
    if(N2132) begin
      \nz.mem_777_sv2v_reg  <= data_i[9];
    end 
    if(N2131) begin
      \nz.mem_776_sv2v_reg  <= data_i[8];
    end 
    if(N2130) begin
      \nz.mem_775_sv2v_reg  <= data_i[7];
    end 
    if(N2129) begin
      \nz.mem_774_sv2v_reg  <= data_i[6];
    end 
    if(N2128) begin
      \nz.mem_773_sv2v_reg  <= data_i[5];
    end 
    if(N2127) begin
      \nz.mem_772_sv2v_reg  <= data_i[4];
    end 
    if(N2126) begin
      \nz.mem_771_sv2v_reg  <= data_i[3];
    end 
    if(N2125) begin
      \nz.mem_770_sv2v_reg  <= data_i[2];
    end 
    if(N2124) begin
      \nz.mem_769_sv2v_reg  <= data_i[1];
    end 
    if(N2123) begin
      \nz.mem_768_sv2v_reg  <= data_i[0];
    end 
    if(N2122) begin
      \nz.mem_767_sv2v_reg  <= data_i[15];
    end 
    if(N2121) begin
      \nz.mem_766_sv2v_reg  <= data_i[14];
    end 
    if(N2120) begin
      \nz.mem_765_sv2v_reg  <= data_i[13];
    end 
    if(N2119) begin
      \nz.mem_764_sv2v_reg  <= data_i[12];
    end 
    if(N2118) begin
      \nz.mem_763_sv2v_reg  <= data_i[11];
    end 
    if(N2117) begin
      \nz.mem_762_sv2v_reg  <= data_i[10];
    end 
    if(N2116) begin
      \nz.mem_761_sv2v_reg  <= data_i[9];
    end 
    if(N2115) begin
      \nz.mem_760_sv2v_reg  <= data_i[8];
    end 
    if(N2114) begin
      \nz.mem_759_sv2v_reg  <= data_i[7];
    end 
    if(N2113) begin
      \nz.mem_758_sv2v_reg  <= data_i[6];
    end 
    if(N2112) begin
      \nz.mem_757_sv2v_reg  <= data_i[5];
    end 
    if(N2111) begin
      \nz.mem_756_sv2v_reg  <= data_i[4];
    end 
    if(N2110) begin
      \nz.mem_755_sv2v_reg  <= data_i[3];
    end 
    if(N2109) begin
      \nz.mem_754_sv2v_reg  <= data_i[2];
    end 
    if(N2108) begin
      \nz.mem_753_sv2v_reg  <= data_i[1];
    end 
    if(N2107) begin
      \nz.mem_752_sv2v_reg  <= data_i[0];
    end 
    if(N2106) begin
      \nz.mem_751_sv2v_reg  <= data_i[15];
    end 
    if(N2105) begin
      \nz.mem_750_sv2v_reg  <= data_i[14];
    end 
    if(N2104) begin
      \nz.mem_749_sv2v_reg  <= data_i[13];
    end 
    if(N2103) begin
      \nz.mem_748_sv2v_reg  <= data_i[12];
    end 
    if(N2102) begin
      \nz.mem_747_sv2v_reg  <= data_i[11];
    end 
    if(N2101) begin
      \nz.mem_746_sv2v_reg  <= data_i[10];
    end 
    if(N2100) begin
      \nz.mem_745_sv2v_reg  <= data_i[9];
    end 
    if(N2099) begin
      \nz.mem_744_sv2v_reg  <= data_i[8];
    end 
    if(N2098) begin
      \nz.mem_743_sv2v_reg  <= data_i[7];
    end 
    if(N2097) begin
      \nz.mem_742_sv2v_reg  <= data_i[6];
    end 
    if(N2096) begin
      \nz.mem_741_sv2v_reg  <= data_i[5];
    end 
    if(N2095) begin
      \nz.mem_740_sv2v_reg  <= data_i[4];
    end 
    if(N2094) begin
      \nz.mem_739_sv2v_reg  <= data_i[3];
    end 
    if(N2093) begin
      \nz.mem_738_sv2v_reg  <= data_i[2];
    end 
    if(N2092) begin
      \nz.mem_737_sv2v_reg  <= data_i[1];
    end 
    if(N2091) begin
      \nz.mem_736_sv2v_reg  <= data_i[0];
    end 
    if(N2090) begin
      \nz.mem_735_sv2v_reg  <= data_i[15];
    end 
    if(N2089) begin
      \nz.mem_734_sv2v_reg  <= data_i[14];
    end 
    if(N2088) begin
      \nz.mem_733_sv2v_reg  <= data_i[13];
    end 
    if(N2087) begin
      \nz.mem_732_sv2v_reg  <= data_i[12];
    end 
    if(N2086) begin
      \nz.mem_731_sv2v_reg  <= data_i[11];
    end 
    if(N2085) begin
      \nz.mem_730_sv2v_reg  <= data_i[10];
    end 
    if(N2084) begin
      \nz.mem_729_sv2v_reg  <= data_i[9];
    end 
    if(N2083) begin
      \nz.mem_728_sv2v_reg  <= data_i[8];
    end 
    if(N2082) begin
      \nz.mem_727_sv2v_reg  <= data_i[7];
    end 
    if(N2081) begin
      \nz.mem_726_sv2v_reg  <= data_i[6];
    end 
    if(N2080) begin
      \nz.mem_725_sv2v_reg  <= data_i[5];
    end 
    if(N2079) begin
      \nz.mem_724_sv2v_reg  <= data_i[4];
    end 
    if(N2078) begin
      \nz.mem_723_sv2v_reg  <= data_i[3];
    end 
    if(N2077) begin
      \nz.mem_722_sv2v_reg  <= data_i[2];
    end 
    if(N2076) begin
      \nz.mem_721_sv2v_reg  <= data_i[1];
    end 
    if(N2075) begin
      \nz.mem_720_sv2v_reg  <= data_i[0];
    end 
    if(N2074) begin
      \nz.mem_719_sv2v_reg  <= data_i[15];
    end 
    if(N2073) begin
      \nz.mem_718_sv2v_reg  <= data_i[14];
    end 
    if(N2072) begin
      \nz.mem_717_sv2v_reg  <= data_i[13];
    end 
    if(N2071) begin
      \nz.mem_716_sv2v_reg  <= data_i[12];
    end 
    if(N2070) begin
      \nz.mem_715_sv2v_reg  <= data_i[11];
    end 
    if(N2069) begin
      \nz.mem_714_sv2v_reg  <= data_i[10];
    end 
    if(N2068) begin
      \nz.mem_713_sv2v_reg  <= data_i[9];
    end 
    if(N2067) begin
      \nz.mem_712_sv2v_reg  <= data_i[8];
    end 
    if(N2066) begin
      \nz.mem_711_sv2v_reg  <= data_i[7];
    end 
    if(N2065) begin
      \nz.mem_710_sv2v_reg  <= data_i[6];
    end 
    if(N2064) begin
      \nz.mem_709_sv2v_reg  <= data_i[5];
    end 
    if(N2063) begin
      \nz.mem_708_sv2v_reg  <= data_i[4];
    end 
    if(N2062) begin
      \nz.mem_707_sv2v_reg  <= data_i[3];
    end 
    if(N2061) begin
      \nz.mem_706_sv2v_reg  <= data_i[2];
    end 
    if(N2060) begin
      \nz.mem_705_sv2v_reg  <= data_i[1];
    end 
    if(N2059) begin
      \nz.mem_704_sv2v_reg  <= data_i[0];
    end 
    if(N2058) begin
      \nz.mem_703_sv2v_reg  <= data_i[15];
    end 
    if(N2057) begin
      \nz.mem_702_sv2v_reg  <= data_i[14];
    end 
    if(N2056) begin
      \nz.mem_701_sv2v_reg  <= data_i[13];
    end 
    if(N2055) begin
      \nz.mem_700_sv2v_reg  <= data_i[12];
    end 
    if(N2054) begin
      \nz.mem_699_sv2v_reg  <= data_i[11];
    end 
    if(N2053) begin
      \nz.mem_698_sv2v_reg  <= data_i[10];
    end 
    if(N2052) begin
      \nz.mem_697_sv2v_reg  <= data_i[9];
    end 
    if(N2051) begin
      \nz.mem_696_sv2v_reg  <= data_i[8];
    end 
    if(N2050) begin
      \nz.mem_695_sv2v_reg  <= data_i[7];
    end 
    if(N2049) begin
      \nz.mem_694_sv2v_reg  <= data_i[6];
    end 
    if(N2048) begin
      \nz.mem_693_sv2v_reg  <= data_i[5];
    end 
    if(N2047) begin
      \nz.mem_692_sv2v_reg  <= data_i[4];
    end 
    if(N2046) begin
      \nz.mem_691_sv2v_reg  <= data_i[3];
    end 
    if(N2045) begin
      \nz.mem_690_sv2v_reg  <= data_i[2];
    end 
    if(N2044) begin
      \nz.mem_689_sv2v_reg  <= data_i[1];
    end 
    if(N2043) begin
      \nz.mem_688_sv2v_reg  <= data_i[0];
    end 
    if(N2042) begin
      \nz.mem_687_sv2v_reg  <= data_i[15];
    end 
    if(N2041) begin
      \nz.mem_686_sv2v_reg  <= data_i[14];
    end 
    if(N2040) begin
      \nz.mem_685_sv2v_reg  <= data_i[13];
    end 
    if(N2039) begin
      \nz.mem_684_sv2v_reg  <= data_i[12];
    end 
    if(N2038) begin
      \nz.mem_683_sv2v_reg  <= data_i[11];
    end 
    if(N2037) begin
      \nz.mem_682_sv2v_reg  <= data_i[10];
    end 
    if(N2036) begin
      \nz.mem_681_sv2v_reg  <= data_i[9];
    end 
    if(N2035) begin
      \nz.mem_680_sv2v_reg  <= data_i[8];
    end 
    if(N2034) begin
      \nz.mem_679_sv2v_reg  <= data_i[7];
    end 
    if(N2033) begin
      \nz.mem_678_sv2v_reg  <= data_i[6];
    end 
    if(N2032) begin
      \nz.mem_677_sv2v_reg  <= data_i[5];
    end 
    if(N2031) begin
      \nz.mem_676_sv2v_reg  <= data_i[4];
    end 
    if(N2030) begin
      \nz.mem_675_sv2v_reg  <= data_i[3];
    end 
    if(N2029) begin
      \nz.mem_674_sv2v_reg  <= data_i[2];
    end 
    if(N2028) begin
      \nz.mem_673_sv2v_reg  <= data_i[1];
    end 
    if(N2027) begin
      \nz.mem_672_sv2v_reg  <= data_i[0];
    end 
    if(N2026) begin
      \nz.mem_671_sv2v_reg  <= data_i[15];
    end 
    if(N2025) begin
      \nz.mem_670_sv2v_reg  <= data_i[14];
    end 
    if(N2024) begin
      \nz.mem_669_sv2v_reg  <= data_i[13];
    end 
    if(N2023) begin
      \nz.mem_668_sv2v_reg  <= data_i[12];
    end 
    if(N2022) begin
      \nz.mem_667_sv2v_reg  <= data_i[11];
    end 
    if(N2021) begin
      \nz.mem_666_sv2v_reg  <= data_i[10];
    end 
    if(N2020) begin
      \nz.mem_665_sv2v_reg  <= data_i[9];
    end 
    if(N2019) begin
      \nz.mem_664_sv2v_reg  <= data_i[8];
    end 
    if(N2018) begin
      \nz.mem_663_sv2v_reg  <= data_i[7];
    end 
    if(N2017) begin
      \nz.mem_662_sv2v_reg  <= data_i[6];
    end 
    if(N2016) begin
      \nz.mem_661_sv2v_reg  <= data_i[5];
    end 
    if(N2015) begin
      \nz.mem_660_sv2v_reg  <= data_i[4];
    end 
    if(N2014) begin
      \nz.mem_659_sv2v_reg  <= data_i[3];
    end 
    if(N2013) begin
      \nz.mem_658_sv2v_reg  <= data_i[2];
    end 
    if(N2012) begin
      \nz.mem_657_sv2v_reg  <= data_i[1];
    end 
    if(N2011) begin
      \nz.mem_656_sv2v_reg  <= data_i[0];
    end 
    if(N2010) begin
      \nz.mem_655_sv2v_reg  <= data_i[15];
    end 
    if(N2009) begin
      \nz.mem_654_sv2v_reg  <= data_i[14];
    end 
    if(N2008) begin
      \nz.mem_653_sv2v_reg  <= data_i[13];
    end 
    if(N2007) begin
      \nz.mem_652_sv2v_reg  <= data_i[12];
    end 
    if(N2006) begin
      \nz.mem_651_sv2v_reg  <= data_i[11];
    end 
    if(N2005) begin
      \nz.mem_650_sv2v_reg  <= data_i[10];
    end 
    if(N2004) begin
      \nz.mem_649_sv2v_reg  <= data_i[9];
    end 
    if(N2003) begin
      \nz.mem_648_sv2v_reg  <= data_i[8];
    end 
    if(N2002) begin
      \nz.mem_647_sv2v_reg  <= data_i[7];
    end 
    if(N2001) begin
      \nz.mem_646_sv2v_reg  <= data_i[6];
    end 
    if(N2000) begin
      \nz.mem_645_sv2v_reg  <= data_i[5];
    end 
    if(N1999) begin
      \nz.mem_644_sv2v_reg  <= data_i[4];
    end 
    if(N1998) begin
      \nz.mem_643_sv2v_reg  <= data_i[3];
    end 
    if(N1997) begin
      \nz.mem_642_sv2v_reg  <= data_i[2];
    end 
    if(N1996) begin
      \nz.mem_641_sv2v_reg  <= data_i[1];
    end 
    if(N1995) begin
      \nz.mem_640_sv2v_reg  <= data_i[0];
    end 
    if(N1994) begin
      \nz.mem_639_sv2v_reg  <= data_i[15];
    end 
    if(N1993) begin
      \nz.mem_638_sv2v_reg  <= data_i[14];
    end 
    if(N1992) begin
      \nz.mem_637_sv2v_reg  <= data_i[13];
    end 
    if(N1991) begin
      \nz.mem_636_sv2v_reg  <= data_i[12];
    end 
    if(N1990) begin
      \nz.mem_635_sv2v_reg  <= data_i[11];
    end 
    if(N1989) begin
      \nz.mem_634_sv2v_reg  <= data_i[10];
    end 
    if(N1988) begin
      \nz.mem_633_sv2v_reg  <= data_i[9];
    end 
    if(N1987) begin
      \nz.mem_632_sv2v_reg  <= data_i[8];
    end 
    if(N1986) begin
      \nz.mem_631_sv2v_reg  <= data_i[7];
    end 
    if(N1985) begin
      \nz.mem_630_sv2v_reg  <= data_i[6];
    end 
    if(N1984) begin
      \nz.mem_629_sv2v_reg  <= data_i[5];
    end 
    if(N1983) begin
      \nz.mem_628_sv2v_reg  <= data_i[4];
    end 
    if(N1982) begin
      \nz.mem_627_sv2v_reg  <= data_i[3];
    end 
    if(N1981) begin
      \nz.mem_626_sv2v_reg  <= data_i[2];
    end 
    if(N1980) begin
      \nz.mem_625_sv2v_reg  <= data_i[1];
    end 
    if(N1979) begin
      \nz.mem_624_sv2v_reg  <= data_i[0];
    end 
    if(N1978) begin
      \nz.mem_623_sv2v_reg  <= data_i[15];
    end 
    if(N1977) begin
      \nz.mem_622_sv2v_reg  <= data_i[14];
    end 
    if(N1976) begin
      \nz.mem_621_sv2v_reg  <= data_i[13];
    end 
    if(N1975) begin
      \nz.mem_620_sv2v_reg  <= data_i[12];
    end 
    if(N1974) begin
      \nz.mem_619_sv2v_reg  <= data_i[11];
    end 
    if(N1973) begin
      \nz.mem_618_sv2v_reg  <= data_i[10];
    end 
    if(N1972) begin
      \nz.mem_617_sv2v_reg  <= data_i[9];
    end 
    if(N1971) begin
      \nz.mem_616_sv2v_reg  <= data_i[8];
    end 
    if(N1970) begin
      \nz.mem_615_sv2v_reg  <= data_i[7];
    end 
    if(N1969) begin
      \nz.mem_614_sv2v_reg  <= data_i[6];
    end 
    if(N1968) begin
      \nz.mem_613_sv2v_reg  <= data_i[5];
    end 
    if(N1967) begin
      \nz.mem_612_sv2v_reg  <= data_i[4];
    end 
    if(N1966) begin
      \nz.mem_611_sv2v_reg  <= data_i[3];
    end 
    if(N1965) begin
      \nz.mem_610_sv2v_reg  <= data_i[2];
    end 
    if(N1964) begin
      \nz.mem_609_sv2v_reg  <= data_i[1];
    end 
    if(N1963) begin
      \nz.mem_608_sv2v_reg  <= data_i[0];
    end 
    if(N1962) begin
      \nz.mem_607_sv2v_reg  <= data_i[15];
    end 
    if(N1961) begin
      \nz.mem_606_sv2v_reg  <= data_i[14];
    end 
    if(N1960) begin
      \nz.mem_605_sv2v_reg  <= data_i[13];
    end 
    if(N1959) begin
      \nz.mem_604_sv2v_reg  <= data_i[12];
    end 
    if(N1958) begin
      \nz.mem_603_sv2v_reg  <= data_i[11];
    end 
    if(N1957) begin
      \nz.mem_602_sv2v_reg  <= data_i[10];
    end 
    if(N1956) begin
      \nz.mem_601_sv2v_reg  <= data_i[9];
    end 
    if(N1955) begin
      \nz.mem_600_sv2v_reg  <= data_i[8];
    end 
    if(N1954) begin
      \nz.mem_599_sv2v_reg  <= data_i[7];
    end 
    if(N1953) begin
      \nz.mem_598_sv2v_reg  <= data_i[6];
    end 
    if(N1952) begin
      \nz.mem_597_sv2v_reg  <= data_i[5];
    end 
    if(N1951) begin
      \nz.mem_596_sv2v_reg  <= data_i[4];
    end 
    if(N1950) begin
      \nz.mem_595_sv2v_reg  <= data_i[3];
    end 
    if(N1949) begin
      \nz.mem_594_sv2v_reg  <= data_i[2];
    end 
    if(N1948) begin
      \nz.mem_593_sv2v_reg  <= data_i[1];
    end 
    if(N1947) begin
      \nz.mem_592_sv2v_reg  <= data_i[0];
    end 
    if(N1946) begin
      \nz.mem_591_sv2v_reg  <= data_i[15];
    end 
    if(N1945) begin
      \nz.mem_590_sv2v_reg  <= data_i[14];
    end 
    if(N1944) begin
      \nz.mem_589_sv2v_reg  <= data_i[13];
    end 
    if(N1943) begin
      \nz.mem_588_sv2v_reg  <= data_i[12];
    end 
    if(N1942) begin
      \nz.mem_587_sv2v_reg  <= data_i[11];
    end 
    if(N1941) begin
      \nz.mem_586_sv2v_reg  <= data_i[10];
    end 
    if(N1940) begin
      \nz.mem_585_sv2v_reg  <= data_i[9];
    end 
    if(N1939) begin
      \nz.mem_584_sv2v_reg  <= data_i[8];
    end 
    if(N1938) begin
      \nz.mem_583_sv2v_reg  <= data_i[7];
    end 
    if(N1937) begin
      \nz.mem_582_sv2v_reg  <= data_i[6];
    end 
    if(N1936) begin
      \nz.mem_581_sv2v_reg  <= data_i[5];
    end 
    if(N1935) begin
      \nz.mem_580_sv2v_reg  <= data_i[4];
    end 
    if(N1934) begin
      \nz.mem_579_sv2v_reg  <= data_i[3];
    end 
    if(N1933) begin
      \nz.mem_578_sv2v_reg  <= data_i[2];
    end 
    if(N1932) begin
      \nz.mem_577_sv2v_reg  <= data_i[1];
    end 
    if(N1931) begin
      \nz.mem_576_sv2v_reg  <= data_i[0];
    end 
    if(N1930) begin
      \nz.mem_575_sv2v_reg  <= data_i[15];
    end 
    if(N1929) begin
      \nz.mem_574_sv2v_reg  <= data_i[14];
    end 
    if(N1928) begin
      \nz.mem_573_sv2v_reg  <= data_i[13];
    end 
    if(N1927) begin
      \nz.mem_572_sv2v_reg  <= data_i[12];
    end 
    if(N1926) begin
      \nz.mem_571_sv2v_reg  <= data_i[11];
    end 
    if(N1925) begin
      \nz.mem_570_sv2v_reg  <= data_i[10];
    end 
    if(N1924) begin
      \nz.mem_569_sv2v_reg  <= data_i[9];
    end 
    if(N1923) begin
      \nz.mem_568_sv2v_reg  <= data_i[8];
    end 
    if(N1922) begin
      \nz.mem_567_sv2v_reg  <= data_i[7];
    end 
    if(N1921) begin
      \nz.mem_566_sv2v_reg  <= data_i[6];
    end 
    if(N1920) begin
      \nz.mem_565_sv2v_reg  <= data_i[5];
    end 
    if(N1919) begin
      \nz.mem_564_sv2v_reg  <= data_i[4];
    end 
    if(N1918) begin
      \nz.mem_563_sv2v_reg  <= data_i[3];
    end 
    if(N1917) begin
      \nz.mem_562_sv2v_reg  <= data_i[2];
    end 
    if(N1916) begin
      \nz.mem_561_sv2v_reg  <= data_i[1];
    end 
    if(N1915) begin
      \nz.mem_560_sv2v_reg  <= data_i[0];
    end 
    if(N1914) begin
      \nz.mem_559_sv2v_reg  <= data_i[15];
    end 
    if(N1913) begin
      \nz.mem_558_sv2v_reg  <= data_i[14];
    end 
    if(N1912) begin
      \nz.mem_557_sv2v_reg  <= data_i[13];
    end 
    if(N1911) begin
      \nz.mem_556_sv2v_reg  <= data_i[12];
    end 
    if(N1910) begin
      \nz.mem_555_sv2v_reg  <= data_i[11];
    end 
    if(N1909) begin
      \nz.mem_554_sv2v_reg  <= data_i[10];
    end 
    if(N1908) begin
      \nz.mem_553_sv2v_reg  <= data_i[9];
    end 
    if(N1907) begin
      \nz.mem_552_sv2v_reg  <= data_i[8];
    end 
    if(N1906) begin
      \nz.mem_551_sv2v_reg  <= data_i[7];
    end 
    if(N1905) begin
      \nz.mem_550_sv2v_reg  <= data_i[6];
    end 
    if(N1904) begin
      \nz.mem_549_sv2v_reg  <= data_i[5];
    end 
    if(N1903) begin
      \nz.mem_548_sv2v_reg  <= data_i[4];
    end 
    if(N1902) begin
      \nz.mem_547_sv2v_reg  <= data_i[3];
    end 
    if(N1901) begin
      \nz.mem_546_sv2v_reg  <= data_i[2];
    end 
    if(N1900) begin
      \nz.mem_545_sv2v_reg  <= data_i[1];
    end 
    if(N1899) begin
      \nz.mem_544_sv2v_reg  <= data_i[0];
    end 
    if(N1898) begin
      \nz.mem_543_sv2v_reg  <= data_i[15];
    end 
    if(N1897) begin
      \nz.mem_542_sv2v_reg  <= data_i[14];
    end 
    if(N1896) begin
      \nz.mem_541_sv2v_reg  <= data_i[13];
    end 
    if(N1895) begin
      \nz.mem_540_sv2v_reg  <= data_i[12];
    end 
    if(N1894) begin
      \nz.mem_539_sv2v_reg  <= data_i[11];
    end 
    if(N1893) begin
      \nz.mem_538_sv2v_reg  <= data_i[10];
    end 
    if(N1892) begin
      \nz.mem_537_sv2v_reg  <= data_i[9];
    end 
    if(N1891) begin
      \nz.mem_536_sv2v_reg  <= data_i[8];
    end 
    if(N1890) begin
      \nz.mem_535_sv2v_reg  <= data_i[7];
    end 
    if(N1889) begin
      \nz.mem_534_sv2v_reg  <= data_i[6];
    end 
    if(N1888) begin
      \nz.mem_533_sv2v_reg  <= data_i[5];
    end 
    if(N1887) begin
      \nz.mem_532_sv2v_reg  <= data_i[4];
    end 
    if(N1886) begin
      \nz.mem_531_sv2v_reg  <= data_i[3];
    end 
    if(N1885) begin
      \nz.mem_530_sv2v_reg  <= data_i[2];
    end 
    if(N1884) begin
      \nz.mem_529_sv2v_reg  <= data_i[1];
    end 
    if(N1883) begin
      \nz.mem_528_sv2v_reg  <= data_i[0];
    end 
    if(N1882) begin
      \nz.mem_527_sv2v_reg  <= data_i[15];
    end 
    if(N1881) begin
      \nz.mem_526_sv2v_reg  <= data_i[14];
    end 
    if(N1880) begin
      \nz.mem_525_sv2v_reg  <= data_i[13];
    end 
    if(N1879) begin
      \nz.mem_524_sv2v_reg  <= data_i[12];
    end 
    if(N1878) begin
      \nz.mem_523_sv2v_reg  <= data_i[11];
    end 
    if(N1877) begin
      \nz.mem_522_sv2v_reg  <= data_i[10];
    end 
    if(N1876) begin
      \nz.mem_521_sv2v_reg  <= data_i[9];
    end 
    if(N1875) begin
      \nz.mem_520_sv2v_reg  <= data_i[8];
    end 
    if(N1874) begin
      \nz.mem_519_sv2v_reg  <= data_i[7];
    end 
    if(N1873) begin
      \nz.mem_518_sv2v_reg  <= data_i[6];
    end 
    if(N1872) begin
      \nz.mem_517_sv2v_reg  <= data_i[5];
    end 
    if(N1871) begin
      \nz.mem_516_sv2v_reg  <= data_i[4];
    end 
    if(N1870) begin
      \nz.mem_515_sv2v_reg  <= data_i[3];
    end 
    if(N1869) begin
      \nz.mem_514_sv2v_reg  <= data_i[2];
    end 
    if(N1868) begin
      \nz.mem_513_sv2v_reg  <= data_i[1];
    end 
    if(N1867) begin
      \nz.mem_512_sv2v_reg  <= data_i[0];
    end 
    if(N1866) begin
      \nz.mem_511_sv2v_reg  <= data_i[15];
    end 
    if(N1865) begin
      \nz.mem_510_sv2v_reg  <= data_i[14];
    end 
    if(N1864) begin
      \nz.mem_509_sv2v_reg  <= data_i[13];
    end 
    if(N1863) begin
      \nz.mem_508_sv2v_reg  <= data_i[12];
    end 
    if(N1862) begin
      \nz.mem_507_sv2v_reg  <= data_i[11];
    end 
    if(N1861) begin
      \nz.mem_506_sv2v_reg  <= data_i[10];
    end 
    if(N1860) begin
      \nz.mem_505_sv2v_reg  <= data_i[9];
    end 
    if(N1859) begin
      \nz.mem_504_sv2v_reg  <= data_i[8];
    end 
    if(N1858) begin
      \nz.mem_503_sv2v_reg  <= data_i[7];
    end 
    if(N1857) begin
      \nz.mem_502_sv2v_reg  <= data_i[6];
    end 
    if(N1856) begin
      \nz.mem_501_sv2v_reg  <= data_i[5];
    end 
    if(N1855) begin
      \nz.mem_500_sv2v_reg  <= data_i[4];
    end 
    if(N1854) begin
      \nz.mem_499_sv2v_reg  <= data_i[3];
    end 
    if(N1853) begin
      \nz.mem_498_sv2v_reg  <= data_i[2];
    end 
    if(N1852) begin
      \nz.mem_497_sv2v_reg  <= data_i[1];
    end 
    if(N1851) begin
      \nz.mem_496_sv2v_reg  <= data_i[0];
    end 
    if(N1850) begin
      \nz.mem_495_sv2v_reg  <= data_i[15];
    end 
    if(N1849) begin
      \nz.mem_494_sv2v_reg  <= data_i[14];
    end 
    if(N1848) begin
      \nz.mem_493_sv2v_reg  <= data_i[13];
    end 
    if(N1847) begin
      \nz.mem_492_sv2v_reg  <= data_i[12];
    end 
    if(N1846) begin
      \nz.mem_491_sv2v_reg  <= data_i[11];
    end 
    if(N1845) begin
      \nz.mem_490_sv2v_reg  <= data_i[10];
    end 
    if(N1844) begin
      \nz.mem_489_sv2v_reg  <= data_i[9];
    end 
    if(N1843) begin
      \nz.mem_488_sv2v_reg  <= data_i[8];
    end 
    if(N1842) begin
      \nz.mem_487_sv2v_reg  <= data_i[7];
    end 
    if(N1841) begin
      \nz.mem_486_sv2v_reg  <= data_i[6];
    end 
    if(N1840) begin
      \nz.mem_485_sv2v_reg  <= data_i[5];
    end 
    if(N1839) begin
      \nz.mem_484_sv2v_reg  <= data_i[4];
    end 
    if(N1838) begin
      \nz.mem_483_sv2v_reg  <= data_i[3];
    end 
    if(N1837) begin
      \nz.mem_482_sv2v_reg  <= data_i[2];
    end 
    if(N1836) begin
      \nz.mem_481_sv2v_reg  <= data_i[1];
    end 
    if(N1835) begin
      \nz.mem_480_sv2v_reg  <= data_i[0];
    end 
    if(N1834) begin
      \nz.mem_479_sv2v_reg  <= data_i[15];
    end 
    if(N1833) begin
      \nz.mem_478_sv2v_reg  <= data_i[14];
    end 
    if(N1832) begin
      \nz.mem_477_sv2v_reg  <= data_i[13];
    end 
    if(N1831) begin
      \nz.mem_476_sv2v_reg  <= data_i[12];
    end 
    if(N1830) begin
      \nz.mem_475_sv2v_reg  <= data_i[11];
    end 
    if(N1829) begin
      \nz.mem_474_sv2v_reg  <= data_i[10];
    end 
    if(N1828) begin
      \nz.mem_473_sv2v_reg  <= data_i[9];
    end 
    if(N1827) begin
      \nz.mem_472_sv2v_reg  <= data_i[8];
    end 
    if(N1826) begin
      \nz.mem_471_sv2v_reg  <= data_i[7];
    end 
    if(N1825) begin
      \nz.mem_470_sv2v_reg  <= data_i[6];
    end 
    if(N1824) begin
      \nz.mem_469_sv2v_reg  <= data_i[5];
    end 
    if(N1823) begin
      \nz.mem_468_sv2v_reg  <= data_i[4];
    end 
    if(N1822) begin
      \nz.mem_467_sv2v_reg  <= data_i[3];
    end 
    if(N1821) begin
      \nz.mem_466_sv2v_reg  <= data_i[2];
    end 
    if(N1820) begin
      \nz.mem_465_sv2v_reg  <= data_i[1];
    end 
    if(N1819) begin
      \nz.mem_464_sv2v_reg  <= data_i[0];
    end 
    if(N1818) begin
      \nz.mem_463_sv2v_reg  <= data_i[15];
    end 
    if(N1817) begin
      \nz.mem_462_sv2v_reg  <= data_i[14];
    end 
    if(N1816) begin
      \nz.mem_461_sv2v_reg  <= data_i[13];
    end 
    if(N1815) begin
      \nz.mem_460_sv2v_reg  <= data_i[12];
    end 
    if(N1814) begin
      \nz.mem_459_sv2v_reg  <= data_i[11];
    end 
    if(N1813) begin
      \nz.mem_458_sv2v_reg  <= data_i[10];
    end 
    if(N1812) begin
      \nz.mem_457_sv2v_reg  <= data_i[9];
    end 
    if(N1811) begin
      \nz.mem_456_sv2v_reg  <= data_i[8];
    end 
    if(N1810) begin
      \nz.mem_455_sv2v_reg  <= data_i[7];
    end 
    if(N1809) begin
      \nz.mem_454_sv2v_reg  <= data_i[6];
    end 
    if(N1808) begin
      \nz.mem_453_sv2v_reg  <= data_i[5];
    end 
    if(N1807) begin
      \nz.mem_452_sv2v_reg  <= data_i[4];
    end 
    if(N1806) begin
      \nz.mem_451_sv2v_reg  <= data_i[3];
    end 
    if(N1805) begin
      \nz.mem_450_sv2v_reg  <= data_i[2];
    end 
    if(N1804) begin
      \nz.mem_449_sv2v_reg  <= data_i[1];
    end 
    if(N1803) begin
      \nz.mem_448_sv2v_reg  <= data_i[0];
    end 
    if(N1802) begin
      \nz.mem_447_sv2v_reg  <= data_i[15];
    end 
    if(N1801) begin
      \nz.mem_446_sv2v_reg  <= data_i[14];
    end 
    if(N1800) begin
      \nz.mem_445_sv2v_reg  <= data_i[13];
    end 
    if(N1799) begin
      \nz.mem_444_sv2v_reg  <= data_i[12];
    end 
    if(N1798) begin
      \nz.mem_443_sv2v_reg  <= data_i[11];
    end 
    if(N1797) begin
      \nz.mem_442_sv2v_reg  <= data_i[10];
    end 
    if(N1796) begin
      \nz.mem_441_sv2v_reg  <= data_i[9];
    end 
    if(N1795) begin
      \nz.mem_440_sv2v_reg  <= data_i[8];
    end 
    if(N1794) begin
      \nz.mem_439_sv2v_reg  <= data_i[7];
    end 
    if(N1793) begin
      \nz.mem_438_sv2v_reg  <= data_i[6];
    end 
    if(N1792) begin
      \nz.mem_437_sv2v_reg  <= data_i[5];
    end 
    if(N1791) begin
      \nz.mem_436_sv2v_reg  <= data_i[4];
    end 
    if(N1790) begin
      \nz.mem_435_sv2v_reg  <= data_i[3];
    end 
    if(N1789) begin
      \nz.mem_434_sv2v_reg  <= data_i[2];
    end 
    if(N1788) begin
      \nz.mem_433_sv2v_reg  <= data_i[1];
    end 
    if(N1787) begin
      \nz.mem_432_sv2v_reg  <= data_i[0];
    end 
    if(N1786) begin
      \nz.mem_431_sv2v_reg  <= data_i[15];
    end 
    if(N1785) begin
      \nz.mem_430_sv2v_reg  <= data_i[14];
    end 
    if(N1784) begin
      \nz.mem_429_sv2v_reg  <= data_i[13];
    end 
    if(N1783) begin
      \nz.mem_428_sv2v_reg  <= data_i[12];
    end 
    if(N1782) begin
      \nz.mem_427_sv2v_reg  <= data_i[11];
    end 
    if(N1781) begin
      \nz.mem_426_sv2v_reg  <= data_i[10];
    end 
    if(N1780) begin
      \nz.mem_425_sv2v_reg  <= data_i[9];
    end 
    if(N1779) begin
      \nz.mem_424_sv2v_reg  <= data_i[8];
    end 
    if(N1778) begin
      \nz.mem_423_sv2v_reg  <= data_i[7];
    end 
    if(N1777) begin
      \nz.mem_422_sv2v_reg  <= data_i[6];
    end 
    if(N1776) begin
      \nz.mem_421_sv2v_reg  <= data_i[5];
    end 
    if(N1775) begin
      \nz.mem_420_sv2v_reg  <= data_i[4];
    end 
    if(N1774) begin
      \nz.mem_419_sv2v_reg  <= data_i[3];
    end 
    if(N1773) begin
      \nz.mem_418_sv2v_reg  <= data_i[2];
    end 
    if(N1772) begin
      \nz.mem_417_sv2v_reg  <= data_i[1];
    end 
    if(N1771) begin
      \nz.mem_416_sv2v_reg  <= data_i[0];
    end 
    if(N1770) begin
      \nz.mem_415_sv2v_reg  <= data_i[15];
    end 
    if(N1769) begin
      \nz.mem_414_sv2v_reg  <= data_i[14];
    end 
    if(N1768) begin
      \nz.mem_413_sv2v_reg  <= data_i[13];
    end 
    if(N1767) begin
      \nz.mem_412_sv2v_reg  <= data_i[12];
    end 
    if(N1766) begin
      \nz.mem_411_sv2v_reg  <= data_i[11];
    end 
    if(N1765) begin
      \nz.mem_410_sv2v_reg  <= data_i[10];
    end 
    if(N1764) begin
      \nz.mem_409_sv2v_reg  <= data_i[9];
    end 
    if(N1763) begin
      \nz.mem_408_sv2v_reg  <= data_i[8];
    end 
    if(N1762) begin
      \nz.mem_407_sv2v_reg  <= data_i[7];
    end 
    if(N1761) begin
      \nz.mem_406_sv2v_reg  <= data_i[6];
    end 
    if(N1760) begin
      \nz.mem_405_sv2v_reg  <= data_i[5];
    end 
    if(N1759) begin
      \nz.mem_404_sv2v_reg  <= data_i[4];
    end 
    if(N1758) begin
      \nz.mem_403_sv2v_reg  <= data_i[3];
    end 
    if(N1757) begin
      \nz.mem_402_sv2v_reg  <= data_i[2];
    end 
    if(N1756) begin
      \nz.mem_401_sv2v_reg  <= data_i[1];
    end 
    if(N1755) begin
      \nz.mem_400_sv2v_reg  <= data_i[0];
    end 
    if(N1754) begin
      \nz.mem_399_sv2v_reg  <= data_i[15];
    end 
    if(N1753) begin
      \nz.mem_398_sv2v_reg  <= data_i[14];
    end 
    if(N1752) begin
      \nz.mem_397_sv2v_reg  <= data_i[13];
    end 
    if(N1751) begin
      \nz.mem_396_sv2v_reg  <= data_i[12];
    end 
    if(N1750) begin
      \nz.mem_395_sv2v_reg  <= data_i[11];
    end 
    if(N1749) begin
      \nz.mem_394_sv2v_reg  <= data_i[10];
    end 
    if(N1748) begin
      \nz.mem_393_sv2v_reg  <= data_i[9];
    end 
    if(N1747) begin
      \nz.mem_392_sv2v_reg  <= data_i[8];
    end 
    if(N1746) begin
      \nz.mem_391_sv2v_reg  <= data_i[7];
    end 
    if(N1745) begin
      \nz.mem_390_sv2v_reg  <= data_i[6];
    end 
    if(N1744) begin
      \nz.mem_389_sv2v_reg  <= data_i[5];
    end 
    if(N1743) begin
      \nz.mem_388_sv2v_reg  <= data_i[4];
    end 
    if(N1742) begin
      \nz.mem_387_sv2v_reg  <= data_i[3];
    end 
    if(N1741) begin
      \nz.mem_386_sv2v_reg  <= data_i[2];
    end 
    if(N1740) begin
      \nz.mem_385_sv2v_reg  <= data_i[1];
    end 
    if(N1739) begin
      \nz.mem_384_sv2v_reg  <= data_i[0];
    end 
    if(N1738) begin
      \nz.mem_383_sv2v_reg  <= data_i[15];
    end 
    if(N1737) begin
      \nz.mem_382_sv2v_reg  <= data_i[14];
    end 
    if(N1736) begin
      \nz.mem_381_sv2v_reg  <= data_i[13];
    end 
    if(N1735) begin
      \nz.mem_380_sv2v_reg  <= data_i[12];
    end 
    if(N1734) begin
      \nz.mem_379_sv2v_reg  <= data_i[11];
    end 
    if(N1733) begin
      \nz.mem_378_sv2v_reg  <= data_i[10];
    end 
    if(N1732) begin
      \nz.mem_377_sv2v_reg  <= data_i[9];
    end 
    if(N1731) begin
      \nz.mem_376_sv2v_reg  <= data_i[8];
    end 
    if(N1730) begin
      \nz.mem_375_sv2v_reg  <= data_i[7];
    end 
    if(N1729) begin
      \nz.mem_374_sv2v_reg  <= data_i[6];
    end 
    if(N1728) begin
      \nz.mem_373_sv2v_reg  <= data_i[5];
    end 
    if(N1727) begin
      \nz.mem_372_sv2v_reg  <= data_i[4];
    end 
    if(N1726) begin
      \nz.mem_371_sv2v_reg  <= data_i[3];
    end 
    if(N1725) begin
      \nz.mem_370_sv2v_reg  <= data_i[2];
    end 
    if(N1724) begin
      \nz.mem_369_sv2v_reg  <= data_i[1];
    end 
    if(N1723) begin
      \nz.mem_368_sv2v_reg  <= data_i[0];
    end 
    if(N1722) begin
      \nz.mem_367_sv2v_reg  <= data_i[15];
    end 
    if(N1721) begin
      \nz.mem_366_sv2v_reg  <= data_i[14];
    end 
    if(N1720) begin
      \nz.mem_365_sv2v_reg  <= data_i[13];
    end 
    if(N1719) begin
      \nz.mem_364_sv2v_reg  <= data_i[12];
    end 
    if(N1718) begin
      \nz.mem_363_sv2v_reg  <= data_i[11];
    end 
    if(N1717) begin
      \nz.mem_362_sv2v_reg  <= data_i[10];
    end 
    if(N1716) begin
      \nz.mem_361_sv2v_reg  <= data_i[9];
    end 
    if(N1715) begin
      \nz.mem_360_sv2v_reg  <= data_i[8];
    end 
    if(N1714) begin
      \nz.mem_359_sv2v_reg  <= data_i[7];
    end 
    if(N1713) begin
      \nz.mem_358_sv2v_reg  <= data_i[6];
    end 
    if(N1712) begin
      \nz.mem_357_sv2v_reg  <= data_i[5];
    end 
    if(N1711) begin
      \nz.mem_356_sv2v_reg  <= data_i[4];
    end 
    if(N1710) begin
      \nz.mem_355_sv2v_reg  <= data_i[3];
    end 
    if(N1709) begin
      \nz.mem_354_sv2v_reg  <= data_i[2];
    end 
    if(N1708) begin
      \nz.mem_353_sv2v_reg  <= data_i[1];
    end 
    if(N1707) begin
      \nz.mem_352_sv2v_reg  <= data_i[0];
    end 
    if(N1706) begin
      \nz.mem_351_sv2v_reg  <= data_i[15];
    end 
    if(N1705) begin
      \nz.mem_350_sv2v_reg  <= data_i[14];
    end 
    if(N1704) begin
      \nz.mem_349_sv2v_reg  <= data_i[13];
    end 
    if(N1703) begin
      \nz.mem_348_sv2v_reg  <= data_i[12];
    end 
    if(N1702) begin
      \nz.mem_347_sv2v_reg  <= data_i[11];
    end 
    if(N1701) begin
      \nz.mem_346_sv2v_reg  <= data_i[10];
    end 
    if(N1700) begin
      \nz.mem_345_sv2v_reg  <= data_i[9];
    end 
    if(N1699) begin
      \nz.mem_344_sv2v_reg  <= data_i[8];
    end 
    if(N1698) begin
      \nz.mem_343_sv2v_reg  <= data_i[7];
    end 
    if(N1697) begin
      \nz.mem_342_sv2v_reg  <= data_i[6];
    end 
    if(N1696) begin
      \nz.mem_341_sv2v_reg  <= data_i[5];
    end 
    if(N1695) begin
      \nz.mem_340_sv2v_reg  <= data_i[4];
    end 
    if(N1694) begin
      \nz.mem_339_sv2v_reg  <= data_i[3];
    end 
    if(N1693) begin
      \nz.mem_338_sv2v_reg  <= data_i[2];
    end 
    if(N1692) begin
      \nz.mem_337_sv2v_reg  <= data_i[1];
    end 
    if(N1691) begin
      \nz.mem_336_sv2v_reg  <= data_i[0];
    end 
    if(N1690) begin
      \nz.mem_335_sv2v_reg  <= data_i[15];
    end 
    if(N1689) begin
      \nz.mem_334_sv2v_reg  <= data_i[14];
    end 
    if(N1688) begin
      \nz.mem_333_sv2v_reg  <= data_i[13];
    end 
    if(N1687) begin
      \nz.mem_332_sv2v_reg  <= data_i[12];
    end 
    if(N1686) begin
      \nz.mem_331_sv2v_reg  <= data_i[11];
    end 
    if(N1685) begin
      \nz.mem_330_sv2v_reg  <= data_i[10];
    end 
    if(N1684) begin
      \nz.mem_329_sv2v_reg  <= data_i[9];
    end 
    if(N1683) begin
      \nz.mem_328_sv2v_reg  <= data_i[8];
    end 
    if(N1682) begin
      \nz.mem_327_sv2v_reg  <= data_i[7];
    end 
    if(N1681) begin
      \nz.mem_326_sv2v_reg  <= data_i[6];
    end 
    if(N1680) begin
      \nz.mem_325_sv2v_reg  <= data_i[5];
    end 
    if(N1679) begin
      \nz.mem_324_sv2v_reg  <= data_i[4];
    end 
    if(N1678) begin
      \nz.mem_323_sv2v_reg  <= data_i[3];
    end 
    if(N1677) begin
      \nz.mem_322_sv2v_reg  <= data_i[2];
    end 
    if(N1676) begin
      \nz.mem_321_sv2v_reg  <= data_i[1];
    end 
    if(N1675) begin
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N1674) begin
      \nz.mem_319_sv2v_reg  <= data_i[15];
    end 
    if(N1673) begin
      \nz.mem_318_sv2v_reg  <= data_i[14];
    end 
    if(N1672) begin
      \nz.mem_317_sv2v_reg  <= data_i[13];
    end 
    if(N1671) begin
      \nz.mem_316_sv2v_reg  <= data_i[12];
    end 
    if(N1670) begin
      \nz.mem_315_sv2v_reg  <= data_i[11];
    end 
    if(N1669) begin
      \nz.mem_314_sv2v_reg  <= data_i[10];
    end 
    if(N1668) begin
      \nz.mem_313_sv2v_reg  <= data_i[9];
    end 
    if(N1667) begin
      \nz.mem_312_sv2v_reg  <= data_i[8];
    end 
    if(N1666) begin
      \nz.mem_311_sv2v_reg  <= data_i[7];
    end 
    if(N1665) begin
      \nz.mem_310_sv2v_reg  <= data_i[6];
    end 
    if(N1664) begin
      \nz.mem_309_sv2v_reg  <= data_i[5];
    end 
    if(N1663) begin
      \nz.mem_308_sv2v_reg  <= data_i[4];
    end 
    if(N1662) begin
      \nz.mem_307_sv2v_reg  <= data_i[3];
    end 
    if(N1661) begin
      \nz.mem_306_sv2v_reg  <= data_i[2];
    end 
    if(N1660) begin
      \nz.mem_305_sv2v_reg  <= data_i[1];
    end 
    if(N1659) begin
      \nz.mem_304_sv2v_reg  <= data_i[0];
    end 
    if(N1658) begin
      \nz.mem_303_sv2v_reg  <= data_i[15];
    end 
    if(N1657) begin
      \nz.mem_302_sv2v_reg  <= data_i[14];
    end 
    if(N1656) begin
      \nz.mem_301_sv2v_reg  <= data_i[13];
    end 
    if(N1655) begin
      \nz.mem_300_sv2v_reg  <= data_i[12];
    end 
    if(N1654) begin
      \nz.mem_299_sv2v_reg  <= data_i[11];
    end 
    if(N1653) begin
      \nz.mem_298_sv2v_reg  <= data_i[10];
    end 
    if(N1652) begin
      \nz.mem_297_sv2v_reg  <= data_i[9];
    end 
    if(N1651) begin
      \nz.mem_296_sv2v_reg  <= data_i[8];
    end 
    if(N1650) begin
      \nz.mem_295_sv2v_reg  <= data_i[7];
    end 
    if(N1649) begin
      \nz.mem_294_sv2v_reg  <= data_i[6];
    end 
    if(N1648) begin
      \nz.mem_293_sv2v_reg  <= data_i[5];
    end 
    if(N1647) begin
      \nz.mem_292_sv2v_reg  <= data_i[4];
    end 
    if(N1646) begin
      \nz.mem_291_sv2v_reg  <= data_i[3];
    end 
    if(N1645) begin
      \nz.mem_290_sv2v_reg  <= data_i[2];
    end 
    if(N1644) begin
      \nz.mem_289_sv2v_reg  <= data_i[1];
    end 
    if(N1643) begin
      \nz.mem_288_sv2v_reg  <= data_i[0];
    end 
    if(N1642) begin
      \nz.mem_287_sv2v_reg  <= data_i[15];
    end 
    if(N1641) begin
      \nz.mem_286_sv2v_reg  <= data_i[14];
    end 
    if(N1640) begin
      \nz.mem_285_sv2v_reg  <= data_i[13];
    end 
    if(N1639) begin
      \nz.mem_284_sv2v_reg  <= data_i[12];
    end 
    if(N1638) begin
      \nz.mem_283_sv2v_reg  <= data_i[11];
    end 
    if(N1637) begin
      \nz.mem_282_sv2v_reg  <= data_i[10];
    end 
    if(N1636) begin
      \nz.mem_281_sv2v_reg  <= data_i[9];
    end 
    if(N1635) begin
      \nz.mem_280_sv2v_reg  <= data_i[8];
    end 
    if(N1634) begin
      \nz.mem_279_sv2v_reg  <= data_i[7];
    end 
    if(N1633) begin
      \nz.mem_278_sv2v_reg  <= data_i[6];
    end 
    if(N1632) begin
      \nz.mem_277_sv2v_reg  <= data_i[5];
    end 
    if(N1631) begin
      \nz.mem_276_sv2v_reg  <= data_i[4];
    end 
    if(N1630) begin
      \nz.mem_275_sv2v_reg  <= data_i[3];
    end 
    if(N1629) begin
      \nz.mem_274_sv2v_reg  <= data_i[2];
    end 
    if(N1628) begin
      \nz.mem_273_sv2v_reg  <= data_i[1];
    end 
    if(N1627) begin
      \nz.mem_272_sv2v_reg  <= data_i[0];
    end 
    if(N1626) begin
      \nz.mem_271_sv2v_reg  <= data_i[15];
    end 
    if(N1625) begin
      \nz.mem_270_sv2v_reg  <= data_i[14];
    end 
    if(N1624) begin
      \nz.mem_269_sv2v_reg  <= data_i[13];
    end 
    if(N1623) begin
      \nz.mem_268_sv2v_reg  <= data_i[12];
    end 
    if(N1622) begin
      \nz.mem_267_sv2v_reg  <= data_i[11];
    end 
    if(N1621) begin
      \nz.mem_266_sv2v_reg  <= data_i[10];
    end 
    if(N1620) begin
      \nz.mem_265_sv2v_reg  <= data_i[9];
    end 
    if(N1619) begin
      \nz.mem_264_sv2v_reg  <= data_i[8];
    end 
    if(N1618) begin
      \nz.mem_263_sv2v_reg  <= data_i[7];
    end 
    if(N1617) begin
      \nz.mem_262_sv2v_reg  <= data_i[6];
    end 
    if(N1616) begin
      \nz.mem_261_sv2v_reg  <= data_i[5];
    end 
    if(N1615) begin
      \nz.mem_260_sv2v_reg  <= data_i[4];
    end 
    if(N1614) begin
      \nz.mem_259_sv2v_reg  <= data_i[3];
    end 
    if(N1613) begin
      \nz.mem_258_sv2v_reg  <= data_i[2];
    end 
    if(N1612) begin
      \nz.mem_257_sv2v_reg  <= data_i[1];
    end 
    if(N1611) begin
      \nz.mem_256_sv2v_reg  <= data_i[0];
    end 
    if(N1610) begin
      \nz.mem_255_sv2v_reg  <= data_i[15];
    end 
    if(N1609) begin
      \nz.mem_254_sv2v_reg  <= data_i[14];
    end 
    if(N1608) begin
      \nz.mem_253_sv2v_reg  <= data_i[13];
    end 
    if(N1607) begin
      \nz.mem_252_sv2v_reg  <= data_i[12];
    end 
    if(N1606) begin
      \nz.mem_251_sv2v_reg  <= data_i[11];
    end 
    if(N1605) begin
      \nz.mem_250_sv2v_reg  <= data_i[10];
    end 
    if(N1604) begin
      \nz.mem_249_sv2v_reg  <= data_i[9];
    end 
    if(N1603) begin
      \nz.mem_248_sv2v_reg  <= data_i[8];
    end 
    if(N1602) begin
      \nz.mem_247_sv2v_reg  <= data_i[7];
    end 
    if(N1601) begin
      \nz.mem_246_sv2v_reg  <= data_i[6];
    end 
    if(N1600) begin
      \nz.mem_245_sv2v_reg  <= data_i[5];
    end 
    if(N1599) begin
      \nz.mem_244_sv2v_reg  <= data_i[4];
    end 
    if(N1598) begin
      \nz.mem_243_sv2v_reg  <= data_i[3];
    end 
    if(N1597) begin
      \nz.mem_242_sv2v_reg  <= data_i[2];
    end 
    if(N1596) begin
      \nz.mem_241_sv2v_reg  <= data_i[1];
    end 
    if(N1595) begin
      \nz.mem_240_sv2v_reg  <= data_i[0];
    end 
    if(N1594) begin
      \nz.mem_239_sv2v_reg  <= data_i[15];
    end 
    if(N1593) begin
      \nz.mem_238_sv2v_reg  <= data_i[14];
    end 
    if(N1592) begin
      \nz.mem_237_sv2v_reg  <= data_i[13];
    end 
    if(N1591) begin
      \nz.mem_236_sv2v_reg  <= data_i[12];
    end 
    if(N1590) begin
      \nz.mem_235_sv2v_reg  <= data_i[11];
    end 
    if(N1589) begin
      \nz.mem_234_sv2v_reg  <= data_i[10];
    end 
    if(N1588) begin
      \nz.mem_233_sv2v_reg  <= data_i[9];
    end 
    if(N1587) begin
      \nz.mem_232_sv2v_reg  <= data_i[8];
    end 
    if(N1586) begin
      \nz.mem_231_sv2v_reg  <= data_i[7];
    end 
    if(N1585) begin
      \nz.mem_230_sv2v_reg  <= data_i[6];
    end 
    if(N1584) begin
      \nz.mem_229_sv2v_reg  <= data_i[5];
    end 
    if(N1583) begin
      \nz.mem_228_sv2v_reg  <= data_i[4];
    end 
    if(N1582) begin
      \nz.mem_227_sv2v_reg  <= data_i[3];
    end 
    if(N1581) begin
      \nz.mem_226_sv2v_reg  <= data_i[2];
    end 
    if(N1580) begin
      \nz.mem_225_sv2v_reg  <= data_i[1];
    end 
    if(N1579) begin
      \nz.mem_224_sv2v_reg  <= data_i[0];
    end 
    if(N1578) begin
      \nz.mem_223_sv2v_reg  <= data_i[15];
    end 
    if(N1577) begin
      \nz.mem_222_sv2v_reg  <= data_i[14];
    end 
    if(N1576) begin
      \nz.mem_221_sv2v_reg  <= data_i[13];
    end 
    if(N1575) begin
      \nz.mem_220_sv2v_reg  <= data_i[12];
    end 
    if(N1574) begin
      \nz.mem_219_sv2v_reg  <= data_i[11];
    end 
    if(N1573) begin
      \nz.mem_218_sv2v_reg  <= data_i[10];
    end 
    if(N1572) begin
      \nz.mem_217_sv2v_reg  <= data_i[9];
    end 
    if(N1571) begin
      \nz.mem_216_sv2v_reg  <= data_i[8];
    end 
    if(N1570) begin
      \nz.mem_215_sv2v_reg  <= data_i[7];
    end 
    if(N1569) begin
      \nz.mem_214_sv2v_reg  <= data_i[6];
    end 
    if(N1568) begin
      \nz.mem_213_sv2v_reg  <= data_i[5];
    end 
    if(N1567) begin
      \nz.mem_212_sv2v_reg  <= data_i[4];
    end 
    if(N1566) begin
      \nz.mem_211_sv2v_reg  <= data_i[3];
    end 
    if(N1565) begin
      \nz.mem_210_sv2v_reg  <= data_i[2];
    end 
    if(N1564) begin
      \nz.mem_209_sv2v_reg  <= data_i[1];
    end 
    if(N1563) begin
      \nz.mem_208_sv2v_reg  <= data_i[0];
    end 
    if(N1562) begin
      \nz.mem_207_sv2v_reg  <= data_i[15];
    end 
    if(N1561) begin
      \nz.mem_206_sv2v_reg  <= data_i[14];
    end 
    if(N1560) begin
      \nz.mem_205_sv2v_reg  <= data_i[13];
    end 
    if(N1559) begin
      \nz.mem_204_sv2v_reg  <= data_i[12];
    end 
    if(N1558) begin
      \nz.mem_203_sv2v_reg  <= data_i[11];
    end 
    if(N1557) begin
      \nz.mem_202_sv2v_reg  <= data_i[10];
    end 
    if(N1556) begin
      \nz.mem_201_sv2v_reg  <= data_i[9];
    end 
    if(N1555) begin
      \nz.mem_200_sv2v_reg  <= data_i[8];
    end 
    if(N1554) begin
      \nz.mem_199_sv2v_reg  <= data_i[7];
    end 
    if(N1553) begin
      \nz.mem_198_sv2v_reg  <= data_i[6];
    end 
    if(N1552) begin
      \nz.mem_197_sv2v_reg  <= data_i[5];
    end 
    if(N1551) begin
      \nz.mem_196_sv2v_reg  <= data_i[4];
    end 
    if(N1550) begin
      \nz.mem_195_sv2v_reg  <= data_i[3];
    end 
    if(N1549) begin
      \nz.mem_194_sv2v_reg  <= data_i[2];
    end 
    if(N1548) begin
      \nz.mem_193_sv2v_reg  <= data_i[1];
    end 
    if(N1547) begin
      \nz.mem_192_sv2v_reg  <= data_i[0];
    end 
    if(N1546) begin
      \nz.mem_191_sv2v_reg  <= data_i[15];
    end 
    if(N1545) begin
      \nz.mem_190_sv2v_reg  <= data_i[14];
    end 
    if(N1544) begin
      \nz.mem_189_sv2v_reg  <= data_i[13];
    end 
    if(N1543) begin
      \nz.mem_188_sv2v_reg  <= data_i[12];
    end 
    if(N1542) begin
      \nz.mem_187_sv2v_reg  <= data_i[11];
    end 
    if(N1541) begin
      \nz.mem_186_sv2v_reg  <= data_i[10];
    end 
    if(N1540) begin
      \nz.mem_185_sv2v_reg  <= data_i[9];
    end 
    if(N1539) begin
      \nz.mem_184_sv2v_reg  <= data_i[8];
    end 
    if(N1538) begin
      \nz.mem_183_sv2v_reg  <= data_i[7];
    end 
    if(N1537) begin
      \nz.mem_182_sv2v_reg  <= data_i[6];
    end 
    if(N1536) begin
      \nz.mem_181_sv2v_reg  <= data_i[5];
    end 
    if(N1535) begin
      \nz.mem_180_sv2v_reg  <= data_i[4];
    end 
    if(N1534) begin
      \nz.mem_179_sv2v_reg  <= data_i[3];
    end 
    if(N1533) begin
      \nz.mem_178_sv2v_reg  <= data_i[2];
    end 
    if(N1532) begin
      \nz.mem_177_sv2v_reg  <= data_i[1];
    end 
    if(N1531) begin
      \nz.mem_176_sv2v_reg  <= data_i[0];
    end 
    if(N1530) begin
      \nz.mem_175_sv2v_reg  <= data_i[15];
    end 
    if(N1529) begin
      \nz.mem_174_sv2v_reg  <= data_i[14];
    end 
    if(N1528) begin
      \nz.mem_173_sv2v_reg  <= data_i[13];
    end 
    if(N1527) begin
      \nz.mem_172_sv2v_reg  <= data_i[12];
    end 
    if(N1526) begin
      \nz.mem_171_sv2v_reg  <= data_i[11];
    end 
    if(N1525) begin
      \nz.mem_170_sv2v_reg  <= data_i[10];
    end 
    if(N1524) begin
      \nz.mem_169_sv2v_reg  <= data_i[9];
    end 
    if(N1523) begin
      \nz.mem_168_sv2v_reg  <= data_i[8];
    end 
    if(N1522) begin
      \nz.mem_167_sv2v_reg  <= data_i[7];
    end 
    if(N1521) begin
      \nz.mem_166_sv2v_reg  <= data_i[6];
    end 
    if(N1520) begin
      \nz.mem_165_sv2v_reg  <= data_i[5];
    end 
    if(N1519) begin
      \nz.mem_164_sv2v_reg  <= data_i[4];
    end 
    if(N1518) begin
      \nz.mem_163_sv2v_reg  <= data_i[3];
    end 
    if(N1517) begin
      \nz.mem_162_sv2v_reg  <= data_i[2];
    end 
    if(N1516) begin
      \nz.mem_161_sv2v_reg  <= data_i[1];
    end 
    if(N1515) begin
      \nz.mem_160_sv2v_reg  <= data_i[0];
    end 
    if(N1514) begin
      \nz.mem_159_sv2v_reg  <= data_i[15];
    end 
    if(N1513) begin
      \nz.mem_158_sv2v_reg  <= data_i[14];
    end 
    if(N1512) begin
      \nz.mem_157_sv2v_reg  <= data_i[13];
    end 
    if(N1511) begin
      \nz.mem_156_sv2v_reg  <= data_i[12];
    end 
    if(N1510) begin
      \nz.mem_155_sv2v_reg  <= data_i[11];
    end 
    if(N1509) begin
      \nz.mem_154_sv2v_reg  <= data_i[10];
    end 
    if(N1508) begin
      \nz.mem_153_sv2v_reg  <= data_i[9];
    end 
    if(N1507) begin
      \nz.mem_152_sv2v_reg  <= data_i[8];
    end 
    if(N1506) begin
      \nz.mem_151_sv2v_reg  <= data_i[7];
    end 
    if(N1505) begin
      \nz.mem_150_sv2v_reg  <= data_i[6];
    end 
    if(N1504) begin
      \nz.mem_149_sv2v_reg  <= data_i[5];
    end 
    if(N1503) begin
      \nz.mem_148_sv2v_reg  <= data_i[4];
    end 
    if(N1502) begin
      \nz.mem_147_sv2v_reg  <= data_i[3];
    end 
    if(N1501) begin
      \nz.mem_146_sv2v_reg  <= data_i[2];
    end 
    if(N1500) begin
      \nz.mem_145_sv2v_reg  <= data_i[1];
    end 
    if(N1499) begin
      \nz.mem_144_sv2v_reg  <= data_i[0];
    end 
    if(N1498) begin
      \nz.mem_143_sv2v_reg  <= data_i[15];
    end 
    if(N1497) begin
      \nz.mem_142_sv2v_reg  <= data_i[14];
    end 
    if(N1496) begin
      \nz.mem_141_sv2v_reg  <= data_i[13];
    end 
    if(N1495) begin
      \nz.mem_140_sv2v_reg  <= data_i[12];
    end 
    if(N1494) begin
      \nz.mem_139_sv2v_reg  <= data_i[11];
    end 
    if(N1493) begin
      \nz.mem_138_sv2v_reg  <= data_i[10];
    end 
    if(N1492) begin
      \nz.mem_137_sv2v_reg  <= data_i[9];
    end 
    if(N1491) begin
      \nz.mem_136_sv2v_reg  <= data_i[8];
    end 
    if(N1490) begin
      \nz.mem_135_sv2v_reg  <= data_i[7];
    end 
    if(N1489) begin
      \nz.mem_134_sv2v_reg  <= data_i[6];
    end 
    if(N1488) begin
      \nz.mem_133_sv2v_reg  <= data_i[5];
    end 
    if(N1487) begin
      \nz.mem_132_sv2v_reg  <= data_i[4];
    end 
    if(N1486) begin
      \nz.mem_131_sv2v_reg  <= data_i[3];
    end 
    if(N1485) begin
      \nz.mem_130_sv2v_reg  <= data_i[2];
    end 
    if(N1484) begin
      \nz.mem_129_sv2v_reg  <= data_i[1];
    end 
    if(N1483) begin
      \nz.mem_128_sv2v_reg  <= data_i[0];
    end 
    if(N1482) begin
      \nz.mem_127_sv2v_reg  <= data_i[15];
    end 
    if(N1481) begin
      \nz.mem_126_sv2v_reg  <= data_i[14];
    end 
    if(N1480) begin
      \nz.mem_125_sv2v_reg  <= data_i[13];
    end 
    if(N1479) begin
      \nz.mem_124_sv2v_reg  <= data_i[12];
    end 
    if(N1478) begin
      \nz.mem_123_sv2v_reg  <= data_i[11];
    end 
    if(N1477) begin
      \nz.mem_122_sv2v_reg  <= data_i[10];
    end 
    if(N1476) begin
      \nz.mem_121_sv2v_reg  <= data_i[9];
    end 
    if(N1475) begin
      \nz.mem_120_sv2v_reg  <= data_i[8];
    end 
    if(N1474) begin
      \nz.mem_119_sv2v_reg  <= data_i[7];
    end 
    if(N1473) begin
      \nz.mem_118_sv2v_reg  <= data_i[6];
    end 
    if(N1472) begin
      \nz.mem_117_sv2v_reg  <= data_i[5];
    end 
    if(N1471) begin
      \nz.mem_116_sv2v_reg  <= data_i[4];
    end 
    if(N1470) begin
      \nz.mem_115_sv2v_reg  <= data_i[3];
    end 
    if(N1469) begin
      \nz.mem_114_sv2v_reg  <= data_i[2];
    end 
    if(N1468) begin
      \nz.mem_113_sv2v_reg  <= data_i[1];
    end 
    if(N1467) begin
      \nz.mem_112_sv2v_reg  <= data_i[0];
    end 
    if(N1466) begin
      \nz.mem_111_sv2v_reg  <= data_i[15];
    end 
    if(N1465) begin
      \nz.mem_110_sv2v_reg  <= data_i[14];
    end 
    if(N1464) begin
      \nz.mem_109_sv2v_reg  <= data_i[13];
    end 
    if(N1463) begin
      \nz.mem_108_sv2v_reg  <= data_i[12];
    end 
    if(N1462) begin
      \nz.mem_107_sv2v_reg  <= data_i[11];
    end 
    if(N1461) begin
      \nz.mem_106_sv2v_reg  <= data_i[10];
    end 
    if(N1460) begin
      \nz.mem_105_sv2v_reg  <= data_i[9];
    end 
    if(N1459) begin
      \nz.mem_104_sv2v_reg  <= data_i[8];
    end 
    if(N1458) begin
      \nz.mem_103_sv2v_reg  <= data_i[7];
    end 
    if(N1457) begin
      \nz.mem_102_sv2v_reg  <= data_i[6];
    end 
    if(N1456) begin
      \nz.mem_101_sv2v_reg  <= data_i[5];
    end 
    if(N1455) begin
      \nz.mem_100_sv2v_reg  <= data_i[4];
    end 
    if(N1454) begin
      \nz.mem_99_sv2v_reg  <= data_i[3];
    end 
    if(N1453) begin
      \nz.mem_98_sv2v_reg  <= data_i[2];
    end 
    if(N1452) begin
      \nz.mem_97_sv2v_reg  <= data_i[1];
    end 
    if(N1451) begin
      \nz.mem_96_sv2v_reg  <= data_i[0];
    end 
    if(N1450) begin
      \nz.mem_95_sv2v_reg  <= data_i[15];
    end 
    if(N1449) begin
      \nz.mem_94_sv2v_reg  <= data_i[14];
    end 
    if(N1448) begin
      \nz.mem_93_sv2v_reg  <= data_i[13];
    end 
    if(N1447) begin
      \nz.mem_92_sv2v_reg  <= data_i[12];
    end 
    if(N1446) begin
      \nz.mem_91_sv2v_reg  <= data_i[11];
    end 
    if(N1445) begin
      \nz.mem_90_sv2v_reg  <= data_i[10];
    end 
    if(N1444) begin
      \nz.mem_89_sv2v_reg  <= data_i[9];
    end 
    if(N1443) begin
      \nz.mem_88_sv2v_reg  <= data_i[8];
    end 
    if(N1442) begin
      \nz.mem_87_sv2v_reg  <= data_i[7];
    end 
    if(N1441) begin
      \nz.mem_86_sv2v_reg  <= data_i[6];
    end 
    if(N1440) begin
      \nz.mem_85_sv2v_reg  <= data_i[5];
    end 
    if(N1439) begin
      \nz.mem_84_sv2v_reg  <= data_i[4];
    end 
    if(N1438) begin
      \nz.mem_83_sv2v_reg  <= data_i[3];
    end 
    if(N1437) begin
      \nz.mem_82_sv2v_reg  <= data_i[2];
    end 
    if(N1436) begin
      \nz.mem_81_sv2v_reg  <= data_i[1];
    end 
    if(N1435) begin
      \nz.mem_80_sv2v_reg  <= data_i[0];
    end 
    if(N1434) begin
      \nz.mem_79_sv2v_reg  <= data_i[15];
    end 
    if(N1433) begin
      \nz.mem_78_sv2v_reg  <= data_i[14];
    end 
    if(N1432) begin
      \nz.mem_77_sv2v_reg  <= data_i[13];
    end 
    if(N1431) begin
      \nz.mem_76_sv2v_reg  <= data_i[12];
    end 
    if(N1430) begin
      \nz.mem_75_sv2v_reg  <= data_i[11];
    end 
    if(N1429) begin
      \nz.mem_74_sv2v_reg  <= data_i[10];
    end 
    if(N1428) begin
      \nz.mem_73_sv2v_reg  <= data_i[9];
    end 
    if(N1427) begin
      \nz.mem_72_sv2v_reg  <= data_i[8];
    end 
    if(N1426) begin
      \nz.mem_71_sv2v_reg  <= data_i[7];
    end 
    if(N1425) begin
      \nz.mem_70_sv2v_reg  <= data_i[6];
    end 
    if(N1424) begin
      \nz.mem_69_sv2v_reg  <= data_i[5];
    end 
    if(N1423) begin
      \nz.mem_68_sv2v_reg  <= data_i[4];
    end 
    if(N1422) begin
      \nz.mem_67_sv2v_reg  <= data_i[3];
    end 
    if(N1421) begin
      \nz.mem_66_sv2v_reg  <= data_i[2];
    end 
    if(N1420) begin
      \nz.mem_65_sv2v_reg  <= data_i[1];
    end 
    if(N1419) begin
      \nz.mem_64_sv2v_reg  <= data_i[0];
    end 
    if(N1418) begin
      \nz.mem_63_sv2v_reg  <= data_i[15];
    end 
    if(N1417) begin
      \nz.mem_62_sv2v_reg  <= data_i[14];
    end 
    if(N1416) begin
      \nz.mem_61_sv2v_reg  <= data_i[13];
    end 
    if(N1415) begin
      \nz.mem_60_sv2v_reg  <= data_i[12];
    end 
    if(N1414) begin
      \nz.mem_59_sv2v_reg  <= data_i[11];
    end 
    if(N1413) begin
      \nz.mem_58_sv2v_reg  <= data_i[10];
    end 
    if(N1412) begin
      \nz.mem_57_sv2v_reg  <= data_i[9];
    end 
    if(N1411) begin
      \nz.mem_56_sv2v_reg  <= data_i[8];
    end 
    if(N1410) begin
      \nz.mem_55_sv2v_reg  <= data_i[7];
    end 
    if(N1409) begin
      \nz.mem_54_sv2v_reg  <= data_i[6];
    end 
    if(N1408) begin
      \nz.mem_53_sv2v_reg  <= data_i[5];
    end 
    if(N1407) begin
      \nz.mem_52_sv2v_reg  <= data_i[4];
    end 
    if(N1406) begin
      \nz.mem_51_sv2v_reg  <= data_i[3];
    end 
    if(N1405) begin
      \nz.mem_50_sv2v_reg  <= data_i[2];
    end 
    if(N1404) begin
      \nz.mem_49_sv2v_reg  <= data_i[1];
    end 
    if(N1403) begin
      \nz.mem_48_sv2v_reg  <= data_i[0];
    end 
    if(N1402) begin
      \nz.mem_47_sv2v_reg  <= data_i[15];
    end 
    if(N1401) begin
      \nz.mem_46_sv2v_reg  <= data_i[14];
    end 
    if(N1400) begin
      \nz.mem_45_sv2v_reg  <= data_i[13];
    end 
    if(N1399) begin
      \nz.mem_44_sv2v_reg  <= data_i[12];
    end 
    if(N1398) begin
      \nz.mem_43_sv2v_reg  <= data_i[11];
    end 
    if(N1397) begin
      \nz.mem_42_sv2v_reg  <= data_i[10];
    end 
    if(N1396) begin
      \nz.mem_41_sv2v_reg  <= data_i[9];
    end 
    if(N1395) begin
      \nz.mem_40_sv2v_reg  <= data_i[8];
    end 
    if(N1394) begin
      \nz.mem_39_sv2v_reg  <= data_i[7];
    end 
    if(N1393) begin
      \nz.mem_38_sv2v_reg  <= data_i[6];
    end 
    if(N1392) begin
      \nz.mem_37_sv2v_reg  <= data_i[5];
    end 
    if(N1391) begin
      \nz.mem_36_sv2v_reg  <= data_i[4];
    end 
    if(N1390) begin
      \nz.mem_35_sv2v_reg  <= data_i[3];
    end 
    if(N1389) begin
      \nz.mem_34_sv2v_reg  <= data_i[2];
    end 
    if(N1388) begin
      \nz.mem_33_sv2v_reg  <= data_i[1];
    end 
    if(N1387) begin
      \nz.mem_32_sv2v_reg  <= data_i[0];
    end 
    if(N1386) begin
      \nz.mem_31_sv2v_reg  <= data_i[15];
    end 
    if(N1385) begin
      \nz.mem_30_sv2v_reg  <= data_i[14];
    end 
    if(N1384) begin
      \nz.mem_29_sv2v_reg  <= data_i[13];
    end 
    if(N1383) begin
      \nz.mem_28_sv2v_reg  <= data_i[12];
    end 
    if(N1382) begin
      \nz.mem_27_sv2v_reg  <= data_i[11];
    end 
    if(N1381) begin
      \nz.mem_26_sv2v_reg  <= data_i[10];
    end 
    if(N1380) begin
      \nz.mem_25_sv2v_reg  <= data_i[9];
    end 
    if(N1379) begin
      \nz.mem_24_sv2v_reg  <= data_i[8];
    end 
    if(N1378) begin
      \nz.mem_23_sv2v_reg  <= data_i[7];
    end 
    if(N1377) begin
      \nz.mem_22_sv2v_reg  <= data_i[6];
    end 
    if(N1376) begin
      \nz.mem_21_sv2v_reg  <= data_i[5];
    end 
    if(N1375) begin
      \nz.mem_20_sv2v_reg  <= data_i[4];
    end 
    if(N1374) begin
      \nz.mem_19_sv2v_reg  <= data_i[3];
    end 
    if(N1373) begin
      \nz.mem_18_sv2v_reg  <= data_i[2];
    end 
    if(N1372) begin
      \nz.mem_17_sv2v_reg  <= data_i[1];
    end 
    if(N1371) begin
      \nz.mem_16_sv2v_reg  <= data_i[0];
    end 
    if(N1370) begin
      \nz.mem_15_sv2v_reg  <= data_i[15];
    end 
    if(N1369) begin
      \nz.mem_14_sv2v_reg  <= data_i[14];
    end 
    if(N1368) begin
      \nz.mem_13_sv2v_reg  <= data_i[13];
    end 
    if(N1367) begin
      \nz.mem_12_sv2v_reg  <= data_i[12];
    end 
    if(N1366) begin
      \nz.mem_11_sv2v_reg  <= data_i[11];
    end 
    if(N1365) begin
      \nz.mem_10_sv2v_reg  <= data_i[10];
    end 
    if(N1364) begin
      \nz.mem_9_sv2v_reg  <= data_i[9];
    end 
    if(N1363) begin
      \nz.mem_8_sv2v_reg  <= data_i[8];
    end 
    if(N1362) begin
      \nz.mem_7_sv2v_reg  <= data_i[7];
    end 
    if(N1361) begin
      \nz.mem_6_sv2v_reg  <= data_i[6];
    end 
    if(N1360) begin
      \nz.mem_5_sv2v_reg  <= data_i[5];
    end 
    if(N1359) begin
      \nz.mem_4_sv2v_reg  <= data_i[4];
    end 
    if(N1358) begin
      \nz.mem_3_sv2v_reg  <= data_i[3];
    end 
    if(N1357) begin
      \nz.mem_2_sv2v_reg  <= data_i[2];
    end 
    if(N1356) begin
      \nz.mem_1_sv2v_reg  <= data_i[1];
    end 
    if(N1355) begin
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p16_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [15:0] data_i;
  input [5:0] addr_i;
  input [15:0] w_mask_i;
  output [15:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [15:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p16_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p4_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [3:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire t_1__3_,t_1__2_,t_1__1_,t_1__0_;
  assign t_1__3_ = i[0] | 1'b0;
  assign t_1__2_ = i[1] | i[0];
  assign t_1__1_ = i[2] | i[1];
  assign t_1__0_ = i[3] | i[2];
  assign o[0] = t_1__3_ | 1'b0;
  assign o[1] = t_1__2_ | 1'b0;
  assign o[2] = t_1__1_ | t_1__3_;
  assign o[3] = t_1__0_ | t_1__2_;

endmodule



module bsg_priority_encode_one_hot_out_width_p4_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [3:0] i;
  output [3:0] o;
  output v_o;
  wire [3:0] o;
  wire v_o,N0,N1,N2;
  wire [2:1] scan_lo;

  bsg_scan_width_p4_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, scan_lo, o[0:0] })
  );

  assign o[3] = v_o & N0;
  assign N0 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N1;
  assign N1 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N2;
  assign N2 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p4_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o;
  wire v_o,v_1__0_;
  assign v_1__0_ = i[1] | i[0];
  assign addr_o[1] = i[3] | i[2];
  assign v_o = addr_o[1] | v_1__0_;
  assign addr_o[0] = i[1] | i[3];

endmodule



module bsg_priority_encode_width_p4_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o;
  wire v_o;
  wire [3:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p4_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p4_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o)
  );


endmodule



module bsg_dff_en_width_p7_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  input en_i;
  wire [6:0] data_o;
  reg data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,
  data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p7
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [6:0] data_i;
  output [6:0] data_o;
  input clk_i;
  input en_i;
  wire [6:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p7_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p7_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,\nz.read_en ,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,
  \nz.llr.read_en_r ,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141;
  wire [5:0] \nz.addr_r ;
  wire [447:0] \nz.mem ;
  reg \nz.addr_r_5_sv2v_reg ,\nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,
  \nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,\nz.mem_447_sv2v_reg ,
  \nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,
  \nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,
  \nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,
  \nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,
  \nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,
  \nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,
  \nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,
  \nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,
  \nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,
  \nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,
  \nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,
  \nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,
  \nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,
  \nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,
  \nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,
  \nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,
  \nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,
  \nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,
  \nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,
  \nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,
  \nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,
  \nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,
  \nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,
  \nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,
  \nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,
  \nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,
  \nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,
  \nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,
  \nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,
  \nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,
  \nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,
  \nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,
  \nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,
  \nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,
  \nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,
  \nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,
  \nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,
  \nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,
  \nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,
  \nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,
  \nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,
  \nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,
  \nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,
  \nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,
  \nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,
  \nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,
  \nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,
  \nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,
  \nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,
  \nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,
  \nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,
  \nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,
  \nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,
  \nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,
  \nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,
  \nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,
  \nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,
  \nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,
  \nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,
  \nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,
  \nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,
  \nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,
  \nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,
  \nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,
  \nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,
  \nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,
  \nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,
  \nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,
  \nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,
  \nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,
  \nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,
  \nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,
  \nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,
  \nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,
  \nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,
  \nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,
  \nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,
  \nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,
  \nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,
  \nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,
  \nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,
  \nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,
  \nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,
  \nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,
  \nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,
  \nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,
  \nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,
  \nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,
  \nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,
  \nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,
  \nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,
  \nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,
  \nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,
  \nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,
  \nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,
  \nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,
  \nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,
  \nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,
  \nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,
  \nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,
  \nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,
  \nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,
  \nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,
  \nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,
  \nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,
  \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,
  \nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,
  \nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,
  \nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,
  \nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,
  \nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,
  \nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,
  \nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [6] = (N82)? \nz.mem [6] : 
                            (N84)? \nz.mem [13] : 
                            (N86)? \nz.mem [20] : 
                            (N88)? \nz.mem [27] : 
                            (N90)? \nz.mem [34] : 
                            (N92)? \nz.mem [41] : 
                            (N94)? \nz.mem [48] : 
                            (N96)? \nz.mem [55] : 
                            (N98)? \nz.mem [62] : 
                            (N100)? \nz.mem [69] : 
                            (N102)? \nz.mem [76] : 
                            (N104)? \nz.mem [83] : 
                            (N106)? \nz.mem [90] : 
                            (N108)? \nz.mem [97] : 
                            (N110)? \nz.mem [104] : 
                            (N112)? \nz.mem [111] : 
                            (N114)? \nz.mem [118] : 
                            (N116)? \nz.mem [125] : 
                            (N118)? \nz.mem [132] : 
                            (N120)? \nz.mem [139] : 
                            (N122)? \nz.mem [146] : 
                            (N124)? \nz.mem [153] : 
                            (N126)? \nz.mem [160] : 
                            (N128)? \nz.mem [167] : 
                            (N130)? \nz.mem [174] : 
                            (N132)? \nz.mem [181] : 
                            (N134)? \nz.mem [188] : 
                            (N136)? \nz.mem [195] : 
                            (N138)? \nz.mem [202] : 
                            (N140)? \nz.mem [209] : 
                            (N142)? \nz.mem [216] : 
                            (N144)? \nz.mem [223] : 
                            (N83)? \nz.mem [230] : 
                            (N85)? \nz.mem [237] : 
                            (N87)? \nz.mem [244] : 
                            (N89)? \nz.mem [251] : 
                            (N91)? \nz.mem [258] : 
                            (N93)? \nz.mem [265] : 
                            (N95)? \nz.mem [272] : 
                            (N97)? \nz.mem [279] : 
                            (N99)? \nz.mem [286] : 
                            (N101)? \nz.mem [293] : 
                            (N103)? \nz.mem [300] : 
                            (N105)? \nz.mem [307] : 
                            (N107)? \nz.mem [314] : 
                            (N109)? \nz.mem [321] : 
                            (N111)? \nz.mem [328] : 
                            (N113)? \nz.mem [335] : 
                            (N115)? \nz.mem [342] : 
                            (N117)? \nz.mem [349] : 
                            (N119)? \nz.mem [356] : 
                            (N121)? \nz.mem [363] : 
                            (N123)? \nz.mem [370] : 
                            (N125)? \nz.mem [377] : 
                            (N127)? \nz.mem [384] : 
                            (N129)? \nz.mem [391] : 
                            (N131)? \nz.mem [398] : 
                            (N133)? \nz.mem [405] : 
                            (N135)? \nz.mem [412] : 
                            (N137)? \nz.mem [419] : 
                            (N139)? \nz.mem [426] : 
                            (N141)? \nz.mem [433] : 
                            (N143)? \nz.mem [440] : 
                            (N145)? \nz.mem [447] : 1'b0;
  assign \nz.data_out [5] = (N82)? \nz.mem [5] : 
                            (N84)? \nz.mem [12] : 
                            (N86)? \nz.mem [19] : 
                            (N88)? \nz.mem [26] : 
                            (N90)? \nz.mem [33] : 
                            (N92)? \nz.mem [40] : 
                            (N94)? \nz.mem [47] : 
                            (N96)? \nz.mem [54] : 
                            (N98)? \nz.mem [61] : 
                            (N100)? \nz.mem [68] : 
                            (N102)? \nz.mem [75] : 
                            (N104)? \nz.mem [82] : 
                            (N106)? \nz.mem [89] : 
                            (N108)? \nz.mem [96] : 
                            (N110)? \nz.mem [103] : 
                            (N112)? \nz.mem [110] : 
                            (N114)? \nz.mem [117] : 
                            (N116)? \nz.mem [124] : 
                            (N118)? \nz.mem [131] : 
                            (N120)? \nz.mem [138] : 
                            (N122)? \nz.mem [145] : 
                            (N124)? \nz.mem [152] : 
                            (N126)? \nz.mem [159] : 
                            (N128)? \nz.mem [166] : 
                            (N130)? \nz.mem [173] : 
                            (N132)? \nz.mem [180] : 
                            (N134)? \nz.mem [187] : 
                            (N136)? \nz.mem [194] : 
                            (N138)? \nz.mem [201] : 
                            (N140)? \nz.mem [208] : 
                            (N142)? \nz.mem [215] : 
                            (N144)? \nz.mem [222] : 
                            (N83)? \nz.mem [229] : 
                            (N85)? \nz.mem [236] : 
                            (N87)? \nz.mem [243] : 
                            (N89)? \nz.mem [250] : 
                            (N91)? \nz.mem [257] : 
                            (N93)? \nz.mem [264] : 
                            (N95)? \nz.mem [271] : 
                            (N97)? \nz.mem [278] : 
                            (N99)? \nz.mem [285] : 
                            (N101)? \nz.mem [292] : 
                            (N103)? \nz.mem [299] : 
                            (N105)? \nz.mem [306] : 
                            (N107)? \nz.mem [313] : 
                            (N109)? \nz.mem [320] : 
                            (N111)? \nz.mem [327] : 
                            (N113)? \nz.mem [334] : 
                            (N115)? \nz.mem [341] : 
                            (N117)? \nz.mem [348] : 
                            (N119)? \nz.mem [355] : 
                            (N121)? \nz.mem [362] : 
                            (N123)? \nz.mem [369] : 
                            (N125)? \nz.mem [376] : 
                            (N127)? \nz.mem [383] : 
                            (N129)? \nz.mem [390] : 
                            (N131)? \nz.mem [397] : 
                            (N133)? \nz.mem [404] : 
                            (N135)? \nz.mem [411] : 
                            (N137)? \nz.mem [418] : 
                            (N139)? \nz.mem [425] : 
                            (N141)? \nz.mem [432] : 
                            (N143)? \nz.mem [439] : 
                            (N145)? \nz.mem [446] : 1'b0;
  assign \nz.data_out [4] = (N82)? \nz.mem [4] : 
                            (N84)? \nz.mem [11] : 
                            (N86)? \nz.mem [18] : 
                            (N88)? \nz.mem [25] : 
                            (N90)? \nz.mem [32] : 
                            (N92)? \nz.mem [39] : 
                            (N94)? \nz.mem [46] : 
                            (N96)? \nz.mem [53] : 
                            (N98)? \nz.mem [60] : 
                            (N100)? \nz.mem [67] : 
                            (N102)? \nz.mem [74] : 
                            (N104)? \nz.mem [81] : 
                            (N106)? \nz.mem [88] : 
                            (N108)? \nz.mem [95] : 
                            (N110)? \nz.mem [102] : 
                            (N112)? \nz.mem [109] : 
                            (N114)? \nz.mem [116] : 
                            (N116)? \nz.mem [123] : 
                            (N118)? \nz.mem [130] : 
                            (N120)? \nz.mem [137] : 
                            (N122)? \nz.mem [144] : 
                            (N124)? \nz.mem [151] : 
                            (N126)? \nz.mem [158] : 
                            (N128)? \nz.mem [165] : 
                            (N130)? \nz.mem [172] : 
                            (N132)? \nz.mem [179] : 
                            (N134)? \nz.mem [186] : 
                            (N136)? \nz.mem [193] : 
                            (N138)? \nz.mem [200] : 
                            (N140)? \nz.mem [207] : 
                            (N142)? \nz.mem [214] : 
                            (N144)? \nz.mem [221] : 
                            (N83)? \nz.mem [228] : 
                            (N85)? \nz.mem [235] : 
                            (N87)? \nz.mem [242] : 
                            (N89)? \nz.mem [249] : 
                            (N91)? \nz.mem [256] : 
                            (N93)? \nz.mem [263] : 
                            (N95)? \nz.mem [270] : 
                            (N97)? \nz.mem [277] : 
                            (N99)? \nz.mem [284] : 
                            (N101)? \nz.mem [291] : 
                            (N103)? \nz.mem [298] : 
                            (N105)? \nz.mem [305] : 
                            (N107)? \nz.mem [312] : 
                            (N109)? \nz.mem [319] : 
                            (N111)? \nz.mem [326] : 
                            (N113)? \nz.mem [333] : 
                            (N115)? \nz.mem [340] : 
                            (N117)? \nz.mem [347] : 
                            (N119)? \nz.mem [354] : 
                            (N121)? \nz.mem [361] : 
                            (N123)? \nz.mem [368] : 
                            (N125)? \nz.mem [375] : 
                            (N127)? \nz.mem [382] : 
                            (N129)? \nz.mem [389] : 
                            (N131)? \nz.mem [396] : 
                            (N133)? \nz.mem [403] : 
                            (N135)? \nz.mem [410] : 
                            (N137)? \nz.mem [417] : 
                            (N139)? \nz.mem [424] : 
                            (N141)? \nz.mem [431] : 
                            (N143)? \nz.mem [438] : 
                            (N145)? \nz.mem [445] : 1'b0;
  assign \nz.data_out [3] = (N82)? \nz.mem [3] : 
                            (N84)? \nz.mem [10] : 
                            (N86)? \nz.mem [17] : 
                            (N88)? \nz.mem [24] : 
                            (N90)? \nz.mem [31] : 
                            (N92)? \nz.mem [38] : 
                            (N94)? \nz.mem [45] : 
                            (N96)? \nz.mem [52] : 
                            (N98)? \nz.mem [59] : 
                            (N100)? \nz.mem [66] : 
                            (N102)? \nz.mem [73] : 
                            (N104)? \nz.mem [80] : 
                            (N106)? \nz.mem [87] : 
                            (N108)? \nz.mem [94] : 
                            (N110)? \nz.mem [101] : 
                            (N112)? \nz.mem [108] : 
                            (N114)? \nz.mem [115] : 
                            (N116)? \nz.mem [122] : 
                            (N118)? \nz.mem [129] : 
                            (N120)? \nz.mem [136] : 
                            (N122)? \nz.mem [143] : 
                            (N124)? \nz.mem [150] : 
                            (N126)? \nz.mem [157] : 
                            (N128)? \nz.mem [164] : 
                            (N130)? \nz.mem [171] : 
                            (N132)? \nz.mem [178] : 
                            (N134)? \nz.mem [185] : 
                            (N136)? \nz.mem [192] : 
                            (N138)? \nz.mem [199] : 
                            (N140)? \nz.mem [206] : 
                            (N142)? \nz.mem [213] : 
                            (N144)? \nz.mem [220] : 
                            (N83)? \nz.mem [227] : 
                            (N85)? \nz.mem [234] : 
                            (N87)? \nz.mem [241] : 
                            (N89)? \nz.mem [248] : 
                            (N91)? \nz.mem [255] : 
                            (N93)? \nz.mem [262] : 
                            (N95)? \nz.mem [269] : 
                            (N97)? \nz.mem [276] : 
                            (N99)? \nz.mem [283] : 
                            (N101)? \nz.mem [290] : 
                            (N103)? \nz.mem [297] : 
                            (N105)? \nz.mem [304] : 
                            (N107)? \nz.mem [311] : 
                            (N109)? \nz.mem [318] : 
                            (N111)? \nz.mem [325] : 
                            (N113)? \nz.mem [332] : 
                            (N115)? \nz.mem [339] : 
                            (N117)? \nz.mem [346] : 
                            (N119)? \nz.mem [353] : 
                            (N121)? \nz.mem [360] : 
                            (N123)? \nz.mem [367] : 
                            (N125)? \nz.mem [374] : 
                            (N127)? \nz.mem [381] : 
                            (N129)? \nz.mem [388] : 
                            (N131)? \nz.mem [395] : 
                            (N133)? \nz.mem [402] : 
                            (N135)? \nz.mem [409] : 
                            (N137)? \nz.mem [416] : 
                            (N139)? \nz.mem [423] : 
                            (N141)? \nz.mem [430] : 
                            (N143)? \nz.mem [437] : 
                            (N145)? \nz.mem [444] : 1'b0;
  assign \nz.data_out [2] = (N82)? \nz.mem [2] : 
                            (N84)? \nz.mem [9] : 
                            (N86)? \nz.mem [16] : 
                            (N88)? \nz.mem [23] : 
                            (N90)? \nz.mem [30] : 
                            (N92)? \nz.mem [37] : 
                            (N94)? \nz.mem [44] : 
                            (N96)? \nz.mem [51] : 
                            (N98)? \nz.mem [58] : 
                            (N100)? \nz.mem [65] : 
                            (N102)? \nz.mem [72] : 
                            (N104)? \nz.mem [79] : 
                            (N106)? \nz.mem [86] : 
                            (N108)? \nz.mem [93] : 
                            (N110)? \nz.mem [100] : 
                            (N112)? \nz.mem [107] : 
                            (N114)? \nz.mem [114] : 
                            (N116)? \nz.mem [121] : 
                            (N118)? \nz.mem [128] : 
                            (N120)? \nz.mem [135] : 
                            (N122)? \nz.mem [142] : 
                            (N124)? \nz.mem [149] : 
                            (N126)? \nz.mem [156] : 
                            (N128)? \nz.mem [163] : 
                            (N130)? \nz.mem [170] : 
                            (N132)? \nz.mem [177] : 
                            (N134)? \nz.mem [184] : 
                            (N136)? \nz.mem [191] : 
                            (N138)? \nz.mem [198] : 
                            (N140)? \nz.mem [205] : 
                            (N142)? \nz.mem [212] : 
                            (N144)? \nz.mem [219] : 
                            (N83)? \nz.mem [226] : 
                            (N85)? \nz.mem [233] : 
                            (N87)? \nz.mem [240] : 
                            (N89)? \nz.mem [247] : 
                            (N91)? \nz.mem [254] : 
                            (N93)? \nz.mem [261] : 
                            (N95)? \nz.mem [268] : 
                            (N97)? \nz.mem [275] : 
                            (N99)? \nz.mem [282] : 
                            (N101)? \nz.mem [289] : 
                            (N103)? \nz.mem [296] : 
                            (N105)? \nz.mem [303] : 
                            (N107)? \nz.mem [310] : 
                            (N109)? \nz.mem [317] : 
                            (N111)? \nz.mem [324] : 
                            (N113)? \nz.mem [331] : 
                            (N115)? \nz.mem [338] : 
                            (N117)? \nz.mem [345] : 
                            (N119)? \nz.mem [352] : 
                            (N121)? \nz.mem [359] : 
                            (N123)? \nz.mem [366] : 
                            (N125)? \nz.mem [373] : 
                            (N127)? \nz.mem [380] : 
                            (N129)? \nz.mem [387] : 
                            (N131)? \nz.mem [394] : 
                            (N133)? \nz.mem [401] : 
                            (N135)? \nz.mem [408] : 
                            (N137)? \nz.mem [415] : 
                            (N139)? \nz.mem [422] : 
                            (N141)? \nz.mem [429] : 
                            (N143)? \nz.mem [436] : 
                            (N145)? \nz.mem [443] : 1'b0;
  assign \nz.data_out [1] = (N82)? \nz.mem [1] : 
                            (N84)? \nz.mem [8] : 
                            (N86)? \nz.mem [15] : 
                            (N88)? \nz.mem [22] : 
                            (N90)? \nz.mem [29] : 
                            (N92)? \nz.mem [36] : 
                            (N94)? \nz.mem [43] : 
                            (N96)? \nz.mem [50] : 
                            (N98)? \nz.mem [57] : 
                            (N100)? \nz.mem [64] : 
                            (N102)? \nz.mem [71] : 
                            (N104)? \nz.mem [78] : 
                            (N106)? \nz.mem [85] : 
                            (N108)? \nz.mem [92] : 
                            (N110)? \nz.mem [99] : 
                            (N112)? \nz.mem [106] : 
                            (N114)? \nz.mem [113] : 
                            (N116)? \nz.mem [120] : 
                            (N118)? \nz.mem [127] : 
                            (N120)? \nz.mem [134] : 
                            (N122)? \nz.mem [141] : 
                            (N124)? \nz.mem [148] : 
                            (N126)? \nz.mem [155] : 
                            (N128)? \nz.mem [162] : 
                            (N130)? \nz.mem [169] : 
                            (N132)? \nz.mem [176] : 
                            (N134)? \nz.mem [183] : 
                            (N136)? \nz.mem [190] : 
                            (N138)? \nz.mem [197] : 
                            (N140)? \nz.mem [204] : 
                            (N142)? \nz.mem [211] : 
                            (N144)? \nz.mem [218] : 
                            (N83)? \nz.mem [225] : 
                            (N85)? \nz.mem [232] : 
                            (N87)? \nz.mem [239] : 
                            (N89)? \nz.mem [246] : 
                            (N91)? \nz.mem [253] : 
                            (N93)? \nz.mem [260] : 
                            (N95)? \nz.mem [267] : 
                            (N97)? \nz.mem [274] : 
                            (N99)? \nz.mem [281] : 
                            (N101)? \nz.mem [288] : 
                            (N103)? \nz.mem [295] : 
                            (N105)? \nz.mem [302] : 
                            (N107)? \nz.mem [309] : 
                            (N109)? \nz.mem [316] : 
                            (N111)? \nz.mem [323] : 
                            (N113)? \nz.mem [330] : 
                            (N115)? \nz.mem [337] : 
                            (N117)? \nz.mem [344] : 
                            (N119)? \nz.mem [351] : 
                            (N121)? \nz.mem [358] : 
                            (N123)? \nz.mem [365] : 
                            (N125)? \nz.mem [372] : 
                            (N127)? \nz.mem [379] : 
                            (N129)? \nz.mem [386] : 
                            (N131)? \nz.mem [393] : 
                            (N133)? \nz.mem [400] : 
                            (N135)? \nz.mem [407] : 
                            (N137)? \nz.mem [414] : 
                            (N139)? \nz.mem [421] : 
                            (N141)? \nz.mem [428] : 
                            (N143)? \nz.mem [435] : 
                            (N145)? \nz.mem [442] : 1'b0;
  assign \nz.data_out [0] = (N82)? \nz.mem [0] : 
                            (N84)? \nz.mem [7] : 
                            (N86)? \nz.mem [14] : 
                            (N88)? \nz.mem [21] : 
                            (N90)? \nz.mem [28] : 
                            (N92)? \nz.mem [35] : 
                            (N94)? \nz.mem [42] : 
                            (N96)? \nz.mem [49] : 
                            (N98)? \nz.mem [56] : 
                            (N100)? \nz.mem [63] : 
                            (N102)? \nz.mem [70] : 
                            (N104)? \nz.mem [77] : 
                            (N106)? \nz.mem [84] : 
                            (N108)? \nz.mem [91] : 
                            (N110)? \nz.mem [98] : 
                            (N112)? \nz.mem [105] : 
                            (N114)? \nz.mem [112] : 
                            (N116)? \nz.mem [119] : 
                            (N118)? \nz.mem [126] : 
                            (N120)? \nz.mem [133] : 
                            (N122)? \nz.mem [140] : 
                            (N124)? \nz.mem [147] : 
                            (N126)? \nz.mem [154] : 
                            (N128)? \nz.mem [161] : 
                            (N130)? \nz.mem [168] : 
                            (N132)? \nz.mem [175] : 
                            (N134)? \nz.mem [182] : 
                            (N136)? \nz.mem [189] : 
                            (N138)? \nz.mem [196] : 
                            (N140)? \nz.mem [203] : 
                            (N142)? \nz.mem [210] : 
                            (N144)? \nz.mem [217] : 
                            (N83)? \nz.mem [224] : 
                            (N85)? \nz.mem [231] : 
                            (N87)? \nz.mem [238] : 
                            (N89)? \nz.mem [245] : 
                            (N91)? \nz.mem [252] : 
                            (N93)? \nz.mem [259] : 
                            (N95)? \nz.mem [266] : 
                            (N97)? \nz.mem [273] : 
                            (N99)? \nz.mem [280] : 
                            (N101)? \nz.mem [287] : 
                            (N103)? \nz.mem [294] : 
                            (N105)? \nz.mem [301] : 
                            (N107)? \nz.mem [308] : 
                            (N109)? \nz.mem [315] : 
                            (N111)? \nz.mem [322] : 
                            (N113)? \nz.mem [329] : 
                            (N115)? \nz.mem [336] : 
                            (N117)? \nz.mem [343] : 
                            (N119)? \nz.mem [350] : 
                            (N121)? \nz.mem [357] : 
                            (N123)? \nz.mem [364] : 
                            (N125)? \nz.mem [371] : 
                            (N127)? \nz.mem [378] : 
                            (N129)? \nz.mem [385] : 
                            (N131)? \nz.mem [392] : 
                            (N133)? \nz.mem [399] : 
                            (N135)? \nz.mem [406] : 
                            (N137)? \nz.mem [413] : 
                            (N139)? \nz.mem [420] : 
                            (N141)? \nz.mem [427] : 
                            (N143)? \nz.mem [434] : 
                            (N145)? \nz.mem [441] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p7
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N1115 = ~addr_i[5];
  assign N1116 = addr_i[3] & addr_i[4];
  assign N1117 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N1118 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N1119 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N1120 = addr_i[5] & N1116;
  assign N1121 = addr_i[5] & N1117;
  assign N1122 = addr_i[5] & N1118;
  assign N1123 = addr_i[5] & N1119;
  assign N1124 = N1115 & N1116;
  assign N1125 = N1115 & N1117;
  assign N1126 = N1115 & N1118;
  assign N1127 = N1115 & N1119;
  assign N1128 = ~addr_i[2];
  assign N1129 = addr_i[0] & addr_i[1];
  assign N1130 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N1131 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N1132 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N1133 = addr_i[2] & N1129;
  assign N1134 = addr_i[2] & N1130;
  assign N1135 = addr_i[2] & N1131;
  assign N1136 = addr_i[2] & N1132;
  assign N1137 = N1128 & N1129;
  assign N1138 = N1128 & N1130;
  assign N1139 = N1128 & N1131;
  assign N1140 = N1128 & N1132;
  assign N602 = N1120 & N1133;
  assign N601 = N1120 & N1134;
  assign N600 = N1120 & N1135;
  assign N599 = N1120 & N1136;
  assign N598 = N1120 & N1137;
  assign N597 = N1120 & N1138;
  assign N596 = N1120 & N1139;
  assign N595 = N1120 & N1140;
  assign N594 = N1121 & N1133;
  assign N593 = N1121 & N1134;
  assign N592 = N1121 & N1135;
  assign N591 = N1121 & N1136;
  assign N590 = N1121 & N1137;
  assign N589 = N1121 & N1138;
  assign N588 = N1121 & N1139;
  assign N587 = N1121 & N1140;
  assign N586 = N1122 & N1133;
  assign N585 = N1122 & N1134;
  assign N584 = N1122 & N1135;
  assign N583 = N1122 & N1136;
  assign N582 = N1122 & N1137;
  assign N581 = N1122 & N1138;
  assign N580 = N1122 & N1139;
  assign N579 = N1122 & N1140;
  assign N578 = N1123 & N1133;
  assign N577 = N1123 & N1134;
  assign N576 = N1123 & N1135;
  assign N575 = N1123 & N1136;
  assign N574 = N1123 & N1137;
  assign N573 = N1123 & N1138;
  assign N572 = N1123 & N1139;
  assign N571 = N1123 & N1140;
  assign N570 = N1124 & N1133;
  assign N569 = N1124 & N1134;
  assign N568 = N1124 & N1135;
  assign N567 = N1124 & N1136;
  assign N566 = N1124 & N1137;
  assign N565 = N1124 & N1138;
  assign N564 = N1124 & N1139;
  assign N563 = N1124 & N1140;
  assign N562 = N1125 & N1133;
  assign N561 = N1125 & N1134;
  assign N560 = N1125 & N1135;
  assign N559 = N1125 & N1136;
  assign N558 = N1125 & N1137;
  assign N557 = N1125 & N1138;
  assign N556 = N1125 & N1139;
  assign N555 = N1125 & N1140;
  assign N554 = N1126 & N1133;
  assign N553 = N1126 & N1134;
  assign N552 = N1126 & N1135;
  assign N551 = N1126 & N1136;
  assign N550 = N1126 & N1137;
  assign N549 = N1126 & N1138;
  assign N548 = N1126 & N1139;
  assign N547 = N1126 & N1140;
  assign N546 = N1127 & N1133;
  assign N545 = N1127 & N1134;
  assign N544 = N1127 & N1135;
  assign N543 = N1127 & N1136;
  assign N542 = N1127 & N1137;
  assign N541 = N1127 & N1138;
  assign N540 = N1127 & N1139;
  assign N539 = N1127 & N1140;
  assign { N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149 } = (N8)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N148)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214 } = (N9)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N213)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 } = (N10)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N278)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344 } = (N11)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N343)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409 } = (N12)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N408)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474 } = (N13)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N473)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603 } = (N14)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N538)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667 } = (N15)? { N666, N537, N472, N407, N342, N277, N212, N665, N536, N471, N406, N341, N276, N211, N664, N535, N470, N405, N340, N275, N210, N663, N534, N469, N404, N339, N274, N209, N662, N533, N468, N403, N338, N273, N208, N661, N532, N467, N402, N337, N272, N207, N660, N531, N466, N401, N336, N271, N206, N659, N530, N465, N400, N335, N270, N205, N658, N529, N464, N399, N334, N269, N204, N657, N528, N463, N398, N333, N268, N203, N656, N527, N462, N397, N332, N267, N202, N655, N526, N461, N396, N331, N266, N201, N654, N525, N460, N395, N330, N265, N200, N653, N524, N459, N394, N329, N264, N199, N652, N523, N458, N393, N328, N263, N198, N651, N522, N457, N392, N327, N262, N197, N650, N521, N456, N391, N326, N261, N196, N649, N520, N455, N390, N325, N260, N195, N648, N519, N454, N389, N324, N259, N194, N647, N518, N453, N388, N323, N258, N193, N646, N517, N452, N387, N322, N257, N192, N645, N516, N451, N386, N321, N256, N191, N644, N515, N450, N385, N320, N255, N190, N643, N514, N449, N384, N319, N254, N189, N642, N513, N448, N383, N318, N253, N188, N641, N512, N447, N382, N317, N252, N187, N640, N511, N446, N381, N316, N251, N186, N639, N510, N445, N380, N315, N250, N185, N638, N509, N444, N379, N314, N249, N184, N637, N508, N443, N378, N313, N248, N183, N636, N507, N442, N377, N312, N247, N182, N635, N506, N441, N376, N311, N246, N181, N634, N505, N440, N375, N310, N245, N180, N633, N504, N439, N374, N309, N244, N179, N632, N503, N438, N373, N308, N243, N178, N631, N502, N437, N372, N307, N242, N177, N630, N501, N436, N371, N306, N241, N176, N629, N500, N435, N370, N305, N240, N175, N628, N499, N434, N369, N304, N239, N174, N627, N498, N433, N368, N303, N238, N173, N626, N497, N432, N367, N302, N237, N172, N625, N496, N431, N366, N301, N236, N171, N624, N495, N430, N365, N300, N235, N170, N623, N494, N429, N364, N299, N234, N169, N622, N493, N428, N363, N298, N233, N168, N621, N492, N427, N362, N297, N232, N167, N620, N491, N426, N361, N296, N231, N166, N619, N490, N425, N360, N295, N230, N165, N618, N489, N424, N359, N294, N229, N164, N617, N488, N423, N358, N293, N228, N163, N616, N487, N422, N357, N292, N227, N162, N615, N486, N421, N356, N291, N226, N161, N614, N485, N420, N355, N290, N225, N160, N613, N484, N419, N354, N289, N224, N159, N612, N483, N418, N353, N288, N223, N158, N611, N482, N417, N352, N287, N222, N157, N610, N481, N416, N351, N286, N221, N156, N609, N480, N415, N350, N285, N220, N155, N608, N479, N414, N349, N284, N219, N154, N607, N478, N413, N348, N283, N218, N153, N606, N477, N412, N347, N282, N217, N152, N605, N476, N411, N346, N281, N216, N151, N604, N475, N410, N345, N280, N215, N150, N603, N474, N409, N344, N279, N214, N149 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 (N147)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N146;
  assign \nz.read_en  = v_i & N1141;
  assign N1141 = ~w_i;
  assign N16 = ~\nz.addr_r [0];
  assign N17 = ~\nz.addr_r [1];
  assign N18 = N16 & N17;
  assign N19 = N16 & \nz.addr_r [1];
  assign N20 = \nz.addr_r [0] & N17;
  assign N21 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N22 = ~\nz.addr_r [2];
  assign N23 = N18 & N22;
  assign N24 = N18 & \nz.addr_r [2];
  assign N25 = N20 & N22;
  assign N26 = N20 & \nz.addr_r [2];
  assign N27 = N19 & N22;
  assign N28 = N19 & \nz.addr_r [2];
  assign N29 = N21 & N22;
  assign N30 = N21 & \nz.addr_r [2];
  assign N31 = ~\nz.addr_r [3];
  assign N32 = N23 & N31;
  assign N33 = N23 & \nz.addr_r [3];
  assign N34 = N25 & N31;
  assign N35 = N25 & \nz.addr_r [3];
  assign N36 = N27 & N31;
  assign N37 = N27 & \nz.addr_r [3];
  assign N38 = N29 & N31;
  assign N39 = N29 & \nz.addr_r [3];
  assign N40 = N24 & N31;
  assign N41 = N24 & \nz.addr_r [3];
  assign N42 = N26 & N31;
  assign N43 = N26 & \nz.addr_r [3];
  assign N44 = N28 & N31;
  assign N45 = N28 & \nz.addr_r [3];
  assign N46 = N30 & N31;
  assign N47 = N30 & \nz.addr_r [3];
  assign N48 = ~\nz.addr_r [4];
  assign N49 = N32 & N48;
  assign N50 = N32 & \nz.addr_r [4];
  assign N51 = N34 & N48;
  assign N52 = N34 & \nz.addr_r [4];
  assign N53 = N36 & N48;
  assign N54 = N36 & \nz.addr_r [4];
  assign N55 = N38 & N48;
  assign N56 = N38 & \nz.addr_r [4];
  assign N57 = N40 & N48;
  assign N58 = N40 & \nz.addr_r [4];
  assign N59 = N42 & N48;
  assign N60 = N42 & \nz.addr_r [4];
  assign N61 = N44 & N48;
  assign N62 = N44 & \nz.addr_r [4];
  assign N63 = N46 & N48;
  assign N64 = N46 & \nz.addr_r [4];
  assign N65 = N33 & N48;
  assign N66 = N33 & \nz.addr_r [4];
  assign N67 = N35 & N48;
  assign N68 = N35 & \nz.addr_r [4];
  assign N69 = N37 & N48;
  assign N70 = N37 & \nz.addr_r [4];
  assign N71 = N39 & N48;
  assign N72 = N39 & \nz.addr_r [4];
  assign N73 = N41 & N48;
  assign N74 = N41 & \nz.addr_r [4];
  assign N75 = N43 & N48;
  assign N76 = N43 & \nz.addr_r [4];
  assign N77 = N45 & N48;
  assign N78 = N45 & \nz.addr_r [4];
  assign N79 = N47 & N48;
  assign N80 = N47 & \nz.addr_r [4];
  assign N81 = ~\nz.addr_r [5];
  assign N82 = N49 & N81;
  assign N83 = N49 & \nz.addr_r [5];
  assign N84 = N51 & N81;
  assign N85 = N51 & \nz.addr_r [5];
  assign N86 = N53 & N81;
  assign N87 = N53 & \nz.addr_r [5];
  assign N88 = N55 & N81;
  assign N89 = N55 & \nz.addr_r [5];
  assign N90 = N57 & N81;
  assign N91 = N57 & \nz.addr_r [5];
  assign N92 = N59 & N81;
  assign N93 = N59 & \nz.addr_r [5];
  assign N94 = N61 & N81;
  assign N95 = N61 & \nz.addr_r [5];
  assign N96 = N63 & N81;
  assign N97 = N63 & \nz.addr_r [5];
  assign N98 = N65 & N81;
  assign N99 = N65 & \nz.addr_r [5];
  assign N100 = N67 & N81;
  assign N101 = N67 & \nz.addr_r [5];
  assign N102 = N69 & N81;
  assign N103 = N69 & \nz.addr_r [5];
  assign N104 = N71 & N81;
  assign N105 = N71 & \nz.addr_r [5];
  assign N106 = N73 & N81;
  assign N107 = N73 & \nz.addr_r [5];
  assign N108 = N75 & N81;
  assign N109 = N75 & \nz.addr_r [5];
  assign N110 = N77 & N81;
  assign N111 = N77 & \nz.addr_r [5];
  assign N112 = N79 & N81;
  assign N113 = N79 & \nz.addr_r [5];
  assign N114 = N50 & N81;
  assign N115 = N50 & \nz.addr_r [5];
  assign N116 = N52 & N81;
  assign N117 = N52 & \nz.addr_r [5];
  assign N118 = N54 & N81;
  assign N119 = N54 & \nz.addr_r [5];
  assign N120 = N56 & N81;
  assign N121 = N56 & \nz.addr_r [5];
  assign N122 = N58 & N81;
  assign N123 = N58 & \nz.addr_r [5];
  assign N124 = N60 & N81;
  assign N125 = N60 & \nz.addr_r [5];
  assign N126 = N62 & N81;
  assign N127 = N62 & \nz.addr_r [5];
  assign N128 = N64 & N81;
  assign N129 = N64 & \nz.addr_r [5];
  assign N130 = N66 & N81;
  assign N131 = N66 & \nz.addr_r [5];
  assign N132 = N68 & N81;
  assign N133 = N68 & \nz.addr_r [5];
  assign N134 = N70 & N81;
  assign N135 = N70 & \nz.addr_r [5];
  assign N136 = N72 & N81;
  assign N137 = N72 & \nz.addr_r [5];
  assign N138 = N74 & N81;
  assign N139 = N74 & \nz.addr_r [5];
  assign N140 = N76 & N81;
  assign N141 = N76 & \nz.addr_r [5];
  assign N142 = N78 & N81;
  assign N143 = N78 & \nz.addr_r [5];
  assign N144 = N80 & N81;
  assign N145 = N80 & \nz.addr_r [5];
  assign N146 = v_i & w_i;
  assign N147 = ~N146;
  assign N148 = ~w_mask_i[0];
  assign N213 = ~w_mask_i[1];
  assign N278 = ~w_mask_i[2];
  assign N343 = ~w_mask_i[3];
  assign N408 = ~w_mask_i[4];
  assign N473 = ~w_mask_i[5];
  assign N538 = ~w_mask_i[6];

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N1114) begin
      \nz.mem_447_sv2v_reg  <= data_i[6];
    end 
    if(N1113) begin
      \nz.mem_446_sv2v_reg  <= data_i[5];
    end 
    if(N1112) begin
      \nz.mem_445_sv2v_reg  <= data_i[4];
    end 
    if(N1111) begin
      \nz.mem_444_sv2v_reg  <= data_i[3];
    end 
    if(N1110) begin
      \nz.mem_443_sv2v_reg  <= data_i[2];
    end 
    if(N1109) begin
      \nz.mem_442_sv2v_reg  <= data_i[1];
    end 
    if(N1108) begin
      \nz.mem_441_sv2v_reg  <= data_i[0];
    end 
    if(N1107) begin
      \nz.mem_440_sv2v_reg  <= data_i[6];
    end 
    if(N1106) begin
      \nz.mem_439_sv2v_reg  <= data_i[5];
    end 
    if(N1105) begin
      \nz.mem_438_sv2v_reg  <= data_i[4];
    end 
    if(N1104) begin
      \nz.mem_437_sv2v_reg  <= data_i[3];
    end 
    if(N1103) begin
      \nz.mem_436_sv2v_reg  <= data_i[2];
    end 
    if(N1102) begin
      \nz.mem_435_sv2v_reg  <= data_i[1];
    end 
    if(N1101) begin
      \nz.mem_434_sv2v_reg  <= data_i[0];
    end 
    if(N1100) begin
      \nz.mem_433_sv2v_reg  <= data_i[6];
    end 
    if(N1099) begin
      \nz.mem_432_sv2v_reg  <= data_i[5];
    end 
    if(N1098) begin
      \nz.mem_431_sv2v_reg  <= data_i[4];
    end 
    if(N1097) begin
      \nz.mem_430_sv2v_reg  <= data_i[3];
    end 
    if(N1096) begin
      \nz.mem_429_sv2v_reg  <= data_i[2];
    end 
    if(N1095) begin
      \nz.mem_428_sv2v_reg  <= data_i[1];
    end 
    if(N1094) begin
      \nz.mem_427_sv2v_reg  <= data_i[0];
    end 
    if(N1093) begin
      \nz.mem_426_sv2v_reg  <= data_i[6];
    end 
    if(N1092) begin
      \nz.mem_425_sv2v_reg  <= data_i[5];
    end 
    if(N1091) begin
      \nz.mem_424_sv2v_reg  <= data_i[4];
    end 
    if(N1090) begin
      \nz.mem_423_sv2v_reg  <= data_i[3];
    end 
    if(N1089) begin
      \nz.mem_422_sv2v_reg  <= data_i[2];
    end 
    if(N1088) begin
      \nz.mem_421_sv2v_reg  <= data_i[1];
    end 
    if(N1087) begin
      \nz.mem_420_sv2v_reg  <= data_i[0];
    end 
    if(N1086) begin
      \nz.mem_419_sv2v_reg  <= data_i[6];
    end 
    if(N1085) begin
      \nz.mem_418_sv2v_reg  <= data_i[5];
    end 
    if(N1084) begin
      \nz.mem_417_sv2v_reg  <= data_i[4];
    end 
    if(N1083) begin
      \nz.mem_416_sv2v_reg  <= data_i[3];
    end 
    if(N1082) begin
      \nz.mem_415_sv2v_reg  <= data_i[2];
    end 
    if(N1081) begin
      \nz.mem_414_sv2v_reg  <= data_i[1];
    end 
    if(N1080) begin
      \nz.mem_413_sv2v_reg  <= data_i[0];
    end 
    if(N1079) begin
      \nz.mem_412_sv2v_reg  <= data_i[6];
    end 
    if(N1078) begin
      \nz.mem_411_sv2v_reg  <= data_i[5];
    end 
    if(N1077) begin
      \nz.mem_410_sv2v_reg  <= data_i[4];
    end 
    if(N1076) begin
      \nz.mem_409_sv2v_reg  <= data_i[3];
    end 
    if(N1075) begin
      \nz.mem_408_sv2v_reg  <= data_i[2];
    end 
    if(N1074) begin
      \nz.mem_407_sv2v_reg  <= data_i[1];
    end 
    if(N1073) begin
      \nz.mem_406_sv2v_reg  <= data_i[0];
    end 
    if(N1072) begin
      \nz.mem_405_sv2v_reg  <= data_i[6];
    end 
    if(N1071) begin
      \nz.mem_404_sv2v_reg  <= data_i[5];
    end 
    if(N1070) begin
      \nz.mem_403_sv2v_reg  <= data_i[4];
    end 
    if(N1069) begin
      \nz.mem_402_sv2v_reg  <= data_i[3];
    end 
    if(N1068) begin
      \nz.mem_401_sv2v_reg  <= data_i[2];
    end 
    if(N1067) begin
      \nz.mem_400_sv2v_reg  <= data_i[1];
    end 
    if(N1066) begin
      \nz.mem_399_sv2v_reg  <= data_i[0];
    end 
    if(N1065) begin
      \nz.mem_398_sv2v_reg  <= data_i[6];
    end 
    if(N1064) begin
      \nz.mem_397_sv2v_reg  <= data_i[5];
    end 
    if(N1063) begin
      \nz.mem_396_sv2v_reg  <= data_i[4];
    end 
    if(N1062) begin
      \nz.mem_395_sv2v_reg  <= data_i[3];
    end 
    if(N1061) begin
      \nz.mem_394_sv2v_reg  <= data_i[2];
    end 
    if(N1060) begin
      \nz.mem_393_sv2v_reg  <= data_i[1];
    end 
    if(N1059) begin
      \nz.mem_392_sv2v_reg  <= data_i[0];
    end 
    if(N1058) begin
      \nz.mem_391_sv2v_reg  <= data_i[6];
    end 
    if(N1057) begin
      \nz.mem_390_sv2v_reg  <= data_i[5];
    end 
    if(N1056) begin
      \nz.mem_389_sv2v_reg  <= data_i[4];
    end 
    if(N1055) begin
      \nz.mem_388_sv2v_reg  <= data_i[3];
    end 
    if(N1054) begin
      \nz.mem_387_sv2v_reg  <= data_i[2];
    end 
    if(N1053) begin
      \nz.mem_386_sv2v_reg  <= data_i[1];
    end 
    if(N1052) begin
      \nz.mem_385_sv2v_reg  <= data_i[0];
    end 
    if(N1051) begin
      \nz.mem_384_sv2v_reg  <= data_i[6];
    end 
    if(N1050) begin
      \nz.mem_383_sv2v_reg  <= data_i[5];
    end 
    if(N1049) begin
      \nz.mem_382_sv2v_reg  <= data_i[4];
    end 
    if(N1048) begin
      \nz.mem_381_sv2v_reg  <= data_i[3];
    end 
    if(N1047) begin
      \nz.mem_380_sv2v_reg  <= data_i[2];
    end 
    if(N1046) begin
      \nz.mem_379_sv2v_reg  <= data_i[1];
    end 
    if(N1045) begin
      \nz.mem_378_sv2v_reg  <= data_i[0];
    end 
    if(N1044) begin
      \nz.mem_377_sv2v_reg  <= data_i[6];
    end 
    if(N1043) begin
      \nz.mem_376_sv2v_reg  <= data_i[5];
    end 
    if(N1042) begin
      \nz.mem_375_sv2v_reg  <= data_i[4];
    end 
    if(N1041) begin
      \nz.mem_374_sv2v_reg  <= data_i[3];
    end 
    if(N1040) begin
      \nz.mem_373_sv2v_reg  <= data_i[2];
    end 
    if(N1039) begin
      \nz.mem_372_sv2v_reg  <= data_i[1];
    end 
    if(N1038) begin
      \nz.mem_371_sv2v_reg  <= data_i[0];
    end 
    if(N1037) begin
      \nz.mem_370_sv2v_reg  <= data_i[6];
    end 
    if(N1036) begin
      \nz.mem_369_sv2v_reg  <= data_i[5];
    end 
    if(N1035) begin
      \nz.mem_368_sv2v_reg  <= data_i[4];
    end 
    if(N1034) begin
      \nz.mem_367_sv2v_reg  <= data_i[3];
    end 
    if(N1033) begin
      \nz.mem_366_sv2v_reg  <= data_i[2];
    end 
    if(N1032) begin
      \nz.mem_365_sv2v_reg  <= data_i[1];
    end 
    if(N1031) begin
      \nz.mem_364_sv2v_reg  <= data_i[0];
    end 
    if(N1030) begin
      \nz.mem_363_sv2v_reg  <= data_i[6];
    end 
    if(N1029) begin
      \nz.mem_362_sv2v_reg  <= data_i[5];
    end 
    if(N1028) begin
      \nz.mem_361_sv2v_reg  <= data_i[4];
    end 
    if(N1027) begin
      \nz.mem_360_sv2v_reg  <= data_i[3];
    end 
    if(N1026) begin
      \nz.mem_359_sv2v_reg  <= data_i[2];
    end 
    if(N1025) begin
      \nz.mem_358_sv2v_reg  <= data_i[1];
    end 
    if(N1024) begin
      \nz.mem_357_sv2v_reg  <= data_i[0];
    end 
    if(N1023) begin
      \nz.mem_356_sv2v_reg  <= data_i[6];
    end 
    if(N1022) begin
      \nz.mem_355_sv2v_reg  <= data_i[5];
    end 
    if(N1021) begin
      \nz.mem_354_sv2v_reg  <= data_i[4];
    end 
    if(N1020) begin
      \nz.mem_353_sv2v_reg  <= data_i[3];
    end 
    if(N1019) begin
      \nz.mem_352_sv2v_reg  <= data_i[2];
    end 
    if(N1018) begin
      \nz.mem_351_sv2v_reg  <= data_i[1];
    end 
    if(N1017) begin
      \nz.mem_350_sv2v_reg  <= data_i[0];
    end 
    if(N1016) begin
      \nz.mem_349_sv2v_reg  <= data_i[6];
    end 
    if(N1015) begin
      \nz.mem_348_sv2v_reg  <= data_i[5];
    end 
    if(N1014) begin
      \nz.mem_347_sv2v_reg  <= data_i[4];
    end 
    if(N1013) begin
      \nz.mem_346_sv2v_reg  <= data_i[3];
    end 
    if(N1012) begin
      \nz.mem_345_sv2v_reg  <= data_i[2];
    end 
    if(N1011) begin
      \nz.mem_344_sv2v_reg  <= data_i[1];
    end 
    if(N1010) begin
      \nz.mem_343_sv2v_reg  <= data_i[0];
    end 
    if(N1009) begin
      \nz.mem_342_sv2v_reg  <= data_i[6];
    end 
    if(N1008) begin
      \nz.mem_341_sv2v_reg  <= data_i[5];
    end 
    if(N1007) begin
      \nz.mem_340_sv2v_reg  <= data_i[4];
    end 
    if(N1006) begin
      \nz.mem_339_sv2v_reg  <= data_i[3];
    end 
    if(N1005) begin
      \nz.mem_338_sv2v_reg  <= data_i[2];
    end 
    if(N1004) begin
      \nz.mem_337_sv2v_reg  <= data_i[1];
    end 
    if(N1003) begin
      \nz.mem_336_sv2v_reg  <= data_i[0];
    end 
    if(N1002) begin
      \nz.mem_335_sv2v_reg  <= data_i[6];
    end 
    if(N1001) begin
      \nz.mem_334_sv2v_reg  <= data_i[5];
    end 
    if(N1000) begin
      \nz.mem_333_sv2v_reg  <= data_i[4];
    end 
    if(N999) begin
      \nz.mem_332_sv2v_reg  <= data_i[3];
    end 
    if(N998) begin
      \nz.mem_331_sv2v_reg  <= data_i[2];
    end 
    if(N997) begin
      \nz.mem_330_sv2v_reg  <= data_i[1];
    end 
    if(N996) begin
      \nz.mem_329_sv2v_reg  <= data_i[0];
    end 
    if(N995) begin
      \nz.mem_328_sv2v_reg  <= data_i[6];
    end 
    if(N994) begin
      \nz.mem_327_sv2v_reg  <= data_i[5];
    end 
    if(N993) begin
      \nz.mem_326_sv2v_reg  <= data_i[4];
    end 
    if(N992) begin
      \nz.mem_325_sv2v_reg  <= data_i[3];
    end 
    if(N991) begin
      \nz.mem_324_sv2v_reg  <= data_i[2];
    end 
    if(N990) begin
      \nz.mem_323_sv2v_reg  <= data_i[1];
    end 
    if(N989) begin
      \nz.mem_322_sv2v_reg  <= data_i[0];
    end 
    if(N988) begin
      \nz.mem_321_sv2v_reg  <= data_i[6];
    end 
    if(N987) begin
      \nz.mem_320_sv2v_reg  <= data_i[5];
    end 
    if(N986) begin
      \nz.mem_319_sv2v_reg  <= data_i[4];
    end 
    if(N985) begin
      \nz.mem_318_sv2v_reg  <= data_i[3];
    end 
    if(N984) begin
      \nz.mem_317_sv2v_reg  <= data_i[2];
    end 
    if(N983) begin
      \nz.mem_316_sv2v_reg  <= data_i[1];
    end 
    if(N982) begin
      \nz.mem_315_sv2v_reg  <= data_i[0];
    end 
    if(N981) begin
      \nz.mem_314_sv2v_reg  <= data_i[6];
    end 
    if(N980) begin
      \nz.mem_313_sv2v_reg  <= data_i[5];
    end 
    if(N979) begin
      \nz.mem_312_sv2v_reg  <= data_i[4];
    end 
    if(N978) begin
      \nz.mem_311_sv2v_reg  <= data_i[3];
    end 
    if(N977) begin
      \nz.mem_310_sv2v_reg  <= data_i[2];
    end 
    if(N976) begin
      \nz.mem_309_sv2v_reg  <= data_i[1];
    end 
    if(N975) begin
      \nz.mem_308_sv2v_reg  <= data_i[0];
    end 
    if(N974) begin
      \nz.mem_307_sv2v_reg  <= data_i[6];
    end 
    if(N973) begin
      \nz.mem_306_sv2v_reg  <= data_i[5];
    end 
    if(N972) begin
      \nz.mem_305_sv2v_reg  <= data_i[4];
    end 
    if(N971) begin
      \nz.mem_304_sv2v_reg  <= data_i[3];
    end 
    if(N970) begin
      \nz.mem_303_sv2v_reg  <= data_i[2];
    end 
    if(N969) begin
      \nz.mem_302_sv2v_reg  <= data_i[1];
    end 
    if(N968) begin
      \nz.mem_301_sv2v_reg  <= data_i[0];
    end 
    if(N967) begin
      \nz.mem_300_sv2v_reg  <= data_i[6];
    end 
    if(N966) begin
      \nz.mem_299_sv2v_reg  <= data_i[5];
    end 
    if(N965) begin
      \nz.mem_298_sv2v_reg  <= data_i[4];
    end 
    if(N964) begin
      \nz.mem_297_sv2v_reg  <= data_i[3];
    end 
    if(N963) begin
      \nz.mem_296_sv2v_reg  <= data_i[2];
    end 
    if(N962) begin
      \nz.mem_295_sv2v_reg  <= data_i[1];
    end 
    if(N961) begin
      \nz.mem_294_sv2v_reg  <= data_i[0];
    end 
    if(N960) begin
      \nz.mem_293_sv2v_reg  <= data_i[6];
    end 
    if(N959) begin
      \nz.mem_292_sv2v_reg  <= data_i[5];
    end 
    if(N958) begin
      \nz.mem_291_sv2v_reg  <= data_i[4];
    end 
    if(N957) begin
      \nz.mem_290_sv2v_reg  <= data_i[3];
    end 
    if(N956) begin
      \nz.mem_289_sv2v_reg  <= data_i[2];
    end 
    if(N955) begin
      \nz.mem_288_sv2v_reg  <= data_i[1];
    end 
    if(N954) begin
      \nz.mem_287_sv2v_reg  <= data_i[0];
    end 
    if(N953) begin
      \nz.mem_286_sv2v_reg  <= data_i[6];
    end 
    if(N952) begin
      \nz.mem_285_sv2v_reg  <= data_i[5];
    end 
    if(N951) begin
      \nz.mem_284_sv2v_reg  <= data_i[4];
    end 
    if(N950) begin
      \nz.mem_283_sv2v_reg  <= data_i[3];
    end 
    if(N949) begin
      \nz.mem_282_sv2v_reg  <= data_i[2];
    end 
    if(N948) begin
      \nz.mem_281_sv2v_reg  <= data_i[1];
    end 
    if(N947) begin
      \nz.mem_280_sv2v_reg  <= data_i[0];
    end 
    if(N946) begin
      \nz.mem_279_sv2v_reg  <= data_i[6];
    end 
    if(N945) begin
      \nz.mem_278_sv2v_reg  <= data_i[5];
    end 
    if(N944) begin
      \nz.mem_277_sv2v_reg  <= data_i[4];
    end 
    if(N943) begin
      \nz.mem_276_sv2v_reg  <= data_i[3];
    end 
    if(N942) begin
      \nz.mem_275_sv2v_reg  <= data_i[2];
    end 
    if(N941) begin
      \nz.mem_274_sv2v_reg  <= data_i[1];
    end 
    if(N940) begin
      \nz.mem_273_sv2v_reg  <= data_i[0];
    end 
    if(N939) begin
      \nz.mem_272_sv2v_reg  <= data_i[6];
    end 
    if(N938) begin
      \nz.mem_271_sv2v_reg  <= data_i[5];
    end 
    if(N937) begin
      \nz.mem_270_sv2v_reg  <= data_i[4];
    end 
    if(N936) begin
      \nz.mem_269_sv2v_reg  <= data_i[3];
    end 
    if(N935) begin
      \nz.mem_268_sv2v_reg  <= data_i[2];
    end 
    if(N934) begin
      \nz.mem_267_sv2v_reg  <= data_i[1];
    end 
    if(N933) begin
      \nz.mem_266_sv2v_reg  <= data_i[0];
    end 
    if(N932) begin
      \nz.mem_265_sv2v_reg  <= data_i[6];
    end 
    if(N931) begin
      \nz.mem_264_sv2v_reg  <= data_i[5];
    end 
    if(N930) begin
      \nz.mem_263_sv2v_reg  <= data_i[4];
    end 
    if(N929) begin
      \nz.mem_262_sv2v_reg  <= data_i[3];
    end 
    if(N928) begin
      \nz.mem_261_sv2v_reg  <= data_i[2];
    end 
    if(N927) begin
      \nz.mem_260_sv2v_reg  <= data_i[1];
    end 
    if(N926) begin
      \nz.mem_259_sv2v_reg  <= data_i[0];
    end 
    if(N925) begin
      \nz.mem_258_sv2v_reg  <= data_i[6];
    end 
    if(N924) begin
      \nz.mem_257_sv2v_reg  <= data_i[5];
    end 
    if(N923) begin
      \nz.mem_256_sv2v_reg  <= data_i[4];
    end 
    if(N922) begin
      \nz.mem_255_sv2v_reg  <= data_i[3];
    end 
    if(N921) begin
      \nz.mem_254_sv2v_reg  <= data_i[2];
    end 
    if(N920) begin
      \nz.mem_253_sv2v_reg  <= data_i[1];
    end 
    if(N919) begin
      \nz.mem_252_sv2v_reg  <= data_i[0];
    end 
    if(N918) begin
      \nz.mem_251_sv2v_reg  <= data_i[6];
    end 
    if(N917) begin
      \nz.mem_250_sv2v_reg  <= data_i[5];
    end 
    if(N916) begin
      \nz.mem_249_sv2v_reg  <= data_i[4];
    end 
    if(N915) begin
      \nz.mem_248_sv2v_reg  <= data_i[3];
    end 
    if(N914) begin
      \nz.mem_247_sv2v_reg  <= data_i[2];
    end 
    if(N913) begin
      \nz.mem_246_sv2v_reg  <= data_i[1];
    end 
    if(N912) begin
      \nz.mem_245_sv2v_reg  <= data_i[0];
    end 
    if(N911) begin
      \nz.mem_244_sv2v_reg  <= data_i[6];
    end 
    if(N910) begin
      \nz.mem_243_sv2v_reg  <= data_i[5];
    end 
    if(N909) begin
      \nz.mem_242_sv2v_reg  <= data_i[4];
    end 
    if(N908) begin
      \nz.mem_241_sv2v_reg  <= data_i[3];
    end 
    if(N907) begin
      \nz.mem_240_sv2v_reg  <= data_i[2];
    end 
    if(N906) begin
      \nz.mem_239_sv2v_reg  <= data_i[1];
    end 
    if(N905) begin
      \nz.mem_238_sv2v_reg  <= data_i[0];
    end 
    if(N904) begin
      \nz.mem_237_sv2v_reg  <= data_i[6];
    end 
    if(N903) begin
      \nz.mem_236_sv2v_reg  <= data_i[5];
    end 
    if(N902) begin
      \nz.mem_235_sv2v_reg  <= data_i[4];
    end 
    if(N901) begin
      \nz.mem_234_sv2v_reg  <= data_i[3];
    end 
    if(N900) begin
      \nz.mem_233_sv2v_reg  <= data_i[2];
    end 
    if(N899) begin
      \nz.mem_232_sv2v_reg  <= data_i[1];
    end 
    if(N898) begin
      \nz.mem_231_sv2v_reg  <= data_i[0];
    end 
    if(N897) begin
      \nz.mem_230_sv2v_reg  <= data_i[6];
    end 
    if(N896) begin
      \nz.mem_229_sv2v_reg  <= data_i[5];
    end 
    if(N895) begin
      \nz.mem_228_sv2v_reg  <= data_i[4];
    end 
    if(N894) begin
      \nz.mem_227_sv2v_reg  <= data_i[3];
    end 
    if(N893) begin
      \nz.mem_226_sv2v_reg  <= data_i[2];
    end 
    if(N892) begin
      \nz.mem_225_sv2v_reg  <= data_i[1];
    end 
    if(N891) begin
      \nz.mem_224_sv2v_reg  <= data_i[0];
    end 
    if(N890) begin
      \nz.mem_223_sv2v_reg  <= data_i[6];
    end 
    if(N889) begin
      \nz.mem_222_sv2v_reg  <= data_i[5];
    end 
    if(N888) begin
      \nz.mem_221_sv2v_reg  <= data_i[4];
    end 
    if(N887) begin
      \nz.mem_220_sv2v_reg  <= data_i[3];
    end 
    if(N886) begin
      \nz.mem_219_sv2v_reg  <= data_i[2];
    end 
    if(N885) begin
      \nz.mem_218_sv2v_reg  <= data_i[1];
    end 
    if(N884) begin
      \nz.mem_217_sv2v_reg  <= data_i[0];
    end 
    if(N883) begin
      \nz.mem_216_sv2v_reg  <= data_i[6];
    end 
    if(N882) begin
      \nz.mem_215_sv2v_reg  <= data_i[5];
    end 
    if(N881) begin
      \nz.mem_214_sv2v_reg  <= data_i[4];
    end 
    if(N880) begin
      \nz.mem_213_sv2v_reg  <= data_i[3];
    end 
    if(N879) begin
      \nz.mem_212_sv2v_reg  <= data_i[2];
    end 
    if(N878) begin
      \nz.mem_211_sv2v_reg  <= data_i[1];
    end 
    if(N877) begin
      \nz.mem_210_sv2v_reg  <= data_i[0];
    end 
    if(N876) begin
      \nz.mem_209_sv2v_reg  <= data_i[6];
    end 
    if(N875) begin
      \nz.mem_208_sv2v_reg  <= data_i[5];
    end 
    if(N874) begin
      \nz.mem_207_sv2v_reg  <= data_i[4];
    end 
    if(N873) begin
      \nz.mem_206_sv2v_reg  <= data_i[3];
    end 
    if(N872) begin
      \nz.mem_205_sv2v_reg  <= data_i[2];
    end 
    if(N871) begin
      \nz.mem_204_sv2v_reg  <= data_i[1];
    end 
    if(N870) begin
      \nz.mem_203_sv2v_reg  <= data_i[0];
    end 
    if(N869) begin
      \nz.mem_202_sv2v_reg  <= data_i[6];
    end 
    if(N868) begin
      \nz.mem_201_sv2v_reg  <= data_i[5];
    end 
    if(N867) begin
      \nz.mem_200_sv2v_reg  <= data_i[4];
    end 
    if(N866) begin
      \nz.mem_199_sv2v_reg  <= data_i[3];
    end 
    if(N865) begin
      \nz.mem_198_sv2v_reg  <= data_i[2];
    end 
    if(N864) begin
      \nz.mem_197_sv2v_reg  <= data_i[1];
    end 
    if(N863) begin
      \nz.mem_196_sv2v_reg  <= data_i[0];
    end 
    if(N862) begin
      \nz.mem_195_sv2v_reg  <= data_i[6];
    end 
    if(N861) begin
      \nz.mem_194_sv2v_reg  <= data_i[5];
    end 
    if(N860) begin
      \nz.mem_193_sv2v_reg  <= data_i[4];
    end 
    if(N859) begin
      \nz.mem_192_sv2v_reg  <= data_i[3];
    end 
    if(N858) begin
      \nz.mem_191_sv2v_reg  <= data_i[2];
    end 
    if(N857) begin
      \nz.mem_190_sv2v_reg  <= data_i[1];
    end 
    if(N856) begin
      \nz.mem_189_sv2v_reg  <= data_i[0];
    end 
    if(N855) begin
      \nz.mem_188_sv2v_reg  <= data_i[6];
    end 
    if(N854) begin
      \nz.mem_187_sv2v_reg  <= data_i[5];
    end 
    if(N853) begin
      \nz.mem_186_sv2v_reg  <= data_i[4];
    end 
    if(N852) begin
      \nz.mem_185_sv2v_reg  <= data_i[3];
    end 
    if(N851) begin
      \nz.mem_184_sv2v_reg  <= data_i[2];
    end 
    if(N850) begin
      \nz.mem_183_sv2v_reg  <= data_i[1];
    end 
    if(N849) begin
      \nz.mem_182_sv2v_reg  <= data_i[0];
    end 
    if(N848) begin
      \nz.mem_181_sv2v_reg  <= data_i[6];
    end 
    if(N847) begin
      \nz.mem_180_sv2v_reg  <= data_i[5];
    end 
    if(N846) begin
      \nz.mem_179_sv2v_reg  <= data_i[4];
    end 
    if(N845) begin
      \nz.mem_178_sv2v_reg  <= data_i[3];
    end 
    if(N844) begin
      \nz.mem_177_sv2v_reg  <= data_i[2];
    end 
    if(N843) begin
      \nz.mem_176_sv2v_reg  <= data_i[1];
    end 
    if(N842) begin
      \nz.mem_175_sv2v_reg  <= data_i[0];
    end 
    if(N841) begin
      \nz.mem_174_sv2v_reg  <= data_i[6];
    end 
    if(N840) begin
      \nz.mem_173_sv2v_reg  <= data_i[5];
    end 
    if(N839) begin
      \nz.mem_172_sv2v_reg  <= data_i[4];
    end 
    if(N838) begin
      \nz.mem_171_sv2v_reg  <= data_i[3];
    end 
    if(N837) begin
      \nz.mem_170_sv2v_reg  <= data_i[2];
    end 
    if(N836) begin
      \nz.mem_169_sv2v_reg  <= data_i[1];
    end 
    if(N835) begin
      \nz.mem_168_sv2v_reg  <= data_i[0];
    end 
    if(N834) begin
      \nz.mem_167_sv2v_reg  <= data_i[6];
    end 
    if(N833) begin
      \nz.mem_166_sv2v_reg  <= data_i[5];
    end 
    if(N832) begin
      \nz.mem_165_sv2v_reg  <= data_i[4];
    end 
    if(N831) begin
      \nz.mem_164_sv2v_reg  <= data_i[3];
    end 
    if(N830) begin
      \nz.mem_163_sv2v_reg  <= data_i[2];
    end 
    if(N829) begin
      \nz.mem_162_sv2v_reg  <= data_i[1];
    end 
    if(N828) begin
      \nz.mem_161_sv2v_reg  <= data_i[0];
    end 
    if(N827) begin
      \nz.mem_160_sv2v_reg  <= data_i[6];
    end 
    if(N826) begin
      \nz.mem_159_sv2v_reg  <= data_i[5];
    end 
    if(N825) begin
      \nz.mem_158_sv2v_reg  <= data_i[4];
    end 
    if(N824) begin
      \nz.mem_157_sv2v_reg  <= data_i[3];
    end 
    if(N823) begin
      \nz.mem_156_sv2v_reg  <= data_i[2];
    end 
    if(N822) begin
      \nz.mem_155_sv2v_reg  <= data_i[1];
    end 
    if(N821) begin
      \nz.mem_154_sv2v_reg  <= data_i[0];
    end 
    if(N820) begin
      \nz.mem_153_sv2v_reg  <= data_i[6];
    end 
    if(N819) begin
      \nz.mem_152_sv2v_reg  <= data_i[5];
    end 
    if(N818) begin
      \nz.mem_151_sv2v_reg  <= data_i[4];
    end 
    if(N817) begin
      \nz.mem_150_sv2v_reg  <= data_i[3];
    end 
    if(N816) begin
      \nz.mem_149_sv2v_reg  <= data_i[2];
    end 
    if(N815) begin
      \nz.mem_148_sv2v_reg  <= data_i[1];
    end 
    if(N814) begin
      \nz.mem_147_sv2v_reg  <= data_i[0];
    end 
    if(N813) begin
      \nz.mem_146_sv2v_reg  <= data_i[6];
    end 
    if(N812) begin
      \nz.mem_145_sv2v_reg  <= data_i[5];
    end 
    if(N811) begin
      \nz.mem_144_sv2v_reg  <= data_i[4];
    end 
    if(N810) begin
      \nz.mem_143_sv2v_reg  <= data_i[3];
    end 
    if(N809) begin
      \nz.mem_142_sv2v_reg  <= data_i[2];
    end 
    if(N808) begin
      \nz.mem_141_sv2v_reg  <= data_i[1];
    end 
    if(N807) begin
      \nz.mem_140_sv2v_reg  <= data_i[0];
    end 
    if(N806) begin
      \nz.mem_139_sv2v_reg  <= data_i[6];
    end 
    if(N805) begin
      \nz.mem_138_sv2v_reg  <= data_i[5];
    end 
    if(N804) begin
      \nz.mem_137_sv2v_reg  <= data_i[4];
    end 
    if(N803) begin
      \nz.mem_136_sv2v_reg  <= data_i[3];
    end 
    if(N802) begin
      \nz.mem_135_sv2v_reg  <= data_i[2];
    end 
    if(N801) begin
      \nz.mem_134_sv2v_reg  <= data_i[1];
    end 
    if(N800) begin
      \nz.mem_133_sv2v_reg  <= data_i[0];
    end 
    if(N799) begin
      \nz.mem_132_sv2v_reg  <= data_i[6];
    end 
    if(N798) begin
      \nz.mem_131_sv2v_reg  <= data_i[5];
    end 
    if(N797) begin
      \nz.mem_130_sv2v_reg  <= data_i[4];
    end 
    if(N796) begin
      \nz.mem_129_sv2v_reg  <= data_i[3];
    end 
    if(N795) begin
      \nz.mem_128_sv2v_reg  <= data_i[2];
    end 
    if(N794) begin
      \nz.mem_127_sv2v_reg  <= data_i[1];
    end 
    if(N793) begin
      \nz.mem_126_sv2v_reg  <= data_i[0];
    end 
    if(N792) begin
      \nz.mem_125_sv2v_reg  <= data_i[6];
    end 
    if(N791) begin
      \nz.mem_124_sv2v_reg  <= data_i[5];
    end 
    if(N790) begin
      \nz.mem_123_sv2v_reg  <= data_i[4];
    end 
    if(N789) begin
      \nz.mem_122_sv2v_reg  <= data_i[3];
    end 
    if(N788) begin
      \nz.mem_121_sv2v_reg  <= data_i[2];
    end 
    if(N787) begin
      \nz.mem_120_sv2v_reg  <= data_i[1];
    end 
    if(N786) begin
      \nz.mem_119_sv2v_reg  <= data_i[0];
    end 
    if(N785) begin
      \nz.mem_118_sv2v_reg  <= data_i[6];
    end 
    if(N784) begin
      \nz.mem_117_sv2v_reg  <= data_i[5];
    end 
    if(N783) begin
      \nz.mem_116_sv2v_reg  <= data_i[4];
    end 
    if(N782) begin
      \nz.mem_115_sv2v_reg  <= data_i[3];
    end 
    if(N781) begin
      \nz.mem_114_sv2v_reg  <= data_i[2];
    end 
    if(N780) begin
      \nz.mem_113_sv2v_reg  <= data_i[1];
    end 
    if(N779) begin
      \nz.mem_112_sv2v_reg  <= data_i[0];
    end 
    if(N778) begin
      \nz.mem_111_sv2v_reg  <= data_i[6];
    end 
    if(N777) begin
      \nz.mem_110_sv2v_reg  <= data_i[5];
    end 
    if(N776) begin
      \nz.mem_109_sv2v_reg  <= data_i[4];
    end 
    if(N775) begin
      \nz.mem_108_sv2v_reg  <= data_i[3];
    end 
    if(N774) begin
      \nz.mem_107_sv2v_reg  <= data_i[2];
    end 
    if(N773) begin
      \nz.mem_106_sv2v_reg  <= data_i[1];
    end 
    if(N772) begin
      \nz.mem_105_sv2v_reg  <= data_i[0];
    end 
    if(N771) begin
      \nz.mem_104_sv2v_reg  <= data_i[6];
    end 
    if(N770) begin
      \nz.mem_103_sv2v_reg  <= data_i[5];
    end 
    if(N769) begin
      \nz.mem_102_sv2v_reg  <= data_i[4];
    end 
    if(N768) begin
      \nz.mem_101_sv2v_reg  <= data_i[3];
    end 
    if(N767) begin
      \nz.mem_100_sv2v_reg  <= data_i[2];
    end 
    if(N766) begin
      \nz.mem_99_sv2v_reg  <= data_i[1];
    end 
    if(N765) begin
      \nz.mem_98_sv2v_reg  <= data_i[0];
    end 
    if(N764) begin
      \nz.mem_97_sv2v_reg  <= data_i[6];
    end 
    if(N763) begin
      \nz.mem_96_sv2v_reg  <= data_i[5];
    end 
    if(N762) begin
      \nz.mem_95_sv2v_reg  <= data_i[4];
    end 
    if(N761) begin
      \nz.mem_94_sv2v_reg  <= data_i[3];
    end 
    if(N760) begin
      \nz.mem_93_sv2v_reg  <= data_i[2];
    end 
    if(N759) begin
      \nz.mem_92_sv2v_reg  <= data_i[1];
    end 
    if(N758) begin
      \nz.mem_91_sv2v_reg  <= data_i[0];
    end 
    if(N757) begin
      \nz.mem_90_sv2v_reg  <= data_i[6];
    end 
    if(N756) begin
      \nz.mem_89_sv2v_reg  <= data_i[5];
    end 
    if(N755) begin
      \nz.mem_88_sv2v_reg  <= data_i[4];
    end 
    if(N754) begin
      \nz.mem_87_sv2v_reg  <= data_i[3];
    end 
    if(N753) begin
      \nz.mem_86_sv2v_reg  <= data_i[2];
    end 
    if(N752) begin
      \nz.mem_85_sv2v_reg  <= data_i[1];
    end 
    if(N751) begin
      \nz.mem_84_sv2v_reg  <= data_i[0];
    end 
    if(N750) begin
      \nz.mem_83_sv2v_reg  <= data_i[6];
    end 
    if(N749) begin
      \nz.mem_82_sv2v_reg  <= data_i[5];
    end 
    if(N748) begin
      \nz.mem_81_sv2v_reg  <= data_i[4];
    end 
    if(N747) begin
      \nz.mem_80_sv2v_reg  <= data_i[3];
    end 
    if(N746) begin
      \nz.mem_79_sv2v_reg  <= data_i[2];
    end 
    if(N745) begin
      \nz.mem_78_sv2v_reg  <= data_i[1];
    end 
    if(N744) begin
      \nz.mem_77_sv2v_reg  <= data_i[0];
    end 
    if(N743) begin
      \nz.mem_76_sv2v_reg  <= data_i[6];
    end 
    if(N742) begin
      \nz.mem_75_sv2v_reg  <= data_i[5];
    end 
    if(N741) begin
      \nz.mem_74_sv2v_reg  <= data_i[4];
    end 
    if(N740) begin
      \nz.mem_73_sv2v_reg  <= data_i[3];
    end 
    if(N739) begin
      \nz.mem_72_sv2v_reg  <= data_i[2];
    end 
    if(N738) begin
      \nz.mem_71_sv2v_reg  <= data_i[1];
    end 
    if(N737) begin
      \nz.mem_70_sv2v_reg  <= data_i[0];
    end 
    if(N736) begin
      \nz.mem_69_sv2v_reg  <= data_i[6];
    end 
    if(N735) begin
      \nz.mem_68_sv2v_reg  <= data_i[5];
    end 
    if(N734) begin
      \nz.mem_67_sv2v_reg  <= data_i[4];
    end 
    if(N733) begin
      \nz.mem_66_sv2v_reg  <= data_i[3];
    end 
    if(N732) begin
      \nz.mem_65_sv2v_reg  <= data_i[2];
    end 
    if(N731) begin
      \nz.mem_64_sv2v_reg  <= data_i[1];
    end 
    if(N730) begin
      \nz.mem_63_sv2v_reg  <= data_i[0];
    end 
    if(N729) begin
      \nz.mem_62_sv2v_reg  <= data_i[6];
    end 
    if(N728) begin
      \nz.mem_61_sv2v_reg  <= data_i[5];
    end 
    if(N727) begin
      \nz.mem_60_sv2v_reg  <= data_i[4];
    end 
    if(N726) begin
      \nz.mem_59_sv2v_reg  <= data_i[3];
    end 
    if(N725) begin
      \nz.mem_58_sv2v_reg  <= data_i[2];
    end 
    if(N724) begin
      \nz.mem_57_sv2v_reg  <= data_i[1];
    end 
    if(N723) begin
      \nz.mem_56_sv2v_reg  <= data_i[0];
    end 
    if(N722) begin
      \nz.mem_55_sv2v_reg  <= data_i[6];
    end 
    if(N721) begin
      \nz.mem_54_sv2v_reg  <= data_i[5];
    end 
    if(N720) begin
      \nz.mem_53_sv2v_reg  <= data_i[4];
    end 
    if(N719) begin
      \nz.mem_52_sv2v_reg  <= data_i[3];
    end 
    if(N718) begin
      \nz.mem_51_sv2v_reg  <= data_i[2];
    end 
    if(N717) begin
      \nz.mem_50_sv2v_reg  <= data_i[1];
    end 
    if(N716) begin
      \nz.mem_49_sv2v_reg  <= data_i[0];
    end 
    if(N715) begin
      \nz.mem_48_sv2v_reg  <= data_i[6];
    end 
    if(N714) begin
      \nz.mem_47_sv2v_reg  <= data_i[5];
    end 
    if(N713) begin
      \nz.mem_46_sv2v_reg  <= data_i[4];
    end 
    if(N712) begin
      \nz.mem_45_sv2v_reg  <= data_i[3];
    end 
    if(N711) begin
      \nz.mem_44_sv2v_reg  <= data_i[2];
    end 
    if(N710) begin
      \nz.mem_43_sv2v_reg  <= data_i[1];
    end 
    if(N709) begin
      \nz.mem_42_sv2v_reg  <= data_i[0];
    end 
    if(N708) begin
      \nz.mem_41_sv2v_reg  <= data_i[6];
    end 
    if(N707) begin
      \nz.mem_40_sv2v_reg  <= data_i[5];
    end 
    if(N706) begin
      \nz.mem_39_sv2v_reg  <= data_i[4];
    end 
    if(N705) begin
      \nz.mem_38_sv2v_reg  <= data_i[3];
    end 
    if(N704) begin
      \nz.mem_37_sv2v_reg  <= data_i[2];
    end 
    if(N703) begin
      \nz.mem_36_sv2v_reg  <= data_i[1];
    end 
    if(N702) begin
      \nz.mem_35_sv2v_reg  <= data_i[0];
    end 
    if(N701) begin
      \nz.mem_34_sv2v_reg  <= data_i[6];
    end 
    if(N700) begin
      \nz.mem_33_sv2v_reg  <= data_i[5];
    end 
    if(N699) begin
      \nz.mem_32_sv2v_reg  <= data_i[4];
    end 
    if(N698) begin
      \nz.mem_31_sv2v_reg  <= data_i[3];
    end 
    if(N697) begin
      \nz.mem_30_sv2v_reg  <= data_i[2];
    end 
    if(N696) begin
      \nz.mem_29_sv2v_reg  <= data_i[1];
    end 
    if(N695) begin
      \nz.mem_28_sv2v_reg  <= data_i[0];
    end 
    if(N694) begin
      \nz.mem_27_sv2v_reg  <= data_i[6];
    end 
    if(N693) begin
      \nz.mem_26_sv2v_reg  <= data_i[5];
    end 
    if(N692) begin
      \nz.mem_25_sv2v_reg  <= data_i[4];
    end 
    if(N691) begin
      \nz.mem_24_sv2v_reg  <= data_i[3];
    end 
    if(N690) begin
      \nz.mem_23_sv2v_reg  <= data_i[2];
    end 
    if(N689) begin
      \nz.mem_22_sv2v_reg  <= data_i[1];
    end 
    if(N688) begin
      \nz.mem_21_sv2v_reg  <= data_i[0];
    end 
    if(N687) begin
      \nz.mem_20_sv2v_reg  <= data_i[6];
    end 
    if(N686) begin
      \nz.mem_19_sv2v_reg  <= data_i[5];
    end 
    if(N685) begin
      \nz.mem_18_sv2v_reg  <= data_i[4];
    end 
    if(N684) begin
      \nz.mem_17_sv2v_reg  <= data_i[3];
    end 
    if(N683) begin
      \nz.mem_16_sv2v_reg  <= data_i[2];
    end 
    if(N682) begin
      \nz.mem_15_sv2v_reg  <= data_i[1];
    end 
    if(N681) begin
      \nz.mem_14_sv2v_reg  <= data_i[0];
    end 
    if(N680) begin
      \nz.mem_13_sv2v_reg  <= data_i[6];
    end 
    if(N679) begin
      \nz.mem_12_sv2v_reg  <= data_i[5];
    end 
    if(N678) begin
      \nz.mem_11_sv2v_reg  <= data_i[4];
    end 
    if(N677) begin
      \nz.mem_10_sv2v_reg  <= data_i[3];
    end 
    if(N676) begin
      \nz.mem_9_sv2v_reg  <= data_i[2];
    end 
    if(N675) begin
      \nz.mem_8_sv2v_reg  <= data_i[1];
    end 
    if(N674) begin
      \nz.mem_7_sv2v_reg  <= data_i[0];
    end 
    if(N673) begin
      \nz.mem_6_sv2v_reg  <= data_i[6];
    end 
    if(N672) begin
      \nz.mem_5_sv2v_reg  <= data_i[5];
    end 
    if(N671) begin
      \nz.mem_4_sv2v_reg  <= data_i[4];
    end 
    if(N670) begin
      \nz.mem_3_sv2v_reg  <= data_i[3];
    end 
    if(N669) begin
      \nz.mem_2_sv2v_reg  <= data_i[2];
    end 
    if(N668) begin
      \nz.mem_1_sv2v_reg  <= data_i[1];
    end 
    if(N667) begin
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p7_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_lru_pseudo_tree_decode_ways_p4
(
  way_id_i,
  data_o,
  mask_o
);

  input [1:0] way_id_i;
  output [2:0] data_o;
  output [2:0] mask_o;
  wire [2:0] data_o,mask_o;
  wire N0,N1;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[1];
  assign mask_o[1] = 1'b1 & N0;
  assign data_o[1] = mask_o[1] & N1;
  assign N1 = ~way_id_i[0];
  assign mask_o[2] = 1'b1 & way_id_i[1];
  assign data_o[2] = mask_o[2] & N1;

endmodule



module bsg_mux_width_p1_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [1:0] data_i;
  input [0:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[1] : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = ~sel_i[0];

endmodule



module bsg_lru_pseudo_tree_encode_ways_p4
(
  lru_i,
  way_id_o
);

  input [2:0] lru_i;
  output [1:0] way_id_o;
  wire [1:0] way_id_o;
  wire way_id_o_1_;
  assign way_id_o_1_ = lru_i[0];
  assign way_id_o[1] = way_id_o_1_;

  bsg_mux_width_p1_els_p2
  \lru.rank_1_.nz.mux 
  (
    .data_i(lru_i[2:1]),
    .sel_i(way_id_o_1_),
    .data_o(way_id_o[0])
  );


endmodule



module bsg_decode_num_out_p4
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4_word_tracking_p1
(
  clk_i,
  reset_i,
  miss_v_i,
  track_miss_i,
  decode_v_i,
  addr_v_i,
  mask_v_i,
  tag_v_i,
  valid_v_i,
  lock_v_i,
  tag_hit_v_i,
  tag_hit_way_id_i,
  tag_hit_found_i,
  sbuf_empty_i,
  tbuf_empty_i,
  dma_cmd_o,
  dma_way_o,
  dma_addr_o,
  dma_done_i,
  track_data_we_o,
  stat_info_i,
  stat_mem_v_o,
  stat_mem_w_o,
  stat_mem_addr_o,
  stat_mem_data_o,
  stat_mem_w_mask_o,
  tag_mem_v_o,
  tag_mem_w_o,
  tag_mem_addr_o,
  tag_mem_data_o,
  tag_mem_w_mask_o,
  track_mem_v_o,
  track_mem_w_o,
  track_mem_addr_o,
  track_mem_w_mask_o,
  track_mem_data_o,
  done_o,
  recover_o,
  chosen_way_o,
  select_snoop_data_r_o,
  ack_i
);

  input [20:0] decode_v_i;
  input [27:0] addr_v_i;
  input [3:0] mask_v_i;
  input [71:0] tag_v_i;
  input [3:0] valid_v_i;
  input [3:0] lock_v_i;
  input [3:0] tag_hit_v_i;
  input [1:0] tag_hit_way_id_i;
  output [3:0] dma_cmd_o;
  output [1:0] dma_way_o;
  output [27:0] dma_addr_o;
  input [6:0] stat_info_i;
  output [5:0] stat_mem_addr_o;
  output [6:0] stat_mem_data_o;
  output [6:0] stat_mem_w_mask_o;
  output [5:0] tag_mem_addr_o;
  output [79:0] tag_mem_data_o;
  output [79:0] tag_mem_w_mask_o;
  output [5:0] track_mem_addr_o;
  output [15:0] track_mem_w_mask_o;
  output [15:0] track_mem_data_o;
  output [1:0] chosen_way_o;
  input clk_i;
  input reset_i;
  input miss_v_i;
  input track_miss_i;
  input tag_hit_found_i;
  input sbuf_empty_i;
  input tbuf_empty_i;
  input dma_done_i;
  input ack_i;
  output track_data_we_o;
  output stat_mem_v_o;
  output stat_mem_w_o;
  output tag_mem_v_o;
  output tag_mem_w_o;
  output track_mem_v_o;
  output track_mem_w_o;
  output done_o;
  output recover_o;
  output select_snoop_data_r_o;
  wire [3:0] dma_cmd_o,chosen_way_decode,addr_way_v_decode,flush_way_decode,miss_state_r,
  miss_state_n;
  wire [1:0] dma_way_o,chosen_way_o,invalid_way_id,flush_way_r,lru_way_id,chosen_way_n;
  wire [27:0] dma_addr_o;
  wire [5:0] stat_mem_addr_o,tag_mem_addr_o,track_mem_addr_o;
  wire [6:0] stat_mem_data_o,stat_mem_w_mask_o;
  wire [79:0] tag_mem_data_o,tag_mem_w_mask_o;
  wire [15:0] track_mem_w_mask_o,track_mem_data_o;
  wire track_data_we_o,stat_mem_v_o,stat_mem_w_o,tag_mem_v_o,tag_mem_w_o,track_mem_v_o,
  track_mem_w_o,done_o,recover_o,select_snoop_data_r_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,track_mem_data_o_3__3_,
  _0_net__3_,_0_net__2_,_0_net__1_,_0_net__0_,invalid_exist,goto_flush_op,
  goto_lock_op,N23,N24,full_word_op,st_tag_miss_op,N25,N26,select_snoop_data_n,N27,N28,N29,
  N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,
  N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,
  N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,
  N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,
  N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,
  N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,
  N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264;
  wire [2:0] chosen_way_lru_data,chosen_way_lru_mask,modify_mask_lo,modify_data_lo,
  modified_lru_bits;
  reg track_data_we_o_sv2v_reg,miss_state_r_3_sv2v_reg,miss_state_r_2_sv2v_reg,
  miss_state_r_1_sv2v_reg,miss_state_r_0_sv2v_reg,chosen_way_o_1_sv2v_reg,
  chosen_way_o_0_sv2v_reg,flush_way_r_1_sv2v_reg,flush_way_r_0_sv2v_reg,
  select_snoop_data_r_o_sv2v_reg;
  assign track_data_we_o = track_data_we_o_sv2v_reg;
  assign miss_state_r[3] = miss_state_r_3_sv2v_reg;
  assign miss_state_r[2] = miss_state_r_2_sv2v_reg;
  assign miss_state_r[1] = miss_state_r_1_sv2v_reg;
  assign miss_state_r[0] = miss_state_r_0_sv2v_reg;
  assign chosen_way_o[1] = chosen_way_o_1_sv2v_reg;
  assign chosen_way_o[0] = chosen_way_o_0_sv2v_reg;
  assign flush_way_r[1] = flush_way_r_1_sv2v_reg;
  assign flush_way_r[0] = flush_way_r_0_sv2v_reg;
  assign select_snoop_data_r_o = select_snoop_data_r_o_sv2v_reg;
  assign dma_addr_o[0] = 1'b0;
  assign dma_addr_o[1] = 1'b0;
  assign stat_mem_addr_o[5] = addr_v_i[9];
  assign track_mem_addr_o[5] = stat_mem_addr_o[5];
  assign tag_mem_addr_o[5] = stat_mem_addr_o[5];
  assign stat_mem_addr_o[4] = addr_v_i[8];
  assign track_mem_addr_o[4] = stat_mem_addr_o[4];
  assign tag_mem_addr_o[4] = stat_mem_addr_o[4];
  assign stat_mem_addr_o[3] = addr_v_i[7];
  assign track_mem_addr_o[3] = stat_mem_addr_o[3];
  assign tag_mem_addr_o[3] = stat_mem_addr_o[3];
  assign stat_mem_addr_o[2] = addr_v_i[6];
  assign track_mem_addr_o[2] = stat_mem_addr_o[2];
  assign tag_mem_addr_o[2] = stat_mem_addr_o[2];
  assign stat_mem_addr_o[1] = addr_v_i[5];
  assign track_mem_addr_o[1] = stat_mem_addr_o[1];
  assign tag_mem_addr_o[1] = stat_mem_addr_o[1];
  assign stat_mem_addr_o[0] = addr_v_i[4];
  assign track_mem_addr_o[0] = stat_mem_addr_o[0];
  assign tag_mem_addr_o[0] = stat_mem_addr_o[0];
  assign dma_cmd_o[2] = track_mem_data_o_3__3_;
  assign track_mem_data_o[0] = track_mem_data_o_3__3_;
  assign track_mem_data_o[1] = track_mem_data_o_3__3_;
  assign track_mem_data_o[2] = track_mem_data_o_3__3_;
  assign track_mem_data_o[3] = track_mem_data_o_3__3_;
  assign track_mem_data_o[4] = track_mem_data_o_3__3_;
  assign track_mem_data_o[5] = track_mem_data_o_3__3_;
  assign track_mem_data_o[6] = track_mem_data_o_3__3_;
  assign track_mem_data_o[7] = track_mem_data_o_3__3_;
  assign track_mem_data_o[8] = track_mem_data_o_3__3_;
  assign track_mem_data_o[9] = track_mem_data_o_3__3_;
  assign track_mem_data_o[10] = track_mem_data_o_3__3_;
  assign track_mem_data_o[11] = track_mem_data_o_3__3_;
  assign track_mem_data_o[12] = track_mem_data_o_3__3_;
  assign track_mem_data_o[13] = track_mem_data_o_3__3_;
  assign track_mem_data_o[14] = track_mem_data_o_3__3_;
  assign track_mem_data_o[15] = track_mem_data_o_3__3_;

  bsg_priority_encode_width_p4_lo_to_hi_p1
  invalid_way_pe
  (
    .i({ _0_net__3_, _0_net__2_, _0_net__1_, _0_net__0_ }),
    .addr_o(invalid_way_id),
    .v_o(invalid_exist)
  );


  bsg_lru_pseudo_tree_decode_ways_p4
  chosen_way_lru_decode
  (
    .way_id_i(chosen_way_o),
    .data_o(chosen_way_lru_data),
    .mask_o(chosen_way_lru_mask)
  );


  bsg_lru_pseudo_tree_backup
  backup_lru
  (
    .disabled_ways_i(lock_v_i),
    .modify_mask_o(modify_mask_lo),
    .modify_data_o(modify_data_lo)
  );


  bsg_mux_bitwise
  lru_bit_mux
  (
    .data0_i(stat_info_i[2:0]),
    .data1_i(modify_data_lo),
    .sel_i(modify_mask_lo),
    .data_o(modified_lru_bits)
  );


  bsg_lru_pseudo_tree_encode_ways_p4
  lru_encode
  (
    .lru_i(modified_lru_bits),
    .way_id_o(lru_way_id)
  );


  bsg_decode_num_out_p4
  chosen_way_demux
  (
    .i(chosen_way_n),
    .o(chosen_way_decode)
  );


  bsg_decode_num_out_p4
  addr_way_v_demux
  (
    .i(addr_v_i[11:10]),
    .o(addr_way_v_decode)
  );

  assign N31 = N27 & N28;
  assign N32 = N29 & N30;
  assign N33 = N31 & N32;
  assign N34 = miss_state_r[3] | N28;
  assign N35 = miss_state_r[1] | miss_state_r[0];
  assign N36 = N34 | N35;
  assign N38 = miss_state_r[3] | miss_state_r[2];
  assign N39 = miss_state_r[1] | N30;
  assign N40 = N38 | N39;
  assign N42 = miss_state_r[3] | miss_state_r[2];
  assign N43 = N29 | miss_state_r[0];
  assign N44 = N42 | N43;
  assign N46 = miss_state_r[3] | miss_state_r[2];
  assign N47 = N29 | N30;
  assign N48 = N46 | N47;
  assign N50 = miss_state_r[3] | N28;
  assign N51 = miss_state_r[1] | N30;
  assign N52 = N50 | N51;
  assign N54 = miss_state_r[3] | N28;
  assign N55 = N29 | miss_state_r[0];
  assign N56 = N54 | N55;
  assign N58 = miss_state_r[3] | N28;
  assign N59 = N29 | N30;
  assign N60 = N58 | N59;
  assign N62 = N27 | miss_state_r[2];
  assign N63 = miss_state_r[1] | miss_state_r[0];
  assign N64 = N62 | N63;
  assign N66 = N27 | miss_state_r[2];
  assign N67 = miss_state_r[1] | N30;
  assign N68 = N66 | N67;
  assign N70 = N27 | miss_state_r[2];
  assign N71 = N29 | miss_state_r[0];
  assign N72 = N70 | N71;
  assign N74 = miss_state_r[3] & miss_state_r[1];
  assign N75 = N74 & miss_state_r[0];
  assign N76 = miss_state_r[3] & miss_state_r[2];
  assign N99 = (N95)? stat_info_i[3] : 
               (N97)? stat_info_i[4] : 
               (N96)? stat_info_i[5] : 
               (N98)? stat_info_i[6] : 1'b0;
  assign N100 = (N95)? valid_v_i[0] : 
                (N97)? valid_v_i[1] : 
                (N96)? valid_v_i[2] : 
                (N98)? valid_v_i[3] : 1'b0;
  assign N121 = (N117)? stat_info_i[3] : 
                (N119)? stat_info_i[4] : 
                (N118)? stat_info_i[5] : 
                (N120)? stat_info_i[6] : 1'b0;
  assign N122 = (N117)? valid_v_i[0] : 
                (N119)? valid_v_i[1] : 
                (N118)? valid_v_i[2] : 
                (N120)? valid_v_i[3] : 1'b0;
  assign N131 = (N127)? tag_v_i[17] : 
                (N129)? tag_v_i[35] : 
                (N128)? tag_v_i[53] : 
                (N130)? tag_v_i[71] : 1'b0;
  assign N132 = (N127)? tag_v_i[16] : 
                (N129)? tag_v_i[34] : 
                (N128)? tag_v_i[52] : 
                (N130)? tag_v_i[70] : 1'b0;
  assign N133 = (N127)? tag_v_i[15] : 
                (N129)? tag_v_i[33] : 
                (N128)? tag_v_i[51] : 
                (N130)? tag_v_i[69] : 1'b0;
  assign N134 = (N127)? tag_v_i[14] : 
                (N129)? tag_v_i[32] : 
                (N128)? tag_v_i[50] : 
                (N130)? tag_v_i[68] : 1'b0;
  assign N135 = (N127)? tag_v_i[13] : 
                (N129)? tag_v_i[31] : 
                (N128)? tag_v_i[49] : 
                (N130)? tag_v_i[67] : 1'b0;
  assign N136 = (N127)? tag_v_i[12] : 
                (N129)? tag_v_i[30] : 
                (N128)? tag_v_i[48] : 
                (N130)? tag_v_i[66] : 1'b0;
  assign N137 = (N127)? tag_v_i[11] : 
                (N129)? tag_v_i[29] : 
                (N128)? tag_v_i[47] : 
                (N130)? tag_v_i[65] : 1'b0;
  assign N138 = (N127)? tag_v_i[10] : 
                (N129)? tag_v_i[28] : 
                (N128)? tag_v_i[46] : 
                (N130)? tag_v_i[64] : 1'b0;
  assign N139 = (N127)? tag_v_i[9] : 
                (N129)? tag_v_i[27] : 
                (N128)? tag_v_i[45] : 
                (N130)? tag_v_i[63] : 1'b0;
  assign N140 = (N127)? tag_v_i[8] : 
                (N129)? tag_v_i[26] : 
                (N128)? tag_v_i[44] : 
                (N130)? tag_v_i[62] : 1'b0;
  assign N141 = (N127)? tag_v_i[7] : 
                (N129)? tag_v_i[25] : 
                (N128)? tag_v_i[43] : 
                (N130)? tag_v_i[61] : 1'b0;
  assign N142 = (N127)? tag_v_i[6] : 
                (N129)? tag_v_i[24] : 
                (N128)? tag_v_i[42] : 
                (N130)? tag_v_i[60] : 1'b0;
  assign N143 = (N127)? tag_v_i[5] : 
                (N129)? tag_v_i[23] : 
                (N128)? tag_v_i[41] : 
                (N130)? tag_v_i[59] : 1'b0;
  assign N144 = (N127)? tag_v_i[4] : 
                (N129)? tag_v_i[22] : 
                (N128)? tag_v_i[40] : 
                (N130)? tag_v_i[58] : 1'b0;
  assign N145 = (N127)? tag_v_i[3] : 
                (N129)? tag_v_i[21] : 
                (N128)? tag_v_i[39] : 
                (N130)? tag_v_i[57] : 1'b0;
  assign N146 = (N127)? tag_v_i[2] : 
                (N129)? tag_v_i[20] : 
                (N128)? tag_v_i[38] : 
                (N130)? tag_v_i[56] : 1'b0;
  assign N147 = (N127)? tag_v_i[1] : 
                (N129)? tag_v_i[19] : 
                (N128)? tag_v_i[37] : 
                (N130)? tag_v_i[55] : 1'b0;
  assign N148 = (N127)? tag_v_i[0] : 
                (N129)? tag_v_i[18] : 
                (N128)? tag_v_i[36] : 
                (N130)? tag_v_i[54] : 1'b0;
  assign N154 = (N150)? tag_v_i[17] : 
                (N152)? tag_v_i[35] : 
                (N151)? tag_v_i[53] : 
                (N153)? tag_v_i[71] : 1'b0;
  assign N155 = (N150)? tag_v_i[16] : 
                (N152)? tag_v_i[34] : 
                (N151)? tag_v_i[52] : 
                (N153)? tag_v_i[70] : 1'b0;
  assign N156 = (N150)? tag_v_i[15] : 
                (N152)? tag_v_i[33] : 
                (N151)? tag_v_i[51] : 
                (N153)? tag_v_i[69] : 1'b0;
  assign N157 = (N150)? tag_v_i[14] : 
                (N152)? tag_v_i[32] : 
                (N151)? tag_v_i[50] : 
                (N153)? tag_v_i[68] : 1'b0;
  assign N158 = (N150)? tag_v_i[13] : 
                (N152)? tag_v_i[31] : 
                (N151)? tag_v_i[49] : 
                (N153)? tag_v_i[67] : 1'b0;
  assign N159 = (N150)? tag_v_i[12] : 
                (N152)? tag_v_i[30] : 
                (N151)? tag_v_i[48] : 
                (N153)? tag_v_i[66] : 1'b0;
  assign N160 = (N150)? tag_v_i[11] : 
                (N152)? tag_v_i[29] : 
                (N151)? tag_v_i[47] : 
                (N153)? tag_v_i[65] : 1'b0;
  assign N161 = (N150)? tag_v_i[10] : 
                (N152)? tag_v_i[28] : 
                (N151)? tag_v_i[46] : 
                (N153)? tag_v_i[64] : 1'b0;
  assign N162 = (N150)? tag_v_i[9] : 
                (N152)? tag_v_i[27] : 
                (N151)? tag_v_i[45] : 
                (N153)? tag_v_i[63] : 1'b0;
  assign N163 = (N150)? tag_v_i[8] : 
                (N152)? tag_v_i[26] : 
                (N151)? tag_v_i[44] : 
                (N153)? tag_v_i[62] : 1'b0;
  assign N164 = (N150)? tag_v_i[7] : 
                (N152)? tag_v_i[25] : 
                (N151)? tag_v_i[43] : 
                (N153)? tag_v_i[61] : 1'b0;
  assign N165 = (N150)? tag_v_i[6] : 
                (N152)? tag_v_i[24] : 
                (N151)? tag_v_i[42] : 
                (N153)? tag_v_i[60] : 1'b0;
  assign N166 = (N150)? tag_v_i[5] : 
                (N152)? tag_v_i[23] : 
                (N151)? tag_v_i[41] : 
                (N153)? tag_v_i[59] : 1'b0;
  assign N167 = (N150)? tag_v_i[4] : 
                (N152)? tag_v_i[22] : 
                (N151)? tag_v_i[40] : 
                (N153)? tag_v_i[58] : 1'b0;
  assign N168 = (N150)? tag_v_i[3] : 
                (N152)? tag_v_i[21] : 
                (N151)? tag_v_i[39] : 
                (N153)? tag_v_i[57] : 1'b0;
  assign N169 = (N150)? tag_v_i[2] : 
                (N152)? tag_v_i[20] : 
                (N151)? tag_v_i[38] : 
                (N153)? tag_v_i[56] : 1'b0;
  assign N170 = (N150)? tag_v_i[1] : 
                (N152)? tag_v_i[19] : 
                (N151)? tag_v_i[37] : 
                (N153)? tag_v_i[55] : 1'b0;
  assign N171 = (N150)? tag_v_i[0] : 
                (N152)? tag_v_i[18] : 
                (N151)? tag_v_i[36] : 
                (N153)? tag_v_i[54] : 1'b0;
  assign N195 = (N191)? stat_info_i[3] : 
                (N193)? stat_info_i[4] : 
                (N192)? stat_info_i[5] : 
                (N194)? stat_info_i[6] : 1'b0;
  assign N196 = (N191)? valid_v_i[0] : 
                (N193)? valid_v_i[1] : 
                (N192)? valid_v_i[2] : 
                (N194)? valid_v_i[3] : 1'b0;
  assign full_word_op = (N0)? N24 : 
                        (N23)? decode_v_i[20] : 1'b0;
  assign N0 = decode_v_i[17];
  assign dma_way_o = (N1)? flush_way_r : 
                     (N2)? chosen_way_o : 1'b0;
  assign N1 = goto_flush_op;
  assign N2 = N25;
  assign flush_way_decode = (N3)? addr_way_v_decode : 
                            (N26)? tag_hit_v_i : 1'b0;
  assign N3 = decode_v_i[13];
  assign { N85, N84, N83 } = (N1)? { 1'b0, 1'b0, 1'b1 } : 
                             (N203)? { 1'b0, 1'b1, 1'b0 } : 
                             (N206)? { 1'b1, 1'b1, 1'b1 } : 
                             (N82)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign { N88, N87, N86 } = (N4)? { N85, N84, N83 } : 
                             (N79)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = N78;
  assign { N92, N91 } = (N5)? tag_hit_way_id_i : 
                        (N208)? invalid_way_id : 
                        (N90)? lru_way_id : 1'b0;
  assign N5 = track_miss_i;
  assign N102 = ~N101;
  assign { N104, N103 } = (N6)? { N102, N101 } : 
                          (N7)? { 1'b1, 1'b0 } : 1'b0;
  assign N6 = dma_done_i;
  assign N7 = N149;
  assign { N106, N105 } = (N3)? addr_v_i[11:10] : 
                          (N26)? tag_hit_way_id_i : 1'b0;
  assign N124 = ~N123;
  assign N176 = ~N175;
  assign { N180, N179, N178, N177 } = (N6)? { N175, N176, N176, N175 } : 
                                      (N7)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign { N185, N184, N183, N182 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N8)? chosen_way_decode : 1'b0;
  assign N8 = N250;
  assign { N188, N187 } = (N9)? invalid_way_id : 
                          (N10)? lru_way_id : 1'b0;
  assign N9 = invalid_exist;
  assign N10 = N186;
  assign N198 = ~N197;
  assign stat_mem_v_o = (N11)? N78 : 
                        (N12)? 1'b0 : 
                        (N13)? 1'b1 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? N172 : 
                        (N17)? dma_done_i : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b1 : 
                        (N20)? 1'b0 : 
                        (N21)? 1'b0 : 
                        (N22)? 1'b0 : 1'b0;
  assign N11 = N33;
  assign N12 = dma_cmd_o[0];
  assign N13 = N41;
  assign N14 = N45;
  assign N15 = dma_cmd_o[1];
  assign N16 = dma_cmd_o[3];
  assign N17 = track_mem_data_o_3__3_;
  assign N18 = N61;
  assign N19 = N65;
  assign N20 = N69;
  assign N21 = N73;
  assign N22 = N77;
  assign track_mem_v_o = (N11)? N78 : 
                         (N12)? 1'b0 : 
                         (N13)? 1'b0 : 
                         (N14)? 1'b0 : 
                         (N15)? 1'b0 : 
                         (N16)? N174 : 
                         (N17)? dma_done_i : 
                         (N18)? 1'b0 : 
                         (N19)? 1'b1 : 
                         (N20)? 1'b0 : 
                         (N21)? 1'b0 : 
                         (N22)? 1'b0 : 1'b0;
  assign miss_state_n = (N11)? { 1'b0, N88, N87, N86 } : 
                        (N12)? { 1'b0, N104, dma_done_i, N103 } : 
                        (N13)? { N124, 1'b0, N123, 1'b1 } : 
                        (N14)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                        (N15)? { 1'b0, dma_done_i, N149, 1'b1 } : 
                        (N16)? { N180, N179, N178, N177 } : 
                        (N17)? { dma_done_i, N149, N149, dma_done_i } : 
                        (N18)? { N198, 1'b0, N197, N197 } : 
                        (N19)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                        (N20)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                        (N21)? { N199, 1'b0, N199, 1'b0 } : 
                        (N22)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign chosen_way_n = (N11)? chosen_way_o : 
                        (N12)? { N92, N91 } : 
                        (N13)? chosen_way_o : 
                        (N14)? chosen_way_o : 
                        (N15)? chosen_way_o : 
                        (N16)? chosen_way_o : 
                        (N17)? chosen_way_o : 
                        (N18)? { N188, N187 } : 
                        (N19)? chosen_way_o : 
                        (N20)? chosen_way_o : 
                        (N21)? chosen_way_o : 
                        (N22)? chosen_way_o : 1'b0;
  assign dma_addr_o[3:2] = (N17)? addr_v_i[3:2] : 
                           (N201)? { 1'b0, 1'b0 } : 1'b0;
  assign dma_addr_o[27:4] = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N12)? { addr_v_i[27:10], stat_mem_addr_o } : 
                            (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N15)? { N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, stat_mem_addr_o } : 
                            (N16)? { N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, stat_mem_addr_o } : 
                            (N17)? { addr_v_i[27:10], stat_mem_addr_o } : 
                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_o = (N11)? 1'b0 : 
                        (N12)? 1'b0 : 
                        (N13)? 1'b1 : 
                        (N14)? 1'b0 : 
                        (N15)? 1'b0 : 
                        (N16)? 1'b1 : 
                        (N17)? 1'b1 : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b1 : 
                        (N20)? 1'b0 : 
                        (N21)? 1'b0 : 
                        (N22)? 1'b0 : 1'b0;
  assign stat_mem_data_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, chosen_way_lru_data } : 
                           (N17)? { N181, N181, N181, N181, chosen_way_lru_data } : 
                           (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N19)? { 1'b1, 1'b1, 1'b1, 1'b1, chosen_way_lru_data } : 
                           (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                           (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N13)? { flush_way_decode, 1'b0, 1'b0, 1'b0 } : 
                             (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N16)? { chosen_way_decode, chosen_way_lru_mask } : 
                             (N17)? { N185, N184, N183, N182, chosen_way_lru_mask } : 
                             (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N19)? { chosen_way_decode, chosen_way_lru_mask } : 
                             (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_v_o = (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b1 : 
                       (N14)? 1'b1 : 
                       (N15)? 1'b0 : 
                       (N16)? N173 : 
                       (N17)? dma_done_i : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b1 : 
                       (N20)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 1'b0;
  assign tag_mem_w_o = (N11)? 1'b0 : 
                       (N12)? 1'b0 : 
                       (N13)? 1'b1 : 
                       (N14)? 1'b1 : 
                       (N15)? 1'b0 : 
                       (N16)? 1'b1 : 
                       (N17)? 1'b1 : 
                       (N18)? 1'b0 : 
                       (N19)? 1'b1 : 
                       (N20)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 1'b0;
  assign tag_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N13)? { N113, N114, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N111, N112, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N109, N110, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N107, N108, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N14)? { 1'b0, tag_hit_v_i[3:3], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[2:2], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N16)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N17)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_data_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N14)? { 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N16)? { 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10] } : 
                          (N17)? { 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10] } : 
                          (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N19)? { 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10] } : 
                          (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign track_mem_w_o = (N11)? 1'b0 : 
                         (N12)? 1'b0 : 
                         (N13)? 1'b0 : 
                         (N14)? 1'b0 : 
                         (N15)? 1'b0 : 
                         (N16)? 1'b1 : 
                         (N17)? 1'b1 : 
                         (N18)? 1'b0 : 
                         (N19)? 1'b1 : 
                         (N20)? 1'b0 : 
                         (N21)? 1'b0 : 
                         (N22)? 1'b0 : 1'b0;
  assign track_mem_w_mask_o = (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N16)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N17)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N19)? { chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:3], chosen_way_decode[3:2], chosen_way_decode[2:2], chosen_way_decode[2:2], chosen_way_decode[2:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N20)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign select_snoop_data_n = (N17)? 1'b1 : 
                               (N21)? 1'b0 : 1'b0;
  assign recover_o = (N11)? 1'b0 : 
                     (N12)? 1'b0 : 
                     (N13)? 1'b0 : 
                     (N14)? 1'b0 : 
                     (N15)? 1'b0 : 
                     (N16)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N20)? 1'b1 : 
                     (N21)? 1'b0 : 
                     (N22)? 1'b0 : 1'b0;
  assign done_o = (N11)? 1'b0 : 
                  (N12)? 1'b0 : 
                  (N13)? 1'b0 : 
                  (N14)? 1'b0 : 
                  (N15)? 1'b0 : 
                  (N16)? 1'b0 : 
                  (N17)? 1'b0 : 
                  (N18)? 1'b0 : 
                  (N19)? 1'b0 : 
                  (N20)? 1'b0 : 
                  (N21)? 1'b1 : 
                  (N22)? 1'b0 : 1'b0;
  assign _0_net__3_ = N234 & N235;
  assign N234 = ~valid_v_i[3];
  assign N235 = ~lock_v_i[3];
  assign _0_net__2_ = N236 & N237;
  assign N236 = ~valid_v_i[2];
  assign N237 = ~lock_v_i[2];
  assign _0_net__1_ = N238 & N239;
  assign N238 = ~valid_v_i[1];
  assign N239 = ~lock_v_i[1];
  assign _0_net__0_ = N240 & N241;
  assign N240 = ~valid_v_i[0];
  assign N241 = ~lock_v_i[0];
  assign goto_flush_op = N243 | decode_v_i[9];
  assign N243 = N242 | decode_v_i[10];
  assign N242 = decode_v_i[13] | decode_v_i[8];
  assign goto_lock_op = decode_v_i[6] | N244;
  assign N244 = decode_v_i[7] & tag_hit_found_i;
  assign N23 = ~decode_v_i[17];
  assign N24 = N246 & mask_v_i[0];
  assign N246 = N245 & mask_v_i[1];
  assign N245 = mask_v_i[3] & mask_v_i[2];
  assign st_tag_miss_op = N247 & N248;
  assign N247 = decode_v_i[15] & full_word_op;
  assign N248 = ~tag_hit_found_i;
  assign N25 = ~goto_flush_op;
  assign N26 = ~decode_v_i[13];
  assign N27 = ~miss_state_r[3];
  assign N28 = ~miss_state_r[2];
  assign N29 = ~miss_state_r[1];
  assign N30 = ~miss_state_r[0];
  assign N37 = ~N36;
  assign N41 = ~N40;
  assign N45 = ~N44;
  assign N49 = ~N48;
  assign N53 = ~N52;
  assign N57 = ~N56;
  assign N61 = ~N60;
  assign N65 = ~N64;
  assign N69 = ~N68;
  assign N73 = ~N72;
  assign N77 = N75 | N76;
  assign dma_cmd_o[0] = N37;
  assign dma_cmd_o[1] = N49;
  assign dma_cmd_o[3] = N53;
  assign track_mem_data_o_3__3_ = N57;
  assign N78 = N249 & tbuf_empty_i;
  assign N249 = miss_v_i & sbuf_empty_i;
  assign N79 = ~N78;
  assign N80 = goto_lock_op | goto_flush_op;
  assign N81 = st_tag_miss_op | N80;
  assign N82 = ~N81;
  assign N89 = invalid_exist | track_miss_i;
  assign N90 = ~N89;
  assign N93 = ~N91;
  assign N94 = ~N92;
  assign N95 = N93 & N94;
  assign N96 = N93 & N92;
  assign N97 = N91 & N94;
  assign N98 = N91 & N92;
  assign N101 = N251 & N100;
  assign N251 = N250 & N99;
  assign N250 = ~track_miss_i;
  assign N107 = N252 & flush_way_decode[0];
  assign N252 = decode_v_i[8] | decode_v_i[9];
  assign N108 = N253 & flush_way_decode[0];
  assign N253 = decode_v_i[8] | decode_v_i[9];
  assign N109 = N254 & flush_way_decode[1];
  assign N254 = decode_v_i[8] | decode_v_i[9];
  assign N110 = N255 & flush_way_decode[1];
  assign N255 = decode_v_i[8] | decode_v_i[9];
  assign N111 = N256 & flush_way_decode[2];
  assign N256 = decode_v_i[8] | decode_v_i[9];
  assign N112 = N257 & flush_way_decode[2];
  assign N257 = decode_v_i[8] | decode_v_i[9];
  assign N113 = N258 & flush_way_decode[3];
  assign N258 = decode_v_i[8] | decode_v_i[9];
  assign N114 = N259 & flush_way_decode[3];
  assign N259 = decode_v_i[8] | decode_v_i[9];
  assign N115 = ~N105;
  assign N116 = ~N106;
  assign N117 = N115 & N116;
  assign N118 = N115 & N106;
  assign N119 = N105 & N116;
  assign N120 = N105 & N106;
  assign N123 = N261 & N122;
  assign N261 = N260 & N121;
  assign N260 = ~decode_v_i[8];
  assign N125 = ~dma_way_o[0];
  assign N126 = ~dma_way_o[1];
  assign N127 = N125 & N126;
  assign N128 = N125 & dma_way_o[1];
  assign N129 = dma_way_o[0] & N126;
  assign N130 = dma_way_o[0] & dma_way_o[1];
  assign N149 = ~dma_done_i;
  assign N150 = N125 & N126;
  assign N151 = N125 & dma_way_o[1];
  assign N152 = dma_way_o[0] & N126;
  assign N153 = dma_way_o[0] & dma_way_o[1];
  assign N172 = dma_done_i & st_tag_miss_op;
  assign N173 = dma_done_i & st_tag_miss_op;
  assign N174 = dma_done_i & st_tag_miss_op;
  assign N175 = N263 | st_tag_miss_op;
  assign N263 = N262 | decode_v_i[10];
  assign N262 = decode_v_i[13] | decode_v_i[9];
  assign N181 = decode_v_i[15] | decode_v_i[4];
  assign N186 = ~invalid_exist;
  assign N189 = ~N187;
  assign N190 = ~N188;
  assign N191 = N189 & N190;
  assign N192 = N189 & N188;
  assign N193 = N187 & N190;
  assign N194 = N187 & N188;
  assign N197 = N195 & N196;
  assign N199 = ~ack_i;
  assign N200 = ~track_mem_data_o_3__3_;
  assign N201 = N200;
  assign N202 = ~goto_flush_op;
  assign N203 = goto_lock_op & N202;
  assign N204 = ~goto_lock_op;
  assign N205 = N202 & N204;
  assign N206 = st_tag_miss_op & N205;
  assign N207 = ~track_miss_i;
  assign N208 = invalid_exist & N207;
  assign N209 = track_mem_v_o & N264;
  assign N264 = ~track_mem_w_o;
  assign N210 = N33 | dma_cmd_o[0];
  assign N211 = N210 | N45;
  assign N212 = N211 | dma_cmd_o[1];
  assign N213 = N212 | dma_cmd_o[3];
  assign N214 = N213 | track_mem_data_o_3__3_;
  assign N215 = N214 | N61;
  assign N216 = N215 | N65;
  assign N217 = N216 | N69;
  assign N218 = N217 | N73;
  assign N219 = N218 | N77;
  assign N220 = ~N219;
  assign N221 = N210 | N41;
  assign N222 = N221 | N45;
  assign N223 = N222 | dma_cmd_o[1];
  assign N224 = N223 | dma_cmd_o[3];
  assign N225 = N149 & track_mem_data_o_3__3_;
  assign N226 = N224 | N225;
  assign N227 = N226 | N61;
  assign N228 = N227 | N65;
  assign N229 = N228 | N69;
  assign N230 = N199 & N73;
  assign N231 = N229 | N230;
  assign N232 = N231 | N77;
  assign N233 = ~N232;

  always @(posedge clk_i) begin
    if(reset_i) begin
      track_data_we_o_sv2v_reg <= 1'b0;
      miss_state_r_3_sv2v_reg <= 1'b0;
      miss_state_r_2_sv2v_reg <= 1'b0;
      miss_state_r_1_sv2v_reg <= 1'b0;
      miss_state_r_0_sv2v_reg <= 1'b0;
      chosen_way_o_1_sv2v_reg <= 1'b0;
      chosen_way_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      track_data_we_o_sv2v_reg <= N209;
      miss_state_r_3_sv2v_reg <= miss_state_n[3];
      miss_state_r_2_sv2v_reg <= miss_state_n[2];
      miss_state_r_1_sv2v_reg <= miss_state_n[1];
      miss_state_r_0_sv2v_reg <= miss_state_n[0];
      chosen_way_o_1_sv2v_reg <= chosen_way_n[1];
      chosen_way_o_0_sv2v_reg <= chosen_way_n[0];
    end 
    if(reset_i) begin
      flush_way_r_1_sv2v_reg <= 1'b0;
      flush_way_r_0_sv2v_reg <= 1'b0;
    end else if(N220) begin
      flush_way_r_1_sv2v_reg <= N106;
      flush_way_r_0_sv2v_reg <= N105;
    end 
    if(reset_i) begin
      select_snoop_data_r_o_sv2v_reg <= 1'b0;
    end else if(N233) begin
      select_snoop_data_r_o_sv2v_reg <= select_snoop_data_n;
    end 
  end


endmodule



module bsg_counter_clear_up_4_0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [2:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [2:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N2,N3,N7,N30,N16;
  reg count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N16 = reset_i | clear_i;
  assign { N8, N6, N5 } = count_o + 1'b1;
  assign N9 = (N0)? 1'b1 : 
              (N7)? 1'b1 : 
              (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N11 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N10 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N15;
  assign N12 = ~reset_i;
  assign N13 = ~clear_i;
  assign N14 = N12 & N13;
  assign N15 = up_i & N14;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N13;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N16) begin
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N11) begin
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N9) begin
      count_o_0_sv2v_reg <= N10;
    end 
  end


endmodule



module bsg_circular_ptr_slots_p4_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1  = o + 1'b1;
  assign n_o = (N0)? \genblk1.genblk1.ptr_r_p1  : 
               (N1)? o : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p4
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p4_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p4_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;
  wire [127:0] \nz.mem ;
  reg \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,
  \nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,
  \nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N8)? \nz.mem [31] : 
                        (N10)? \nz.mem [63] : 
                        (N9)? \nz.mem [95] : 
                        (N11)? \nz.mem [127] : 1'b0;
  assign r_data_o[30] = (N8)? \nz.mem [30] : 
                        (N10)? \nz.mem [62] : 
                        (N9)? \nz.mem [94] : 
                        (N11)? \nz.mem [126] : 1'b0;
  assign r_data_o[29] = (N8)? \nz.mem [29] : 
                        (N10)? \nz.mem [61] : 
                        (N9)? \nz.mem [93] : 
                        (N11)? \nz.mem [125] : 1'b0;
  assign r_data_o[28] = (N8)? \nz.mem [28] : 
                        (N10)? \nz.mem [60] : 
                        (N9)? \nz.mem [92] : 
                        (N11)? \nz.mem [124] : 1'b0;
  assign r_data_o[27] = (N8)? \nz.mem [27] : 
                        (N10)? \nz.mem [59] : 
                        (N9)? \nz.mem [91] : 
                        (N11)? \nz.mem [123] : 1'b0;
  assign r_data_o[26] = (N8)? \nz.mem [26] : 
                        (N10)? \nz.mem [58] : 
                        (N9)? \nz.mem [90] : 
                        (N11)? \nz.mem [122] : 1'b0;
  assign r_data_o[25] = (N8)? \nz.mem [25] : 
                        (N10)? \nz.mem [57] : 
                        (N9)? \nz.mem [89] : 
                        (N11)? \nz.mem [121] : 1'b0;
  assign r_data_o[24] = (N8)? \nz.mem [24] : 
                        (N10)? \nz.mem [56] : 
                        (N9)? \nz.mem [88] : 
                        (N11)? \nz.mem [120] : 1'b0;
  assign r_data_o[23] = (N8)? \nz.mem [23] : 
                        (N10)? \nz.mem [55] : 
                        (N9)? \nz.mem [87] : 
                        (N11)? \nz.mem [119] : 1'b0;
  assign r_data_o[22] = (N8)? \nz.mem [22] : 
                        (N10)? \nz.mem [54] : 
                        (N9)? \nz.mem [86] : 
                        (N11)? \nz.mem [118] : 1'b0;
  assign r_data_o[21] = (N8)? \nz.mem [21] : 
                        (N10)? \nz.mem [53] : 
                        (N9)? \nz.mem [85] : 
                        (N11)? \nz.mem [117] : 1'b0;
  assign r_data_o[20] = (N8)? \nz.mem [20] : 
                        (N10)? \nz.mem [52] : 
                        (N9)? \nz.mem [84] : 
                        (N11)? \nz.mem [116] : 1'b0;
  assign r_data_o[19] = (N8)? \nz.mem [19] : 
                        (N10)? \nz.mem [51] : 
                        (N9)? \nz.mem [83] : 
                        (N11)? \nz.mem [115] : 1'b0;
  assign r_data_o[18] = (N8)? \nz.mem [18] : 
                        (N10)? \nz.mem [50] : 
                        (N9)? \nz.mem [82] : 
                        (N11)? \nz.mem [114] : 1'b0;
  assign r_data_o[17] = (N8)? \nz.mem [17] : 
                        (N10)? \nz.mem [49] : 
                        (N9)? \nz.mem [81] : 
                        (N11)? \nz.mem [113] : 1'b0;
  assign r_data_o[16] = (N8)? \nz.mem [16] : 
                        (N10)? \nz.mem [48] : 
                        (N9)? \nz.mem [80] : 
                        (N11)? \nz.mem [112] : 1'b0;
  assign r_data_o[15] = (N8)? \nz.mem [15] : 
                        (N10)? \nz.mem [47] : 
                        (N9)? \nz.mem [79] : 
                        (N11)? \nz.mem [111] : 1'b0;
  assign r_data_o[14] = (N8)? \nz.mem [14] : 
                        (N10)? \nz.mem [46] : 
                        (N9)? \nz.mem [78] : 
                        (N11)? \nz.mem [110] : 1'b0;
  assign r_data_o[13] = (N8)? \nz.mem [13] : 
                        (N10)? \nz.mem [45] : 
                        (N9)? \nz.mem [77] : 
                        (N11)? \nz.mem [109] : 1'b0;
  assign r_data_o[12] = (N8)? \nz.mem [12] : 
                        (N10)? \nz.mem [44] : 
                        (N9)? \nz.mem [76] : 
                        (N11)? \nz.mem [108] : 1'b0;
  assign r_data_o[11] = (N8)? \nz.mem [11] : 
                        (N10)? \nz.mem [43] : 
                        (N9)? \nz.mem [75] : 
                        (N11)? \nz.mem [107] : 1'b0;
  assign r_data_o[10] = (N8)? \nz.mem [10] : 
                        (N10)? \nz.mem [42] : 
                        (N9)? \nz.mem [74] : 
                        (N11)? \nz.mem [106] : 1'b0;
  assign r_data_o[9] = (N8)? \nz.mem [9] : 
                       (N10)? \nz.mem [41] : 
                       (N9)? \nz.mem [73] : 
                       (N11)? \nz.mem [105] : 1'b0;
  assign r_data_o[8] = (N8)? \nz.mem [8] : 
                       (N10)? \nz.mem [40] : 
                       (N9)? \nz.mem [72] : 
                       (N11)? \nz.mem [104] : 1'b0;
  assign r_data_o[7] = (N8)? \nz.mem [7] : 
                       (N10)? \nz.mem [39] : 
                       (N9)? \nz.mem [71] : 
                       (N11)? \nz.mem [103] : 1'b0;
  assign r_data_o[6] = (N8)? \nz.mem [6] : 
                       (N10)? \nz.mem [38] : 
                       (N9)? \nz.mem [70] : 
                       (N11)? \nz.mem [102] : 1'b0;
  assign r_data_o[5] = (N8)? \nz.mem [5] : 
                       (N10)? \nz.mem [37] : 
                       (N9)? \nz.mem [69] : 
                       (N11)? \nz.mem [101] : 1'b0;
  assign r_data_o[4] = (N8)? \nz.mem [4] : 
                       (N10)? \nz.mem [36] : 
                       (N9)? \nz.mem [68] : 
                       (N11)? \nz.mem [100] : 1'b0;
  assign r_data_o[3] = (N8)? \nz.mem [3] : 
                       (N10)? \nz.mem [35] : 
                       (N9)? \nz.mem [67] : 
                       (N11)? \nz.mem [99] : 1'b0;
  assign r_data_o[2] = (N8)? \nz.mem [2] : 
                       (N10)? \nz.mem [34] : 
                       (N9)? \nz.mem [66] : 
                       (N11)? \nz.mem [98] : 1'b0;
  assign r_data_o[1] = (N8)? \nz.mem [1] : 
                       (N10)? \nz.mem [33] : 
                       (N9)? \nz.mem [65] : 
                       (N11)? \nz.mem [97] : 1'b0;
  assign r_data_o[0] = (N8)? \nz.mem [0] : 
                       (N10)? \nz.mem [32] : 
                       (N9)? \nz.mem [64] : 
                       (N11)? \nz.mem [96] : 1'b0;
  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N20, N19, N18, N17 } = (N4)? { N16, N15, N14, N13 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N20) begin
      \nz.mem_127_sv2v_reg  <= w_data_i[31];
      \nz.mem_126_sv2v_reg  <= w_data_i[30];
      \nz.mem_125_sv2v_reg  <= w_data_i[29];
      \nz.mem_124_sv2v_reg  <= w_data_i[28];
      \nz.mem_123_sv2v_reg  <= w_data_i[27];
      \nz.mem_122_sv2v_reg  <= w_data_i[26];
      \nz.mem_121_sv2v_reg  <= w_data_i[25];
      \nz.mem_120_sv2v_reg  <= w_data_i[24];
      \nz.mem_119_sv2v_reg  <= w_data_i[23];
      \nz.mem_118_sv2v_reg  <= w_data_i[22];
      \nz.mem_117_sv2v_reg  <= w_data_i[21];
      \nz.mem_116_sv2v_reg  <= w_data_i[20];
      \nz.mem_115_sv2v_reg  <= w_data_i[19];
      \nz.mem_114_sv2v_reg  <= w_data_i[18];
      \nz.mem_113_sv2v_reg  <= w_data_i[17];
      \nz.mem_112_sv2v_reg  <= w_data_i[16];
      \nz.mem_111_sv2v_reg  <= w_data_i[15];
      \nz.mem_110_sv2v_reg  <= w_data_i[14];
      \nz.mem_109_sv2v_reg  <= w_data_i[13];
      \nz.mem_108_sv2v_reg  <= w_data_i[12];
      \nz.mem_107_sv2v_reg  <= w_data_i[11];
      \nz.mem_106_sv2v_reg  <= w_data_i[10];
      \nz.mem_105_sv2v_reg  <= w_data_i[9];
      \nz.mem_104_sv2v_reg  <= w_data_i[8];
      \nz.mem_103_sv2v_reg  <= w_data_i[7];
      \nz.mem_102_sv2v_reg  <= w_data_i[6];
      \nz.mem_101_sv2v_reg  <= w_data_i[5];
      \nz.mem_100_sv2v_reg  <= w_data_i[4];
      \nz.mem_99_sv2v_reg  <= w_data_i[3];
      \nz.mem_98_sv2v_reg  <= w_data_i[2];
      \nz.mem_97_sv2v_reg  <= w_data_i[1];
      \nz.mem_96_sv2v_reg  <= w_data_i[0];
    end 
    if(N19) begin
      \nz.mem_95_sv2v_reg  <= w_data_i[31];
      \nz.mem_94_sv2v_reg  <= w_data_i[30];
      \nz.mem_93_sv2v_reg  <= w_data_i[29];
      \nz.mem_92_sv2v_reg  <= w_data_i[28];
      \nz.mem_91_sv2v_reg  <= w_data_i[27];
      \nz.mem_90_sv2v_reg  <= w_data_i[26];
      \nz.mem_89_sv2v_reg  <= w_data_i[25];
      \nz.mem_88_sv2v_reg  <= w_data_i[24];
      \nz.mem_87_sv2v_reg  <= w_data_i[23];
      \nz.mem_86_sv2v_reg  <= w_data_i[22];
      \nz.mem_85_sv2v_reg  <= w_data_i[21];
      \nz.mem_84_sv2v_reg  <= w_data_i[20];
      \nz.mem_83_sv2v_reg  <= w_data_i[19];
      \nz.mem_82_sv2v_reg  <= w_data_i[18];
      \nz.mem_81_sv2v_reg  <= w_data_i[17];
      \nz.mem_80_sv2v_reg  <= w_data_i[16];
      \nz.mem_79_sv2v_reg  <= w_data_i[15];
      \nz.mem_78_sv2v_reg  <= w_data_i[14];
      \nz.mem_77_sv2v_reg  <= w_data_i[13];
      \nz.mem_76_sv2v_reg  <= w_data_i[12];
      \nz.mem_75_sv2v_reg  <= w_data_i[11];
      \nz.mem_74_sv2v_reg  <= w_data_i[10];
      \nz.mem_73_sv2v_reg  <= w_data_i[9];
      \nz.mem_72_sv2v_reg  <= w_data_i[8];
      \nz.mem_71_sv2v_reg  <= w_data_i[7];
      \nz.mem_70_sv2v_reg  <= w_data_i[6];
      \nz.mem_69_sv2v_reg  <= w_data_i[5];
      \nz.mem_68_sv2v_reg  <= w_data_i[4];
      \nz.mem_67_sv2v_reg  <= w_data_i[3];
      \nz.mem_66_sv2v_reg  <= w_data_i[2];
      \nz.mem_65_sv2v_reg  <= w_data_i[1];
      \nz.mem_64_sv2v_reg  <= w_data_i[0];
    end 
    if(N18) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N17) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p4
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p32_els_p4
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [63:0] \nz.mem ;
  reg \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [53] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [52] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [51] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [50] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [49] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [48] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [47] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [46] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [45] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [44] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [43] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [42] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [41] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [40] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [39] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [38] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [37] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [36] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [35] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [34] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [33] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_mux_width_p4_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [15:0] data_i;
  input [1:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[7] : 
                     (N3)? data_i[11] : 
                     (N5)? data_i[15] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[6] : 
                     (N3)? data_i[10] : 
                     (N5)? data_i[14] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[5] : 
                     (N3)? data_i[9] : 
                     (N5)? data_i[13] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[4] : 
                     (N3)? data_i[8] : 
                     (N5)? data_i[12] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p1_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [3:0] data_i;
  input [1:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[1] : 
                     (N3)? data_i[2] : 
                     (N5)? data_i[3] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p32_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [127:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[31] = (N2)? data_i[31] : 
                      (N4)? data_i[63] : 
                      (N3)? data_i[95] : 
                      (N5)? data_i[127] : 1'b0;
  assign data_o[30] = (N2)? data_i[30] : 
                      (N4)? data_i[62] : 
                      (N3)? data_i[94] : 
                      (N5)? data_i[126] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N4)? data_i[61] : 
                      (N3)? data_i[93] : 
                      (N5)? data_i[125] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N4)? data_i[60] : 
                      (N3)? data_i[92] : 
                      (N5)? data_i[124] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N4)? data_i[59] : 
                      (N3)? data_i[91] : 
                      (N5)? data_i[123] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N4)? data_i[58] : 
                      (N3)? data_i[90] : 
                      (N5)? data_i[122] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N4)? data_i[57] : 
                      (N3)? data_i[89] : 
                      (N5)? data_i[121] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N4)? data_i[56] : 
                      (N3)? data_i[88] : 
                      (N5)? data_i[120] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N4)? data_i[55] : 
                      (N3)? data_i[87] : 
                      (N5)? data_i[119] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N4)? data_i[54] : 
                      (N3)? data_i[86] : 
                      (N5)? data_i[118] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N4)? data_i[53] : 
                      (N3)? data_i[85] : 
                      (N5)? data_i[117] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N4)? data_i[52] : 
                      (N3)? data_i[84] : 
                      (N5)? data_i[116] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N4)? data_i[51] : 
                      (N3)? data_i[83] : 
                      (N5)? data_i[115] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N4)? data_i[50] : 
                      (N3)? data_i[82] : 
                      (N5)? data_i[114] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N4)? data_i[49] : 
                      (N3)? data_i[81] : 
                      (N5)? data_i[113] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N4)? data_i[48] : 
                      (N3)? data_i[80] : 
                      (N5)? data_i[112] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N4)? data_i[47] : 
                      (N3)? data_i[79] : 
                      (N5)? data_i[111] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N4)? data_i[46] : 
                      (N3)? data_i[78] : 
                      (N5)? data_i[110] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N4)? data_i[45] : 
                      (N3)? data_i[77] : 
                      (N5)? data_i[109] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N4)? data_i[44] : 
                      (N3)? data_i[76] : 
                      (N5)? data_i[108] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N4)? data_i[43] : 
                      (N3)? data_i[75] : 
                      (N5)? data_i[107] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N4)? data_i[42] : 
                      (N3)? data_i[74] : 
                      (N5)? data_i[106] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N4)? data_i[41] : 
                     (N3)? data_i[73] : 
                     (N5)? data_i[105] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N4)? data_i[40] : 
                     (N3)? data_i[72] : 
                     (N5)? data_i[104] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[39] : 
                     (N3)? data_i[71] : 
                     (N5)? data_i[103] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[38] : 
                     (N3)? data_i[70] : 
                     (N5)? data_i[102] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[37] : 
                     (N3)? data_i[69] : 
                     (N5)? data_i[101] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[36] : 
                     (N3)? data_i[68] : 
                     (N5)? data_i[100] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[35] : 
                     (N3)? data_i[67] : 
                     (N5)? data_i[99] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[34] : 
                     (N3)? data_i[66] : 
                     (N5)? data_i[98] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[33] : 
                     (N3)? data_i[65] : 
                     (N5)? data_i[97] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[32] : 
                     (N3)? data_i[64] : 
                     (N5)? data_i[96] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p32_els_p1
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4_word_tracking_p1_dma_data_width_p32_debug_p0
(
  clk_i,
  reset_i,
  dma_cmd_i,
  dma_way_i,
  dma_addr_i,
  done_o,
  track_data_we_i,
  snoop_word_o,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  data_mem_v_o,
  data_mem_w_o,
  data_mem_addr_o,
  data_mem_w_mask_o,
  data_mem_data_o,
  data_mem_data_i,
  track_miss_i,
  track_mem_data_i,
  dma_evict_o
);

  input [3:0] dma_cmd_i;
  input [1:0] dma_way_i;
  input [27:0] dma_addr_i;
  output [31:0] snoop_word_o;
  output [32:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  output [7:0] data_mem_addr_o;
  output [15:0] data_mem_w_mask_o;
  output [127:0] data_mem_data_o;
  input [127:0] data_mem_data_i;
  input [15:0] track_mem_data_i;
  input clk_i;
  input reset_i;
  input track_data_we_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  input track_miss_i;
  output done_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output data_mem_v_o;
  output data_mem_w_o;
  output dma_evict_o;
  wire [31:0] snoop_word_o,dma_data_o,out_fifo_data_li,snoop_word_n;
  wire [32:0] dma_pkt_o;
  wire [7:0] data_mem_addr_o;
  wire [15:0] data_mem_w_mask_o,dma_way_mask_expanded,track_mem_data_r;
  wire [127:0] data_mem_data_o;
  wire done_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,data_mem_v_o,data_mem_w_o,
  dma_evict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,dma_pkt_o_31_,dma_pkt_o_30_,
  dma_pkt_o_29_,dma_pkt_o_28_,dma_pkt_o_27_,dma_pkt_o_26_,dma_pkt_o_25_,dma_pkt_o_24_,
  dma_pkt_o_23_,dma_pkt_o_22_,dma_pkt_o_21_,dma_pkt_o_20_,dma_pkt_o_19_,
  dma_pkt_o_18_,dma_pkt_o_17_,dma_pkt_o_16_,dma_pkt_o_15_,dma_pkt_o_14_,data_mem_addr_o_7_,
  data_mem_addr_o_6_,data_mem_addr_o_5_,data_mem_addr_o_4_,data_mem_addr_o_3_,
  data_mem_addr_o_2_,data_mem_data_o_3__31_,data_mem_data_o_3__30_,data_mem_data_o_3__29_,
  data_mem_data_o_3__28_,data_mem_data_o_3__27_,data_mem_data_o_3__26_,
  data_mem_data_o_3__25_,data_mem_data_o_3__24_,data_mem_data_o_3__23_,
  data_mem_data_o_3__22_,data_mem_data_o_3__21_,data_mem_data_o_3__20_,data_mem_data_o_3__19_,
  data_mem_data_o_3__18_,data_mem_data_o_3__17_,data_mem_data_o_3__16_,
  data_mem_data_o_3__15_,data_mem_data_o_3__14_,data_mem_data_o_3__13_,data_mem_data_o_3__12_,
  data_mem_data_o_3__11_,data_mem_data_o_3__10_,data_mem_data_o_3__9_,
  data_mem_data_o_3__8_,data_mem_data_o_3__7_,data_mem_data_o_3__6_,data_mem_data_o_3__5_,
  data_mem_data_o_3__4_,data_mem_data_o_3__3_,data_mem_data_o_3__2_,data_mem_data_o_3__1_,
  data_mem_data_o_3__0_,counter_clear,counter_up,in_fifo_v_lo,in_fifo_yumi_li,
  out_fifo_v_li,out_fifo_ready_lo,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,
  N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  N66,N67,N68,N69,N70,N71,snoop_word_we,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89;
  wire [2:2] counter_r;
  wire [3:0] dma_way_mask,track_data_way_picked,track_bits_offset_picked_expanded,
  data_mem_w_mask_way_picked;
  wire [0:0] track_bits_offset_picked;
  wire [1:0] dma_state_r,dma_state_n;
  reg track_mem_data_r_15_sv2v_reg,track_mem_data_r_14_sv2v_reg,
  track_mem_data_r_13_sv2v_reg,track_mem_data_r_12_sv2v_reg,track_mem_data_r_11_sv2v_reg,
  track_mem_data_r_10_sv2v_reg,track_mem_data_r_9_sv2v_reg,track_mem_data_r_8_sv2v_reg,
  track_mem_data_r_7_sv2v_reg,track_mem_data_r_6_sv2v_reg,track_mem_data_r_5_sv2v_reg,
  track_mem_data_r_4_sv2v_reg,track_mem_data_r_3_sv2v_reg,track_mem_data_r_2_sv2v_reg,
  track_mem_data_r_1_sv2v_reg,track_mem_data_r_0_sv2v_reg,dma_state_r_1_sv2v_reg,
  dma_state_r_0_sv2v_reg,snoop_word_o_31_sv2v_reg,snoop_word_o_30_sv2v_reg,
  snoop_word_o_29_sv2v_reg,snoop_word_o_28_sv2v_reg,snoop_word_o_27_sv2v_reg,
  snoop_word_o_26_sv2v_reg,snoop_word_o_25_sv2v_reg,snoop_word_o_24_sv2v_reg,
  snoop_word_o_23_sv2v_reg,snoop_word_o_22_sv2v_reg,snoop_word_o_21_sv2v_reg,snoop_word_o_20_sv2v_reg,
  snoop_word_o_19_sv2v_reg,snoop_word_o_18_sv2v_reg,snoop_word_o_17_sv2v_reg,
  snoop_word_o_16_sv2v_reg,snoop_word_o_15_sv2v_reg,snoop_word_o_14_sv2v_reg,
  snoop_word_o_13_sv2v_reg,snoop_word_o_12_sv2v_reg,snoop_word_o_11_sv2v_reg,
  snoop_word_o_10_sv2v_reg,snoop_word_o_9_sv2v_reg,snoop_word_o_8_sv2v_reg,
  snoop_word_o_7_sv2v_reg,snoop_word_o_6_sv2v_reg,snoop_word_o_5_sv2v_reg,snoop_word_o_4_sv2v_reg,
  snoop_word_o_3_sv2v_reg,snoop_word_o_2_sv2v_reg,snoop_word_o_1_sv2v_reg,
  snoop_word_o_0_sv2v_reg;
  assign track_mem_data_r[15] = track_mem_data_r_15_sv2v_reg;
  assign track_mem_data_r[14] = track_mem_data_r_14_sv2v_reg;
  assign track_mem_data_r[13] = track_mem_data_r_13_sv2v_reg;
  assign track_mem_data_r[12] = track_mem_data_r_12_sv2v_reg;
  assign track_mem_data_r[11] = track_mem_data_r_11_sv2v_reg;
  assign track_mem_data_r[10] = track_mem_data_r_10_sv2v_reg;
  assign track_mem_data_r[9] = track_mem_data_r_9_sv2v_reg;
  assign track_mem_data_r[8] = track_mem_data_r_8_sv2v_reg;
  assign track_mem_data_r[7] = track_mem_data_r_7_sv2v_reg;
  assign track_mem_data_r[6] = track_mem_data_r_6_sv2v_reg;
  assign track_mem_data_r[5] = track_mem_data_r_5_sv2v_reg;
  assign track_mem_data_r[4] = track_mem_data_r_4_sv2v_reg;
  assign track_mem_data_r[3] = track_mem_data_r_3_sv2v_reg;
  assign track_mem_data_r[2] = track_mem_data_r_2_sv2v_reg;
  assign track_mem_data_r[1] = track_mem_data_r_1_sv2v_reg;
  assign track_mem_data_r[0] = track_mem_data_r_0_sv2v_reg;
  assign dma_state_r[1] = dma_state_r_1_sv2v_reg;
  assign dma_state_r[0] = dma_state_r_0_sv2v_reg;
  assign snoop_word_o[31] = snoop_word_o_31_sv2v_reg;
  assign snoop_word_o[30] = snoop_word_o_30_sv2v_reg;
  assign snoop_word_o[29] = snoop_word_o_29_sv2v_reg;
  assign snoop_word_o[28] = snoop_word_o_28_sv2v_reg;
  assign snoop_word_o[27] = snoop_word_o_27_sv2v_reg;
  assign snoop_word_o[26] = snoop_word_o_26_sv2v_reg;
  assign snoop_word_o[25] = snoop_word_o_25_sv2v_reg;
  assign snoop_word_o[24] = snoop_word_o_24_sv2v_reg;
  assign snoop_word_o[23] = snoop_word_o_23_sv2v_reg;
  assign snoop_word_o[22] = snoop_word_o_22_sv2v_reg;
  assign snoop_word_o[21] = snoop_word_o_21_sv2v_reg;
  assign snoop_word_o[20] = snoop_word_o_20_sv2v_reg;
  assign snoop_word_o[19] = snoop_word_o_19_sv2v_reg;
  assign snoop_word_o[18] = snoop_word_o_18_sv2v_reg;
  assign snoop_word_o[17] = snoop_word_o_17_sv2v_reg;
  assign snoop_word_o[16] = snoop_word_o_16_sv2v_reg;
  assign snoop_word_o[15] = snoop_word_o_15_sv2v_reg;
  assign snoop_word_o[14] = snoop_word_o_14_sv2v_reg;
  assign snoop_word_o[13] = snoop_word_o_13_sv2v_reg;
  assign snoop_word_o[12] = snoop_word_o_12_sv2v_reg;
  assign snoop_word_o[11] = snoop_word_o_11_sv2v_reg;
  assign snoop_word_o[10] = snoop_word_o_10_sv2v_reg;
  assign snoop_word_o[9] = snoop_word_o_9_sv2v_reg;
  assign snoop_word_o[8] = snoop_word_o_8_sv2v_reg;
  assign snoop_word_o[7] = snoop_word_o_7_sv2v_reg;
  assign snoop_word_o[6] = snoop_word_o_6_sv2v_reg;
  assign snoop_word_o[5] = snoop_word_o_5_sv2v_reg;
  assign snoop_word_o[4] = snoop_word_o_4_sv2v_reg;
  assign snoop_word_o[3] = snoop_word_o_3_sv2v_reg;
  assign snoop_word_o[2] = snoop_word_o_2_sv2v_reg;
  assign snoop_word_o[1] = snoop_word_o_1_sv2v_reg;
  assign snoop_word_o[0] = snoop_word_o_0_sv2v_reg;
  assign dma_pkt_o[4] = 1'b0;
  assign dma_pkt_o[5] = 1'b0;
  assign dma_pkt_o[6] = 1'b0;
  assign dma_pkt_o[7] = 1'b0;
  assign dma_pkt_o_31_ = dma_addr_i[27];
  assign dma_pkt_o[31] = dma_pkt_o_31_;
  assign dma_pkt_o_30_ = dma_addr_i[26];
  assign dma_pkt_o[30] = dma_pkt_o_30_;
  assign dma_pkt_o_29_ = dma_addr_i[25];
  assign dma_pkt_o[29] = dma_pkt_o_29_;
  assign dma_pkt_o_28_ = dma_addr_i[24];
  assign dma_pkt_o[28] = dma_pkt_o_28_;
  assign dma_pkt_o_27_ = dma_addr_i[23];
  assign dma_pkt_o[27] = dma_pkt_o_27_;
  assign dma_pkt_o_26_ = dma_addr_i[22];
  assign dma_pkt_o[26] = dma_pkt_o_26_;
  assign dma_pkt_o_25_ = dma_addr_i[21];
  assign dma_pkt_o[25] = dma_pkt_o_25_;
  assign dma_pkt_o_24_ = dma_addr_i[20];
  assign dma_pkt_o[24] = dma_pkt_o_24_;
  assign dma_pkt_o_23_ = dma_addr_i[19];
  assign dma_pkt_o[23] = dma_pkt_o_23_;
  assign dma_pkt_o_22_ = dma_addr_i[18];
  assign dma_pkt_o[22] = dma_pkt_o_22_;
  assign dma_pkt_o_21_ = dma_addr_i[17];
  assign dma_pkt_o[21] = dma_pkt_o_21_;
  assign dma_pkt_o_20_ = dma_addr_i[16];
  assign dma_pkt_o[20] = dma_pkt_o_20_;
  assign dma_pkt_o_19_ = dma_addr_i[15];
  assign dma_pkt_o[19] = dma_pkt_o_19_;
  assign dma_pkt_o_18_ = dma_addr_i[14];
  assign dma_pkt_o[18] = dma_pkt_o_18_;
  assign dma_pkt_o_17_ = dma_addr_i[13];
  assign dma_pkt_o[17] = dma_pkt_o_17_;
  assign dma_pkt_o_16_ = dma_addr_i[12];
  assign dma_pkt_o[16] = dma_pkt_o_16_;
  assign dma_pkt_o_15_ = dma_addr_i[11];
  assign dma_pkt_o[15] = dma_pkt_o_15_;
  assign dma_pkt_o_14_ = dma_addr_i[10];
  assign dma_pkt_o[14] = dma_pkt_o_14_;
  assign data_mem_addr_o_7_ = dma_addr_i[9];
  assign dma_pkt_o[13] = data_mem_addr_o_7_;
  assign data_mem_addr_o[7] = data_mem_addr_o_7_;
  assign data_mem_addr_o_6_ = dma_addr_i[8];
  assign dma_pkt_o[12] = data_mem_addr_o_6_;
  assign data_mem_addr_o[6] = data_mem_addr_o_6_;
  assign data_mem_addr_o_5_ = dma_addr_i[7];
  assign dma_pkt_o[11] = data_mem_addr_o_5_;
  assign data_mem_addr_o[5] = data_mem_addr_o_5_;
  assign data_mem_addr_o_4_ = dma_addr_i[6];
  assign dma_pkt_o[10] = data_mem_addr_o_4_;
  assign data_mem_addr_o[4] = data_mem_addr_o_4_;
  assign data_mem_addr_o_3_ = dma_addr_i[5];
  assign dma_pkt_o[9] = data_mem_addr_o_3_;
  assign data_mem_addr_o[3] = data_mem_addr_o_3_;
  assign data_mem_addr_o_2_ = dma_addr_i[4];
  assign dma_pkt_o[8] = data_mem_addr_o_2_;
  assign data_mem_addr_o[2] = data_mem_addr_o_2_;
  assign data_mem_data_o[31] = data_mem_data_o_3__31_;
  assign data_mem_data_o[63] = data_mem_data_o_3__31_;
  assign data_mem_data_o[95] = data_mem_data_o_3__31_;
  assign data_mem_data_o[127] = data_mem_data_o_3__31_;
  assign data_mem_data_o[30] = data_mem_data_o_3__30_;
  assign data_mem_data_o[62] = data_mem_data_o_3__30_;
  assign data_mem_data_o[94] = data_mem_data_o_3__30_;
  assign data_mem_data_o[126] = data_mem_data_o_3__30_;
  assign data_mem_data_o[29] = data_mem_data_o_3__29_;
  assign data_mem_data_o[61] = data_mem_data_o_3__29_;
  assign data_mem_data_o[93] = data_mem_data_o_3__29_;
  assign data_mem_data_o[125] = data_mem_data_o_3__29_;
  assign data_mem_data_o[28] = data_mem_data_o_3__28_;
  assign data_mem_data_o[60] = data_mem_data_o_3__28_;
  assign data_mem_data_o[92] = data_mem_data_o_3__28_;
  assign data_mem_data_o[124] = data_mem_data_o_3__28_;
  assign data_mem_data_o[27] = data_mem_data_o_3__27_;
  assign data_mem_data_o[59] = data_mem_data_o_3__27_;
  assign data_mem_data_o[91] = data_mem_data_o_3__27_;
  assign data_mem_data_o[123] = data_mem_data_o_3__27_;
  assign data_mem_data_o[26] = data_mem_data_o_3__26_;
  assign data_mem_data_o[58] = data_mem_data_o_3__26_;
  assign data_mem_data_o[90] = data_mem_data_o_3__26_;
  assign data_mem_data_o[122] = data_mem_data_o_3__26_;
  assign data_mem_data_o[25] = data_mem_data_o_3__25_;
  assign data_mem_data_o[57] = data_mem_data_o_3__25_;
  assign data_mem_data_o[89] = data_mem_data_o_3__25_;
  assign data_mem_data_o[121] = data_mem_data_o_3__25_;
  assign data_mem_data_o[24] = data_mem_data_o_3__24_;
  assign data_mem_data_o[56] = data_mem_data_o_3__24_;
  assign data_mem_data_o[88] = data_mem_data_o_3__24_;
  assign data_mem_data_o[120] = data_mem_data_o_3__24_;
  assign data_mem_data_o[23] = data_mem_data_o_3__23_;
  assign data_mem_data_o[55] = data_mem_data_o_3__23_;
  assign data_mem_data_o[87] = data_mem_data_o_3__23_;
  assign data_mem_data_o[119] = data_mem_data_o_3__23_;
  assign data_mem_data_o[22] = data_mem_data_o_3__22_;
  assign data_mem_data_o[54] = data_mem_data_o_3__22_;
  assign data_mem_data_o[86] = data_mem_data_o_3__22_;
  assign data_mem_data_o[118] = data_mem_data_o_3__22_;
  assign data_mem_data_o[21] = data_mem_data_o_3__21_;
  assign data_mem_data_o[53] = data_mem_data_o_3__21_;
  assign data_mem_data_o[85] = data_mem_data_o_3__21_;
  assign data_mem_data_o[117] = data_mem_data_o_3__21_;
  assign data_mem_data_o[20] = data_mem_data_o_3__20_;
  assign data_mem_data_o[52] = data_mem_data_o_3__20_;
  assign data_mem_data_o[84] = data_mem_data_o_3__20_;
  assign data_mem_data_o[116] = data_mem_data_o_3__20_;
  assign data_mem_data_o[19] = data_mem_data_o_3__19_;
  assign data_mem_data_o[51] = data_mem_data_o_3__19_;
  assign data_mem_data_o[83] = data_mem_data_o_3__19_;
  assign data_mem_data_o[115] = data_mem_data_o_3__19_;
  assign data_mem_data_o[18] = data_mem_data_o_3__18_;
  assign data_mem_data_o[50] = data_mem_data_o_3__18_;
  assign data_mem_data_o[82] = data_mem_data_o_3__18_;
  assign data_mem_data_o[114] = data_mem_data_o_3__18_;
  assign data_mem_data_o[17] = data_mem_data_o_3__17_;
  assign data_mem_data_o[49] = data_mem_data_o_3__17_;
  assign data_mem_data_o[81] = data_mem_data_o_3__17_;
  assign data_mem_data_o[113] = data_mem_data_o_3__17_;
  assign data_mem_data_o[16] = data_mem_data_o_3__16_;
  assign data_mem_data_o[48] = data_mem_data_o_3__16_;
  assign data_mem_data_o[80] = data_mem_data_o_3__16_;
  assign data_mem_data_o[112] = data_mem_data_o_3__16_;
  assign data_mem_data_o[15] = data_mem_data_o_3__15_;
  assign data_mem_data_o[47] = data_mem_data_o_3__15_;
  assign data_mem_data_o[79] = data_mem_data_o_3__15_;
  assign data_mem_data_o[111] = data_mem_data_o_3__15_;
  assign data_mem_data_o[14] = data_mem_data_o_3__14_;
  assign data_mem_data_o[46] = data_mem_data_o_3__14_;
  assign data_mem_data_o[78] = data_mem_data_o_3__14_;
  assign data_mem_data_o[110] = data_mem_data_o_3__14_;
  assign data_mem_data_o[13] = data_mem_data_o_3__13_;
  assign data_mem_data_o[45] = data_mem_data_o_3__13_;
  assign data_mem_data_o[77] = data_mem_data_o_3__13_;
  assign data_mem_data_o[109] = data_mem_data_o_3__13_;
  assign data_mem_data_o[12] = data_mem_data_o_3__12_;
  assign data_mem_data_o[44] = data_mem_data_o_3__12_;
  assign data_mem_data_o[76] = data_mem_data_o_3__12_;
  assign data_mem_data_o[108] = data_mem_data_o_3__12_;
  assign data_mem_data_o[11] = data_mem_data_o_3__11_;
  assign data_mem_data_o[43] = data_mem_data_o_3__11_;
  assign data_mem_data_o[75] = data_mem_data_o_3__11_;
  assign data_mem_data_o[107] = data_mem_data_o_3__11_;
  assign data_mem_data_o[10] = data_mem_data_o_3__10_;
  assign data_mem_data_o[42] = data_mem_data_o_3__10_;
  assign data_mem_data_o[74] = data_mem_data_o_3__10_;
  assign data_mem_data_o[106] = data_mem_data_o_3__10_;
  assign data_mem_data_o[9] = data_mem_data_o_3__9_;
  assign data_mem_data_o[41] = data_mem_data_o_3__9_;
  assign data_mem_data_o[73] = data_mem_data_o_3__9_;
  assign data_mem_data_o[105] = data_mem_data_o_3__9_;
  assign data_mem_data_o[8] = data_mem_data_o_3__8_;
  assign data_mem_data_o[40] = data_mem_data_o_3__8_;
  assign data_mem_data_o[72] = data_mem_data_o_3__8_;
  assign data_mem_data_o[104] = data_mem_data_o_3__8_;
  assign data_mem_data_o[7] = data_mem_data_o_3__7_;
  assign data_mem_data_o[39] = data_mem_data_o_3__7_;
  assign data_mem_data_o[71] = data_mem_data_o_3__7_;
  assign data_mem_data_o[103] = data_mem_data_o_3__7_;
  assign data_mem_data_o[6] = data_mem_data_o_3__6_;
  assign data_mem_data_o[38] = data_mem_data_o_3__6_;
  assign data_mem_data_o[70] = data_mem_data_o_3__6_;
  assign data_mem_data_o[102] = data_mem_data_o_3__6_;
  assign data_mem_data_o[5] = data_mem_data_o_3__5_;
  assign data_mem_data_o[37] = data_mem_data_o_3__5_;
  assign data_mem_data_o[69] = data_mem_data_o_3__5_;
  assign data_mem_data_o[101] = data_mem_data_o_3__5_;
  assign data_mem_data_o[4] = data_mem_data_o_3__4_;
  assign data_mem_data_o[36] = data_mem_data_o_3__4_;
  assign data_mem_data_o[68] = data_mem_data_o_3__4_;
  assign data_mem_data_o[100] = data_mem_data_o_3__4_;
  assign data_mem_data_o[3] = data_mem_data_o_3__3_;
  assign data_mem_data_o[35] = data_mem_data_o_3__3_;
  assign data_mem_data_o[67] = data_mem_data_o_3__3_;
  assign data_mem_data_o[99] = data_mem_data_o_3__3_;
  assign data_mem_data_o[2] = data_mem_data_o_3__2_;
  assign data_mem_data_o[34] = data_mem_data_o_3__2_;
  assign data_mem_data_o[66] = data_mem_data_o_3__2_;
  assign data_mem_data_o[98] = data_mem_data_o_3__2_;
  assign data_mem_data_o[1] = data_mem_data_o_3__1_;
  assign data_mem_data_o[33] = data_mem_data_o_3__1_;
  assign data_mem_data_o[65] = data_mem_data_o_3__1_;
  assign data_mem_data_o[97] = data_mem_data_o_3__1_;
  assign data_mem_data_o[0] = data_mem_data_o_3__0_;
  assign data_mem_data_o[32] = data_mem_data_o_3__0_;
  assign data_mem_data_o[64] = data_mem_data_o_3__0_;
  assign data_mem_data_o[96] = data_mem_data_o_3__0_;

  bsg_counter_clear_up_4_0
  dma_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(counter_clear),
    .up_i(counter_up),
    .count_o({ counter_r[2:2], data_mem_addr_o[1:0] })
  );


  bsg_fifo_1r1w_small_width_p32_els_p4
  in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(dma_data_v_i),
    .ready_o(dma_data_ready_o),
    .data_i(dma_data_i),
    .v_o(in_fifo_v_lo),
    .data_o({ data_mem_data_o_3__31_, data_mem_data_o_3__30_, data_mem_data_o_3__29_, data_mem_data_o_3__28_, data_mem_data_o_3__27_, data_mem_data_o_3__26_, data_mem_data_o_3__25_, data_mem_data_o_3__24_, data_mem_data_o_3__23_, data_mem_data_o_3__22_, data_mem_data_o_3__21_, data_mem_data_o_3__20_, data_mem_data_o_3__19_, data_mem_data_o_3__18_, data_mem_data_o_3__17_, data_mem_data_o_3__16_, data_mem_data_o_3__15_, data_mem_data_o_3__14_, data_mem_data_o_3__13_, data_mem_data_o_3__12_, data_mem_data_o_3__11_, data_mem_data_o_3__10_, data_mem_data_o_3__9_, data_mem_data_o_3__8_, data_mem_data_o_3__7_, data_mem_data_o_3__6_, data_mem_data_o_3__5_, data_mem_data_o_3__4_, data_mem_data_o_3__3_, data_mem_data_o_3__2_, data_mem_data_o_3__1_, data_mem_data_o_3__0_ }),
    .yumi_i(in_fifo_yumi_li)
  );


  bsg_two_fifo_width_p32
  out_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(out_fifo_ready_lo),
    .data_i(out_fifo_data_li),
    .v_i(out_fifo_v_li),
    .v_o(dma_data_v_o),
    .data_o(dma_data_o),
    .yumi_i(dma_data_yumi_i)
  );


  bsg_decode_num_out_p4
  dma_way_demux
  (
    .i(dma_way_i),
    .o(dma_way_mask)
  );


  bsg_expand_bitmask
  expand0
  (
    .i(dma_way_mask),
    .o(dma_way_mask_expanded)
  );


  bsg_mux_width_p4_els_p4
  track_way_mux
  (
    .data_i(track_mem_data_r),
    .sel_i(dma_way_i),
    .data_o(track_data_way_picked)
  );


  bsg_mux_width_p1_els_p4
  track_offset_mux
  (
    .data_i(track_data_way_picked),
    .sel_i(data_mem_addr_o[1:0]),
    .data_o(track_bits_offset_picked[0])
  );


  bsg_expand_bitmask
  expand1
  (
    .i(track_bits_offset_picked[0]),
    .o(track_bits_offset_picked_expanded)
  );


  bsg_mux_width_p32_els_p4
  write_data_mux
  (
    .data_i(data_mem_data_i),
    .sel_i(dma_way_i),
    .data_o(out_fifo_data_li)
  );

  assign N18 = N17 & N85;
  assign N19 = dma_state_r[1] | N85;
  assign N21 = N17 | dma_state_r[0];
  assign N23 = dma_state_r[1] & dma_state_r[0];
  assign N24 = dma_cmd_i[1] | N41;
  assign N25 = N27 | N24;
  assign N27 = dma_cmd_i[3] | dma_cmd_i[2];
  assign N28 = N40 | dma_cmd_i[0];
  assign N29 = N27 | N28;
  assign N31 = dma_cmd_i[3] | N39;
  assign N32 = N31 | N35;
  assign N34 = N38 | dma_cmd_i[2];
  assign N35 = dma_cmd_i[1] | dma_cmd_i[0];
  assign N36 = N34 | N35;
  assign N42 = N38 & N39;
  assign N43 = N40 & N41;
  assign N44 = N42 & N43;
  assign N71 = data_mem_addr_o[1:0] == dma_addr_i[3:2];

  bsg_mux_width_p32_els_p1
  snoop_mux0
  (
    .data_i({ data_mem_data_o_3__31_, data_mem_data_o_3__30_, data_mem_data_o_3__29_, data_mem_data_o_3__28_, data_mem_data_o_3__27_, data_mem_data_o_3__26_, data_mem_data_o_3__25_, data_mem_data_o_3__24_, data_mem_data_o_3__23_, data_mem_data_o_3__22_, data_mem_data_o_3__21_, data_mem_data_o_3__20_, data_mem_data_o_3__19_, data_mem_data_o_3__18_, data_mem_data_o_3__17_, data_mem_data_o_3__16_, data_mem_data_o_3__15_, data_mem_data_o_3__14_, data_mem_data_o_3__13_, data_mem_data_o_3__12_, data_mem_data_o_3__11_, data_mem_data_o_3__10_, data_mem_data_o_3__9_, data_mem_data_o_3__8_, data_mem_data_o_3__7_, data_mem_data_o_3__6_, data_mem_data_o_3__5_, data_mem_data_o_3__4_, data_mem_data_o_3__3_, data_mem_data_o_3__2_, data_mem_data_o_3__1_, data_mem_data_o_3__0_ }),
    .sel_i(dma_addr_i[2]),
    .data_o(snoop_word_n)
  );

  assign N76 = ~counter_r[2];
  assign N77 = data_mem_addr_o[1] | N76;
  assign N78 = data_mem_addr_o[0] | N77;
  assign N79 = ~N78;
  assign N80 = ~data_mem_addr_o[1];
  assign N81 = ~data_mem_addr_o[0];
  assign N82 = N80 | counter_r[2];
  assign N83 = N81 | N82;
  assign N84 = ~N83;
  assign N85 = ~dma_state_r[0];
  assign N86 = N85 | dma_state_r[1];
  assign N87 = ~N86;
  assign data_mem_w_mask_way_picked = (N0)? { N13, N14, N15, N16 } : 
                                      (N12)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N0 = track_miss_i;
  assign N50 = (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N1 = N26;
  assign N2 = N30;
  assign N3 = N33;
  assign N4 = N37;
  assign N5 = N44;
  assign { N55, N54, N53, N52, N51 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N2)? { 1'b1, track_data_way_picked } : 
                                       (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N49)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = (N1)? dma_pkt_yumi_i : 
               (N2)? dma_pkt_yumi_i : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N57 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b1 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N58 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N59 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? track_bits_offset_picked[0] : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N61 = ~N60;
  assign N66 = ~N65;
  assign counter_clear = (N6)? N57 : 
                         (N7)? N63 : 
                         (N8)? N68 : 
                         (N9)? 1'b0 : 1'b0;
  assign N6 = N18;
  assign N7 = N20;
  assign N8 = N22;
  assign N9 = N23;
  assign counter_up = (N6)? N58 : 
                      (N7)? N62 : 
                      (N8)? N67 : 
                      (N9)? 1'b0 : 1'b0;
  assign data_mem_v_o = (N6)? N59 : 
                        (N7)? in_fifo_v_lo : 
                        (N8)? N69 : 
                        (N9)? 1'b0 : 1'b0;
  assign dma_pkt_v_o = (N6)? N50 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b0 : 
                       (N9)? 1'b0 : 1'b0;
  assign { dma_pkt_o[32:32], dma_pkt_o[3:0] } = (N6)? { N55, N54, N53, N52, N51 } : 
                                                (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign done_o = (N6)? N56 : 
                  (N7)? N64 : 
                  (N8)? N70 : 
                  (N9)? 1'b0 : 1'b0;
  assign dma_state_n = (N6)? { N37, N33 } : 
                       (N7)? { 1'b0, N61 } : 
                       (N8)? { N66, 1'b0 } : 
                       (N9)? { 1'b0, 1'b0 } : 1'b0;
  assign data_mem_w_o = (N6)? 1'b0 : 
                        (N7)? in_fifo_v_lo : 
                        (N8)? 1'b0 : 
                        (N9)? 1'b0 : 1'b0;
  assign in_fifo_yumi_li = (N6)? 1'b0 : 
                           (N7)? in_fifo_v_lo : 
                           (N8)? 1'b0 : 
                           (N9)? 1'b0 : 1'b0;
  assign out_fifo_v_li = (N6)? 1'b0 : 
                         (N7)? 1'b0 : 
                         (N8)? 1'b1 : 
                         (N9)? 1'b0 : 1'b0;
  assign dma_evict_o = (N6)? 1'b0 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b1 : 
                       (N9)? 1'b0 : 1'b0;
  assign N74 = (N10)? 1'b0 : 
               (N11)? snoop_word_we : 1'b0;
  assign N10 = N73;
  assign N11 = N72;
  assign N75 = (N10)? 1'b0 : 
               (N11)? track_data_we_i : 1'b0;
  assign N12 = ~track_miss_i;
  assign N13 = ~track_bits_offset_picked_expanded[3];
  assign N14 = ~track_bits_offset_picked_expanded[2];
  assign N15 = ~track_bits_offset_picked_expanded[1];
  assign N16 = ~track_bits_offset_picked_expanded[0];
  assign data_mem_w_mask_o[15] = dma_way_mask_expanded[15] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[14] = dma_way_mask_expanded[14] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[13] = dma_way_mask_expanded[13] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[12] = dma_way_mask_expanded[12] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[11] = dma_way_mask_expanded[11] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[10] = dma_way_mask_expanded[10] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[9] = dma_way_mask_expanded[9] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[8] = dma_way_mask_expanded[8] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[7] = dma_way_mask_expanded[7] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[6] = dma_way_mask_expanded[6] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[5] = dma_way_mask_expanded[5] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[4] = dma_way_mask_expanded[4] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[3] = dma_way_mask_expanded[3] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[2] = dma_way_mask_expanded[2] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[1] = dma_way_mask_expanded[1] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[0] = dma_way_mask_expanded[0] & data_mem_w_mask_way_picked[0];
  assign N17 = ~dma_state_r[1];
  assign N20 = ~N19;
  assign N22 = ~N21;
  assign N26 = ~N25;
  assign N30 = ~N29;
  assign N33 = ~N32;
  assign N37 = ~N36;
  assign N38 = ~dma_cmd_i[3];
  assign N39 = ~dma_cmd_i[2];
  assign N40 = ~dma_cmd_i[1];
  assign N41 = ~dma_cmd_i[0];
  assign N45 = N30 | N26;
  assign N46 = N33 | N45;
  assign N47 = N37 | N46;
  assign N48 = N44 | N47;
  assign N49 = ~N48;
  assign N60 = N84 & in_fifo_v_lo;
  assign N62 = in_fifo_v_lo & N83;
  assign N63 = in_fifo_v_lo & N84;
  assign N64 = N84 & in_fifo_v_lo;
  assign N65 = N79 & out_fifo_ready_lo;
  assign N67 = out_fifo_ready_lo & N78;
  assign N68 = out_fifo_ready_lo & N79;
  assign N69 = N88 & track_bits_offset_picked[0];
  assign N88 = out_fifo_ready_lo & N78;
  assign N70 = N79 & out_fifo_ready_lo;
  assign snoop_word_we = N89 & N71;
  assign N89 = N87 & in_fifo_v_lo;
  assign N72 = ~reset_i;
  assign N73 = reset_i;

  always @(posedge clk_i) begin
    if(N75) begin
      track_mem_data_r_15_sv2v_reg <= track_mem_data_i[15];
      track_mem_data_r_14_sv2v_reg <= track_mem_data_i[14];
      track_mem_data_r_13_sv2v_reg <= track_mem_data_i[13];
      track_mem_data_r_12_sv2v_reg <= track_mem_data_i[12];
      track_mem_data_r_11_sv2v_reg <= track_mem_data_i[11];
      track_mem_data_r_10_sv2v_reg <= track_mem_data_i[10];
      track_mem_data_r_9_sv2v_reg <= track_mem_data_i[9];
      track_mem_data_r_8_sv2v_reg <= track_mem_data_i[8];
      track_mem_data_r_7_sv2v_reg <= track_mem_data_i[7];
      track_mem_data_r_6_sv2v_reg <= track_mem_data_i[6];
      track_mem_data_r_5_sv2v_reg <= track_mem_data_i[5];
      track_mem_data_r_4_sv2v_reg <= track_mem_data_i[4];
      track_mem_data_r_3_sv2v_reg <= track_mem_data_i[3];
      track_mem_data_r_2_sv2v_reg <= track_mem_data_i[2];
      track_mem_data_r_1_sv2v_reg <= track_mem_data_i[1];
      track_mem_data_r_0_sv2v_reg <= track_mem_data_i[0];
    end 
    if(reset_i) begin
      dma_state_r_1_sv2v_reg <= 1'b0;
      dma_state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      dma_state_r_1_sv2v_reg <= dma_state_n[1];
      dma_state_r_0_sv2v_reg <= dma_state_n[0];
    end 
    if(N74) begin
      snoop_word_o_31_sv2v_reg <= snoop_word_n[31];
      snoop_word_o_30_sv2v_reg <= snoop_word_n[30];
      snoop_word_o_29_sv2v_reg <= snoop_word_n[29];
      snoop_word_o_28_sv2v_reg <= snoop_word_n[28];
      snoop_word_o_27_sv2v_reg <= snoop_word_n[27];
      snoop_word_o_26_sv2v_reg <= snoop_word_n[26];
      snoop_word_o_25_sv2v_reg <= snoop_word_n[25];
      snoop_word_o_24_sv2v_reg <= snoop_word_n[24];
      snoop_word_o_23_sv2v_reg <= snoop_word_n[23];
      snoop_word_o_22_sv2v_reg <= snoop_word_n[22];
      snoop_word_o_21_sv2v_reg <= snoop_word_n[21];
      snoop_word_o_20_sv2v_reg <= snoop_word_n[20];
      snoop_word_o_19_sv2v_reg <= snoop_word_n[19];
      snoop_word_o_18_sv2v_reg <= snoop_word_n[18];
      snoop_word_o_17_sv2v_reg <= snoop_word_n[17];
      snoop_word_o_16_sv2v_reg <= snoop_word_n[16];
      snoop_word_o_15_sv2v_reg <= snoop_word_n[15];
      snoop_word_o_14_sv2v_reg <= snoop_word_n[14];
      snoop_word_o_13_sv2v_reg <= snoop_word_n[13];
      snoop_word_o_12_sv2v_reg <= snoop_word_n[12];
      snoop_word_o_11_sv2v_reg <= snoop_word_n[11];
      snoop_word_o_10_sv2v_reg <= snoop_word_n[10];
      snoop_word_o_9_sv2v_reg <= snoop_word_n[9];
      snoop_word_o_8_sv2v_reg <= snoop_word_n[8];
      snoop_word_o_7_sv2v_reg <= snoop_word_n[7];
      snoop_word_o_6_sv2v_reg <= snoop_word_n[6];
      snoop_word_o_5_sv2v_reg <= snoop_word_n[5];
      snoop_word_o_4_sv2v_reg <= snoop_word_n[4];
      snoop_word_o_3_sv2v_reg <= snoop_word_n[3];
      snoop_word_o_2_sv2v_reg <= snoop_word_n[2];
      snoop_word_o_1_sv2v_reg <= snoop_word_n[1];
      snoop_word_o_0_sv2v_reg <= snoop_word_n[0];
    end 
  end


endmodule



module bsg_cache_buffer_queue_width_p66
(
  clk_i,
  reset_i,
  v_i,
  data_i,
  v_o,
  data_o,
  yumi_i,
  el0_valid_o,
  el1_valid_o,
  el0_snoop_o,
  el1_snoop_o,
  empty_o,
  full_o
);

  input [65:0] data_i;
  output [65:0] data_o;
  output [65:0] el0_snoop_o;
  output [65:0] el1_snoop_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output v_o;
  output el0_valid_o;
  output el1_valid_o;
  output empty_o;
  output full_o;
  wire [65:0] data_o,el0_snoop_o,el1_snoop_o;
  wire v_o,el0_valid_o,el1_valid_o,empty_o,full_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,el0_enable,el1_enable,mux0_sel,mux1_sel,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92;
  wire [1:0] num_els_r;
  reg num_els_r_1_sv2v_reg,num_els_r_0_sv2v_reg,el0_snoop_o_65_sv2v_reg,
  el0_snoop_o_64_sv2v_reg,el0_snoop_o_63_sv2v_reg,el0_snoop_o_62_sv2v_reg,
  el0_snoop_o_61_sv2v_reg,el0_snoop_o_60_sv2v_reg,el0_snoop_o_59_sv2v_reg,el0_snoop_o_58_sv2v_reg,
  el0_snoop_o_57_sv2v_reg,el0_snoop_o_56_sv2v_reg,el0_snoop_o_55_sv2v_reg,
  el0_snoop_o_54_sv2v_reg,el0_snoop_o_53_sv2v_reg,el0_snoop_o_52_sv2v_reg,
  el0_snoop_o_51_sv2v_reg,el0_snoop_o_50_sv2v_reg,el0_snoop_o_49_sv2v_reg,el0_snoop_o_48_sv2v_reg,
  el0_snoop_o_47_sv2v_reg,el0_snoop_o_46_sv2v_reg,el0_snoop_o_45_sv2v_reg,
  el0_snoop_o_44_sv2v_reg,el0_snoop_o_43_sv2v_reg,el0_snoop_o_42_sv2v_reg,
  el0_snoop_o_41_sv2v_reg,el0_snoop_o_40_sv2v_reg,el0_snoop_o_39_sv2v_reg,el0_snoop_o_38_sv2v_reg,
  el0_snoop_o_37_sv2v_reg,el0_snoop_o_36_sv2v_reg,el0_snoop_o_35_sv2v_reg,
  el0_snoop_o_34_sv2v_reg,el0_snoop_o_33_sv2v_reg,el0_snoop_o_32_sv2v_reg,
  el0_snoop_o_31_sv2v_reg,el0_snoop_o_30_sv2v_reg,el0_snoop_o_29_sv2v_reg,el0_snoop_o_28_sv2v_reg,
  el0_snoop_o_27_sv2v_reg,el0_snoop_o_26_sv2v_reg,el0_snoop_o_25_sv2v_reg,
  el0_snoop_o_24_sv2v_reg,el0_snoop_o_23_sv2v_reg,el0_snoop_o_22_sv2v_reg,
  el0_snoop_o_21_sv2v_reg,el0_snoop_o_20_sv2v_reg,el0_snoop_o_19_sv2v_reg,el0_snoop_o_18_sv2v_reg,
  el0_snoop_o_17_sv2v_reg,el0_snoop_o_16_sv2v_reg,el0_snoop_o_15_sv2v_reg,
  el0_snoop_o_14_sv2v_reg,el0_snoop_o_13_sv2v_reg,el0_snoop_o_12_sv2v_reg,
  el0_snoop_o_11_sv2v_reg,el0_snoop_o_10_sv2v_reg,el0_snoop_o_9_sv2v_reg,el0_snoop_o_8_sv2v_reg,
  el0_snoop_o_7_sv2v_reg,el0_snoop_o_6_sv2v_reg,el0_snoop_o_5_sv2v_reg,
  el0_snoop_o_4_sv2v_reg,el0_snoop_o_3_sv2v_reg,el0_snoop_o_2_sv2v_reg,el0_snoop_o_1_sv2v_reg,
  el0_snoop_o_0_sv2v_reg,el1_snoop_o_65_sv2v_reg,el1_snoop_o_64_sv2v_reg,
  el1_snoop_o_63_sv2v_reg,el1_snoop_o_62_sv2v_reg,el1_snoop_o_61_sv2v_reg,el1_snoop_o_60_sv2v_reg,
  el1_snoop_o_59_sv2v_reg,el1_snoop_o_58_sv2v_reg,el1_snoop_o_57_sv2v_reg,
  el1_snoop_o_56_sv2v_reg,el1_snoop_o_55_sv2v_reg,el1_snoop_o_54_sv2v_reg,
  el1_snoop_o_53_sv2v_reg,el1_snoop_o_52_sv2v_reg,el1_snoop_o_51_sv2v_reg,el1_snoop_o_50_sv2v_reg,
  el1_snoop_o_49_sv2v_reg,el1_snoop_o_48_sv2v_reg,el1_snoop_o_47_sv2v_reg,
  el1_snoop_o_46_sv2v_reg,el1_snoop_o_45_sv2v_reg,el1_snoop_o_44_sv2v_reg,
  el1_snoop_o_43_sv2v_reg,el1_snoop_o_42_sv2v_reg,el1_snoop_o_41_sv2v_reg,el1_snoop_o_40_sv2v_reg,
  el1_snoop_o_39_sv2v_reg,el1_snoop_o_38_sv2v_reg,el1_snoop_o_37_sv2v_reg,
  el1_snoop_o_36_sv2v_reg,el1_snoop_o_35_sv2v_reg,el1_snoop_o_34_sv2v_reg,
  el1_snoop_o_33_sv2v_reg,el1_snoop_o_32_sv2v_reg,el1_snoop_o_31_sv2v_reg,el1_snoop_o_30_sv2v_reg,
  el1_snoop_o_29_sv2v_reg,el1_snoop_o_28_sv2v_reg,el1_snoop_o_27_sv2v_reg,
  el1_snoop_o_26_sv2v_reg,el1_snoop_o_25_sv2v_reg,el1_snoop_o_24_sv2v_reg,
  el1_snoop_o_23_sv2v_reg,el1_snoop_o_22_sv2v_reg,el1_snoop_o_21_sv2v_reg,el1_snoop_o_20_sv2v_reg,
  el1_snoop_o_19_sv2v_reg,el1_snoop_o_18_sv2v_reg,el1_snoop_o_17_sv2v_reg,
  el1_snoop_o_16_sv2v_reg,el1_snoop_o_15_sv2v_reg,el1_snoop_o_14_sv2v_reg,
  el1_snoop_o_13_sv2v_reg,el1_snoop_o_12_sv2v_reg,el1_snoop_o_11_sv2v_reg,el1_snoop_o_10_sv2v_reg,
  el1_snoop_o_9_sv2v_reg,el1_snoop_o_8_sv2v_reg,el1_snoop_o_7_sv2v_reg,
  el1_snoop_o_6_sv2v_reg,el1_snoop_o_5_sv2v_reg,el1_snoop_o_4_sv2v_reg,
  el1_snoop_o_3_sv2v_reg,el1_snoop_o_2_sv2v_reg,el1_snoop_o_1_sv2v_reg,el1_snoop_o_0_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign el0_snoop_o[65] = el0_snoop_o_65_sv2v_reg;
  assign el0_snoop_o[64] = el0_snoop_o_64_sv2v_reg;
  assign el0_snoop_o[63] = el0_snoop_o_63_sv2v_reg;
  assign el0_snoop_o[62] = el0_snoop_o_62_sv2v_reg;
  assign el0_snoop_o[61] = el0_snoop_o_61_sv2v_reg;
  assign el0_snoop_o[60] = el0_snoop_o_60_sv2v_reg;
  assign el0_snoop_o[59] = el0_snoop_o_59_sv2v_reg;
  assign el0_snoop_o[58] = el0_snoop_o_58_sv2v_reg;
  assign el0_snoop_o[57] = el0_snoop_o_57_sv2v_reg;
  assign el0_snoop_o[56] = el0_snoop_o_56_sv2v_reg;
  assign el0_snoop_o[55] = el0_snoop_o_55_sv2v_reg;
  assign el0_snoop_o[54] = el0_snoop_o_54_sv2v_reg;
  assign el0_snoop_o[53] = el0_snoop_o_53_sv2v_reg;
  assign el0_snoop_o[52] = el0_snoop_o_52_sv2v_reg;
  assign el0_snoop_o[51] = el0_snoop_o_51_sv2v_reg;
  assign el0_snoop_o[50] = el0_snoop_o_50_sv2v_reg;
  assign el0_snoop_o[49] = el0_snoop_o_49_sv2v_reg;
  assign el0_snoop_o[48] = el0_snoop_o_48_sv2v_reg;
  assign el0_snoop_o[47] = el0_snoop_o_47_sv2v_reg;
  assign el0_snoop_o[46] = el0_snoop_o_46_sv2v_reg;
  assign el0_snoop_o[45] = el0_snoop_o_45_sv2v_reg;
  assign el0_snoop_o[44] = el0_snoop_o_44_sv2v_reg;
  assign el0_snoop_o[43] = el0_snoop_o_43_sv2v_reg;
  assign el0_snoop_o[42] = el0_snoop_o_42_sv2v_reg;
  assign el0_snoop_o[41] = el0_snoop_o_41_sv2v_reg;
  assign el0_snoop_o[40] = el0_snoop_o_40_sv2v_reg;
  assign el0_snoop_o[39] = el0_snoop_o_39_sv2v_reg;
  assign el0_snoop_o[38] = el0_snoop_o_38_sv2v_reg;
  assign el0_snoop_o[37] = el0_snoop_o_37_sv2v_reg;
  assign el0_snoop_o[36] = el0_snoop_o_36_sv2v_reg;
  assign el0_snoop_o[35] = el0_snoop_o_35_sv2v_reg;
  assign el0_snoop_o[34] = el0_snoop_o_34_sv2v_reg;
  assign el0_snoop_o[33] = el0_snoop_o_33_sv2v_reg;
  assign el0_snoop_o[32] = el0_snoop_o_32_sv2v_reg;
  assign el0_snoop_o[31] = el0_snoop_o_31_sv2v_reg;
  assign el0_snoop_o[30] = el0_snoop_o_30_sv2v_reg;
  assign el0_snoop_o[29] = el0_snoop_o_29_sv2v_reg;
  assign el0_snoop_o[28] = el0_snoop_o_28_sv2v_reg;
  assign el0_snoop_o[27] = el0_snoop_o_27_sv2v_reg;
  assign el0_snoop_o[26] = el0_snoop_o_26_sv2v_reg;
  assign el0_snoop_o[25] = el0_snoop_o_25_sv2v_reg;
  assign el0_snoop_o[24] = el0_snoop_o_24_sv2v_reg;
  assign el0_snoop_o[23] = el0_snoop_o_23_sv2v_reg;
  assign el0_snoop_o[22] = el0_snoop_o_22_sv2v_reg;
  assign el0_snoop_o[21] = el0_snoop_o_21_sv2v_reg;
  assign el0_snoop_o[20] = el0_snoop_o_20_sv2v_reg;
  assign el0_snoop_o[19] = el0_snoop_o_19_sv2v_reg;
  assign el0_snoop_o[18] = el0_snoop_o_18_sv2v_reg;
  assign el0_snoop_o[17] = el0_snoop_o_17_sv2v_reg;
  assign el0_snoop_o[16] = el0_snoop_o_16_sv2v_reg;
  assign el0_snoop_o[15] = el0_snoop_o_15_sv2v_reg;
  assign el0_snoop_o[14] = el0_snoop_o_14_sv2v_reg;
  assign el0_snoop_o[13] = el0_snoop_o_13_sv2v_reg;
  assign el0_snoop_o[12] = el0_snoop_o_12_sv2v_reg;
  assign el0_snoop_o[11] = el0_snoop_o_11_sv2v_reg;
  assign el0_snoop_o[10] = el0_snoop_o_10_sv2v_reg;
  assign el0_snoop_o[9] = el0_snoop_o_9_sv2v_reg;
  assign el0_snoop_o[8] = el0_snoop_o_8_sv2v_reg;
  assign el0_snoop_o[7] = el0_snoop_o_7_sv2v_reg;
  assign el0_snoop_o[6] = el0_snoop_o_6_sv2v_reg;
  assign el0_snoop_o[5] = el0_snoop_o_5_sv2v_reg;
  assign el0_snoop_o[4] = el0_snoop_o_4_sv2v_reg;
  assign el0_snoop_o[3] = el0_snoop_o_3_sv2v_reg;
  assign el0_snoop_o[2] = el0_snoop_o_2_sv2v_reg;
  assign el0_snoop_o[1] = el0_snoop_o_1_sv2v_reg;
  assign el0_snoop_o[0] = el0_snoop_o_0_sv2v_reg;
  assign el1_snoop_o[65] = el1_snoop_o_65_sv2v_reg;
  assign el1_snoop_o[64] = el1_snoop_o_64_sv2v_reg;
  assign el1_snoop_o[63] = el1_snoop_o_63_sv2v_reg;
  assign el1_snoop_o[62] = el1_snoop_o_62_sv2v_reg;
  assign el1_snoop_o[61] = el1_snoop_o_61_sv2v_reg;
  assign el1_snoop_o[60] = el1_snoop_o_60_sv2v_reg;
  assign el1_snoop_o[59] = el1_snoop_o_59_sv2v_reg;
  assign el1_snoop_o[58] = el1_snoop_o_58_sv2v_reg;
  assign el1_snoop_o[57] = el1_snoop_o_57_sv2v_reg;
  assign el1_snoop_o[56] = el1_snoop_o_56_sv2v_reg;
  assign el1_snoop_o[55] = el1_snoop_o_55_sv2v_reg;
  assign el1_snoop_o[54] = el1_snoop_o_54_sv2v_reg;
  assign el1_snoop_o[53] = el1_snoop_o_53_sv2v_reg;
  assign el1_snoop_o[52] = el1_snoop_o_52_sv2v_reg;
  assign el1_snoop_o[51] = el1_snoop_o_51_sv2v_reg;
  assign el1_snoop_o[50] = el1_snoop_o_50_sv2v_reg;
  assign el1_snoop_o[49] = el1_snoop_o_49_sv2v_reg;
  assign el1_snoop_o[48] = el1_snoop_o_48_sv2v_reg;
  assign el1_snoop_o[47] = el1_snoop_o_47_sv2v_reg;
  assign el1_snoop_o[46] = el1_snoop_o_46_sv2v_reg;
  assign el1_snoop_o[45] = el1_snoop_o_45_sv2v_reg;
  assign el1_snoop_o[44] = el1_snoop_o_44_sv2v_reg;
  assign el1_snoop_o[43] = el1_snoop_o_43_sv2v_reg;
  assign el1_snoop_o[42] = el1_snoop_o_42_sv2v_reg;
  assign el1_snoop_o[41] = el1_snoop_o_41_sv2v_reg;
  assign el1_snoop_o[40] = el1_snoop_o_40_sv2v_reg;
  assign el1_snoop_o[39] = el1_snoop_o_39_sv2v_reg;
  assign el1_snoop_o[38] = el1_snoop_o_38_sv2v_reg;
  assign el1_snoop_o[37] = el1_snoop_o_37_sv2v_reg;
  assign el1_snoop_o[36] = el1_snoop_o_36_sv2v_reg;
  assign el1_snoop_o[35] = el1_snoop_o_35_sv2v_reg;
  assign el1_snoop_o[34] = el1_snoop_o_34_sv2v_reg;
  assign el1_snoop_o[33] = el1_snoop_o_33_sv2v_reg;
  assign el1_snoop_o[32] = el1_snoop_o_32_sv2v_reg;
  assign el1_snoop_o[31] = el1_snoop_o_31_sv2v_reg;
  assign el1_snoop_o[30] = el1_snoop_o_30_sv2v_reg;
  assign el1_snoop_o[29] = el1_snoop_o_29_sv2v_reg;
  assign el1_snoop_o[28] = el1_snoop_o_28_sv2v_reg;
  assign el1_snoop_o[27] = el1_snoop_o_27_sv2v_reg;
  assign el1_snoop_o[26] = el1_snoop_o_26_sv2v_reg;
  assign el1_snoop_o[25] = el1_snoop_o_25_sv2v_reg;
  assign el1_snoop_o[24] = el1_snoop_o_24_sv2v_reg;
  assign el1_snoop_o[23] = el1_snoop_o_23_sv2v_reg;
  assign el1_snoop_o[22] = el1_snoop_o_22_sv2v_reg;
  assign el1_snoop_o[21] = el1_snoop_o_21_sv2v_reg;
  assign el1_snoop_o[20] = el1_snoop_o_20_sv2v_reg;
  assign el1_snoop_o[19] = el1_snoop_o_19_sv2v_reg;
  assign el1_snoop_o[18] = el1_snoop_o_18_sv2v_reg;
  assign el1_snoop_o[17] = el1_snoop_o_17_sv2v_reg;
  assign el1_snoop_o[16] = el1_snoop_o_16_sv2v_reg;
  assign el1_snoop_o[15] = el1_snoop_o_15_sv2v_reg;
  assign el1_snoop_o[14] = el1_snoop_o_14_sv2v_reg;
  assign el1_snoop_o[13] = el1_snoop_o_13_sv2v_reg;
  assign el1_snoop_o[12] = el1_snoop_o_12_sv2v_reg;
  assign el1_snoop_o[11] = el1_snoop_o_11_sv2v_reg;
  assign el1_snoop_o[10] = el1_snoop_o_10_sv2v_reg;
  assign el1_snoop_o[9] = el1_snoop_o_9_sv2v_reg;
  assign el1_snoop_o[8] = el1_snoop_o_8_sv2v_reg;
  assign el1_snoop_o[7] = el1_snoop_o_7_sv2v_reg;
  assign el1_snoop_o[6] = el1_snoop_o_6_sv2v_reg;
  assign el1_snoop_o[5] = el1_snoop_o_5_sv2v_reg;
  assign el1_snoop_o[4] = el1_snoop_o_4_sv2v_reg;
  assign el1_snoop_o[3] = el1_snoop_o_3_sv2v_reg;
  assign el1_snoop_o[2] = el1_snoop_o_2_sv2v_reg;
  assign el1_snoop_o[1] = el1_snoop_o_1_sv2v_reg;
  assign el1_snoop_o[0] = el1_snoop_o_0_sv2v_reg;
  assign N10 = N8 & N9;
  assign N11 = num_els_r[1] | N9;
  assign N13 = N8 | num_els_r[0];
  assign N15 = num_els_r[1] & num_els_r[0];
  assign { N20, N19 } = num_els_r + v_i;
  assign { N23, N22 } = { N20, N19 } - N21;
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N10;
  assign N1 = N12;
  assign N2 = N14;
  assign N3 = N15;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign full_o = (N0)? 1'b0 : 
                  (N1)? 1'b0 : 
                  (N2)? 1'b1 : 
                  (N3)? 1'b0 : 1'b0;
  assign el0_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b0 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el1_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b1 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N16 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N16 : 
                      (N1)? N17 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25 } = (N4)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                                        (N5)? data_i : 1'b0;
  assign N4 = mux0_sel;
  assign N5 = N24;
  assign data_o = (N6)? el1_snoop_o : 
                  (N7)? data_i : 1'b0;
  assign N6 = mux1_sel;
  assign N7 = N91;
  assign N8 = ~num_els_r[1];
  assign N9 = ~num_els_r[0];
  assign N12 = ~N11;
  assign N14 = ~N13;
  assign N16 = v_i & N92;
  assign N92 = ~yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N21 = v_o & yumi_i;
  assign N24 = ~mux0_sel;
  assign N91 = ~mux1_sel;

  always @(posedge clk_i) begin
    if(reset_i) begin
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      num_els_r_1_sv2v_reg <= N23;
      num_els_r_0_sv2v_reg <= N22;
    end 
    if(el0_enable) begin
      el0_snoop_o_65_sv2v_reg <= data_i[65];
      el0_snoop_o_64_sv2v_reg <= data_i[64];
      el0_snoop_o_63_sv2v_reg <= data_i[63];
      el0_snoop_o_62_sv2v_reg <= data_i[62];
      el0_snoop_o_61_sv2v_reg <= data_i[61];
      el0_snoop_o_60_sv2v_reg <= data_i[60];
      el0_snoop_o_59_sv2v_reg <= data_i[59];
      el0_snoop_o_58_sv2v_reg <= data_i[58];
      el0_snoop_o_57_sv2v_reg <= data_i[57];
      el0_snoop_o_56_sv2v_reg <= data_i[56];
      el0_snoop_o_55_sv2v_reg <= data_i[55];
      el0_snoop_o_54_sv2v_reg <= data_i[54];
      el0_snoop_o_53_sv2v_reg <= data_i[53];
      el0_snoop_o_52_sv2v_reg <= data_i[52];
      el0_snoop_o_51_sv2v_reg <= data_i[51];
      el0_snoop_o_50_sv2v_reg <= data_i[50];
      el0_snoop_o_49_sv2v_reg <= data_i[49];
      el0_snoop_o_48_sv2v_reg <= data_i[48];
      el0_snoop_o_47_sv2v_reg <= data_i[47];
      el0_snoop_o_46_sv2v_reg <= data_i[46];
      el0_snoop_o_45_sv2v_reg <= data_i[45];
      el0_snoop_o_44_sv2v_reg <= data_i[44];
      el0_snoop_o_43_sv2v_reg <= data_i[43];
      el0_snoop_o_42_sv2v_reg <= data_i[42];
      el0_snoop_o_41_sv2v_reg <= data_i[41];
      el0_snoop_o_40_sv2v_reg <= data_i[40];
      el0_snoop_o_39_sv2v_reg <= data_i[39];
      el0_snoop_o_38_sv2v_reg <= data_i[38];
      el0_snoop_o_37_sv2v_reg <= data_i[37];
      el0_snoop_o_36_sv2v_reg <= data_i[36];
      el0_snoop_o_35_sv2v_reg <= data_i[35];
      el0_snoop_o_34_sv2v_reg <= data_i[34];
      el0_snoop_o_33_sv2v_reg <= data_i[33];
      el0_snoop_o_32_sv2v_reg <= data_i[32];
      el0_snoop_o_31_sv2v_reg <= data_i[31];
      el0_snoop_o_30_sv2v_reg <= data_i[30];
      el0_snoop_o_29_sv2v_reg <= data_i[29];
      el0_snoop_o_28_sv2v_reg <= data_i[28];
      el0_snoop_o_27_sv2v_reg <= data_i[27];
      el0_snoop_o_26_sv2v_reg <= data_i[26];
      el0_snoop_o_25_sv2v_reg <= data_i[25];
      el0_snoop_o_24_sv2v_reg <= data_i[24];
      el0_snoop_o_23_sv2v_reg <= data_i[23];
      el0_snoop_o_22_sv2v_reg <= data_i[22];
      el0_snoop_o_21_sv2v_reg <= data_i[21];
      el0_snoop_o_20_sv2v_reg <= data_i[20];
      el0_snoop_o_19_sv2v_reg <= data_i[19];
      el0_snoop_o_18_sv2v_reg <= data_i[18];
      el0_snoop_o_17_sv2v_reg <= data_i[17];
      el0_snoop_o_16_sv2v_reg <= data_i[16];
      el0_snoop_o_15_sv2v_reg <= data_i[15];
      el0_snoop_o_14_sv2v_reg <= data_i[14];
      el0_snoop_o_13_sv2v_reg <= data_i[13];
      el0_snoop_o_12_sv2v_reg <= data_i[12];
      el0_snoop_o_11_sv2v_reg <= data_i[11];
      el0_snoop_o_10_sv2v_reg <= data_i[10];
      el0_snoop_o_9_sv2v_reg <= data_i[9];
      el0_snoop_o_8_sv2v_reg <= data_i[8];
      el0_snoop_o_7_sv2v_reg <= data_i[7];
      el0_snoop_o_6_sv2v_reg <= data_i[6];
      el0_snoop_o_5_sv2v_reg <= data_i[5];
      el0_snoop_o_4_sv2v_reg <= data_i[4];
      el0_snoop_o_3_sv2v_reg <= data_i[3];
      el0_snoop_o_2_sv2v_reg <= data_i[2];
      el0_snoop_o_1_sv2v_reg <= data_i[1];
      el0_snoop_o_0_sv2v_reg <= data_i[0];
    end 
    if(el1_enable) begin
      el1_snoop_o_65_sv2v_reg <= N90;
      el1_snoop_o_64_sv2v_reg <= N89;
      el1_snoop_o_63_sv2v_reg <= N88;
      el1_snoop_o_62_sv2v_reg <= N87;
      el1_snoop_o_61_sv2v_reg <= N86;
      el1_snoop_o_60_sv2v_reg <= N85;
      el1_snoop_o_59_sv2v_reg <= N84;
      el1_snoop_o_58_sv2v_reg <= N83;
      el1_snoop_o_57_sv2v_reg <= N82;
      el1_snoop_o_56_sv2v_reg <= N81;
      el1_snoop_o_55_sv2v_reg <= N80;
      el1_snoop_o_54_sv2v_reg <= N79;
      el1_snoop_o_53_sv2v_reg <= N78;
      el1_snoop_o_52_sv2v_reg <= N77;
      el1_snoop_o_51_sv2v_reg <= N76;
      el1_snoop_o_50_sv2v_reg <= N75;
      el1_snoop_o_49_sv2v_reg <= N74;
      el1_snoop_o_48_sv2v_reg <= N73;
      el1_snoop_o_47_sv2v_reg <= N72;
      el1_snoop_o_46_sv2v_reg <= N71;
      el1_snoop_o_45_sv2v_reg <= N70;
      el1_snoop_o_44_sv2v_reg <= N69;
      el1_snoop_o_43_sv2v_reg <= N68;
      el1_snoop_o_42_sv2v_reg <= N67;
      el1_snoop_o_41_sv2v_reg <= N66;
      el1_snoop_o_40_sv2v_reg <= N65;
      el1_snoop_o_39_sv2v_reg <= N64;
      el1_snoop_o_38_sv2v_reg <= N63;
      el1_snoop_o_37_sv2v_reg <= N62;
      el1_snoop_o_36_sv2v_reg <= N61;
      el1_snoop_o_35_sv2v_reg <= N60;
      el1_snoop_o_34_sv2v_reg <= N59;
      el1_snoop_o_33_sv2v_reg <= N58;
      el1_snoop_o_32_sv2v_reg <= N57;
      el1_snoop_o_31_sv2v_reg <= N56;
      el1_snoop_o_30_sv2v_reg <= N55;
      el1_snoop_o_29_sv2v_reg <= N54;
      el1_snoop_o_28_sv2v_reg <= N53;
      el1_snoop_o_27_sv2v_reg <= N52;
      el1_snoop_o_26_sv2v_reg <= N51;
      el1_snoop_o_25_sv2v_reg <= N50;
      el1_snoop_o_24_sv2v_reg <= N49;
      el1_snoop_o_23_sv2v_reg <= N48;
      el1_snoop_o_22_sv2v_reg <= N47;
      el1_snoop_o_21_sv2v_reg <= N46;
      el1_snoop_o_20_sv2v_reg <= N45;
      el1_snoop_o_19_sv2v_reg <= N44;
      el1_snoop_o_18_sv2v_reg <= N43;
      el1_snoop_o_17_sv2v_reg <= N42;
      el1_snoop_o_16_sv2v_reg <= N41;
      el1_snoop_o_15_sv2v_reg <= N40;
      el1_snoop_o_14_sv2v_reg <= N39;
      el1_snoop_o_13_sv2v_reg <= N38;
      el1_snoop_o_12_sv2v_reg <= N37;
      el1_snoop_o_11_sv2v_reg <= N36;
      el1_snoop_o_10_sv2v_reg <= N35;
      el1_snoop_o_9_sv2v_reg <= N34;
      el1_snoop_o_8_sv2v_reg <= N33;
      el1_snoop_o_7_sv2v_reg <= N32;
      el1_snoop_o_6_sv2v_reg <= N31;
      el1_snoop_o_5_sv2v_reg <= N30;
      el1_snoop_o_4_sv2v_reg <= N29;
      el1_snoop_o_3_sv2v_reg <= N28;
      el1_snoop_o_2_sv2v_reg <= N27;
      el1_snoop_o_1_sv2v_reg <= N26;
      el1_snoop_o_0_sv2v_reg <= N25;
    end 
  end


endmodule



module bsg_mux_segmented_segments_p4_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [31:0] data0_i;
  input [31:0] data1_i;
  input [3:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N4)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N5)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N6)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N7)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign N4 = ~sel_i[0];
  assign N5 = ~sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = ~sel_i[3];

endmodule



module bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p4
(
  clk_i,
  reset_i,
  sbuf_entry_i,
  v_i,
  sbuf_entry_o,
  v_o,
  yumi_i,
  empty_o,
  full_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o
);

  input [65:0] sbuf_entry_i;
  output [65:0] sbuf_entry_o;
  input [27:0] bypass_addr_i;
  output [31:0] bypass_data_o;
  output [3:0] bypass_mask_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  output full_o;
  wire [65:0] sbuf_entry_o,el0,el1;
  wire [31:0] bypass_data_o,el0or1_data,bypass_data_n;
  wire [3:0] bypass_mask_o,bypass_mask_n;
  wire v_o,empty_o,full_o,N0,el0_valid,el1_valid,tag_hit0_n,tag_hit1_n,tag_hit2_n,
  _2_net__3_,_2_net__2_,_2_net__1_,_2_net__0_,_4_net__3_,_4_net__2_,_4_net__1_,
  _4_net__0_,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  wire [3:3] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  reg bypass_data_o_31_sv2v_reg,bypass_data_o_30_sv2v_reg,bypass_data_o_29_sv2v_reg,
  bypass_data_o_28_sv2v_reg,bypass_data_o_27_sv2v_reg,bypass_data_o_26_sv2v_reg,
  bypass_data_o_25_sv2v_reg,bypass_data_o_24_sv2v_reg,bypass_data_o_23_sv2v_reg,
  bypass_data_o_22_sv2v_reg,bypass_data_o_21_sv2v_reg,bypass_data_o_20_sv2v_reg,
  bypass_data_o_19_sv2v_reg,bypass_data_o_18_sv2v_reg,bypass_data_o_17_sv2v_reg,
  bypass_data_o_16_sv2v_reg,bypass_data_o_15_sv2v_reg,bypass_data_o_14_sv2v_reg,
  bypass_data_o_13_sv2v_reg,bypass_data_o_12_sv2v_reg,bypass_data_o_11_sv2v_reg,
  bypass_data_o_10_sv2v_reg,bypass_data_o_9_sv2v_reg,bypass_data_o_8_sv2v_reg,
  bypass_data_o_7_sv2v_reg,bypass_data_o_6_sv2v_reg,bypass_data_o_5_sv2v_reg,
  bypass_data_o_4_sv2v_reg,bypass_data_o_3_sv2v_reg,bypass_data_o_2_sv2v_reg,bypass_data_o_1_sv2v_reg,
  bypass_data_o_0_sv2v_reg,bypass_mask_o_3_sv2v_reg,bypass_mask_o_2_sv2v_reg,
  bypass_mask_o_1_sv2v_reg,bypass_mask_o_0_sv2v_reg;
  assign bypass_data_o[31] = bypass_data_o_31_sv2v_reg;
  assign bypass_data_o[30] = bypass_data_o_30_sv2v_reg;
  assign bypass_data_o[29] = bypass_data_o_29_sv2v_reg;
  assign bypass_data_o[28] = bypass_data_o_28_sv2v_reg;
  assign bypass_data_o[27] = bypass_data_o_27_sv2v_reg;
  assign bypass_data_o[26] = bypass_data_o_26_sv2v_reg;
  assign bypass_data_o[25] = bypass_data_o_25_sv2v_reg;
  assign bypass_data_o[24] = bypass_data_o_24_sv2v_reg;
  assign bypass_data_o[23] = bypass_data_o_23_sv2v_reg;
  assign bypass_data_o[22] = bypass_data_o_22_sv2v_reg;
  assign bypass_data_o[21] = bypass_data_o_21_sv2v_reg;
  assign bypass_data_o[20] = bypass_data_o_20_sv2v_reg;
  assign bypass_data_o[19] = bypass_data_o_19_sv2v_reg;
  assign bypass_data_o[18] = bypass_data_o_18_sv2v_reg;
  assign bypass_data_o[17] = bypass_data_o_17_sv2v_reg;
  assign bypass_data_o[16] = bypass_data_o_16_sv2v_reg;
  assign bypass_data_o[15] = bypass_data_o_15_sv2v_reg;
  assign bypass_data_o[14] = bypass_data_o_14_sv2v_reg;
  assign bypass_data_o[13] = bypass_data_o_13_sv2v_reg;
  assign bypass_data_o[12] = bypass_data_o_12_sv2v_reg;
  assign bypass_data_o[11] = bypass_data_o_11_sv2v_reg;
  assign bypass_data_o[10] = bypass_data_o_10_sv2v_reg;
  assign bypass_data_o[9] = bypass_data_o_9_sv2v_reg;
  assign bypass_data_o[8] = bypass_data_o_8_sv2v_reg;
  assign bypass_data_o[7] = bypass_data_o_7_sv2v_reg;
  assign bypass_data_o[6] = bypass_data_o_6_sv2v_reg;
  assign bypass_data_o[5] = bypass_data_o_5_sv2v_reg;
  assign bypass_data_o[4] = bypass_data_o_4_sv2v_reg;
  assign bypass_data_o[3] = bypass_data_o_3_sv2v_reg;
  assign bypass_data_o[2] = bypass_data_o_2_sv2v_reg;
  assign bypass_data_o[1] = bypass_data_o_1_sv2v_reg;
  assign bypass_data_o[0] = bypass_data_o_0_sv2v_reg;
  assign bypass_mask_o[3] = bypass_mask_o_3_sv2v_reg;
  assign bypass_mask_o[2] = bypass_mask_o_2_sv2v_reg;
  assign bypass_mask_o[1] = bypass_mask_o_1_sv2v_reg;
  assign bypass_mask_o[0] = bypass_mask_o_0_sv2v_reg;

  bsg_cache_buffer_queue_width_p66
  q0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .data_i(sbuf_entry_i),
    .v_o(v_o),
    .data_o(sbuf_entry_o),
    .yumi_i(yumi_i),
    .el0_valid_o(el0_valid),
    .el1_valid_o(el1_valid),
    .el0_snoop_o(el0),
    .el1_snoop_o(el1),
    .empty_o(empty_o),
    .full_o(full_o)
  );

  assign tag_hit0_n = bypass_addr_i[27:2] == el0[65:40];
  assign tag_hit1_n = bypass_addr_i[27:2] == el1[65:40];
  assign tag_hit2_n = bypass_addr_i[27:2] == sbuf_entry_i[65:40];

  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(el1[37:6]),
    .data1_i(el0[37:6]),
    .sel_i({ _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(sbuf_entry_i[37:6]),
    .sel_i({ _4_net__3_, _4_net__2_, _4_net__1_, _4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = bypass_v_i;
  assign tag_hit0x4[3] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[3] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[3] = tag_hit2_n & v_i;
  assign bypass_mask_n[3] = N5 | N6;
  assign N5 = N3 | N4;
  assign N3 = tag_hit0x4[3] & el0[5];
  assign N4 = tag_hit1x4[3] & el1[5];
  assign N6 = tag_hit2x4[3] & sbuf_entry_i[5];
  assign bypass_mask_n[2] = N9 | N10;
  assign N9 = N7 | N8;
  assign N7 = tag_hit0x4[3] & el0[4];
  assign N8 = tag_hit1x4[3] & el1[4];
  assign N10 = tag_hit2x4[3] & sbuf_entry_i[4];
  assign bypass_mask_n[1] = N13 | N14;
  assign N13 = N11 | N12;
  assign N11 = tag_hit0x4[3] & el0[3];
  assign N12 = tag_hit1x4[3] & el1[3];
  assign N14 = tag_hit2x4[3] & sbuf_entry_i[3];
  assign bypass_mask_n[0] = N17 | N18;
  assign N17 = N15 | N16;
  assign N15 = tag_hit0x4[3] & el0[2];
  assign N16 = tag_hit1x4[3] & el1[2];
  assign N18 = tag_hit2x4[3] & sbuf_entry_i[2];
  assign _2_net__3_ = tag_hit0x4[3] & el0[5];
  assign _2_net__2_ = tag_hit0x4[3] & el0[4];
  assign _2_net__1_ = tag_hit0x4[3] & el0[3];
  assign _2_net__0_ = tag_hit0x4[3] & el0[2];
  assign _4_net__3_ = tag_hit2x4[3] & sbuf_entry_i[5];
  assign _4_net__2_ = tag_hit2x4[3] & sbuf_entry_i[4];
  assign _4_net__1_ = tag_hit2x4[3] & sbuf_entry_i[3];
  assign _4_net__0_ = tag_hit2x4[3] & sbuf_entry_i[2];
  assign N1 = ~bypass_v_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      bypass_data_o_31_sv2v_reg <= 1'b0;
      bypass_data_o_30_sv2v_reg <= 1'b0;
      bypass_data_o_29_sv2v_reg <= 1'b0;
      bypass_data_o_28_sv2v_reg <= 1'b0;
      bypass_data_o_27_sv2v_reg <= 1'b0;
      bypass_data_o_26_sv2v_reg <= 1'b0;
      bypass_data_o_25_sv2v_reg <= 1'b0;
      bypass_data_o_24_sv2v_reg <= 1'b0;
      bypass_data_o_23_sv2v_reg <= 1'b0;
      bypass_data_o_22_sv2v_reg <= 1'b0;
      bypass_data_o_21_sv2v_reg <= 1'b0;
      bypass_data_o_20_sv2v_reg <= 1'b0;
      bypass_data_o_19_sv2v_reg <= 1'b0;
      bypass_data_o_18_sv2v_reg <= 1'b0;
      bypass_data_o_17_sv2v_reg <= 1'b0;
      bypass_data_o_16_sv2v_reg <= 1'b0;
      bypass_data_o_15_sv2v_reg <= 1'b0;
      bypass_data_o_14_sv2v_reg <= 1'b0;
      bypass_data_o_13_sv2v_reg <= 1'b0;
      bypass_data_o_12_sv2v_reg <= 1'b0;
      bypass_data_o_11_sv2v_reg <= 1'b0;
      bypass_data_o_10_sv2v_reg <= 1'b0;
      bypass_data_o_9_sv2v_reg <= 1'b0;
      bypass_data_o_8_sv2v_reg <= 1'b0;
      bypass_data_o_7_sv2v_reg <= 1'b0;
      bypass_data_o_6_sv2v_reg <= 1'b0;
      bypass_data_o_5_sv2v_reg <= 1'b0;
      bypass_data_o_4_sv2v_reg <= 1'b0;
      bypass_data_o_3_sv2v_reg <= 1'b0;
      bypass_data_o_2_sv2v_reg <= 1'b0;
      bypass_data_o_1_sv2v_reg <= 1'b0;
      bypass_data_o_0_sv2v_reg <= 1'b0;
      bypass_mask_o_3_sv2v_reg <= 1'b0;
      bypass_mask_o_2_sv2v_reg <= 1'b0;
      bypass_mask_o_1_sv2v_reg <= 1'b0;
      bypass_mask_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      bypass_data_o_31_sv2v_reg <= bypass_data_n[31];
      bypass_data_o_30_sv2v_reg <= bypass_data_n[30];
      bypass_data_o_29_sv2v_reg <= bypass_data_n[29];
      bypass_data_o_28_sv2v_reg <= bypass_data_n[28];
      bypass_data_o_27_sv2v_reg <= bypass_data_n[27];
      bypass_data_o_26_sv2v_reg <= bypass_data_n[26];
      bypass_data_o_25_sv2v_reg <= bypass_data_n[25];
      bypass_data_o_24_sv2v_reg <= bypass_data_n[24];
      bypass_data_o_23_sv2v_reg <= bypass_data_n[23];
      bypass_data_o_22_sv2v_reg <= bypass_data_n[22];
      bypass_data_o_21_sv2v_reg <= bypass_data_n[21];
      bypass_data_o_20_sv2v_reg <= bypass_data_n[20];
      bypass_data_o_19_sv2v_reg <= bypass_data_n[19];
      bypass_data_o_18_sv2v_reg <= bypass_data_n[18];
      bypass_data_o_17_sv2v_reg <= bypass_data_n[17];
      bypass_data_o_16_sv2v_reg <= bypass_data_n[16];
      bypass_data_o_15_sv2v_reg <= bypass_data_n[15];
      bypass_data_o_14_sv2v_reg <= bypass_data_n[14];
      bypass_data_o_13_sv2v_reg <= bypass_data_n[13];
      bypass_data_o_12_sv2v_reg <= bypass_data_n[12];
      bypass_data_o_11_sv2v_reg <= bypass_data_n[11];
      bypass_data_o_10_sv2v_reg <= bypass_data_n[10];
      bypass_data_o_9_sv2v_reg <= bypass_data_n[9];
      bypass_data_o_8_sv2v_reg <= bypass_data_n[8];
      bypass_data_o_7_sv2v_reg <= bypass_data_n[7];
      bypass_data_o_6_sv2v_reg <= bypass_data_n[6];
      bypass_data_o_5_sv2v_reg <= bypass_data_n[5];
      bypass_data_o_4_sv2v_reg <= bypass_data_n[4];
      bypass_data_o_3_sv2v_reg <= bypass_data_n[3];
      bypass_data_o_2_sv2v_reg <= bypass_data_n[2];
      bypass_data_o_1_sv2v_reg <= bypass_data_n[1];
      bypass_data_o_0_sv2v_reg <= bypass_data_n[0];
      bypass_mask_o_3_sv2v_reg <= bypass_mask_n[3];
      bypass_mask_o_2_sv2v_reg <= bypass_mask_n[2];
      bypass_mask_o_1_sv2v_reg <= bypass_mask_n[1];
      bypass_mask_o_0_sv2v_reg <= bypass_mask_n[0];
    end 
  end


endmodule



module bsg_decode_num_out_p1
(
  i,
  o
);

  input [0:0] i;
  output [0:0] o;
  wire [0:0] o;
  assign o[0] = 1'b1;

endmodule



module bsg_mux_width_p32_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [95:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[31] = (N2)? data_i[31] : 
                      (N3)? data_i[63] : 
                      (N4)? data_i[95] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[30] = (N2)? data_i[30] : 
                      (N3)? data_i[62] : 
                      (N4)? data_i[94] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N3)? data_i[61] : 
                      (N4)? data_i[93] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N3)? data_i[60] : 
                      (N4)? data_i[92] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N3)? data_i[59] : 
                      (N4)? data_i[91] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N3)? data_i[58] : 
                      (N4)? data_i[90] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N3)? data_i[57] : 
                      (N4)? data_i[89] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N3)? data_i[56] : 
                      (N4)? data_i[88] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N3)? data_i[55] : 
                      (N4)? data_i[87] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N3)? data_i[54] : 
                      (N4)? data_i[86] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N3)? data_i[53] : 
                      (N4)? data_i[85] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N3)? data_i[52] : 
                      (N4)? data_i[84] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N3)? data_i[51] : 
                      (N4)? data_i[83] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N3)? data_i[50] : 
                      (N4)? data_i[82] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N3)? data_i[49] : 
                      (N4)? data_i[81] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N3)? data_i[48] : 
                      (N4)? data_i[80] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N3)? data_i[47] : 
                      (N4)? data_i[79] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N3)? data_i[46] : 
                      (N4)? data_i[78] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N3)? data_i[45] : 
                      (N4)? data_i[77] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N3)? data_i[44] : 
                      (N4)? data_i[76] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N3)? data_i[43] : 
                      (N4)? data_i[75] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N3)? data_i[42] : 
                      (N4)? data_i[74] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N3)? data_i[41] : 
                     (N4)? data_i[73] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N3)? data_i[40] : 
                     (N4)? data_i[72] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N3)? data_i[39] : 
                     (N4)? data_i[71] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N3)? data_i[38] : 
                     (N4)? data_i[70] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N3)? data_i[37] : 
                     (N4)? data_i[69] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N3)? data_i[36] : 
                     (N4)? data_i[68] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[35] : 
                     (N4)? data_i[67] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[34] : 
                     (N4)? data_i[66] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[33] : 
                     (N4)? data_i[65] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[32] : 
                     (N4)? data_i[64] : 1'b0;

endmodule



module bsg_mux_width_p4_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [11:0] data_i;
  input [1:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[7] : 
                     (N4)? data_i[11] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[6] : 
                     (N4)? data_i[10] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[5] : 
                     (N4)? data_i[9] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[4] : 
                     (N4)? data_i[8] : 1'b0;

endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_mux_width_p8_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [1:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[15] : 
                     (N3)? data_i[23] : 
                     (N5)? data_i[31] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[14] : 
                     (N3)? data_i[22] : 
                     (N5)? data_i[30] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[13] : 
                     (N3)? data_i[21] : 
                     (N5)? data_i[29] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[12] : 
                     (N3)? data_i[20] : 
                     (N5)? data_i[28] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[11] : 
                     (N3)? data_i[19] : 
                     (N5)? data_i[27] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[10] : 
                     (N3)? data_i[18] : 
                     (N5)? data_i[26] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[9] : 
                     (N3)? data_i[17] : 
                     (N5)? data_i[25] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[8] : 
                     (N3)? data_i[16] : 
                     (N5)? data_i[24] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p16_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[31] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[30] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[29] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[28] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[27] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[26] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[25] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[24] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[23] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[22] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[21] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[20] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[19] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[18] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[17] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[16] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_cache
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  yumi_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [69:0] cache_pkt_i;
  output [31:0] data_o;
  output [32:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output yumi_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;
  wire [31:0] data_o,dma_data_o,data_tl_r,data_v_r,snoop_word_lo,bypass_data_lo,sbuf_data_in,
  atomic_mem_data,atomic_alu_result,\sbuf_in_sel_2_.slice_data ,ld_data_way_picked,
  ld_data_offset_picked,bypass_data_masked,snoop_or_ld_data,expanded_mask_v,
  ld_data_masked,ld_data_final_lo;
  wire [32:0] dma_pkt_o;
  wire yumi_o,v_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,v_we_o,N0,N1,N3,N4,N5,N6,
  N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,
  tl_we,sbuf_hazard,N67,N68,v_tl_r,N69,N70,N71,N72,N73,tag_mem_v_li,tag_mem_w_li,
  data_mem_v_li,data_mem_w_li,track_mem_v_li,track_mem_w_li,N74,N75,N76,v_v_r,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,tag_hit_found,N90,N91,N92,N93,
  partial_st,N94,N95,N96,N97,partial_st_tl,N98,N99,N100,N101,N102,partial_st_v,
  ld_st_amo_tag_miss,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,bypass_track_lo,track_miss,N120,N121,N122,N123,N124,N125,N126,
  tagfl_hit,aflinv_hit,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,
  alock_miss,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,aunlock_hit,miss_v,
  retval_op_v,stat_mem_v_li,stat_mem_w_li,sbuf_empty_lo,tbuf_empty_lo,dma_done_li,
  miss_track_data_we_lo,miss_stat_mem_v_lo,miss_stat_mem_w_lo,miss_tag_mem_v_lo,
  miss_tag_mem_w_lo,miss_track_mem_v_lo,miss_track_mem_w_lo,recover_lo,miss_done_lo,_1_net_,
  select_snoop_data_r_lo,dma_data_mem_v_lo,dma_data_mem_w_lo,dma_evict_lo,
  sbuf_entry_li_data__31_,sbuf_entry_li_data__30_,sbuf_entry_li_data__29_,
  sbuf_entry_li_data__28_,sbuf_entry_li_data__27_,sbuf_entry_li_data__26_,sbuf_entry_li_data__25_,
  sbuf_entry_li_data__24_,sbuf_entry_li_data__23_,sbuf_entry_li_data__22_,
  sbuf_entry_li_data__21_,sbuf_entry_li_data__20_,sbuf_entry_li_data__19_,
  sbuf_entry_li_data__18_,sbuf_entry_li_data__17_,sbuf_entry_li_data__16_,sbuf_entry_li_data__15_,
  sbuf_entry_li_data__14_,sbuf_entry_li_data__13_,sbuf_entry_li_data__12_,
  sbuf_entry_li_data__11_,sbuf_entry_li_data__10_,sbuf_entry_li_data__9_,
  sbuf_entry_li_data__8_,sbuf_entry_li_data__7_,sbuf_entry_li_data__6_,sbuf_entry_li_data__5_,
  sbuf_entry_li_data__4_,sbuf_entry_li_data__3_,sbuf_entry_li_data__2_,
  sbuf_entry_li_data__1_,sbuf_entry_li_data__0_,sbuf_entry_li_mask__3_,sbuf_entry_li_mask__2_,
  sbuf_entry_li_mask__1_,sbuf_entry_li_mask__0_,sbuf_entry_li_way_id__1_,
  sbuf_entry_li_way_id__0_,sbuf_v_li,sbuf_v_lo,sbuf_yumi_li,sbuf_full_lo,sbuf_bypass_v_li,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,ld_data_final_li_1__31_,ld_data_final_li_1__30_,
  ld_data_final_li_1__29_,ld_data_final_li_1__28_,ld_data_final_li_1__27_,ld_data_final_li_1__26_,
  ld_data_final_li_1__25_,ld_data_final_li_1__24_,ld_data_final_li_1__23_,
  ld_data_final_li_1__22_,ld_data_final_li_1__21_,ld_data_final_li_1__20_,
  ld_data_final_li_1__19_,ld_data_final_li_1__18_,ld_data_final_li_1__17_,ld_data_final_li_1__16_,
  ld_data_final_li_0__31_,ld_data_final_li_0__30_,ld_data_final_li_0__29_,
  ld_data_final_li_0__28_,ld_data_final_li_0__27_,ld_data_final_li_0__26_,
  ld_data_final_li_0__25_,ld_data_final_li_0__24_,ld_data_final_li_0__23_,ld_data_final_li_0__22_,
  ld_data_final_li_0__21_,ld_data_final_li_0__20_,ld_data_final_li_0__19_,
  ld_data_final_li_0__18_,ld_data_final_li_0__17_,ld_data_final_li_0__16_,
  ld_data_final_li_0__15_,ld_data_final_li_0__14_,ld_data_final_li_0__13_,ld_data_final_li_0__12_,
  ld_data_final_li_0__11_,ld_data_final_li_0__10_,ld_data_final_li_0__9_,
  ld_data_final_li_0__8_,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,
  N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,
  N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
  N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,
  N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,
  N501,N502,tbuf_v_li,tbuf_v_lo,tbuf_yumi_li,tbuf_full_lo,tbuf_bypass_v_li,N503,N504,
  N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,
  N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,
  N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,
  N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
  N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,
  N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,tl_ready,
  N599,N600,tagst_write_en,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N2,N666,N667,N668,N669,N670,N671,N672,N673,N674,
  N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,
  N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,
  N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,
  N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,
  N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,
  N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,
  N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,
  N787,N788,N789;
  wire [20:0] decode,decode_tl_r,decode_v_r;
  wire [3:0] mask_tl_r,mask_v_r,valid_v_r,lock_v_r,tag_hit_v,dma_cmd_lo,bypass_mask_lo,
  sbuf_way_decode,sbuf_expand_mask,sbuf_mask_in,\sbuf_in_sel_0_.decode_lo ,
  tbuf_way_decode,tbuf_word_offset_decode,addr_way_decode;
  wire [27:0] addr_tl_r,addr_v_r,dma_addr_lo,tbuf_addr_lo;
  wire [5:0] tag_mem_addr_li,track_mem_addr_li,stat_mem_addr_li,miss_stat_mem_addr_lo,
  miss_tag_mem_addr_lo,miss_track_mem_addr_lo;
  wire [79:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo,miss_tag_mem_data_lo,
  miss_tag_mem_w_mask_lo;
  wire [7:0] data_mem_addr_li,dma_data_mem_addr_lo,\ld_data_sel_0_.byte_sel ;
  wire [127:0] data_mem_data_li,data_mem_data_lo,ld_data_v_r,dma_data_mem_data_lo;
  wire [15:0] data_mem_w_mask_li,track_mem_data_li,track_mem_w_mask_li,track_mem_data_lo,
  track_data_v_r,miss_track_mem_w_mask_lo,miss_track_mem_data_lo,
  dma_data_mem_w_mask_lo,sbuf_data_mem_w_mask,tbuf_track_mem_w_mask,\ld_data_sel_1_.byte_sel ;
  wire [71:0] tag_v_r;
  wire [1:0] tag_hit_way_id,dma_way_lo,chosen_way_lo,\sbuf_in_sel_1_.decode_lo ,tbuf_way_li,
  tbuf_way_lo;
  wire [6:0] stat_mem_data_li,stat_mem_w_mask_li,stat_mem_data_lo,miss_stat_mem_data_lo,
  miss_stat_mem_w_mask_lo;
  wire [65:0] sbuf_entry_lo;
  wire [0:0] sbuf_burst_offset_decode,\sbuf_in_sel_2_.decode_lo ;
  wire [11:0] sbuf_mask_in_mux_li;
  wire [2:0] plru_decode_data_lo,plru_decode_mask_lo;
  reg data_tl_r_31_sv2v_reg,data_tl_r_30_sv2v_reg,data_tl_r_29_sv2v_reg,
  data_tl_r_28_sv2v_reg,data_tl_r_27_sv2v_reg,data_tl_r_26_sv2v_reg,data_tl_r_25_sv2v_reg,
  data_tl_r_24_sv2v_reg,data_tl_r_23_sv2v_reg,data_tl_r_22_sv2v_reg,
  data_tl_r_21_sv2v_reg,data_tl_r_20_sv2v_reg,data_tl_r_19_sv2v_reg,data_tl_r_18_sv2v_reg,
  data_tl_r_17_sv2v_reg,data_tl_r_16_sv2v_reg,data_tl_r_15_sv2v_reg,data_tl_r_14_sv2v_reg,
  data_tl_r_13_sv2v_reg,data_tl_r_12_sv2v_reg,data_tl_r_11_sv2v_reg,
  data_tl_r_10_sv2v_reg,data_tl_r_9_sv2v_reg,data_tl_r_8_sv2v_reg,data_tl_r_7_sv2v_reg,
  data_tl_r_6_sv2v_reg,data_tl_r_5_sv2v_reg,data_tl_r_4_sv2v_reg,data_tl_r_3_sv2v_reg,
  data_tl_r_2_sv2v_reg,data_tl_r_1_sv2v_reg,data_tl_r_0_sv2v_reg,v_tl_r_sv2v_reg,
  decode_tl_r_20_sv2v_reg,decode_tl_r_19_sv2v_reg,decode_tl_r_18_sv2v_reg,
  decode_tl_r_17_sv2v_reg,decode_tl_r_16_sv2v_reg,decode_tl_r_15_sv2v_reg,decode_tl_r_14_sv2v_reg,
  decode_tl_r_13_sv2v_reg,decode_tl_r_12_sv2v_reg,decode_tl_r_11_sv2v_reg,
  decode_tl_r_10_sv2v_reg,decode_tl_r_9_sv2v_reg,decode_tl_r_8_sv2v_reg,
  decode_tl_r_7_sv2v_reg,decode_tl_r_6_sv2v_reg,decode_tl_r_5_sv2v_reg,decode_tl_r_4_sv2v_reg,
  decode_tl_r_3_sv2v_reg,decode_tl_r_2_sv2v_reg,decode_tl_r_1_sv2v_reg,
  decode_tl_r_0_sv2v_reg,mask_tl_r_3_sv2v_reg,mask_tl_r_2_sv2v_reg,mask_tl_r_1_sv2v_reg,
  mask_tl_r_0_sv2v_reg,addr_tl_r_27_sv2v_reg,addr_tl_r_26_sv2v_reg,addr_tl_r_25_sv2v_reg,
  addr_tl_r_24_sv2v_reg,addr_tl_r_23_sv2v_reg,addr_tl_r_22_sv2v_reg,
  addr_tl_r_21_sv2v_reg,addr_tl_r_20_sv2v_reg,addr_tl_r_19_sv2v_reg,addr_tl_r_18_sv2v_reg,
  addr_tl_r_17_sv2v_reg,addr_tl_r_16_sv2v_reg,addr_tl_r_15_sv2v_reg,addr_tl_r_14_sv2v_reg,
  addr_tl_r_13_sv2v_reg,addr_tl_r_12_sv2v_reg,addr_tl_r_11_sv2v_reg,
  addr_tl_r_10_sv2v_reg,addr_tl_r_9_sv2v_reg,addr_tl_r_8_sv2v_reg,addr_tl_r_7_sv2v_reg,
  addr_tl_r_6_sv2v_reg,addr_tl_r_5_sv2v_reg,addr_tl_r_4_sv2v_reg,addr_tl_r_3_sv2v_reg,
  addr_tl_r_2_sv2v_reg,addr_tl_r_1_sv2v_reg,addr_tl_r_0_sv2v_reg,ld_data_v_r_127_sv2v_reg,
  ld_data_v_r_126_sv2v_reg,ld_data_v_r_125_sv2v_reg,ld_data_v_r_124_sv2v_reg,
  ld_data_v_r_123_sv2v_reg,ld_data_v_r_122_sv2v_reg,ld_data_v_r_121_sv2v_reg,
  ld_data_v_r_120_sv2v_reg,ld_data_v_r_119_sv2v_reg,ld_data_v_r_118_sv2v_reg,
  ld_data_v_r_117_sv2v_reg,ld_data_v_r_116_sv2v_reg,ld_data_v_r_115_sv2v_reg,
  ld_data_v_r_114_sv2v_reg,ld_data_v_r_113_sv2v_reg,ld_data_v_r_112_sv2v_reg,ld_data_v_r_111_sv2v_reg,
  ld_data_v_r_110_sv2v_reg,ld_data_v_r_109_sv2v_reg,ld_data_v_r_108_sv2v_reg,
  ld_data_v_r_107_sv2v_reg,ld_data_v_r_106_sv2v_reg,ld_data_v_r_105_sv2v_reg,
  ld_data_v_r_104_sv2v_reg,ld_data_v_r_103_sv2v_reg,ld_data_v_r_102_sv2v_reg,
  ld_data_v_r_101_sv2v_reg,ld_data_v_r_100_sv2v_reg,ld_data_v_r_99_sv2v_reg,
  ld_data_v_r_98_sv2v_reg,ld_data_v_r_97_sv2v_reg,ld_data_v_r_96_sv2v_reg,ld_data_v_r_95_sv2v_reg,
  ld_data_v_r_94_sv2v_reg,ld_data_v_r_93_sv2v_reg,ld_data_v_r_92_sv2v_reg,
  ld_data_v_r_91_sv2v_reg,ld_data_v_r_90_sv2v_reg,ld_data_v_r_89_sv2v_reg,
  ld_data_v_r_88_sv2v_reg,ld_data_v_r_87_sv2v_reg,ld_data_v_r_86_sv2v_reg,ld_data_v_r_85_sv2v_reg,
  ld_data_v_r_84_sv2v_reg,ld_data_v_r_83_sv2v_reg,ld_data_v_r_82_sv2v_reg,
  ld_data_v_r_81_sv2v_reg,ld_data_v_r_80_sv2v_reg,ld_data_v_r_79_sv2v_reg,
  ld_data_v_r_78_sv2v_reg,ld_data_v_r_77_sv2v_reg,ld_data_v_r_76_sv2v_reg,ld_data_v_r_75_sv2v_reg,
  ld_data_v_r_74_sv2v_reg,ld_data_v_r_73_sv2v_reg,ld_data_v_r_72_sv2v_reg,
  ld_data_v_r_71_sv2v_reg,ld_data_v_r_70_sv2v_reg,ld_data_v_r_69_sv2v_reg,
  ld_data_v_r_68_sv2v_reg,ld_data_v_r_67_sv2v_reg,ld_data_v_r_66_sv2v_reg,ld_data_v_r_65_sv2v_reg,
  ld_data_v_r_64_sv2v_reg,ld_data_v_r_63_sv2v_reg,ld_data_v_r_62_sv2v_reg,
  ld_data_v_r_61_sv2v_reg,ld_data_v_r_60_sv2v_reg,ld_data_v_r_59_sv2v_reg,
  ld_data_v_r_58_sv2v_reg,ld_data_v_r_57_sv2v_reg,ld_data_v_r_56_sv2v_reg,ld_data_v_r_55_sv2v_reg,
  ld_data_v_r_54_sv2v_reg,ld_data_v_r_53_sv2v_reg,ld_data_v_r_52_sv2v_reg,
  ld_data_v_r_51_sv2v_reg,ld_data_v_r_50_sv2v_reg,ld_data_v_r_49_sv2v_reg,
  ld_data_v_r_48_sv2v_reg,ld_data_v_r_47_sv2v_reg,ld_data_v_r_46_sv2v_reg,ld_data_v_r_45_sv2v_reg,
  ld_data_v_r_44_sv2v_reg,ld_data_v_r_43_sv2v_reg,ld_data_v_r_42_sv2v_reg,
  ld_data_v_r_41_sv2v_reg,ld_data_v_r_40_sv2v_reg,ld_data_v_r_39_sv2v_reg,
  ld_data_v_r_38_sv2v_reg,ld_data_v_r_37_sv2v_reg,ld_data_v_r_36_sv2v_reg,ld_data_v_r_35_sv2v_reg,
  ld_data_v_r_34_sv2v_reg,ld_data_v_r_33_sv2v_reg,ld_data_v_r_32_sv2v_reg,
  ld_data_v_r_31_sv2v_reg,ld_data_v_r_30_sv2v_reg,ld_data_v_r_29_sv2v_reg,
  ld_data_v_r_28_sv2v_reg,ld_data_v_r_27_sv2v_reg,ld_data_v_r_26_sv2v_reg,ld_data_v_r_25_sv2v_reg,
  ld_data_v_r_24_sv2v_reg,ld_data_v_r_23_sv2v_reg,ld_data_v_r_22_sv2v_reg,
  ld_data_v_r_21_sv2v_reg,ld_data_v_r_20_sv2v_reg,ld_data_v_r_19_sv2v_reg,
  ld_data_v_r_18_sv2v_reg,ld_data_v_r_17_sv2v_reg,ld_data_v_r_16_sv2v_reg,ld_data_v_r_15_sv2v_reg,
  ld_data_v_r_14_sv2v_reg,ld_data_v_r_13_sv2v_reg,ld_data_v_r_12_sv2v_reg,
  ld_data_v_r_11_sv2v_reg,ld_data_v_r_10_sv2v_reg,ld_data_v_r_9_sv2v_reg,ld_data_v_r_8_sv2v_reg,
  ld_data_v_r_7_sv2v_reg,ld_data_v_r_6_sv2v_reg,ld_data_v_r_5_sv2v_reg,
  ld_data_v_r_4_sv2v_reg,ld_data_v_r_3_sv2v_reg,ld_data_v_r_2_sv2v_reg,
  ld_data_v_r_1_sv2v_reg,ld_data_v_r_0_sv2v_reg,v_v_r_sv2v_reg,track_data_v_r_15_sv2v_reg,
  track_data_v_r_14_sv2v_reg,track_data_v_r_13_sv2v_reg,track_data_v_r_12_sv2v_reg,
  track_data_v_r_11_sv2v_reg,track_data_v_r_10_sv2v_reg,track_data_v_r_9_sv2v_reg,
  track_data_v_r_8_sv2v_reg,track_data_v_r_7_sv2v_reg,track_data_v_r_6_sv2v_reg,
  track_data_v_r_5_sv2v_reg,track_data_v_r_4_sv2v_reg,track_data_v_r_3_sv2v_reg,
  track_data_v_r_2_sv2v_reg,track_data_v_r_1_sv2v_reg,track_data_v_r_0_sv2v_reg,
  mask_v_r_3_sv2v_reg,mask_v_r_2_sv2v_reg,mask_v_r_1_sv2v_reg,mask_v_r_0_sv2v_reg,
  decode_v_r_20_sv2v_reg,decode_v_r_19_sv2v_reg,decode_v_r_18_sv2v_reg,decode_v_r_17_sv2v_reg,
  decode_v_r_16_sv2v_reg,decode_v_r_15_sv2v_reg,decode_v_r_14_sv2v_reg,
  decode_v_r_13_sv2v_reg,decode_v_r_12_sv2v_reg,decode_v_r_11_sv2v_reg,decode_v_r_10_sv2v_reg,
  decode_v_r_9_sv2v_reg,decode_v_r_8_sv2v_reg,decode_v_r_7_sv2v_reg,
  decode_v_r_6_sv2v_reg,decode_v_r_5_sv2v_reg,decode_v_r_4_sv2v_reg,decode_v_r_3_sv2v_reg,
  decode_v_r_2_sv2v_reg,decode_v_r_1_sv2v_reg,decode_v_r_0_sv2v_reg,addr_v_r_27_sv2v_reg,
  addr_v_r_26_sv2v_reg,addr_v_r_25_sv2v_reg,addr_v_r_24_sv2v_reg,addr_v_r_23_sv2v_reg,
  addr_v_r_22_sv2v_reg,addr_v_r_21_sv2v_reg,addr_v_r_20_sv2v_reg,
  addr_v_r_19_sv2v_reg,addr_v_r_18_sv2v_reg,addr_v_r_17_sv2v_reg,addr_v_r_16_sv2v_reg,
  addr_v_r_15_sv2v_reg,addr_v_r_14_sv2v_reg,addr_v_r_13_sv2v_reg,addr_v_r_12_sv2v_reg,
  addr_v_r_11_sv2v_reg,addr_v_r_10_sv2v_reg,addr_v_r_9_sv2v_reg,addr_v_r_8_sv2v_reg,
  addr_v_r_7_sv2v_reg,addr_v_r_6_sv2v_reg,addr_v_r_5_sv2v_reg,addr_v_r_4_sv2v_reg,
  addr_v_r_3_sv2v_reg,addr_v_r_2_sv2v_reg,addr_v_r_1_sv2v_reg,addr_v_r_0_sv2v_reg,
  data_v_r_31_sv2v_reg,data_v_r_30_sv2v_reg,data_v_r_29_sv2v_reg,data_v_r_28_sv2v_reg,
  data_v_r_27_sv2v_reg,data_v_r_26_sv2v_reg,data_v_r_25_sv2v_reg,data_v_r_24_sv2v_reg,
  data_v_r_23_sv2v_reg,data_v_r_22_sv2v_reg,data_v_r_21_sv2v_reg,
  data_v_r_20_sv2v_reg,data_v_r_19_sv2v_reg,data_v_r_18_sv2v_reg,data_v_r_17_sv2v_reg,
  data_v_r_16_sv2v_reg,data_v_r_15_sv2v_reg,data_v_r_14_sv2v_reg,data_v_r_13_sv2v_reg,
  data_v_r_12_sv2v_reg,data_v_r_11_sv2v_reg,data_v_r_10_sv2v_reg,data_v_r_9_sv2v_reg,
  data_v_r_8_sv2v_reg,data_v_r_7_sv2v_reg,data_v_r_6_sv2v_reg,data_v_r_5_sv2v_reg,
  data_v_r_4_sv2v_reg,data_v_r_3_sv2v_reg,data_v_r_2_sv2v_reg,data_v_r_1_sv2v_reg,
  data_v_r_0_sv2v_reg,valid_v_r_3_sv2v_reg,valid_v_r_2_sv2v_reg,valid_v_r_1_sv2v_reg,
  valid_v_r_0_sv2v_reg,lock_v_r_3_sv2v_reg,lock_v_r_2_sv2v_reg,lock_v_r_1_sv2v_reg,
  lock_v_r_0_sv2v_reg,tag_v_r_71_sv2v_reg,tag_v_r_70_sv2v_reg,tag_v_r_69_sv2v_reg,
  tag_v_r_68_sv2v_reg,tag_v_r_67_sv2v_reg,tag_v_r_66_sv2v_reg,tag_v_r_65_sv2v_reg,
  tag_v_r_64_sv2v_reg,tag_v_r_63_sv2v_reg,tag_v_r_62_sv2v_reg,tag_v_r_61_sv2v_reg,
  tag_v_r_60_sv2v_reg,tag_v_r_59_sv2v_reg,tag_v_r_58_sv2v_reg,tag_v_r_57_sv2v_reg,
  tag_v_r_56_sv2v_reg,tag_v_r_55_sv2v_reg,tag_v_r_54_sv2v_reg,tag_v_r_53_sv2v_reg,
  tag_v_r_52_sv2v_reg,tag_v_r_51_sv2v_reg,tag_v_r_50_sv2v_reg,tag_v_r_49_sv2v_reg,
  tag_v_r_48_sv2v_reg,tag_v_r_47_sv2v_reg,tag_v_r_46_sv2v_reg,tag_v_r_45_sv2v_reg,
  tag_v_r_44_sv2v_reg,tag_v_r_43_sv2v_reg,tag_v_r_42_sv2v_reg,tag_v_r_41_sv2v_reg,
  tag_v_r_40_sv2v_reg,tag_v_r_39_sv2v_reg,tag_v_r_38_sv2v_reg,tag_v_r_37_sv2v_reg,
  tag_v_r_36_sv2v_reg,tag_v_r_35_sv2v_reg,tag_v_r_34_sv2v_reg,tag_v_r_33_sv2v_reg,
  tag_v_r_32_sv2v_reg,tag_v_r_31_sv2v_reg,tag_v_r_30_sv2v_reg,tag_v_r_29_sv2v_reg,
  tag_v_r_28_sv2v_reg,tag_v_r_27_sv2v_reg,tag_v_r_26_sv2v_reg,tag_v_r_25_sv2v_reg,
  tag_v_r_24_sv2v_reg,tag_v_r_23_sv2v_reg,tag_v_r_22_sv2v_reg,tag_v_r_21_sv2v_reg,
  tag_v_r_20_sv2v_reg,tag_v_r_19_sv2v_reg,tag_v_r_18_sv2v_reg,tag_v_r_17_sv2v_reg,
  tag_v_r_16_sv2v_reg,tag_v_r_15_sv2v_reg,tag_v_r_14_sv2v_reg,tag_v_r_13_sv2v_reg,
  tag_v_r_12_sv2v_reg,tag_v_r_11_sv2v_reg,tag_v_r_10_sv2v_reg,tag_v_r_9_sv2v_reg,
  tag_v_r_8_sv2v_reg,tag_v_r_7_sv2v_reg,tag_v_r_6_sv2v_reg,tag_v_r_5_sv2v_reg,
  tag_v_r_4_sv2v_reg,tag_v_r_3_sv2v_reg,tag_v_r_2_sv2v_reg,tag_v_r_1_sv2v_reg,
  tag_v_r_0_sv2v_reg;
  assign data_tl_r[31] = data_tl_r_31_sv2v_reg;
  assign data_tl_r[30] = data_tl_r_30_sv2v_reg;
  assign data_tl_r[29] = data_tl_r_29_sv2v_reg;
  assign data_tl_r[28] = data_tl_r_28_sv2v_reg;
  assign data_tl_r[27] = data_tl_r_27_sv2v_reg;
  assign data_tl_r[26] = data_tl_r_26_sv2v_reg;
  assign data_tl_r[25] = data_tl_r_25_sv2v_reg;
  assign data_tl_r[24] = data_tl_r_24_sv2v_reg;
  assign data_tl_r[23] = data_tl_r_23_sv2v_reg;
  assign data_tl_r[22] = data_tl_r_22_sv2v_reg;
  assign data_tl_r[21] = data_tl_r_21_sv2v_reg;
  assign data_tl_r[20] = data_tl_r_20_sv2v_reg;
  assign data_tl_r[19] = data_tl_r_19_sv2v_reg;
  assign data_tl_r[18] = data_tl_r_18_sv2v_reg;
  assign data_tl_r[17] = data_tl_r_17_sv2v_reg;
  assign data_tl_r[16] = data_tl_r_16_sv2v_reg;
  assign data_tl_r[15] = data_tl_r_15_sv2v_reg;
  assign data_tl_r[14] = data_tl_r_14_sv2v_reg;
  assign data_tl_r[13] = data_tl_r_13_sv2v_reg;
  assign data_tl_r[12] = data_tl_r_12_sv2v_reg;
  assign data_tl_r[11] = data_tl_r_11_sv2v_reg;
  assign data_tl_r[10] = data_tl_r_10_sv2v_reg;
  assign data_tl_r[9] = data_tl_r_9_sv2v_reg;
  assign data_tl_r[8] = data_tl_r_8_sv2v_reg;
  assign data_tl_r[7] = data_tl_r_7_sv2v_reg;
  assign data_tl_r[6] = data_tl_r_6_sv2v_reg;
  assign data_tl_r[5] = data_tl_r_5_sv2v_reg;
  assign data_tl_r[4] = data_tl_r_4_sv2v_reg;
  assign data_tl_r[3] = data_tl_r_3_sv2v_reg;
  assign data_tl_r[2] = data_tl_r_2_sv2v_reg;
  assign data_tl_r[1] = data_tl_r_1_sv2v_reg;
  assign data_tl_r[0] = data_tl_r_0_sv2v_reg;
  assign v_tl_r = v_tl_r_sv2v_reg;
  assign decode_tl_r[20] = decode_tl_r_20_sv2v_reg;
  assign decode_tl_r[19] = decode_tl_r_19_sv2v_reg;
  assign decode_tl_r[18] = decode_tl_r_18_sv2v_reg;
  assign decode_tl_r[17] = decode_tl_r_17_sv2v_reg;
  assign decode_tl_r[16] = decode_tl_r_16_sv2v_reg;
  assign decode_tl_r[15] = decode_tl_r_15_sv2v_reg;
  assign decode_tl_r[14] = decode_tl_r_14_sv2v_reg;
  assign decode_tl_r[13] = decode_tl_r_13_sv2v_reg;
  assign decode_tl_r[12] = decode_tl_r_12_sv2v_reg;
  assign decode_tl_r[11] = decode_tl_r_11_sv2v_reg;
  assign decode_tl_r[10] = decode_tl_r_10_sv2v_reg;
  assign decode_tl_r[9] = decode_tl_r_9_sv2v_reg;
  assign decode_tl_r[8] = decode_tl_r_8_sv2v_reg;
  assign decode_tl_r[7] = decode_tl_r_7_sv2v_reg;
  assign decode_tl_r[6] = decode_tl_r_6_sv2v_reg;
  assign decode_tl_r[5] = decode_tl_r_5_sv2v_reg;
  assign decode_tl_r[4] = decode_tl_r_4_sv2v_reg;
  assign decode_tl_r[3] = decode_tl_r_3_sv2v_reg;
  assign decode_tl_r[2] = decode_tl_r_2_sv2v_reg;
  assign decode_tl_r[1] = decode_tl_r_1_sv2v_reg;
  assign decode_tl_r[0] = decode_tl_r_0_sv2v_reg;
  assign mask_tl_r[3] = mask_tl_r_3_sv2v_reg;
  assign mask_tl_r[2] = mask_tl_r_2_sv2v_reg;
  assign mask_tl_r[1] = mask_tl_r_1_sv2v_reg;
  assign mask_tl_r[0] = mask_tl_r_0_sv2v_reg;
  assign addr_tl_r[27] = addr_tl_r_27_sv2v_reg;
  assign addr_tl_r[26] = addr_tl_r_26_sv2v_reg;
  assign addr_tl_r[25] = addr_tl_r_25_sv2v_reg;
  assign addr_tl_r[24] = addr_tl_r_24_sv2v_reg;
  assign addr_tl_r[23] = addr_tl_r_23_sv2v_reg;
  assign addr_tl_r[22] = addr_tl_r_22_sv2v_reg;
  assign addr_tl_r[21] = addr_tl_r_21_sv2v_reg;
  assign addr_tl_r[20] = addr_tl_r_20_sv2v_reg;
  assign addr_tl_r[19] = addr_tl_r_19_sv2v_reg;
  assign addr_tl_r[18] = addr_tl_r_18_sv2v_reg;
  assign addr_tl_r[17] = addr_tl_r_17_sv2v_reg;
  assign addr_tl_r[16] = addr_tl_r_16_sv2v_reg;
  assign addr_tl_r[15] = addr_tl_r_15_sv2v_reg;
  assign addr_tl_r[14] = addr_tl_r_14_sv2v_reg;
  assign addr_tl_r[13] = addr_tl_r_13_sv2v_reg;
  assign addr_tl_r[12] = addr_tl_r_12_sv2v_reg;
  assign addr_tl_r[11] = addr_tl_r_11_sv2v_reg;
  assign addr_tl_r[10] = addr_tl_r_10_sv2v_reg;
  assign addr_tl_r[9] = addr_tl_r_9_sv2v_reg;
  assign addr_tl_r[8] = addr_tl_r_8_sv2v_reg;
  assign addr_tl_r[7] = addr_tl_r_7_sv2v_reg;
  assign addr_tl_r[6] = addr_tl_r_6_sv2v_reg;
  assign addr_tl_r[5] = addr_tl_r_5_sv2v_reg;
  assign addr_tl_r[4] = addr_tl_r_4_sv2v_reg;
  assign addr_tl_r[3] = addr_tl_r_3_sv2v_reg;
  assign addr_tl_r[2] = addr_tl_r_2_sv2v_reg;
  assign addr_tl_r[1] = addr_tl_r_1_sv2v_reg;
  assign addr_tl_r[0] = addr_tl_r_0_sv2v_reg;
  assign ld_data_v_r[127] = ld_data_v_r_127_sv2v_reg;
  assign ld_data_v_r[126] = ld_data_v_r_126_sv2v_reg;
  assign ld_data_v_r[125] = ld_data_v_r_125_sv2v_reg;
  assign ld_data_v_r[124] = ld_data_v_r_124_sv2v_reg;
  assign ld_data_v_r[123] = ld_data_v_r_123_sv2v_reg;
  assign ld_data_v_r[122] = ld_data_v_r_122_sv2v_reg;
  assign ld_data_v_r[121] = ld_data_v_r_121_sv2v_reg;
  assign ld_data_v_r[120] = ld_data_v_r_120_sv2v_reg;
  assign ld_data_v_r[119] = ld_data_v_r_119_sv2v_reg;
  assign ld_data_v_r[118] = ld_data_v_r_118_sv2v_reg;
  assign ld_data_v_r[117] = ld_data_v_r_117_sv2v_reg;
  assign ld_data_v_r[116] = ld_data_v_r_116_sv2v_reg;
  assign ld_data_v_r[115] = ld_data_v_r_115_sv2v_reg;
  assign ld_data_v_r[114] = ld_data_v_r_114_sv2v_reg;
  assign ld_data_v_r[113] = ld_data_v_r_113_sv2v_reg;
  assign ld_data_v_r[112] = ld_data_v_r_112_sv2v_reg;
  assign ld_data_v_r[111] = ld_data_v_r_111_sv2v_reg;
  assign ld_data_v_r[110] = ld_data_v_r_110_sv2v_reg;
  assign ld_data_v_r[109] = ld_data_v_r_109_sv2v_reg;
  assign ld_data_v_r[108] = ld_data_v_r_108_sv2v_reg;
  assign ld_data_v_r[107] = ld_data_v_r_107_sv2v_reg;
  assign ld_data_v_r[106] = ld_data_v_r_106_sv2v_reg;
  assign ld_data_v_r[105] = ld_data_v_r_105_sv2v_reg;
  assign ld_data_v_r[104] = ld_data_v_r_104_sv2v_reg;
  assign ld_data_v_r[103] = ld_data_v_r_103_sv2v_reg;
  assign ld_data_v_r[102] = ld_data_v_r_102_sv2v_reg;
  assign ld_data_v_r[101] = ld_data_v_r_101_sv2v_reg;
  assign ld_data_v_r[100] = ld_data_v_r_100_sv2v_reg;
  assign ld_data_v_r[99] = ld_data_v_r_99_sv2v_reg;
  assign ld_data_v_r[98] = ld_data_v_r_98_sv2v_reg;
  assign ld_data_v_r[97] = ld_data_v_r_97_sv2v_reg;
  assign ld_data_v_r[96] = ld_data_v_r_96_sv2v_reg;
  assign ld_data_v_r[95] = ld_data_v_r_95_sv2v_reg;
  assign ld_data_v_r[94] = ld_data_v_r_94_sv2v_reg;
  assign ld_data_v_r[93] = ld_data_v_r_93_sv2v_reg;
  assign ld_data_v_r[92] = ld_data_v_r_92_sv2v_reg;
  assign ld_data_v_r[91] = ld_data_v_r_91_sv2v_reg;
  assign ld_data_v_r[90] = ld_data_v_r_90_sv2v_reg;
  assign ld_data_v_r[89] = ld_data_v_r_89_sv2v_reg;
  assign ld_data_v_r[88] = ld_data_v_r_88_sv2v_reg;
  assign ld_data_v_r[87] = ld_data_v_r_87_sv2v_reg;
  assign ld_data_v_r[86] = ld_data_v_r_86_sv2v_reg;
  assign ld_data_v_r[85] = ld_data_v_r_85_sv2v_reg;
  assign ld_data_v_r[84] = ld_data_v_r_84_sv2v_reg;
  assign ld_data_v_r[83] = ld_data_v_r_83_sv2v_reg;
  assign ld_data_v_r[82] = ld_data_v_r_82_sv2v_reg;
  assign ld_data_v_r[81] = ld_data_v_r_81_sv2v_reg;
  assign ld_data_v_r[80] = ld_data_v_r_80_sv2v_reg;
  assign ld_data_v_r[79] = ld_data_v_r_79_sv2v_reg;
  assign ld_data_v_r[78] = ld_data_v_r_78_sv2v_reg;
  assign ld_data_v_r[77] = ld_data_v_r_77_sv2v_reg;
  assign ld_data_v_r[76] = ld_data_v_r_76_sv2v_reg;
  assign ld_data_v_r[75] = ld_data_v_r_75_sv2v_reg;
  assign ld_data_v_r[74] = ld_data_v_r_74_sv2v_reg;
  assign ld_data_v_r[73] = ld_data_v_r_73_sv2v_reg;
  assign ld_data_v_r[72] = ld_data_v_r_72_sv2v_reg;
  assign ld_data_v_r[71] = ld_data_v_r_71_sv2v_reg;
  assign ld_data_v_r[70] = ld_data_v_r_70_sv2v_reg;
  assign ld_data_v_r[69] = ld_data_v_r_69_sv2v_reg;
  assign ld_data_v_r[68] = ld_data_v_r_68_sv2v_reg;
  assign ld_data_v_r[67] = ld_data_v_r_67_sv2v_reg;
  assign ld_data_v_r[66] = ld_data_v_r_66_sv2v_reg;
  assign ld_data_v_r[65] = ld_data_v_r_65_sv2v_reg;
  assign ld_data_v_r[64] = ld_data_v_r_64_sv2v_reg;
  assign ld_data_v_r[63] = ld_data_v_r_63_sv2v_reg;
  assign ld_data_v_r[62] = ld_data_v_r_62_sv2v_reg;
  assign ld_data_v_r[61] = ld_data_v_r_61_sv2v_reg;
  assign ld_data_v_r[60] = ld_data_v_r_60_sv2v_reg;
  assign ld_data_v_r[59] = ld_data_v_r_59_sv2v_reg;
  assign ld_data_v_r[58] = ld_data_v_r_58_sv2v_reg;
  assign ld_data_v_r[57] = ld_data_v_r_57_sv2v_reg;
  assign ld_data_v_r[56] = ld_data_v_r_56_sv2v_reg;
  assign ld_data_v_r[55] = ld_data_v_r_55_sv2v_reg;
  assign ld_data_v_r[54] = ld_data_v_r_54_sv2v_reg;
  assign ld_data_v_r[53] = ld_data_v_r_53_sv2v_reg;
  assign ld_data_v_r[52] = ld_data_v_r_52_sv2v_reg;
  assign ld_data_v_r[51] = ld_data_v_r_51_sv2v_reg;
  assign ld_data_v_r[50] = ld_data_v_r_50_sv2v_reg;
  assign ld_data_v_r[49] = ld_data_v_r_49_sv2v_reg;
  assign ld_data_v_r[48] = ld_data_v_r_48_sv2v_reg;
  assign ld_data_v_r[47] = ld_data_v_r_47_sv2v_reg;
  assign ld_data_v_r[46] = ld_data_v_r_46_sv2v_reg;
  assign ld_data_v_r[45] = ld_data_v_r_45_sv2v_reg;
  assign ld_data_v_r[44] = ld_data_v_r_44_sv2v_reg;
  assign ld_data_v_r[43] = ld_data_v_r_43_sv2v_reg;
  assign ld_data_v_r[42] = ld_data_v_r_42_sv2v_reg;
  assign ld_data_v_r[41] = ld_data_v_r_41_sv2v_reg;
  assign ld_data_v_r[40] = ld_data_v_r_40_sv2v_reg;
  assign ld_data_v_r[39] = ld_data_v_r_39_sv2v_reg;
  assign ld_data_v_r[38] = ld_data_v_r_38_sv2v_reg;
  assign ld_data_v_r[37] = ld_data_v_r_37_sv2v_reg;
  assign ld_data_v_r[36] = ld_data_v_r_36_sv2v_reg;
  assign ld_data_v_r[35] = ld_data_v_r_35_sv2v_reg;
  assign ld_data_v_r[34] = ld_data_v_r_34_sv2v_reg;
  assign ld_data_v_r[33] = ld_data_v_r_33_sv2v_reg;
  assign ld_data_v_r[32] = ld_data_v_r_32_sv2v_reg;
  assign ld_data_v_r[31] = ld_data_v_r_31_sv2v_reg;
  assign ld_data_v_r[30] = ld_data_v_r_30_sv2v_reg;
  assign ld_data_v_r[29] = ld_data_v_r_29_sv2v_reg;
  assign ld_data_v_r[28] = ld_data_v_r_28_sv2v_reg;
  assign ld_data_v_r[27] = ld_data_v_r_27_sv2v_reg;
  assign ld_data_v_r[26] = ld_data_v_r_26_sv2v_reg;
  assign ld_data_v_r[25] = ld_data_v_r_25_sv2v_reg;
  assign ld_data_v_r[24] = ld_data_v_r_24_sv2v_reg;
  assign ld_data_v_r[23] = ld_data_v_r_23_sv2v_reg;
  assign ld_data_v_r[22] = ld_data_v_r_22_sv2v_reg;
  assign ld_data_v_r[21] = ld_data_v_r_21_sv2v_reg;
  assign ld_data_v_r[20] = ld_data_v_r_20_sv2v_reg;
  assign ld_data_v_r[19] = ld_data_v_r_19_sv2v_reg;
  assign ld_data_v_r[18] = ld_data_v_r_18_sv2v_reg;
  assign ld_data_v_r[17] = ld_data_v_r_17_sv2v_reg;
  assign ld_data_v_r[16] = ld_data_v_r_16_sv2v_reg;
  assign ld_data_v_r[15] = ld_data_v_r_15_sv2v_reg;
  assign ld_data_v_r[14] = ld_data_v_r_14_sv2v_reg;
  assign ld_data_v_r[13] = ld_data_v_r_13_sv2v_reg;
  assign ld_data_v_r[12] = ld_data_v_r_12_sv2v_reg;
  assign ld_data_v_r[11] = ld_data_v_r_11_sv2v_reg;
  assign ld_data_v_r[10] = ld_data_v_r_10_sv2v_reg;
  assign ld_data_v_r[9] = ld_data_v_r_9_sv2v_reg;
  assign ld_data_v_r[8] = ld_data_v_r_8_sv2v_reg;
  assign ld_data_v_r[7] = ld_data_v_r_7_sv2v_reg;
  assign ld_data_v_r[6] = ld_data_v_r_6_sv2v_reg;
  assign ld_data_v_r[5] = ld_data_v_r_5_sv2v_reg;
  assign ld_data_v_r[4] = ld_data_v_r_4_sv2v_reg;
  assign ld_data_v_r[3] = ld_data_v_r_3_sv2v_reg;
  assign ld_data_v_r[2] = ld_data_v_r_2_sv2v_reg;
  assign ld_data_v_r[1] = ld_data_v_r_1_sv2v_reg;
  assign ld_data_v_r[0] = ld_data_v_r_0_sv2v_reg;
  assign v_v_r = v_v_r_sv2v_reg;
  assign track_data_v_r[15] = track_data_v_r_15_sv2v_reg;
  assign track_data_v_r[14] = track_data_v_r_14_sv2v_reg;
  assign track_data_v_r[13] = track_data_v_r_13_sv2v_reg;
  assign track_data_v_r[12] = track_data_v_r_12_sv2v_reg;
  assign track_data_v_r[11] = track_data_v_r_11_sv2v_reg;
  assign track_data_v_r[10] = track_data_v_r_10_sv2v_reg;
  assign track_data_v_r[9] = track_data_v_r_9_sv2v_reg;
  assign track_data_v_r[8] = track_data_v_r_8_sv2v_reg;
  assign track_data_v_r[7] = track_data_v_r_7_sv2v_reg;
  assign track_data_v_r[6] = track_data_v_r_6_sv2v_reg;
  assign track_data_v_r[5] = track_data_v_r_5_sv2v_reg;
  assign track_data_v_r[4] = track_data_v_r_4_sv2v_reg;
  assign track_data_v_r[3] = track_data_v_r_3_sv2v_reg;
  assign track_data_v_r[2] = track_data_v_r_2_sv2v_reg;
  assign track_data_v_r[1] = track_data_v_r_1_sv2v_reg;
  assign track_data_v_r[0] = track_data_v_r_0_sv2v_reg;
  assign mask_v_r[3] = mask_v_r_3_sv2v_reg;
  assign mask_v_r[2] = mask_v_r_2_sv2v_reg;
  assign mask_v_r[1] = mask_v_r_1_sv2v_reg;
  assign mask_v_r[0] = mask_v_r_0_sv2v_reg;
  assign decode_v_r[20] = decode_v_r_20_sv2v_reg;
  assign decode_v_r[19] = decode_v_r_19_sv2v_reg;
  assign decode_v_r[18] = decode_v_r_18_sv2v_reg;
  assign decode_v_r[17] = decode_v_r_17_sv2v_reg;
  assign decode_v_r[16] = decode_v_r_16_sv2v_reg;
  assign decode_v_r[15] = decode_v_r_15_sv2v_reg;
  assign decode_v_r[14] = decode_v_r_14_sv2v_reg;
  assign decode_v_r[13] = decode_v_r_13_sv2v_reg;
  assign decode_v_r[12] = decode_v_r_12_sv2v_reg;
  assign decode_v_r[11] = decode_v_r_11_sv2v_reg;
  assign decode_v_r[10] = decode_v_r_10_sv2v_reg;
  assign decode_v_r[9] = decode_v_r_9_sv2v_reg;
  assign decode_v_r[8] = decode_v_r_8_sv2v_reg;
  assign decode_v_r[7] = decode_v_r_7_sv2v_reg;
  assign decode_v_r[6] = decode_v_r_6_sv2v_reg;
  assign decode_v_r[5] = decode_v_r_5_sv2v_reg;
  assign decode_v_r[4] = decode_v_r_4_sv2v_reg;
  assign decode_v_r[3] = decode_v_r_3_sv2v_reg;
  assign decode_v_r[2] = decode_v_r_2_sv2v_reg;
  assign decode_v_r[1] = decode_v_r_1_sv2v_reg;
  assign decode_v_r[0] = decode_v_r_0_sv2v_reg;
  assign addr_v_r[27] = addr_v_r_27_sv2v_reg;
  assign addr_v_r[26] = addr_v_r_26_sv2v_reg;
  assign addr_v_r[25] = addr_v_r_25_sv2v_reg;
  assign addr_v_r[24] = addr_v_r_24_sv2v_reg;
  assign addr_v_r[23] = addr_v_r_23_sv2v_reg;
  assign addr_v_r[22] = addr_v_r_22_sv2v_reg;
  assign addr_v_r[21] = addr_v_r_21_sv2v_reg;
  assign addr_v_r[20] = addr_v_r_20_sv2v_reg;
  assign addr_v_r[19] = addr_v_r_19_sv2v_reg;
  assign addr_v_r[18] = addr_v_r_18_sv2v_reg;
  assign addr_v_r[17] = addr_v_r_17_sv2v_reg;
  assign addr_v_r[16] = addr_v_r_16_sv2v_reg;
  assign addr_v_r[15] = addr_v_r_15_sv2v_reg;
  assign addr_v_r[14] = addr_v_r_14_sv2v_reg;
  assign addr_v_r[13] = addr_v_r_13_sv2v_reg;
  assign addr_v_r[12] = addr_v_r_12_sv2v_reg;
  assign addr_v_r[11] = addr_v_r_11_sv2v_reg;
  assign addr_v_r[10] = addr_v_r_10_sv2v_reg;
  assign addr_v_r[9] = addr_v_r_9_sv2v_reg;
  assign addr_v_r[8] = addr_v_r_8_sv2v_reg;
  assign addr_v_r[7] = addr_v_r_7_sv2v_reg;
  assign addr_v_r[6] = addr_v_r_6_sv2v_reg;
  assign addr_v_r[5] = addr_v_r_5_sv2v_reg;
  assign addr_v_r[4] = addr_v_r_4_sv2v_reg;
  assign addr_v_r[3] = addr_v_r_3_sv2v_reg;
  assign addr_v_r[2] = addr_v_r_2_sv2v_reg;
  assign addr_v_r[1] = addr_v_r_1_sv2v_reg;
  assign addr_v_r[0] = addr_v_r_0_sv2v_reg;
  assign data_v_r[31] = data_v_r_31_sv2v_reg;
  assign data_v_r[30] = data_v_r_30_sv2v_reg;
  assign data_v_r[29] = data_v_r_29_sv2v_reg;
  assign data_v_r[28] = data_v_r_28_sv2v_reg;
  assign data_v_r[27] = data_v_r_27_sv2v_reg;
  assign data_v_r[26] = data_v_r_26_sv2v_reg;
  assign data_v_r[25] = data_v_r_25_sv2v_reg;
  assign data_v_r[24] = data_v_r_24_sv2v_reg;
  assign data_v_r[23] = data_v_r_23_sv2v_reg;
  assign data_v_r[22] = data_v_r_22_sv2v_reg;
  assign data_v_r[21] = data_v_r_21_sv2v_reg;
  assign data_v_r[20] = data_v_r_20_sv2v_reg;
  assign data_v_r[19] = data_v_r_19_sv2v_reg;
  assign data_v_r[18] = data_v_r_18_sv2v_reg;
  assign data_v_r[17] = data_v_r_17_sv2v_reg;
  assign data_v_r[16] = data_v_r_16_sv2v_reg;
  assign data_v_r[15] = data_v_r_15_sv2v_reg;
  assign data_v_r[14] = data_v_r_14_sv2v_reg;
  assign data_v_r[13] = data_v_r_13_sv2v_reg;
  assign data_v_r[12] = data_v_r_12_sv2v_reg;
  assign data_v_r[11] = data_v_r_11_sv2v_reg;
  assign data_v_r[10] = data_v_r_10_sv2v_reg;
  assign data_v_r[9] = data_v_r_9_sv2v_reg;
  assign data_v_r[8] = data_v_r_8_sv2v_reg;
  assign data_v_r[7] = data_v_r_7_sv2v_reg;
  assign data_v_r[6] = data_v_r_6_sv2v_reg;
  assign data_v_r[5] = data_v_r_5_sv2v_reg;
  assign data_v_r[4] = data_v_r_4_sv2v_reg;
  assign data_v_r[3] = data_v_r_3_sv2v_reg;
  assign data_v_r[2] = data_v_r_2_sv2v_reg;
  assign data_v_r[1] = data_v_r_1_sv2v_reg;
  assign data_v_r[0] = data_v_r_0_sv2v_reg;
  assign valid_v_r[3] = valid_v_r_3_sv2v_reg;
  assign valid_v_r[2] = valid_v_r_2_sv2v_reg;
  assign valid_v_r[1] = valid_v_r_1_sv2v_reg;
  assign valid_v_r[0] = valid_v_r_0_sv2v_reg;
  assign lock_v_r[3] = lock_v_r_3_sv2v_reg;
  assign lock_v_r[2] = lock_v_r_2_sv2v_reg;
  assign lock_v_r[1] = lock_v_r_1_sv2v_reg;
  assign lock_v_r[0] = lock_v_r_0_sv2v_reg;
  assign tag_v_r[71] = tag_v_r_71_sv2v_reg;
  assign tag_v_r[70] = tag_v_r_70_sv2v_reg;
  assign tag_v_r[69] = tag_v_r_69_sv2v_reg;
  assign tag_v_r[68] = tag_v_r_68_sv2v_reg;
  assign tag_v_r[67] = tag_v_r_67_sv2v_reg;
  assign tag_v_r[66] = tag_v_r_66_sv2v_reg;
  assign tag_v_r[65] = tag_v_r_65_sv2v_reg;
  assign tag_v_r[64] = tag_v_r_64_sv2v_reg;
  assign tag_v_r[63] = tag_v_r_63_sv2v_reg;
  assign tag_v_r[62] = tag_v_r_62_sv2v_reg;
  assign tag_v_r[61] = tag_v_r_61_sv2v_reg;
  assign tag_v_r[60] = tag_v_r_60_sv2v_reg;
  assign tag_v_r[59] = tag_v_r_59_sv2v_reg;
  assign tag_v_r[58] = tag_v_r_58_sv2v_reg;
  assign tag_v_r[57] = tag_v_r_57_sv2v_reg;
  assign tag_v_r[56] = tag_v_r_56_sv2v_reg;
  assign tag_v_r[55] = tag_v_r_55_sv2v_reg;
  assign tag_v_r[54] = tag_v_r_54_sv2v_reg;
  assign tag_v_r[53] = tag_v_r_53_sv2v_reg;
  assign tag_v_r[52] = tag_v_r_52_sv2v_reg;
  assign tag_v_r[51] = tag_v_r_51_sv2v_reg;
  assign tag_v_r[50] = tag_v_r_50_sv2v_reg;
  assign tag_v_r[49] = tag_v_r_49_sv2v_reg;
  assign tag_v_r[48] = tag_v_r_48_sv2v_reg;
  assign tag_v_r[47] = tag_v_r_47_sv2v_reg;
  assign tag_v_r[46] = tag_v_r_46_sv2v_reg;
  assign tag_v_r[45] = tag_v_r_45_sv2v_reg;
  assign tag_v_r[44] = tag_v_r_44_sv2v_reg;
  assign tag_v_r[43] = tag_v_r_43_sv2v_reg;
  assign tag_v_r[42] = tag_v_r_42_sv2v_reg;
  assign tag_v_r[41] = tag_v_r_41_sv2v_reg;
  assign tag_v_r[40] = tag_v_r_40_sv2v_reg;
  assign tag_v_r[39] = tag_v_r_39_sv2v_reg;
  assign tag_v_r[38] = tag_v_r_38_sv2v_reg;
  assign tag_v_r[37] = tag_v_r_37_sv2v_reg;
  assign tag_v_r[36] = tag_v_r_36_sv2v_reg;
  assign tag_v_r[35] = tag_v_r_35_sv2v_reg;
  assign tag_v_r[34] = tag_v_r_34_sv2v_reg;
  assign tag_v_r[33] = tag_v_r_33_sv2v_reg;
  assign tag_v_r[32] = tag_v_r_32_sv2v_reg;
  assign tag_v_r[31] = tag_v_r_31_sv2v_reg;
  assign tag_v_r[30] = tag_v_r_30_sv2v_reg;
  assign tag_v_r[29] = tag_v_r_29_sv2v_reg;
  assign tag_v_r[28] = tag_v_r_28_sv2v_reg;
  assign tag_v_r[27] = tag_v_r_27_sv2v_reg;
  assign tag_v_r[26] = tag_v_r_26_sv2v_reg;
  assign tag_v_r[25] = tag_v_r_25_sv2v_reg;
  assign tag_v_r[24] = tag_v_r_24_sv2v_reg;
  assign tag_v_r[23] = tag_v_r_23_sv2v_reg;
  assign tag_v_r[22] = tag_v_r_22_sv2v_reg;
  assign tag_v_r[21] = tag_v_r_21_sv2v_reg;
  assign tag_v_r[20] = tag_v_r_20_sv2v_reg;
  assign tag_v_r[19] = tag_v_r_19_sv2v_reg;
  assign tag_v_r[18] = tag_v_r_18_sv2v_reg;
  assign tag_v_r[17] = tag_v_r_17_sv2v_reg;
  assign tag_v_r[16] = tag_v_r_16_sv2v_reg;
  assign tag_v_r[15] = tag_v_r_15_sv2v_reg;
  assign tag_v_r[14] = tag_v_r_14_sv2v_reg;
  assign tag_v_r[13] = tag_v_r_13_sv2v_reg;
  assign tag_v_r[12] = tag_v_r_12_sv2v_reg;
  assign tag_v_r[11] = tag_v_r_11_sv2v_reg;
  assign tag_v_r[10] = tag_v_r_10_sv2v_reg;
  assign tag_v_r[9] = tag_v_r_9_sv2v_reg;
  assign tag_v_r[8] = tag_v_r_8_sv2v_reg;
  assign tag_v_r[7] = tag_v_r_7_sv2v_reg;
  assign tag_v_r[6] = tag_v_r_6_sv2v_reg;
  assign tag_v_r[5] = tag_v_r_5_sv2v_reg;
  assign tag_v_r[4] = tag_v_r_4_sv2v_reg;
  assign tag_v_r[3] = tag_v_r_3_sv2v_reg;
  assign tag_v_r[2] = tag_v_r_2_sv2v_reg;
  assign tag_v_r[1] = tag_v_r_1_sv2v_reg;
  assign tag_v_r[0] = tag_v_r_0_sv2v_reg;

  bsg_cache_decode
  decode0
  (
    .opcode_i(cache_pkt_i[69:64]),
    .decode_o(decode)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p80_els_p64_latch_last_read_p1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p128_latch_last_read_p1
  data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li),
    .data_i(data_mem_data_li),
    .write_mask_i(data_mem_w_mask_li),
    .data_o(data_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p16_els_p64_latch_last_read_p1
  \track_mem_gen.track_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(track_mem_data_li),
    .addr_i(track_mem_addr_li),
    .v_i(track_mem_v_li),
    .w_mask_i(track_mem_w_mask_li),
    .w_i(track_mem_w_li),
    .data_o(track_mem_data_lo)
  );

  assign N86 = addr_v_r[27:10] == tag_v_r[17:0];
  assign N87 = addr_v_r[27:10] == tag_v_r[35:18];
  assign N88 = addr_v_r[27:10] == tag_v_r[53:36];
  assign N89 = addr_v_r[27:10] == tag_v_r[71:54];

  bsg_priority_encode_width_p4_lo_to_hi_p1
  tag_hit_pe
  (
    .i(tag_hit_v),
    .addr_o(tag_hit_way_id),
    .v_o(tag_hit_found)
  );

  assign N109 = (N105)? track_data_v_r[3] : 
                (N107)? track_data_v_r[7] : 
                (N106)? track_data_v_r[11] : 
                (N108)? track_data_v_r[15] : 1'b0;
  assign N110 = (N105)? track_data_v_r[2] : 
                (N107)? track_data_v_r[6] : 
                (N106)? track_data_v_r[10] : 
                (N108)? track_data_v_r[14] : 1'b0;
  assign N111 = (N105)? track_data_v_r[1] : 
                (N107)? track_data_v_r[5] : 
                (N106)? track_data_v_r[9] : 
                (N108)? track_data_v_r[13] : 1'b0;
  assign N112 = (N105)? track_data_v_r[0] : 
                (N107)? track_data_v_r[4] : 
                (N106)? track_data_v_r[8] : 
                (N108)? track_data_v_r[12] : 1'b0;
  assign N119 = (N115)? N112 : 
                (N117)? N111 : 
                (N116)? N110 : 
                (N118)? N109 : 1'b0;
  assign N126 = (N122)? valid_v_r[0] : 
                (N124)? valid_v_r[1] : 
                (N123)? valid_v_r[2] : 
                (N125)? valid_v_r[3] : 1'b0;
  assign N135 = (N131)? lock_v_r[0] : 
                (N133)? lock_v_r[1] : 
                (N132)? lock_v_r[2] : 
                (N134)? lock_v_r[3] : 1'b0;
  assign N146 = (N142)? lock_v_r[0] : 
                (N144)? lock_v_r[1] : 
                (N143)? lock_v_r[2] : 
                (N145)? lock_v_r[3] : 1'b0;

  bsg_mem_1rw_sync_mask_write_bit_width_p7_els_p64_latch_last_read_p1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_w_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4_word_tracking_p1
  miss
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .miss_v_i(miss_v),
    .track_miss_i(track_miss),
    .decode_v_i(decode_v_r),
    .addr_v_i(addr_v_r),
    .mask_v_i(mask_v_r),
    .tag_v_i(tag_v_r),
    .valid_v_i(valid_v_r),
    .lock_v_i(lock_v_r),
    .tag_hit_v_i(tag_hit_v),
    .tag_hit_way_id_i(tag_hit_way_id),
    .tag_hit_found_i(tag_hit_found),
    .sbuf_empty_i(sbuf_empty_lo),
    .tbuf_empty_i(tbuf_empty_lo),
    .dma_cmd_o(dma_cmd_lo),
    .dma_way_o(dma_way_lo),
    .dma_addr_o(dma_addr_lo),
    .dma_done_i(dma_done_li),
    .track_data_we_o(miss_track_data_we_lo),
    .stat_info_i(stat_mem_data_lo),
    .stat_mem_v_o(miss_stat_mem_v_lo),
    .stat_mem_w_o(miss_stat_mem_w_lo),
    .stat_mem_addr_o(miss_stat_mem_addr_lo),
    .stat_mem_data_o(miss_stat_mem_data_lo),
    .stat_mem_w_mask_o(miss_stat_mem_w_mask_lo),
    .tag_mem_v_o(miss_tag_mem_v_lo),
    .tag_mem_w_o(miss_tag_mem_w_lo),
    .tag_mem_addr_o(miss_tag_mem_addr_lo),
    .tag_mem_data_o(miss_tag_mem_data_lo),
    .tag_mem_w_mask_o(miss_tag_mem_w_mask_lo),
    .track_mem_v_o(miss_track_mem_v_lo),
    .track_mem_w_o(miss_track_mem_w_lo),
    .track_mem_addr_o(miss_track_mem_addr_lo),
    .track_mem_w_mask_o(miss_track_mem_w_mask_lo),
    .track_mem_data_o(miss_track_mem_data_lo),
    .done_o(miss_done_lo),
    .recover_o(recover_lo),
    .chosen_way_o(chosen_way_lo),
    .select_snoop_data_r_o(select_snoop_data_r_lo),
    .ack_i(_1_net_)
  );


  bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p4_word_tracking_p1_dma_data_width_p32_debug_p0
  dma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dma_cmd_i(dma_cmd_lo),
    .dma_way_i(dma_way_lo),
    .dma_addr_i(dma_addr_lo),
    .done_o(dma_done_li),
    .track_data_we_i(miss_track_data_we_lo),
    .snoop_word_o(snoop_word_lo),
    .dma_pkt_o(dma_pkt_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_i(dma_data_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_o(dma_data_o),
    .dma_data_v_o(dma_data_v_o),
    .dma_data_yumi_i(dma_data_yumi_i),
    .data_mem_v_o(dma_data_mem_v_lo),
    .data_mem_w_o(dma_data_mem_w_lo),
    .data_mem_addr_o(dma_data_mem_addr_lo),
    .data_mem_w_mask_o(dma_data_mem_w_mask_lo),
    .data_mem_data_o(dma_data_mem_data_lo),
    .data_mem_data_i(data_mem_data_lo),
    .track_miss_i(track_miss),
    .track_mem_data_i(track_mem_data_lo),
    .dma_evict_o(dma_evict_lo)
  );


  bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p4
  sbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .sbuf_entry_i({ addr_v_r, sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_, sbuf_entry_li_way_id__1_, sbuf_entry_li_way_id__0_ }),
    .v_i(sbuf_v_li),
    .sbuf_entry_o(sbuf_entry_lo),
    .v_o(sbuf_v_lo),
    .yumi_i(sbuf_yumi_li),
    .empty_o(sbuf_empty_lo),
    .full_o(sbuf_full_lo),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(sbuf_bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo)
  );


  bsg_decode_num_out_p4
  sbuf_way_demux
  (
    .i(sbuf_entry_lo[1:0]),
    .o(sbuf_way_decode)
  );


  bsg_decode_num_out_p1
  sbuf_bo_demux
  (
    .i(sbuf_entry_lo[40]),
    .o(sbuf_burst_offset_decode[0])
  );


  bsg_expand_bitmask
  expand0
  (
    .i(sbuf_burst_offset_decode[0]),
    .o(sbuf_expand_mask)
  );


  bsg_mux_width_p32_els_p3
  sbuf_data_in_mux
  (
    .data_i({ \sbuf_in_sel_2_.slice_data , data_v_r[15:0], data_v_r[15:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0] }),
    .sel_i(decode_v_r[20:19]),
    .data_o(sbuf_data_in)
  );


  bsg_mux_width_p4_els_p3
  sbuf_mask_in_mux
  (
    .data_i(sbuf_mask_in_mux_li),
    .sel_i(decode_v_r[20:19]),
    .data_o(sbuf_mask_in)
  );

  assign N170 = N169 | decode_v_r[3];
  assign N171 = decode_v_r[2] | decode_v_r[1];
  assign N172 = N170 | N171;
  assign N173 = N172 | decode_v_r[0];
  assign N177 = N169 | decode_v_r[3];
  assign N178 = decode_v_r[2] | N175;
  assign N179 = N177 | N178;
  assign N180 = N179 | N176;
  assign N183 = N169 | decode_v_r[3];
  assign N184 = N182 | decode_v_r[1];
  assign N185 = N183 | N184;
  assign N186 = N185 | decode_v_r[0];
  assign N189 = N169 | decode_v_r[3];
  assign N190 = decode_v_r[2] | N188;
  assign N191 = N189 | N190;
  assign N192 = N191 | decode_v_r[0];
  assign N195 = N169 | decode_v_r[3];
  assign N196 = decode_v_r[2] | decode_v_r[1];
  assign N197 = N195 | N196;
  assign N198 = N197 | N194;
  assign N202 = N169 | decode_v_r[3];
  assign N203 = N200 | decode_v_r[1];
  assign N204 = N202 | N203;
  assign N205 = N204 | N201;
  assign N209 = N169 | decode_v_r[3];
  assign N210 = N207 | N208;
  assign N211 = N209 | N210;
  assign N212 = N211 | decode_v_r[0];
  assign N217 = N169 | decode_v_r[3];
  assign N218 = N214 | N215;
  assign N219 = N217 | N218;
  assign N220 = N219 | N216;
  assign N223 = N169 | N222;
  assign N224 = decode_v_r[2] | decode_v_r[1];
  assign N225 = N223 | N224;
  assign N226 = N225 | decode_v_r[0];
  assign N228 = N168 & decode_v_r[3];
  assign N229 = N228 & decode_v_r[0];
  assign N230 = N168 & decode_v_r[3];
  assign N231 = N230 & decode_v_r[1];
  assign N232 = N168 & decode_v_r[3];
  assign N233 = N232 & decode_v_r[2];
  assign N363 = $signed(data_v_r) < $signed(atomic_mem_data);
  assign N397 = $signed(data_v_r) > $signed(atomic_mem_data);
  assign N431 = data_v_r < atomic_mem_data;
  assign N465 = data_v_r > atomic_mem_data;

  bsg_decode_num_out_p4
  \sbuf_in_sel_0_.dec 
  (
    .i(addr_v_r[1:0]),
    .o(\sbuf_in_sel_0_.decode_lo )
  );


  bsg_expand_bitmask
  \sbuf_in_sel_0_.exp 
  (
    .i(\sbuf_in_sel_0_.decode_lo ),
    .o(sbuf_mask_in_mux_li[3:0])
  );


  bsg_decode_num_out_p2
  \sbuf_in_sel_1_.dec 
  (
    .i(addr_v_r[1]),
    .o(\sbuf_in_sel_1_.decode_lo )
  );


  bsg_expand_bitmask
  \sbuf_in_sel_1_.exp 
  (
    .i(\sbuf_in_sel_1_.decode_lo ),
    .o(sbuf_mask_in_mux_li[7:4])
  );


  bsg_decode_num_out_p1
  \sbuf_in_sel_2_.dec 
  (
    .i(addr_v_r[2]),
    .o(\sbuf_in_sel_2_.decode_lo [0])
  );


  bsg_expand_bitmask
  \sbuf_in_sel_2_.exp 
  (
    .i(\sbuf_in_sel_2_.decode_lo [0]),
    .o(sbuf_mask_in_mux_li[11:8])
  );


  bsg_cache_tbuf
  \tbuf_gen.tbuf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .addr_i(addr_v_r),
    .way_i(tbuf_way_li),
    .v_i(tbuf_v_li),
    .addr_o(tbuf_addr_lo),
    .way_o(tbuf_way_lo),
    .v_o(tbuf_v_lo),
    .yumi_i(tbuf_yumi_li),
    .empty_o(tbuf_empty_lo),
    .full_o(tbuf_full_lo),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(tbuf_bypass_v_li),
    .bypass_track_o(bypass_track_lo)
  );


  bsg_decode_num_out_p4
  tbuf_way_demux
  (
    .i(tbuf_way_lo),
    .o(tbuf_way_decode)
  );


  bsg_decode_num_out_p4
  tbuf_wo_demux
  (
    .i(tbuf_addr_lo[3:2]),
    .o(tbuf_word_offset_decode)
  );


  bsg_mux_width_p32_els_p4
  ld_data_mux
  (
    .data_i(ld_data_v_r),
    .sel_i(tag_hit_way_id),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_width_p32_els_p1
  mux00
  (
    .data_i(ld_data_way_picked),
    .sel_i(addr_v_r[2]),
    .data_o(ld_data_offset_picked)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(ld_data_offset_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_expand_bitmask
  mask_v_expand
  (
    .i(mask_v_r),
    .o(expanded_mask_v)
  );


  bsg_mux_width_p8_els_p4
  \ld_data_sel_0_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1:0]),
    .data_o(\ld_data_sel_0_.byte_sel )
  );


  bsg_mux_width_p16_els_p2
  \ld_data_sel_1_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1]),
    .data_o(\ld_data_sel_1_.byte_sel )
  );


  bsg_mux_width_p32_els_p1
  \ld_data_sel_2_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[2]),
    .data_o(atomic_mem_data)
  );


  bsg_mux_width_p32_els_p3
  ld_data_size_mux
  (
    .data_i({ atomic_mem_data, ld_data_final_li_1__31_, ld_data_final_li_1__30_, ld_data_final_li_1__29_, ld_data_final_li_1__28_, ld_data_final_li_1__27_, ld_data_final_li_1__26_, ld_data_final_li_1__25_, ld_data_final_li_1__24_, ld_data_final_li_1__23_, ld_data_final_li_1__22_, ld_data_final_li_1__21_, ld_data_final_li_1__20_, ld_data_final_li_1__19_, ld_data_final_li_1__18_, ld_data_final_li_1__17_, ld_data_final_li_1__16_, \ld_data_sel_1_.byte_sel , ld_data_final_li_0__31_, ld_data_final_li_0__30_, ld_data_final_li_0__29_, ld_data_final_li_0__28_, ld_data_final_li_0__27_, ld_data_final_li_0__26_, ld_data_final_li_0__25_, ld_data_final_li_0__24_, ld_data_final_li_0__23_, ld_data_final_li_0__22_, ld_data_final_li_0__21_, ld_data_final_li_0__20_, ld_data_final_li_0__19_, ld_data_final_li_0__18_, ld_data_final_li_0__17_, ld_data_final_li_0__16_, ld_data_final_li_0__15_, ld_data_final_li_0__14_, ld_data_final_li_0__13_, ld_data_final_li_0__12_, ld_data_final_li_0__11_, ld_data_final_li_0__10_, ld_data_final_li_0__9_, ld_data_final_li_0__8_, \ld_data_sel_0_.byte_sel  }),
    .sel_i(decode_v_r[20:19]),
    .data_o(ld_data_final_lo)
  );

  assign N521 = (N517)? lock_v_r[0] : 
                (N519)? lock_v_r[1] : 
                (N518)? lock_v_r[2] : 
                (N520)? lock_v_r[3] : 1'b0;
  assign N528 = (N524)? valid_v_r[0] : 
                (N526)? valid_v_r[1] : 
                (N525)? valid_v_r[2] : 
                (N527)? valid_v_r[3] : 1'b0;
  assign N535 = (N531)? tag_v_r[17] : 
                (N533)? tag_v_r[35] : 
                (N532)? tag_v_r[53] : 
                (N534)? tag_v_r[71] : 1'b0;
  assign N536 = (N531)? tag_v_r[16] : 
                (N533)? tag_v_r[34] : 
                (N532)? tag_v_r[52] : 
                (N534)? tag_v_r[70] : 1'b0;
  assign N537 = (N531)? tag_v_r[15] : 
                (N533)? tag_v_r[33] : 
                (N532)? tag_v_r[51] : 
                (N534)? tag_v_r[69] : 1'b0;
  assign N538 = (N531)? tag_v_r[14] : 
                (N533)? tag_v_r[32] : 
                (N532)? tag_v_r[50] : 
                (N534)? tag_v_r[68] : 1'b0;
  assign N539 = (N531)? tag_v_r[13] : 
                (N533)? tag_v_r[31] : 
                (N532)? tag_v_r[49] : 
                (N534)? tag_v_r[67] : 1'b0;
  assign N540 = (N531)? tag_v_r[12] : 
                (N533)? tag_v_r[30] : 
                (N532)? tag_v_r[48] : 
                (N534)? tag_v_r[66] : 1'b0;
  assign N541 = (N531)? tag_v_r[11] : 
                (N533)? tag_v_r[29] : 
                (N532)? tag_v_r[47] : 
                (N534)? tag_v_r[65] : 1'b0;
  assign N542 = (N531)? tag_v_r[10] : 
                (N533)? tag_v_r[28] : 
                (N532)? tag_v_r[46] : 
                (N534)? tag_v_r[64] : 1'b0;
  assign N543 = (N531)? tag_v_r[9] : 
                (N533)? tag_v_r[27] : 
                (N532)? tag_v_r[45] : 
                (N534)? tag_v_r[63] : 1'b0;
  assign N544 = (N531)? tag_v_r[8] : 
                (N533)? tag_v_r[26] : 
                (N532)? tag_v_r[44] : 
                (N534)? tag_v_r[62] : 1'b0;
  assign N545 = (N531)? tag_v_r[7] : 
                (N533)? tag_v_r[25] : 
                (N532)? tag_v_r[43] : 
                (N534)? tag_v_r[61] : 1'b0;
  assign N546 = (N531)? tag_v_r[6] : 
                (N533)? tag_v_r[24] : 
                (N532)? tag_v_r[42] : 
                (N534)? tag_v_r[60] : 1'b0;
  assign N547 = (N531)? tag_v_r[5] : 
                (N533)? tag_v_r[23] : 
                (N532)? tag_v_r[41] : 
                (N534)? tag_v_r[59] : 1'b0;
  assign N548 = (N531)? tag_v_r[4] : 
                (N533)? tag_v_r[22] : 
                (N532)? tag_v_r[40] : 
                (N534)? tag_v_r[58] : 1'b0;
  assign N549 = (N531)? tag_v_r[3] : 
                (N533)? tag_v_r[21] : 
                (N532)? tag_v_r[39] : 
                (N534)? tag_v_r[57] : 1'b0;
  assign N550 = (N531)? tag_v_r[2] : 
                (N533)? tag_v_r[20] : 
                (N532)? tag_v_r[38] : 
                (N534)? tag_v_r[56] : 1'b0;
  assign N551 = (N531)? tag_v_r[1] : 
                (N533)? tag_v_r[19] : 
                (N532)? tag_v_r[37] : 
                (N534)? tag_v_r[55] : 1'b0;
  assign N552 = (N531)? tag_v_r[0] : 
                (N533)? tag_v_r[18] : 
                (N532)? tag_v_r[36] : 
                (N534)? tag_v_r[54] : 1'b0;

  bsg_decode_num_out_p4
  addr_way_demux
  (
    .i(cache_pkt_i[47:46]),
    .o(addr_way_decode)
  );


  bsg_lru_pseudo_tree_decode_ways_p4
  plru_decode
  (
    .way_id_i(tag_hit_way_id),
    .data_o(plru_decode_data_lo),
    .mask_o(plru_decode_mask_lo)
  );

  assign { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331 } = data_v_r + atomic_mem_data;
  assign N69 = (N0)? 1'b1 : 
               (N73)? 1'b1 : 
               (N68)? 1'b0 : 1'b0;
  assign N0 = tl_we;
  assign N70 = (N0)? v_i : 
               (N73)? 1'b0 : 1'b0;
  assign N71 = (N0)? v_i : 
               (N73)? 1'b0 : 
               (N68)? 1'b0 : 1'b0;
  assign N77 = (N1)? 1'b1 : 
               (N2)? 1'b0 : 1'b0;
  assign N1 = v_we_o;
  assign N78 = (N1)? v_tl_r : 
               (N2)? 1'b0 : 1'b0;
  assign { N81, N80, N79 } = (N1)? { v_tl_r, v_tl_r, v_tl_r } : 
                             (N2)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N83, N82 } = (N3)? { 1'b0, 1'b0 } : 
                        (N85)? { v_tl_r, v_tl_r } : 
                        (N76)? { 1'b0, 1'b0 } : 1'b0;
  assign N3 = N74;
  assign N93 = (N4)? N91 : 
               (N90)? N92 : 1'b0;
  assign N4 = decode[17];
  assign N97 = (N5)? N95 : 
               (N94)? N96 : 1'b0;
  assign N5 = decode_tl_r[17];
  assign N102 = (N6)? N100 : 
                (N99)? N101 : 1'b0;
  assign N6 = N98;
  assign N137 = (N7)? N136 : 
                (N8)? 1'b1 : 1'b0;
  assign N7 = N128;
  assign N8 = N127;
  assign N147 = (N9)? N146 : 
                (N10)? 1'b0 : 1'b0;
  assign N9 = N139;
  assign N10 = N138;
  assign sbuf_data_mem_w_mask[3:0] = (N11)? { N149, N150, N151, N152 } : 
                                     (N148)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = sbuf_way_decode[0];
  assign sbuf_data_mem_w_mask[7:4] = (N12)? { N154, N155, N156, N157 } : 
                                     (N153)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = sbuf_way_decode[1];
  assign sbuf_data_mem_w_mask[11:8] = (N13)? { N159, N160, N161, N162 } : 
                                      (N158)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = sbuf_way_decode[2];
  assign sbuf_data_mem_w_mask[15:12] = (N14)? { N164, N165, N166, N167 } : 
                                       (N163)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = sbuf_way_decode[3];
  assign { N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365 } = (N15)? data_v_r : 
                                                                                                                                                                                                              (N364)? atomic_mem_data : 1'b0;
  assign N15 = N363;
  assign { N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399 } = (N16)? data_v_r : 
                                                                                                                                                                                                              (N398)? atomic_mem_data : 1'b0;
  assign N16 = N397;
  assign { N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433 } = (N17)? data_v_r : 
                                                                                                                                                                                                              (N432)? atomic_mem_data : 1'b0;
  assign N17 = N431;
  assign { N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467 } = (N18)? data_v_r : 
                                                                                                                                                                                                              (N466)? atomic_mem_data : 1'b0;
  assign N18 = N465;
  assign atomic_alu_result = (N19)? data_v_r : 
                             (N20)? { N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266 } : 
                             (N21)? { N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298 } : 
                             (N22)? { N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330 } : 
                             (N23)? { N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331 } : 
                             (N24)? { N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365 } : 
                             (N25)? { N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399 } : 
                             (N26)? { N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433 } : 
                             (N27)? { N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467 } : 
                             (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N29)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = N174;
  assign N20 = N181;
  assign N21 = N187;
  assign N22 = N193;
  assign N23 = N199;
  assign N24 = N206;
  assign N25 = N213;
  assign N26 = N221;
  assign N27 = N227;
  assign N28 = N169;
  assign N29 = N234;
  assign \sbuf_in_sel_2_.slice_data  = (N30)? atomic_alu_result : 
                                       (N500)? data_v_r : 1'b0;
  assign N30 = N499;
  assign { sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_ } = (N31)? { data_v_r, mask_v_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N502)? { sbuf_data_in, sbuf_mask_in } : 1'b0;
  assign N31 = N501;
  assign tbuf_track_mem_w_mask[3:0] = (N32)? tbuf_word_offset_decode : 
                                      (N503)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = tbuf_way_decode[0];
  assign tbuf_track_mem_w_mask[7:4] = (N33)? tbuf_word_offset_decode : 
                                      (N504)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = tbuf_way_decode[1];
  assign tbuf_track_mem_w_mask[11:8] = (N34)? tbuf_word_offset_decode : 
                                       (N505)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = tbuf_way_decode[2];
  assign tbuf_track_mem_w_mask[15:12] = (N35)? tbuf_word_offset_decode : 
                                        (N506)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = tbuf_way_decode[3];
  assign snoop_or_ld_data = (N36)? snoop_word_lo : 
                            (N37)? bypass_data_masked : 1'b0;
  assign N36 = select_snoop_data_r_lo;
  assign N37 = N507;
  assign { N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553 } = (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N521, N528 } : 
                                                                                                                                                                                                              (N586)? { 1'b0, 1'b0, 1'b0, 1'b0, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, addr_v_r[9:4], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N589)? ld_data_masked : 
                                                                                                                                                                                                              (N514)? ld_data_final_lo : 1'b0;
  assign N38 = N509;
  assign data_o = (N39)? { N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553 } : 
                  (N40)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N39 = retval_op_v;
  assign N40 = N508;
  assign N592 = (N41)? miss_done_lo : 
                (N42)? 1'b1 : 1'b0;
  assign N41 = N591;
  assign N42 = N590;
  assign v_we_o = (N43)? N594 : 
                  (N44)? 1'b1 : 1'b0;
  assign N43 = v_v_r;
  assign N44 = N593;
  assign N598 = (N45)? N597 : 
                (N46)? 1'b1 : 1'b0;
  assign N45 = N596;
  assign N46 = N595;
  assign N600 = (N47)? v_we_o : 
                (N48)? 1'b1 : 1'b0;
  assign N47 = v_tl_r;
  assign N48 = N599;
  assign tag_mem_w_li = (N49)? N603 : 
                        (N50)? tagst_write_en : 1'b0;
  assign N49 = N602;
  assign N50 = N601;
  assign { N613, N612, N611, N610, N609, N608 } = (N51)? addr_tl_r[9:4] : 
                                                  (N615)? miss_tag_mem_addr_lo : 
                                                  (N607)? cache_pkt_i[45:40] : 1'b0;
  assign N51 = recover_lo;
  assign tag_mem_addr_li = (N52)? { N613, N612, N611, N610, N609, N608 } : 
                           (N53)? cache_pkt_i[45:40] : 1'b0;
  assign N52 = N605;
  assign N53 = N604;
  assign tag_mem_data_li = (N52)? miss_tag_mem_data_lo : 
                           (N53)? { cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4] } : 1'b0;
  assign tag_mem_w_mask_li = (N52)? miss_tag_mem_w_mask_lo : 
                             (N53)? { addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:3], addr_way_decode[3:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:2], addr_way_decode[2:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0] } : 1'b0;
  assign data_mem_data_li = (N54)? dma_data_mem_data_lo : 
                            (N55)? { sbuf_entry_lo[37:6], sbuf_entry_lo[37:6], sbuf_entry_lo[37:6], sbuf_entry_lo[37:6] } : 1'b0;
  assign N54 = dma_data_mem_w_lo;
  assign N55 = N616;
  assign data_mem_addr_li = (N51)? addr_tl_r[9:2] : 
                            (N621)? dma_data_mem_addr_lo : 
                            (N624)? cache_pkt_i[45:38] : 
                            (N620)? sbuf_entry_lo[47:40] : 1'b0;
  assign data_mem_w_mask_li = (N54)? dma_data_mem_w_mask_lo : 
                              (N55)? sbuf_data_mem_w_mask : 1'b0;
  assign track_mem_w_li = (N56)? miss_track_mem_w_lo : 
                          (N57)? N625 : 1'b0;
  assign N56 = miss_track_mem_v_lo;
  assign N57 = N707;
  assign track_mem_data_li = (N56)? miss_track_mem_data_lo : 
                             (N57)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign track_mem_w_mask_li = (N56)? miss_track_mem_w_mask_lo : 
                               (N57)? tbuf_track_mem_w_mask : 1'b0;
  assign track_mem_addr_li = (N51)? addr_tl_r[9:4] : 
                             (N630)? miss_track_mem_addr_lo : 
                             (N633)? cache_pkt_i[45:40] : 
                             (N629)? tbuf_addr_lo[9:4] : 1'b0;
  assign { N654, N653, N652, N651, N650, N649, N648 } = (N58)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N639)? { N640, N641, N642, N643, plru_decode_data_lo } : 1'b0;
  assign N58 = N638;
  assign { N661, N660, N659, N658, N657, N656, N655 } = (N58)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                        (N639)? { N644, N645, N646, N647, plru_decode_mask_lo } : 1'b0;
  assign stat_mem_v_li = (N59)? miss_stat_mem_v_lo : 
                         (N60)? N636 : 1'b0;
  assign N59 = N635;
  assign N60 = N634;
  assign stat_mem_w_li = (N59)? miss_stat_mem_w_lo : 
                         (N60)? N637 : 1'b0;
  assign stat_mem_addr_li = (N59)? miss_stat_mem_addr_lo : 
                            (N60)? addr_v_r[9:4] : 1'b0;
  assign stat_mem_data_li = (N59)? miss_stat_mem_data_lo : 
                            (N60)? { N654, N653, N652, N651, N650, N649, N648 } : 1'b0;
  assign stat_mem_w_mask_li = (N59)? miss_stat_mem_w_mask_lo : 
                              (N60)? { N661, N660, N659, N658, N657, N656, N655 } : 1'b0;
  assign { sbuf_entry_li_way_id__1_, sbuf_entry_li_way_id__0_ } = (N61)? chosen_way_lo : 
                                                                  (N62)? tag_hit_way_id : 1'b0;
  assign N61 = N663;
  assign N62 = N662;
  assign tbuf_way_li = (N63)? chosen_way_lo : 
                       (N64)? tag_hit_way_id : 1'b0;
  assign N63 = N665;
  assign N64 = N664;
  assign N666 = ~decode_v_r[0];
  assign N667 = N65 & N666;
  assign N65 = ~decode_v_r[1];
  assign N168 = N66 & N667;
  assign N66 = ~decode_v_r[3];
  assign N67 = sbuf_hazard | tl_we;
  assign N68 = ~N67;
  assign N72 = ~tl_we;
  assign N73 = sbuf_hazard & N72;
  assign N74 = reset_i;
  assign N75 = v_we_o | N74;
  assign N76 = ~N75;
  assign N84 = ~N74;
  assign N85 = v_we_o & N84;
  assign tag_hit_v[0] = N86 & valid_v_r[0];
  assign tag_hit_v[1] = N87 & valid_v_r[1];
  assign tag_hit_v[2] = N88 & valid_v_r[2];
  assign tag_hit_v[3] = N89 & valid_v_r[3];
  assign N90 = ~decode[17];
  assign N91 = ~N670;
  assign N670 = N669 & cache_pkt_i[0];
  assign N669 = N668 & cache_pkt_i[1];
  assign N668 = cache_pkt_i[3] & cache_pkt_i[2];
  assign N92 = ~decode[20];
  assign partial_st = decode[15] & N93;
  assign N94 = ~decode_tl_r[17];
  assign N95 = ~N673;
  assign N673 = N672 & mask_tl_r[0];
  assign N672 = N671 & mask_tl_r[1];
  assign N671 = mask_tl_r[3] & mask_tl_r[2];
  assign N96 = ~decode_tl_r[20];
  assign partial_st_tl = decode_tl_r[15] & N97;
  assign N98 = decode_v_r[17];
  assign N99 = ~N98;
  assign N100 = ~N676;
  assign N676 = N675 & mask_v_r[0];
  assign N675 = N674 & mask_v_r[1];
  assign N674 = mask_v_r[3] & mask_v_r[2];
  assign N101 = ~decode_v_r[20];
  assign partial_st_v = decode_v_r[15] & N102;
  assign ld_st_amo_tag_miss = N678 & N679;
  assign N678 = N677 | decode_v_r[4];
  assign N677 = decode_v_r[16] | decode_v_r[15];
  assign N679 = ~tag_hit_found;
  assign N103 = ~tag_hit_way_id[0];
  assign N104 = ~tag_hit_way_id[1];
  assign N105 = N103 & N104;
  assign N106 = N103 & tag_hit_way_id[1];
  assign N107 = tag_hit_way_id[0] & N104;
  assign N108 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign N113 = ~addr_v_r[2];
  assign N114 = ~addr_v_r[3];
  assign N115 = N113 & N114;
  assign N116 = N113 & addr_v_r[3];
  assign N117 = addr_v_r[2] & N114;
  assign N118 = addr_v_r[2] & addr_v_r[3];
  assign track_miss = N682 & N684;
  assign N682 = N681 & tag_hit_found;
  assign N681 = N680 | partial_st_v;
  assign N680 = decode_v_r[16] | decode_v_r[4];
  assign N684 = ~N683;
  assign N683 = N119 | bypass_track_lo;
  assign N120 = ~addr_v_r[10];
  assign N121 = ~addr_v_r[11];
  assign N122 = N120 & N121;
  assign N123 = N120 & addr_v_r[11];
  assign N124 = addr_v_r[10] & N121;
  assign N125 = addr_v_r[10] & addr_v_r[11];
  assign tagfl_hit = decode_v_r[13] & N126;
  assign aflinv_hit = N686 & tag_hit_found;
  assign N686 = N685 | decode_v_r[8];
  assign N685 = decode_v_r[10] | decode_v_r[9];
  assign N127 = ~tag_hit_found;
  assign N128 = tag_hit_found;
  assign N129 = ~tag_hit_way_id[0];
  assign N130 = ~tag_hit_way_id[1];
  assign N131 = N129 & N130;
  assign N132 = N129 & tag_hit_way_id[1];
  assign N133 = tag_hit_way_id[0] & N130;
  assign N134 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign N136 = ~N135;
  assign alock_miss = decode_v_r[7] & N137;
  assign N138 = ~tag_hit_found;
  assign N139 = tag_hit_found;
  assign N140 = ~tag_hit_way_id[0];
  assign N141 = ~tag_hit_way_id[1];
  assign N142 = N140 & N141;
  assign N143 = N140 & tag_hit_way_id[1];
  assign N144 = tag_hit_way_id[0] & N141;
  assign N145 = tag_hit_way_id[0] & tag_hit_way_id[1];
  assign aunlock_hit = decode_v_r[6] & N147;
  assign miss_v = N688 & N693;
  assign N688 = N687 & v_v_r;
  assign N687 = ~decode_v_r[14];
  assign N693 = N692 | aunlock_hit;
  assign N692 = N691 | alock_miss;
  assign N691 = N690 | aflinv_hit;
  assign N690 = N689 | tagfl_hit;
  assign N689 = ld_st_amo_tag_miss | track_miss;
  assign retval_op_v = N695 | decode_v_r[4];
  assign N695 = N694 | decode_v_r[11];
  assign N694 = decode_v_r[16] | decode_v_r[12];
  assign _1_net_ = v_o & yumi_i;
  assign N148 = ~sbuf_way_decode[0];
  assign N149 = sbuf_expand_mask[3] & sbuf_entry_lo[5];
  assign N150 = sbuf_expand_mask[2] & sbuf_entry_lo[4];
  assign N151 = sbuf_expand_mask[1] & sbuf_entry_lo[3];
  assign N152 = sbuf_expand_mask[0] & sbuf_entry_lo[2];
  assign N153 = ~sbuf_way_decode[1];
  assign N154 = sbuf_expand_mask[3] & sbuf_entry_lo[5];
  assign N155 = sbuf_expand_mask[2] & sbuf_entry_lo[4];
  assign N156 = sbuf_expand_mask[1] & sbuf_entry_lo[3];
  assign N157 = sbuf_expand_mask[0] & sbuf_entry_lo[2];
  assign N158 = ~sbuf_way_decode[2];
  assign N159 = sbuf_expand_mask[3] & sbuf_entry_lo[5];
  assign N160 = sbuf_expand_mask[2] & sbuf_entry_lo[4];
  assign N161 = sbuf_expand_mask[1] & sbuf_entry_lo[3];
  assign N162 = sbuf_expand_mask[0] & sbuf_entry_lo[2];
  assign N163 = ~sbuf_way_decode[3];
  assign N164 = sbuf_expand_mask[3] & sbuf_entry_lo[5];
  assign N165 = sbuf_expand_mask[2] & sbuf_entry_lo[4];
  assign N166 = sbuf_expand_mask[1] & sbuf_entry_lo[3];
  assign N167 = sbuf_expand_mask[0] & sbuf_entry_lo[2];
  assign N169 = ~N168;
  assign N174 = ~N173;
  assign N175 = ~decode_v_r[1];
  assign N176 = ~decode_v_r[0];
  assign N181 = ~N180;
  assign N182 = ~decode_v_r[2];
  assign N187 = ~N186;
  assign N188 = ~decode_v_r[1];
  assign N193 = ~N192;
  assign N194 = ~decode_v_r[0];
  assign N199 = ~N198;
  assign N200 = ~decode_v_r[2];
  assign N201 = ~decode_v_r[0];
  assign N206 = ~N205;
  assign N207 = ~decode_v_r[2];
  assign N208 = ~decode_v_r[1];
  assign N213 = ~N212;
  assign N214 = ~decode_v_r[2];
  assign N215 = ~decode_v_r[1];
  assign N216 = ~decode_v_r[0];
  assign N221 = ~N220;
  assign N222 = ~decode_v_r[3];
  assign N227 = ~N226;
  assign N234 = N229 | N696;
  assign N696 = N231 | N233;
  assign N235 = data_v_r[31] & atomic_mem_data[31];
  assign N236 = data_v_r[30] & atomic_mem_data[30];
  assign N237 = data_v_r[29] & atomic_mem_data[29];
  assign N238 = data_v_r[28] & atomic_mem_data[28];
  assign N239 = data_v_r[27] & atomic_mem_data[27];
  assign N240 = data_v_r[26] & atomic_mem_data[26];
  assign N241 = data_v_r[25] & atomic_mem_data[25];
  assign N242 = data_v_r[24] & atomic_mem_data[24];
  assign N243 = data_v_r[23] & atomic_mem_data[23];
  assign N244 = data_v_r[22] & atomic_mem_data[22];
  assign N245 = data_v_r[21] & atomic_mem_data[21];
  assign N246 = data_v_r[20] & atomic_mem_data[20];
  assign N247 = data_v_r[19] & atomic_mem_data[19];
  assign N248 = data_v_r[18] & atomic_mem_data[18];
  assign N249 = data_v_r[17] & atomic_mem_data[17];
  assign N250 = data_v_r[16] & atomic_mem_data[16];
  assign N251 = data_v_r[15] & atomic_mem_data[15];
  assign N252 = data_v_r[14] & atomic_mem_data[14];
  assign N253 = data_v_r[13] & atomic_mem_data[13];
  assign N254 = data_v_r[12] & atomic_mem_data[12];
  assign N255 = data_v_r[11] & atomic_mem_data[11];
  assign N256 = data_v_r[10] & atomic_mem_data[10];
  assign N257 = data_v_r[9] & atomic_mem_data[9];
  assign N258 = data_v_r[8] & atomic_mem_data[8];
  assign N259 = data_v_r[7] & atomic_mem_data[7];
  assign N260 = data_v_r[6] & atomic_mem_data[6];
  assign N261 = data_v_r[5] & atomic_mem_data[5];
  assign N262 = data_v_r[4] & atomic_mem_data[4];
  assign N263 = data_v_r[3] & atomic_mem_data[3];
  assign N264 = data_v_r[2] & atomic_mem_data[2];
  assign N265 = data_v_r[1] & atomic_mem_data[1];
  assign N266 = data_v_r[0] & atomic_mem_data[0];
  assign N267 = data_v_r[31] | atomic_mem_data[31];
  assign N268 = data_v_r[30] | atomic_mem_data[30];
  assign N269 = data_v_r[29] | atomic_mem_data[29];
  assign N270 = data_v_r[28] | atomic_mem_data[28];
  assign N271 = data_v_r[27] | atomic_mem_data[27];
  assign N272 = data_v_r[26] | atomic_mem_data[26];
  assign N273 = data_v_r[25] | atomic_mem_data[25];
  assign N274 = data_v_r[24] | atomic_mem_data[24];
  assign N275 = data_v_r[23] | atomic_mem_data[23];
  assign N276 = data_v_r[22] | atomic_mem_data[22];
  assign N277 = data_v_r[21] | atomic_mem_data[21];
  assign N278 = data_v_r[20] | atomic_mem_data[20];
  assign N279 = data_v_r[19] | atomic_mem_data[19];
  assign N280 = data_v_r[18] | atomic_mem_data[18];
  assign N281 = data_v_r[17] | atomic_mem_data[17];
  assign N282 = data_v_r[16] | atomic_mem_data[16];
  assign N283 = data_v_r[15] | atomic_mem_data[15];
  assign N284 = data_v_r[14] | atomic_mem_data[14];
  assign N285 = data_v_r[13] | atomic_mem_data[13];
  assign N286 = data_v_r[12] | atomic_mem_data[12];
  assign N287 = data_v_r[11] | atomic_mem_data[11];
  assign N288 = data_v_r[10] | atomic_mem_data[10];
  assign N289 = data_v_r[9] | atomic_mem_data[9];
  assign N290 = data_v_r[8] | atomic_mem_data[8];
  assign N291 = data_v_r[7] | atomic_mem_data[7];
  assign N292 = data_v_r[6] | atomic_mem_data[6];
  assign N293 = data_v_r[5] | atomic_mem_data[5];
  assign N294 = data_v_r[4] | atomic_mem_data[4];
  assign N295 = data_v_r[3] | atomic_mem_data[3];
  assign N296 = data_v_r[2] | atomic_mem_data[2];
  assign N297 = data_v_r[1] | atomic_mem_data[1];
  assign N298 = data_v_r[0] | atomic_mem_data[0];
  assign N299 = data_v_r[31] ^ atomic_mem_data[31];
  assign N300 = data_v_r[30] ^ atomic_mem_data[30];
  assign N301 = data_v_r[29] ^ atomic_mem_data[29];
  assign N302 = data_v_r[28] ^ atomic_mem_data[28];
  assign N303 = data_v_r[27] ^ atomic_mem_data[27];
  assign N304 = data_v_r[26] ^ atomic_mem_data[26];
  assign N305 = data_v_r[25] ^ atomic_mem_data[25];
  assign N306 = data_v_r[24] ^ atomic_mem_data[24];
  assign N307 = data_v_r[23] ^ atomic_mem_data[23];
  assign N308 = data_v_r[22] ^ atomic_mem_data[22];
  assign N309 = data_v_r[21] ^ atomic_mem_data[21];
  assign N310 = data_v_r[20] ^ atomic_mem_data[20];
  assign N311 = data_v_r[19] ^ atomic_mem_data[19];
  assign N312 = data_v_r[18] ^ atomic_mem_data[18];
  assign N313 = data_v_r[17] ^ atomic_mem_data[17];
  assign N314 = data_v_r[16] ^ atomic_mem_data[16];
  assign N315 = data_v_r[15] ^ atomic_mem_data[15];
  assign N316 = data_v_r[14] ^ atomic_mem_data[14];
  assign N317 = data_v_r[13] ^ atomic_mem_data[13];
  assign N318 = data_v_r[12] ^ atomic_mem_data[12];
  assign N319 = data_v_r[11] ^ atomic_mem_data[11];
  assign N320 = data_v_r[10] ^ atomic_mem_data[10];
  assign N321 = data_v_r[9] ^ atomic_mem_data[9];
  assign N322 = data_v_r[8] ^ atomic_mem_data[8];
  assign N323 = data_v_r[7] ^ atomic_mem_data[7];
  assign N324 = data_v_r[6] ^ atomic_mem_data[6];
  assign N325 = data_v_r[5] ^ atomic_mem_data[5];
  assign N326 = data_v_r[4] ^ atomic_mem_data[4];
  assign N327 = data_v_r[3] ^ atomic_mem_data[3];
  assign N328 = data_v_r[2] ^ atomic_mem_data[2];
  assign N329 = data_v_r[1] ^ atomic_mem_data[1];
  assign N330 = data_v_r[0] ^ atomic_mem_data[0];
  assign N364 = ~N363;
  assign N398 = ~N397;
  assign N432 = ~N431;
  assign N466 = ~N465;
  assign N499 = decode_v_r[4];
  assign N500 = ~N499;
  assign N501 = decode_v_r[17];
  assign N502 = ~N501;
  assign N503 = ~tbuf_way_decode[0];
  assign N504 = ~tbuf_way_decode[1];
  assign N505 = ~tbuf_way_decode[2];
  assign N506 = ~tbuf_way_decode[3];
  assign N507 = ~select_snoop_data_r_lo;
  assign ld_data_masked[31] = snoop_or_ld_data[31] & expanded_mask_v[31];
  assign ld_data_masked[30] = snoop_or_ld_data[30] & expanded_mask_v[30];
  assign ld_data_masked[29] = snoop_or_ld_data[29] & expanded_mask_v[29];
  assign ld_data_masked[28] = snoop_or_ld_data[28] & expanded_mask_v[28];
  assign ld_data_masked[27] = snoop_or_ld_data[27] & expanded_mask_v[27];
  assign ld_data_masked[26] = snoop_or_ld_data[26] & expanded_mask_v[26];
  assign ld_data_masked[25] = snoop_or_ld_data[25] & expanded_mask_v[25];
  assign ld_data_masked[24] = snoop_or_ld_data[24] & expanded_mask_v[24];
  assign ld_data_masked[23] = snoop_or_ld_data[23] & expanded_mask_v[23];
  assign ld_data_masked[22] = snoop_or_ld_data[22] & expanded_mask_v[22];
  assign ld_data_masked[21] = snoop_or_ld_data[21] & expanded_mask_v[21];
  assign ld_data_masked[20] = snoop_or_ld_data[20] & expanded_mask_v[20];
  assign ld_data_masked[19] = snoop_or_ld_data[19] & expanded_mask_v[19];
  assign ld_data_masked[18] = snoop_or_ld_data[18] & expanded_mask_v[18];
  assign ld_data_masked[17] = snoop_or_ld_data[17] & expanded_mask_v[17];
  assign ld_data_masked[16] = snoop_or_ld_data[16] & expanded_mask_v[16];
  assign ld_data_masked[15] = snoop_or_ld_data[15] & expanded_mask_v[15];
  assign ld_data_masked[14] = snoop_or_ld_data[14] & expanded_mask_v[14];
  assign ld_data_masked[13] = snoop_or_ld_data[13] & expanded_mask_v[13];
  assign ld_data_masked[12] = snoop_or_ld_data[12] & expanded_mask_v[12];
  assign ld_data_masked[11] = snoop_or_ld_data[11] & expanded_mask_v[11];
  assign ld_data_masked[10] = snoop_or_ld_data[10] & expanded_mask_v[10];
  assign ld_data_masked[9] = snoop_or_ld_data[9] & expanded_mask_v[9];
  assign ld_data_masked[8] = snoop_or_ld_data[8] & expanded_mask_v[8];
  assign ld_data_masked[7] = snoop_or_ld_data[7] & expanded_mask_v[7];
  assign ld_data_masked[6] = snoop_or_ld_data[6] & expanded_mask_v[6];
  assign ld_data_masked[5] = snoop_or_ld_data[5] & expanded_mask_v[5];
  assign ld_data_masked[4] = snoop_or_ld_data[4] & expanded_mask_v[4];
  assign ld_data_masked[3] = snoop_or_ld_data[3] & expanded_mask_v[3];
  assign ld_data_masked[2] = snoop_or_ld_data[2] & expanded_mask_v[2];
  assign ld_data_masked[1] = snoop_or_ld_data[1] & expanded_mask_v[1];
  assign ld_data_masked[0] = snoop_or_ld_data[0] & expanded_mask_v[0];
  assign ld_data_final_li_0__31_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__30_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__29_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__28_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__27_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__26_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__25_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__24_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__23_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__22_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__21_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__20_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__19_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__18_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__17_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__16_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__15_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__14_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__13_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__12_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__11_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__10_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__9_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__8_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_1__31_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__30_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__29_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__28_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__27_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__26_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__25_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__24_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__23_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__22_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__21_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__20_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__19_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__18_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__17_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__16_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign N508 = ~retval_op_v;
  assign N509 = decode_v_r[12];
  assign N510 = decode_v_r[11];
  assign N511 = decode_v_r[17];
  assign N512 = N510 | N509;
  assign N513 = N511 | N512;
  assign N514 = ~N513;
  assign N515 = ~addr_v_r[10];
  assign N516 = ~addr_v_r[11];
  assign N517 = N515 & N516;
  assign N518 = N515 & addr_v_r[11];
  assign N519 = addr_v_r[10] & N516;
  assign N520 = addr_v_r[10] & addr_v_r[11];
  assign N522 = ~addr_v_r[10];
  assign N523 = ~addr_v_r[11];
  assign N524 = N522 & N523;
  assign N525 = N522 & addr_v_r[11];
  assign N526 = addr_v_r[10] & N523;
  assign N527 = addr_v_r[10] & addr_v_r[11];
  assign N529 = ~addr_v_r[10];
  assign N530 = ~addr_v_r[11];
  assign N531 = N529 & N530;
  assign N532 = N529 & addr_v_r[11];
  assign N533 = addr_v_r[10] & N530;
  assign N534 = addr_v_r[10] & addr_v_r[11];
  assign N585 = ~N509;
  assign N586 = N510 & N585;
  assign N587 = ~N510;
  assign N588 = N585 & N587;
  assign N589 = N511 & N588;
  assign N590 = ~miss_v;
  assign N591 = miss_v;
  assign v_o = v_v_r & N592;
  assign N593 = ~v_v_r;
  assign N594 = v_o & yumi_i;
  assign sbuf_hazard = N700 & N702;
  assign N700 = sbuf_full_lo & N699;
  assign N699 = N697 & N698;
  assign N697 = v_o & yumi_i;
  assign N698 = decode_v_r[15] | decode_v_r[4];
  assign N702 = v_i & N701;
  assign N701 = decode[16] | decode[4];
  assign N595 = ~miss_v;
  assign N596 = miss_v;
  assign N597 = N712 & N713;
  assign N712 = N710 & N711;
  assign N710 = N708 & N709;
  assign N708 = N706 & N707;
  assign N706 = N704 & N705;
  assign N704 = ~N703;
  assign N703 = decode[14] & v_i;
  assign N705 = ~miss_tag_mem_v_lo;
  assign N707 = ~miss_track_mem_v_lo;
  assign N709 = ~dma_data_mem_v_lo;
  assign N711 = ~recover_lo;
  assign N713 = ~dma_evict_lo;
  assign tl_ready = N598 & N714;
  assign N714 = ~sbuf_hazard;
  assign N599 = ~v_tl_r;
  assign tl_we = tl_ready & N600;
  assign yumi_o = v_i & tl_we;
  assign tagst_write_en = decode[14] & yumi_o;
  assign tag_mem_v_li = N719 | N720;
  assign N719 = N718 | miss_tag_mem_v_lo;
  assign N718 = N715 | N717;
  assign N715 = decode[5] & yumi_o;
  assign N717 = N716 & v_tl_r;
  assign N716 = recover_lo & decode_tl_r[5];
  assign N720 = decode[14] & yumi_o;
  assign N601 = ~miss_v;
  assign N602 = miss_v;
  assign N603 = miss_tag_mem_v_lo & miss_tag_mem_w_lo;
  assign N604 = ~miss_v;
  assign N605 = miss_v;
  assign N606 = miss_tag_mem_v_lo | recover_lo;
  assign N607 = ~N606;
  assign N614 = ~recover_lo;
  assign N615 = miss_tag_mem_v_lo & N614;
  assign data_mem_v_li = N727 | N728;
  assign N727 = N726 | dma_data_mem_v_lo;
  assign N726 = N722 | N725;
  assign N722 = yumi_o & N721;
  assign N721 = decode[16] | decode[4];
  assign N725 = N723 & N724;
  assign N723 = v_tl_r & recover_lo;
  assign N724 = decode_tl_r[16] | decode_tl_r[4];
  assign N728 = sbuf_v_lo & sbuf_yumi_li;
  assign data_mem_w_li = dma_data_mem_w_lo | N729;
  assign N729 = sbuf_v_lo & sbuf_yumi_li;
  assign N616 = ~dma_data_mem_w_lo;
  assign N617 = N730 & yumi_o;
  assign N730 = decode[16] | decode[4];
  assign N618 = dma_data_mem_v_lo | recover_lo;
  assign N619 = N617 | N618;
  assign N620 = ~N619;
  assign N621 = dma_data_mem_v_lo & N614;
  assign N622 = ~dma_data_mem_v_lo;
  assign N623 = N614 & N622;
  assign N624 = N617 & N623;
  assign track_mem_v_li = N739 | N740;
  assign N739 = N738 | miss_track_mem_v_lo;
  assign N738 = N733 | N737;
  assign N733 = yumi_o & N732;
  assign N732 = N731 | partial_st;
  assign N731 = decode[16] | decode[4];
  assign N737 = N734 & N736;
  assign N734 = v_tl_r & recover_lo;
  assign N736 = N735 | partial_st_tl;
  assign N735 = decode_tl_r[16] | decode_tl_r[4];
  assign N740 = tbuf_v_lo & tbuf_yumi_li;
  assign N625 = tbuf_v_lo & tbuf_yumi_li;
  assign N626 = N742 & yumi_o;
  assign N742 = N741 | partial_st;
  assign N741 = decode[16] | decode[4];
  assign N627 = miss_track_mem_v_lo | recover_lo;
  assign N628 = N626 | N627;
  assign N629 = ~N628;
  assign N630 = miss_track_mem_v_lo & N614;
  assign N631 = ~miss_track_mem_v_lo;
  assign N632 = N614 & N631;
  assign N633 = N626 & N632;
  assign N634 = ~miss_v;
  assign N635 = miss_v;
  assign N636 = N746 & yumi_i;
  assign N746 = N745 & v_o;
  assign N745 = N744 | decode_v_r[4];
  assign N744 = N743 | decode_v_r[14];
  assign N743 = decode_v_r[15] | decode_v_r[16];
  assign N637 = N750 & yumi_i;
  assign N750 = N749 & v_o;
  assign N749 = N748 | decode_v_r[4];
  assign N748 = N747 | decode_v_r[14];
  assign N747 = decode_v_r[15] | decode_v_r[16];
  assign N638 = decode_v_r[14];
  assign N639 = ~N638;
  assign N640 = decode_v_r[15] | decode_v_r[4];
  assign N641 = decode_v_r[15] | decode_v_r[4];
  assign N642 = decode_v_r[15] | decode_v_r[4];
  assign N643 = decode_v_r[15] | decode_v_r[4];
  assign N644 = N751 & tag_hit_v[3];
  assign N751 = decode_v_r[15] | decode_v_r[4];
  assign N645 = N752 & tag_hit_v[2];
  assign N752 = decode_v_r[15] | decode_v_r[4];
  assign N646 = N753 & tag_hit_v[1];
  assign N753 = decode_v_r[15] | decode_v_r[4];
  assign N647 = N754 & tag_hit_v[0];
  assign N754 = decode_v_r[15] | decode_v_r[4];
  assign sbuf_v_li = N756 & yumi_i;
  assign N756 = N755 & v_o;
  assign N755 = decode_v_r[15] | decode_v_r[4];
  assign N662 = ~miss_v;
  assign N663 = miss_v;
  assign sbuf_yumi_li = N761 & N768;
  assign N761 = N760 & N709;
  assign N760 = sbuf_v_lo & N759;
  assign N759 = ~N758;
  assign N758 = N757 & yumi_o;
  assign N757 = decode[16] | decode[4];
  assign N768 = ~N767;
  assign N767 = N765 & N766;
  assign N765 = N763 & N764;
  assign N763 = v_tl_r & N762;
  assign N762 = decode_tl_r[16] | decode_tl_r[4];
  assign N764 = ~v_we_o;
  assign N766 = ~miss_v;
  assign sbuf_bypass_v_li = N770 & v_we_o;
  assign N770 = N769 & v_tl_r;
  assign N769 = decode_tl_r[16] | decode_tl_r[4];
  assign tbuf_v_li = N773 & yumi_i;
  assign N773 = N772 & v_o;
  assign N772 = decode_v_r[15] & N771;
  assign N771 = ~partial_st_v;
  assign N664 = ~miss_v;
  assign N665 = miss_v;
  assign tbuf_yumi_li = N779 & N786;
  assign N779 = N778 & N707;
  assign N778 = tbuf_v_lo & N777;
  assign N777 = ~N776;
  assign N776 = N775 & yumi_o;
  assign N775 = N774 | partial_st;
  assign N774 = decode[16] | decode[4];
  assign N786 = ~N785;
  assign N785 = N783 & N784;
  assign N783 = N782 & N764;
  assign N782 = v_tl_r & N781;
  assign N781 = N780 | partial_st_tl;
  assign N780 = decode_tl_r[16] | decode_tl_r[4];
  assign N784 = ~miss_v;
  assign tbuf_bypass_v_li = N789 & v_we_o;
  assign N789 = N788 & v_tl_r;
  assign N788 = N787 | partial_st_tl;
  assign N787 = decode_tl_r[16] | decode_tl_r[4];
  assign N2 = ~v_we_o;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_tl_r_31_sv2v_reg <= 1'b0;
      data_tl_r_30_sv2v_reg <= 1'b0;
      data_tl_r_29_sv2v_reg <= 1'b0;
      data_tl_r_28_sv2v_reg <= 1'b0;
      data_tl_r_27_sv2v_reg <= 1'b0;
      data_tl_r_26_sv2v_reg <= 1'b0;
      data_tl_r_25_sv2v_reg <= 1'b0;
      data_tl_r_24_sv2v_reg <= 1'b0;
      data_tl_r_23_sv2v_reg <= 1'b0;
      data_tl_r_22_sv2v_reg <= 1'b0;
      data_tl_r_21_sv2v_reg <= 1'b0;
      data_tl_r_20_sv2v_reg <= 1'b0;
      data_tl_r_19_sv2v_reg <= 1'b0;
      data_tl_r_18_sv2v_reg <= 1'b0;
      data_tl_r_17_sv2v_reg <= 1'b0;
      data_tl_r_16_sv2v_reg <= 1'b0;
      data_tl_r_15_sv2v_reg <= 1'b0;
      data_tl_r_14_sv2v_reg <= 1'b0;
      data_tl_r_13_sv2v_reg <= 1'b0;
      data_tl_r_12_sv2v_reg <= 1'b0;
      data_tl_r_11_sv2v_reg <= 1'b0;
      data_tl_r_10_sv2v_reg <= 1'b0;
      data_tl_r_9_sv2v_reg <= 1'b0;
      data_tl_r_8_sv2v_reg <= 1'b0;
      data_tl_r_7_sv2v_reg <= 1'b0;
      data_tl_r_6_sv2v_reg <= 1'b0;
      data_tl_r_5_sv2v_reg <= 1'b0;
      data_tl_r_4_sv2v_reg <= 1'b0;
      data_tl_r_3_sv2v_reg <= 1'b0;
      data_tl_r_2_sv2v_reg <= 1'b0;
      data_tl_r_1_sv2v_reg <= 1'b0;
      data_tl_r_0_sv2v_reg <= 1'b0;
      decode_tl_r_20_sv2v_reg <= 1'b0;
      decode_tl_r_19_sv2v_reg <= 1'b0;
      decode_tl_r_18_sv2v_reg <= 1'b0;
      decode_tl_r_17_sv2v_reg <= 1'b0;
      decode_tl_r_16_sv2v_reg <= 1'b0;
      decode_tl_r_15_sv2v_reg <= 1'b0;
      decode_tl_r_14_sv2v_reg <= 1'b0;
      decode_tl_r_13_sv2v_reg <= 1'b0;
      decode_tl_r_12_sv2v_reg <= 1'b0;
      decode_tl_r_11_sv2v_reg <= 1'b0;
      decode_tl_r_10_sv2v_reg <= 1'b0;
      decode_tl_r_9_sv2v_reg <= 1'b0;
      decode_tl_r_8_sv2v_reg <= 1'b0;
      decode_tl_r_7_sv2v_reg <= 1'b0;
      decode_tl_r_6_sv2v_reg <= 1'b0;
      decode_tl_r_5_sv2v_reg <= 1'b0;
      decode_tl_r_4_sv2v_reg <= 1'b0;
      decode_tl_r_3_sv2v_reg <= 1'b0;
      decode_tl_r_2_sv2v_reg <= 1'b0;
      decode_tl_r_1_sv2v_reg <= 1'b0;
      decode_tl_r_0_sv2v_reg <= 1'b0;
      mask_tl_r_3_sv2v_reg <= 1'b0;
      mask_tl_r_2_sv2v_reg <= 1'b0;
      mask_tl_r_1_sv2v_reg <= 1'b0;
      mask_tl_r_0_sv2v_reg <= 1'b0;
      addr_tl_r_27_sv2v_reg <= 1'b0;
      addr_tl_r_26_sv2v_reg <= 1'b0;
      addr_tl_r_25_sv2v_reg <= 1'b0;
      addr_tl_r_24_sv2v_reg <= 1'b0;
      addr_tl_r_23_sv2v_reg <= 1'b0;
      addr_tl_r_22_sv2v_reg <= 1'b0;
      addr_tl_r_21_sv2v_reg <= 1'b0;
      addr_tl_r_20_sv2v_reg <= 1'b0;
      addr_tl_r_19_sv2v_reg <= 1'b0;
      addr_tl_r_18_sv2v_reg <= 1'b0;
      addr_tl_r_17_sv2v_reg <= 1'b0;
      addr_tl_r_16_sv2v_reg <= 1'b0;
      addr_tl_r_15_sv2v_reg <= 1'b0;
      addr_tl_r_14_sv2v_reg <= 1'b0;
      addr_tl_r_13_sv2v_reg <= 1'b0;
      addr_tl_r_12_sv2v_reg <= 1'b0;
      addr_tl_r_11_sv2v_reg <= 1'b0;
      addr_tl_r_10_sv2v_reg <= 1'b0;
      addr_tl_r_9_sv2v_reg <= 1'b0;
      addr_tl_r_8_sv2v_reg <= 1'b0;
      addr_tl_r_7_sv2v_reg <= 1'b0;
      addr_tl_r_6_sv2v_reg <= 1'b0;
      addr_tl_r_5_sv2v_reg <= 1'b0;
      addr_tl_r_4_sv2v_reg <= 1'b0;
      addr_tl_r_3_sv2v_reg <= 1'b0;
      addr_tl_r_2_sv2v_reg <= 1'b0;
      addr_tl_r_1_sv2v_reg <= 1'b0;
      addr_tl_r_0_sv2v_reg <= 1'b0;
    end else if(N71) begin
      data_tl_r_31_sv2v_reg <= cache_pkt_i[35];
      data_tl_r_30_sv2v_reg <= cache_pkt_i[34];
      data_tl_r_29_sv2v_reg <= cache_pkt_i[33];
      data_tl_r_28_sv2v_reg <= cache_pkt_i[32];
      data_tl_r_27_sv2v_reg <= cache_pkt_i[31];
      data_tl_r_26_sv2v_reg <= cache_pkt_i[30];
      data_tl_r_25_sv2v_reg <= cache_pkt_i[29];
      data_tl_r_24_sv2v_reg <= cache_pkt_i[28];
      data_tl_r_23_sv2v_reg <= cache_pkt_i[27];
      data_tl_r_22_sv2v_reg <= cache_pkt_i[26];
      data_tl_r_21_sv2v_reg <= cache_pkt_i[25];
      data_tl_r_20_sv2v_reg <= cache_pkt_i[24];
      data_tl_r_19_sv2v_reg <= cache_pkt_i[23];
      data_tl_r_18_sv2v_reg <= cache_pkt_i[22];
      data_tl_r_17_sv2v_reg <= cache_pkt_i[21];
      data_tl_r_16_sv2v_reg <= cache_pkt_i[20];
      data_tl_r_15_sv2v_reg <= cache_pkt_i[19];
      data_tl_r_14_sv2v_reg <= cache_pkt_i[18];
      data_tl_r_13_sv2v_reg <= cache_pkt_i[17];
      data_tl_r_12_sv2v_reg <= cache_pkt_i[16];
      data_tl_r_11_sv2v_reg <= cache_pkt_i[15];
      data_tl_r_10_sv2v_reg <= cache_pkt_i[14];
      data_tl_r_9_sv2v_reg <= cache_pkt_i[13];
      data_tl_r_8_sv2v_reg <= cache_pkt_i[12];
      data_tl_r_7_sv2v_reg <= cache_pkt_i[11];
      data_tl_r_6_sv2v_reg <= cache_pkt_i[10];
      data_tl_r_5_sv2v_reg <= cache_pkt_i[9];
      data_tl_r_4_sv2v_reg <= cache_pkt_i[8];
      data_tl_r_3_sv2v_reg <= cache_pkt_i[7];
      data_tl_r_2_sv2v_reg <= cache_pkt_i[6];
      data_tl_r_1_sv2v_reg <= cache_pkt_i[5];
      data_tl_r_0_sv2v_reg <= cache_pkt_i[4];
      decode_tl_r_20_sv2v_reg <= decode[20];
      decode_tl_r_19_sv2v_reg <= decode[19];
      decode_tl_r_18_sv2v_reg <= decode[18];
      decode_tl_r_17_sv2v_reg <= decode[17];
      decode_tl_r_16_sv2v_reg <= decode[16];
      decode_tl_r_15_sv2v_reg <= decode[15];
      decode_tl_r_14_sv2v_reg <= decode[14];
      decode_tl_r_13_sv2v_reg <= decode[13];
      decode_tl_r_12_sv2v_reg <= decode[12];
      decode_tl_r_11_sv2v_reg <= decode[11];
      decode_tl_r_10_sv2v_reg <= decode[10];
      decode_tl_r_9_sv2v_reg <= decode[9];
      decode_tl_r_8_sv2v_reg <= decode[8];
      decode_tl_r_7_sv2v_reg <= decode[7];
      decode_tl_r_6_sv2v_reg <= decode[6];
      decode_tl_r_5_sv2v_reg <= decode[5];
      decode_tl_r_4_sv2v_reg <= decode[4];
      decode_tl_r_3_sv2v_reg <= decode[3];
      decode_tl_r_2_sv2v_reg <= decode[2];
      decode_tl_r_1_sv2v_reg <= decode[1];
      decode_tl_r_0_sv2v_reg <= decode[0];
      mask_tl_r_3_sv2v_reg <= cache_pkt_i[3];
      mask_tl_r_2_sv2v_reg <= cache_pkt_i[2];
      mask_tl_r_1_sv2v_reg <= cache_pkt_i[1];
      mask_tl_r_0_sv2v_reg <= cache_pkt_i[0];
      addr_tl_r_27_sv2v_reg <= cache_pkt_i[63];
      addr_tl_r_26_sv2v_reg <= cache_pkt_i[62];
      addr_tl_r_25_sv2v_reg <= cache_pkt_i[61];
      addr_tl_r_24_sv2v_reg <= cache_pkt_i[60];
      addr_tl_r_23_sv2v_reg <= cache_pkt_i[59];
      addr_tl_r_22_sv2v_reg <= cache_pkt_i[58];
      addr_tl_r_21_sv2v_reg <= cache_pkt_i[57];
      addr_tl_r_20_sv2v_reg <= cache_pkt_i[56];
      addr_tl_r_19_sv2v_reg <= cache_pkt_i[55];
      addr_tl_r_18_sv2v_reg <= cache_pkt_i[54];
      addr_tl_r_17_sv2v_reg <= cache_pkt_i[53];
      addr_tl_r_16_sv2v_reg <= cache_pkt_i[52];
      addr_tl_r_15_sv2v_reg <= cache_pkt_i[51];
      addr_tl_r_14_sv2v_reg <= cache_pkt_i[50];
      addr_tl_r_13_sv2v_reg <= cache_pkt_i[49];
      addr_tl_r_12_sv2v_reg <= cache_pkt_i[48];
      addr_tl_r_11_sv2v_reg <= cache_pkt_i[47];
      addr_tl_r_10_sv2v_reg <= cache_pkt_i[46];
      addr_tl_r_9_sv2v_reg <= cache_pkt_i[45];
      addr_tl_r_8_sv2v_reg <= cache_pkt_i[44];
      addr_tl_r_7_sv2v_reg <= cache_pkt_i[43];
      addr_tl_r_6_sv2v_reg <= cache_pkt_i[42];
      addr_tl_r_5_sv2v_reg <= cache_pkt_i[41];
      addr_tl_r_4_sv2v_reg <= cache_pkt_i[40];
      addr_tl_r_3_sv2v_reg <= cache_pkt_i[39];
      addr_tl_r_2_sv2v_reg <= cache_pkt_i[38];
      addr_tl_r_1_sv2v_reg <= cache_pkt_i[37];
      addr_tl_r_0_sv2v_reg <= cache_pkt_i[36];
    end 
    if(reset_i) begin
      v_tl_r_sv2v_reg <= 1'b0;
    end else if(N69) begin
      v_tl_r_sv2v_reg <= N70;
    end 
    if(N83) begin
      ld_data_v_r_127_sv2v_reg <= data_mem_data_lo[127];
      ld_data_v_r_126_sv2v_reg <= data_mem_data_lo[126];
      ld_data_v_r_125_sv2v_reg <= data_mem_data_lo[125];
      ld_data_v_r_124_sv2v_reg <= data_mem_data_lo[124];
      ld_data_v_r_123_sv2v_reg <= data_mem_data_lo[123];
      ld_data_v_r_122_sv2v_reg <= data_mem_data_lo[122];
      ld_data_v_r_121_sv2v_reg <= data_mem_data_lo[121];
      ld_data_v_r_120_sv2v_reg <= data_mem_data_lo[120];
      ld_data_v_r_119_sv2v_reg <= data_mem_data_lo[119];
      ld_data_v_r_118_sv2v_reg <= data_mem_data_lo[118];
      ld_data_v_r_117_sv2v_reg <= data_mem_data_lo[117];
      ld_data_v_r_116_sv2v_reg <= data_mem_data_lo[116];
      ld_data_v_r_115_sv2v_reg <= data_mem_data_lo[115];
      ld_data_v_r_114_sv2v_reg <= data_mem_data_lo[114];
      ld_data_v_r_113_sv2v_reg <= data_mem_data_lo[113];
      ld_data_v_r_112_sv2v_reg <= data_mem_data_lo[112];
      ld_data_v_r_111_sv2v_reg <= data_mem_data_lo[111];
      ld_data_v_r_110_sv2v_reg <= data_mem_data_lo[110];
      ld_data_v_r_109_sv2v_reg <= data_mem_data_lo[109];
      ld_data_v_r_108_sv2v_reg <= data_mem_data_lo[108];
      ld_data_v_r_107_sv2v_reg <= data_mem_data_lo[107];
      ld_data_v_r_106_sv2v_reg <= data_mem_data_lo[106];
      ld_data_v_r_105_sv2v_reg <= data_mem_data_lo[105];
      ld_data_v_r_104_sv2v_reg <= data_mem_data_lo[104];
      ld_data_v_r_103_sv2v_reg <= data_mem_data_lo[103];
      ld_data_v_r_102_sv2v_reg <= data_mem_data_lo[102];
      ld_data_v_r_101_sv2v_reg <= data_mem_data_lo[101];
      ld_data_v_r_100_sv2v_reg <= data_mem_data_lo[100];
      ld_data_v_r_99_sv2v_reg <= data_mem_data_lo[99];
      ld_data_v_r_98_sv2v_reg <= data_mem_data_lo[98];
      ld_data_v_r_97_sv2v_reg <= data_mem_data_lo[97];
      ld_data_v_r_96_sv2v_reg <= data_mem_data_lo[96];
      ld_data_v_r_95_sv2v_reg <= data_mem_data_lo[95];
      ld_data_v_r_94_sv2v_reg <= data_mem_data_lo[94];
      ld_data_v_r_93_sv2v_reg <= data_mem_data_lo[93];
      ld_data_v_r_92_sv2v_reg <= data_mem_data_lo[92];
      ld_data_v_r_91_sv2v_reg <= data_mem_data_lo[91];
      ld_data_v_r_90_sv2v_reg <= data_mem_data_lo[90];
      ld_data_v_r_89_sv2v_reg <= data_mem_data_lo[89];
      ld_data_v_r_88_sv2v_reg <= data_mem_data_lo[88];
      ld_data_v_r_87_sv2v_reg <= data_mem_data_lo[87];
      ld_data_v_r_86_sv2v_reg <= data_mem_data_lo[86];
      ld_data_v_r_85_sv2v_reg <= data_mem_data_lo[85];
      ld_data_v_r_84_sv2v_reg <= data_mem_data_lo[84];
      ld_data_v_r_83_sv2v_reg <= data_mem_data_lo[83];
      ld_data_v_r_82_sv2v_reg <= data_mem_data_lo[82];
      ld_data_v_r_81_sv2v_reg <= data_mem_data_lo[81];
      ld_data_v_r_80_sv2v_reg <= data_mem_data_lo[80];
      ld_data_v_r_79_sv2v_reg <= data_mem_data_lo[79];
      ld_data_v_r_78_sv2v_reg <= data_mem_data_lo[78];
      ld_data_v_r_77_sv2v_reg <= data_mem_data_lo[77];
      ld_data_v_r_76_sv2v_reg <= data_mem_data_lo[76];
      ld_data_v_r_75_sv2v_reg <= data_mem_data_lo[75];
      ld_data_v_r_74_sv2v_reg <= data_mem_data_lo[74];
      ld_data_v_r_73_sv2v_reg <= data_mem_data_lo[73];
      ld_data_v_r_72_sv2v_reg <= data_mem_data_lo[72];
      ld_data_v_r_71_sv2v_reg <= data_mem_data_lo[71];
      ld_data_v_r_70_sv2v_reg <= data_mem_data_lo[70];
      ld_data_v_r_69_sv2v_reg <= data_mem_data_lo[69];
      ld_data_v_r_68_sv2v_reg <= data_mem_data_lo[68];
      ld_data_v_r_67_sv2v_reg <= data_mem_data_lo[67];
      ld_data_v_r_66_sv2v_reg <= data_mem_data_lo[66];
      ld_data_v_r_65_sv2v_reg <= data_mem_data_lo[65];
      ld_data_v_r_64_sv2v_reg <= data_mem_data_lo[64];
      ld_data_v_r_63_sv2v_reg <= data_mem_data_lo[63];
      ld_data_v_r_62_sv2v_reg <= data_mem_data_lo[62];
      ld_data_v_r_61_sv2v_reg <= data_mem_data_lo[61];
      ld_data_v_r_60_sv2v_reg <= data_mem_data_lo[60];
      ld_data_v_r_59_sv2v_reg <= data_mem_data_lo[59];
      ld_data_v_r_58_sv2v_reg <= data_mem_data_lo[58];
      ld_data_v_r_57_sv2v_reg <= data_mem_data_lo[57];
      ld_data_v_r_56_sv2v_reg <= data_mem_data_lo[56];
      ld_data_v_r_55_sv2v_reg <= data_mem_data_lo[55];
      ld_data_v_r_54_sv2v_reg <= data_mem_data_lo[54];
      ld_data_v_r_53_sv2v_reg <= data_mem_data_lo[53];
      ld_data_v_r_52_sv2v_reg <= data_mem_data_lo[52];
      ld_data_v_r_51_sv2v_reg <= data_mem_data_lo[51];
      ld_data_v_r_50_sv2v_reg <= data_mem_data_lo[50];
      ld_data_v_r_49_sv2v_reg <= data_mem_data_lo[49];
      ld_data_v_r_48_sv2v_reg <= data_mem_data_lo[48];
      ld_data_v_r_47_sv2v_reg <= data_mem_data_lo[47];
      ld_data_v_r_46_sv2v_reg <= data_mem_data_lo[46];
      ld_data_v_r_45_sv2v_reg <= data_mem_data_lo[45];
    end 
    if(N82) begin
      ld_data_v_r_44_sv2v_reg <= data_mem_data_lo[44];
      ld_data_v_r_43_sv2v_reg <= data_mem_data_lo[43];
      ld_data_v_r_42_sv2v_reg <= data_mem_data_lo[42];
      ld_data_v_r_41_sv2v_reg <= data_mem_data_lo[41];
      ld_data_v_r_40_sv2v_reg <= data_mem_data_lo[40];
      ld_data_v_r_39_sv2v_reg <= data_mem_data_lo[39];
      ld_data_v_r_38_sv2v_reg <= data_mem_data_lo[38];
      ld_data_v_r_37_sv2v_reg <= data_mem_data_lo[37];
      ld_data_v_r_36_sv2v_reg <= data_mem_data_lo[36];
      ld_data_v_r_35_sv2v_reg <= data_mem_data_lo[35];
      ld_data_v_r_34_sv2v_reg <= data_mem_data_lo[34];
      ld_data_v_r_33_sv2v_reg <= data_mem_data_lo[33];
      ld_data_v_r_32_sv2v_reg <= data_mem_data_lo[32];
      ld_data_v_r_31_sv2v_reg <= data_mem_data_lo[31];
      ld_data_v_r_30_sv2v_reg <= data_mem_data_lo[30];
      ld_data_v_r_29_sv2v_reg <= data_mem_data_lo[29];
      ld_data_v_r_28_sv2v_reg <= data_mem_data_lo[28];
      ld_data_v_r_27_sv2v_reg <= data_mem_data_lo[27];
      ld_data_v_r_26_sv2v_reg <= data_mem_data_lo[26];
      ld_data_v_r_25_sv2v_reg <= data_mem_data_lo[25];
      ld_data_v_r_24_sv2v_reg <= data_mem_data_lo[24];
      ld_data_v_r_23_sv2v_reg <= data_mem_data_lo[23];
      ld_data_v_r_22_sv2v_reg <= data_mem_data_lo[22];
      ld_data_v_r_21_sv2v_reg <= data_mem_data_lo[21];
      ld_data_v_r_20_sv2v_reg <= data_mem_data_lo[20];
      ld_data_v_r_19_sv2v_reg <= data_mem_data_lo[19];
      ld_data_v_r_18_sv2v_reg <= data_mem_data_lo[18];
      ld_data_v_r_17_sv2v_reg <= data_mem_data_lo[17];
      ld_data_v_r_16_sv2v_reg <= data_mem_data_lo[16];
      ld_data_v_r_15_sv2v_reg <= data_mem_data_lo[15];
      ld_data_v_r_14_sv2v_reg <= data_mem_data_lo[14];
      ld_data_v_r_13_sv2v_reg <= data_mem_data_lo[13];
      ld_data_v_r_12_sv2v_reg <= data_mem_data_lo[12];
      ld_data_v_r_11_sv2v_reg <= data_mem_data_lo[11];
      ld_data_v_r_10_sv2v_reg <= data_mem_data_lo[10];
      ld_data_v_r_9_sv2v_reg <= data_mem_data_lo[9];
      ld_data_v_r_8_sv2v_reg <= data_mem_data_lo[8];
      ld_data_v_r_7_sv2v_reg <= data_mem_data_lo[7];
      ld_data_v_r_6_sv2v_reg <= data_mem_data_lo[6];
      ld_data_v_r_5_sv2v_reg <= data_mem_data_lo[5];
      ld_data_v_r_4_sv2v_reg <= data_mem_data_lo[4];
      ld_data_v_r_3_sv2v_reg <= data_mem_data_lo[3];
      ld_data_v_r_2_sv2v_reg <= data_mem_data_lo[2];
      ld_data_v_r_1_sv2v_reg <= data_mem_data_lo[1];
      ld_data_v_r_0_sv2v_reg <= data_mem_data_lo[0];
    end 
    if(reset_i) begin
      v_v_r_sv2v_reg <= 1'b0;
    end else if(N77) begin
      v_v_r_sv2v_reg <= v_tl_r;
    end 
    if(reset_i) begin
      track_data_v_r_15_sv2v_reg <= 1'b0;
      track_data_v_r_14_sv2v_reg <= 1'b0;
      track_data_v_r_13_sv2v_reg <= 1'b0;
      track_data_v_r_12_sv2v_reg <= 1'b0;
      track_data_v_r_11_sv2v_reg <= 1'b0;
      track_data_v_r_10_sv2v_reg <= 1'b0;
      track_data_v_r_9_sv2v_reg <= 1'b0;
      track_data_v_r_8_sv2v_reg <= 1'b0;
      track_data_v_r_7_sv2v_reg <= 1'b0;
      track_data_v_r_6_sv2v_reg <= 1'b0;
      track_data_v_r_5_sv2v_reg <= 1'b0;
      track_data_v_r_4_sv2v_reg <= 1'b0;
      track_data_v_r_3_sv2v_reg <= 1'b0;
      track_data_v_r_2_sv2v_reg <= 1'b0;
      track_data_v_r_1_sv2v_reg <= 1'b0;
      track_data_v_r_0_sv2v_reg <= 1'b0;
      mask_v_r_0_sv2v_reg <= 1'b0;
    end else if(N78) begin
      track_data_v_r_15_sv2v_reg <= track_mem_data_lo[15];
      track_data_v_r_14_sv2v_reg <= track_mem_data_lo[14];
      track_data_v_r_13_sv2v_reg <= track_mem_data_lo[13];
      track_data_v_r_12_sv2v_reg <= track_mem_data_lo[12];
      track_data_v_r_11_sv2v_reg <= track_mem_data_lo[11];
      track_data_v_r_10_sv2v_reg <= track_mem_data_lo[10];
      track_data_v_r_9_sv2v_reg <= track_mem_data_lo[9];
      track_data_v_r_8_sv2v_reg <= track_mem_data_lo[8];
      track_data_v_r_7_sv2v_reg <= track_mem_data_lo[7];
      track_data_v_r_6_sv2v_reg <= track_mem_data_lo[6];
      track_data_v_r_5_sv2v_reg <= track_mem_data_lo[5];
      track_data_v_r_4_sv2v_reg <= track_mem_data_lo[4];
      track_data_v_r_3_sv2v_reg <= track_mem_data_lo[3];
      track_data_v_r_2_sv2v_reg <= track_mem_data_lo[2];
      track_data_v_r_1_sv2v_reg <= track_mem_data_lo[1];
      track_data_v_r_0_sv2v_reg <= track_mem_data_lo[0];
      mask_v_r_0_sv2v_reg <= mask_tl_r[0];
    end 
    if(reset_i) begin
      mask_v_r_3_sv2v_reg <= 1'b0;
      decode_v_r_7_sv2v_reg <= 1'b0;
      decode_v_r_6_sv2v_reg <= 1'b0;
      decode_v_r_5_sv2v_reg <= 1'b0;
      decode_v_r_4_sv2v_reg <= 1'b0;
      decode_v_r_3_sv2v_reg <= 1'b0;
      decode_v_r_2_sv2v_reg <= 1'b0;
      decode_v_r_1_sv2v_reg <= 1'b0;
      decode_v_r_0_sv2v_reg <= 1'b0;
    end else if(N81) begin
      mask_v_r_3_sv2v_reg <= mask_tl_r[3];
      decode_v_r_7_sv2v_reg <= decode_tl_r[7];
      decode_v_r_6_sv2v_reg <= decode_tl_r[6];
      decode_v_r_5_sv2v_reg <= decode_tl_r[5];
      decode_v_r_4_sv2v_reg <= decode_tl_r[4];
      decode_v_r_3_sv2v_reg <= decode_tl_r[3];
      decode_v_r_2_sv2v_reg <= decode_tl_r[2];
      decode_v_r_1_sv2v_reg <= decode_tl_r[1];
      decode_v_r_0_sv2v_reg <= decode_tl_r[0];
    end 
    if(reset_i) begin
      mask_v_r_2_sv2v_reg <= 1'b0;
      decode_v_r_20_sv2v_reg <= 1'b0;
      decode_v_r_19_sv2v_reg <= 1'b0;
      decode_v_r_18_sv2v_reg <= 1'b0;
      decode_v_r_17_sv2v_reg <= 1'b0;
      decode_v_r_16_sv2v_reg <= 1'b0;
      decode_v_r_15_sv2v_reg <= 1'b0;
      decode_v_r_14_sv2v_reg <= 1'b0;
      decode_v_r_13_sv2v_reg <= 1'b0;
      decode_v_r_12_sv2v_reg <= 1'b0;
      decode_v_r_11_sv2v_reg <= 1'b0;
      decode_v_r_10_sv2v_reg <= 1'b0;
      decode_v_r_9_sv2v_reg <= 1'b0;
      decode_v_r_8_sv2v_reg <= 1'b0;
      addr_v_r_27_sv2v_reg <= 1'b0;
      addr_v_r_26_sv2v_reg <= 1'b0;
      addr_v_r_25_sv2v_reg <= 1'b0;
      addr_v_r_24_sv2v_reg <= 1'b0;
      addr_v_r_23_sv2v_reg <= 1'b0;
      addr_v_r_22_sv2v_reg <= 1'b0;
      addr_v_r_21_sv2v_reg <= 1'b0;
      addr_v_r_20_sv2v_reg <= 1'b0;
      addr_v_r_19_sv2v_reg <= 1'b0;
      addr_v_r_18_sv2v_reg <= 1'b0;
      addr_v_r_17_sv2v_reg <= 1'b0;
      addr_v_r_16_sv2v_reg <= 1'b0;
      addr_v_r_15_sv2v_reg <= 1'b0;
      addr_v_r_14_sv2v_reg <= 1'b0;
      addr_v_r_13_sv2v_reg <= 1'b0;
      addr_v_r_12_sv2v_reg <= 1'b0;
      addr_v_r_11_sv2v_reg <= 1'b0;
      addr_v_r_10_sv2v_reg <= 1'b0;
      addr_v_r_9_sv2v_reg <= 1'b0;
      addr_v_r_8_sv2v_reg <= 1'b0;
      addr_v_r_7_sv2v_reg <= 1'b0;
      addr_v_r_6_sv2v_reg <= 1'b0;
      addr_v_r_5_sv2v_reg <= 1'b0;
      addr_v_r_4_sv2v_reg <= 1'b0;
      addr_v_r_3_sv2v_reg <= 1'b0;
      addr_v_r_2_sv2v_reg <= 1'b0;
      addr_v_r_1_sv2v_reg <= 1'b0;
      addr_v_r_0_sv2v_reg <= 1'b0;
      data_v_r_31_sv2v_reg <= 1'b0;
      data_v_r_30_sv2v_reg <= 1'b0;
      data_v_r_29_sv2v_reg <= 1'b0;
      data_v_r_28_sv2v_reg <= 1'b0;
      data_v_r_27_sv2v_reg <= 1'b0;
      data_v_r_26_sv2v_reg <= 1'b0;
      data_v_r_25_sv2v_reg <= 1'b0;
      data_v_r_24_sv2v_reg <= 1'b0;
      data_v_r_23_sv2v_reg <= 1'b0;
      data_v_r_22_sv2v_reg <= 1'b0;
      data_v_r_21_sv2v_reg <= 1'b0;
      data_v_r_20_sv2v_reg <= 1'b0;
      data_v_r_19_sv2v_reg <= 1'b0;
      data_v_r_18_sv2v_reg <= 1'b0;
      data_v_r_17_sv2v_reg <= 1'b0;
      data_v_r_16_sv2v_reg <= 1'b0;
      data_v_r_15_sv2v_reg <= 1'b0;
      data_v_r_14_sv2v_reg <= 1'b0;
      data_v_r_13_sv2v_reg <= 1'b0;
      data_v_r_12_sv2v_reg <= 1'b0;
      data_v_r_11_sv2v_reg <= 1'b0;
      data_v_r_10_sv2v_reg <= 1'b0;
      data_v_r_9_sv2v_reg <= 1'b0;
      data_v_r_8_sv2v_reg <= 1'b0;
      data_v_r_7_sv2v_reg <= 1'b0;
      data_v_r_6_sv2v_reg <= 1'b0;
      data_v_r_5_sv2v_reg <= 1'b0;
      data_v_r_4_sv2v_reg <= 1'b0;
      data_v_r_3_sv2v_reg <= 1'b0;
      data_v_r_2_sv2v_reg <= 1'b0;
      data_v_r_1_sv2v_reg <= 1'b0;
      data_v_r_0_sv2v_reg <= 1'b0;
      valid_v_r_3_sv2v_reg <= 1'b0;
      valid_v_r_2_sv2v_reg <= 1'b0;
      valid_v_r_1_sv2v_reg <= 1'b0;
      valid_v_r_0_sv2v_reg <= 1'b0;
      tag_v_r_21_sv2v_reg <= 1'b0;
      tag_v_r_20_sv2v_reg <= 1'b0;
      tag_v_r_19_sv2v_reg <= 1'b0;
      tag_v_r_18_sv2v_reg <= 1'b0;
      tag_v_r_17_sv2v_reg <= 1'b0;
      tag_v_r_16_sv2v_reg <= 1'b0;
      tag_v_r_15_sv2v_reg <= 1'b0;
      tag_v_r_14_sv2v_reg <= 1'b0;
      tag_v_r_13_sv2v_reg <= 1'b0;
      tag_v_r_12_sv2v_reg <= 1'b0;
      tag_v_r_11_sv2v_reg <= 1'b0;
      tag_v_r_10_sv2v_reg <= 1'b0;
      tag_v_r_9_sv2v_reg <= 1'b0;
      tag_v_r_8_sv2v_reg <= 1'b0;
      tag_v_r_7_sv2v_reg <= 1'b0;
      tag_v_r_6_sv2v_reg <= 1'b0;
      tag_v_r_5_sv2v_reg <= 1'b0;
      tag_v_r_4_sv2v_reg <= 1'b0;
      tag_v_r_3_sv2v_reg <= 1'b0;
      tag_v_r_2_sv2v_reg <= 1'b0;
      tag_v_r_1_sv2v_reg <= 1'b0;
      tag_v_r_0_sv2v_reg <= 1'b0;
    end else if(N80) begin
      mask_v_r_2_sv2v_reg <= mask_tl_r[2];
      decode_v_r_20_sv2v_reg <= decode_tl_r[20];
      decode_v_r_19_sv2v_reg <= decode_tl_r[19];
      decode_v_r_18_sv2v_reg <= decode_tl_r[18];
      decode_v_r_17_sv2v_reg <= decode_tl_r[17];
      decode_v_r_16_sv2v_reg <= decode_tl_r[16];
      decode_v_r_15_sv2v_reg <= decode_tl_r[15];
      decode_v_r_14_sv2v_reg <= decode_tl_r[14];
      decode_v_r_13_sv2v_reg <= decode_tl_r[13];
      decode_v_r_12_sv2v_reg <= decode_tl_r[12];
      decode_v_r_11_sv2v_reg <= decode_tl_r[11];
      decode_v_r_10_sv2v_reg <= decode_tl_r[10];
      decode_v_r_9_sv2v_reg <= decode_tl_r[9];
      decode_v_r_8_sv2v_reg <= decode_tl_r[8];
      addr_v_r_27_sv2v_reg <= addr_tl_r[27];
      addr_v_r_26_sv2v_reg <= addr_tl_r[26];
      addr_v_r_25_sv2v_reg <= addr_tl_r[25];
      addr_v_r_24_sv2v_reg <= addr_tl_r[24];
      addr_v_r_23_sv2v_reg <= addr_tl_r[23];
      addr_v_r_22_sv2v_reg <= addr_tl_r[22];
      addr_v_r_21_sv2v_reg <= addr_tl_r[21];
      addr_v_r_20_sv2v_reg <= addr_tl_r[20];
      addr_v_r_19_sv2v_reg <= addr_tl_r[19];
      addr_v_r_18_sv2v_reg <= addr_tl_r[18];
      addr_v_r_17_sv2v_reg <= addr_tl_r[17];
      addr_v_r_16_sv2v_reg <= addr_tl_r[16];
      addr_v_r_15_sv2v_reg <= addr_tl_r[15];
      addr_v_r_14_sv2v_reg <= addr_tl_r[14];
      addr_v_r_13_sv2v_reg <= addr_tl_r[13];
      addr_v_r_12_sv2v_reg <= addr_tl_r[12];
      addr_v_r_11_sv2v_reg <= addr_tl_r[11];
      addr_v_r_10_sv2v_reg <= addr_tl_r[10];
      addr_v_r_9_sv2v_reg <= addr_tl_r[9];
      addr_v_r_8_sv2v_reg <= addr_tl_r[8];
      addr_v_r_7_sv2v_reg <= addr_tl_r[7];
      addr_v_r_6_sv2v_reg <= addr_tl_r[6];
      addr_v_r_5_sv2v_reg <= addr_tl_r[5];
      addr_v_r_4_sv2v_reg <= addr_tl_r[4];
      addr_v_r_3_sv2v_reg <= addr_tl_r[3];
      addr_v_r_2_sv2v_reg <= addr_tl_r[2];
      addr_v_r_1_sv2v_reg <= addr_tl_r[1];
      addr_v_r_0_sv2v_reg <= addr_tl_r[0];
      data_v_r_31_sv2v_reg <= data_tl_r[31];
      data_v_r_30_sv2v_reg <= data_tl_r[30];
      data_v_r_29_sv2v_reg <= data_tl_r[29];
      data_v_r_28_sv2v_reg <= data_tl_r[28];
      data_v_r_27_sv2v_reg <= data_tl_r[27];
      data_v_r_26_sv2v_reg <= data_tl_r[26];
      data_v_r_25_sv2v_reg <= data_tl_r[25];
      data_v_r_24_sv2v_reg <= data_tl_r[24];
      data_v_r_23_sv2v_reg <= data_tl_r[23];
      data_v_r_22_sv2v_reg <= data_tl_r[22];
      data_v_r_21_sv2v_reg <= data_tl_r[21];
      data_v_r_20_sv2v_reg <= data_tl_r[20];
      data_v_r_19_sv2v_reg <= data_tl_r[19];
      data_v_r_18_sv2v_reg <= data_tl_r[18];
      data_v_r_17_sv2v_reg <= data_tl_r[17];
      data_v_r_16_sv2v_reg <= data_tl_r[16];
      data_v_r_15_sv2v_reg <= data_tl_r[15];
      data_v_r_14_sv2v_reg <= data_tl_r[14];
      data_v_r_13_sv2v_reg <= data_tl_r[13];
      data_v_r_12_sv2v_reg <= data_tl_r[12];
      data_v_r_11_sv2v_reg <= data_tl_r[11];
      data_v_r_10_sv2v_reg <= data_tl_r[10];
      data_v_r_9_sv2v_reg <= data_tl_r[9];
      data_v_r_8_sv2v_reg <= data_tl_r[8];
      data_v_r_7_sv2v_reg <= data_tl_r[7];
      data_v_r_6_sv2v_reg <= data_tl_r[6];
      data_v_r_5_sv2v_reg <= data_tl_r[5];
      data_v_r_4_sv2v_reg <= data_tl_r[4];
      data_v_r_3_sv2v_reg <= data_tl_r[3];
      data_v_r_2_sv2v_reg <= data_tl_r[2];
      data_v_r_1_sv2v_reg <= data_tl_r[1];
      data_v_r_0_sv2v_reg <= data_tl_r[0];
      valid_v_r_3_sv2v_reg <= tag_mem_data_lo[79];
      valid_v_r_2_sv2v_reg <= tag_mem_data_lo[59];
      valid_v_r_1_sv2v_reg <= tag_mem_data_lo[39];
      valid_v_r_0_sv2v_reg <= tag_mem_data_lo[19];
      tag_v_r_21_sv2v_reg <= tag_mem_data_lo[23];
      tag_v_r_20_sv2v_reg <= tag_mem_data_lo[22];
      tag_v_r_19_sv2v_reg <= tag_mem_data_lo[21];
      tag_v_r_18_sv2v_reg <= tag_mem_data_lo[20];
      tag_v_r_17_sv2v_reg <= tag_mem_data_lo[17];
      tag_v_r_16_sv2v_reg <= tag_mem_data_lo[16];
      tag_v_r_15_sv2v_reg <= tag_mem_data_lo[15];
      tag_v_r_14_sv2v_reg <= tag_mem_data_lo[14];
      tag_v_r_13_sv2v_reg <= tag_mem_data_lo[13];
      tag_v_r_12_sv2v_reg <= tag_mem_data_lo[12];
      tag_v_r_11_sv2v_reg <= tag_mem_data_lo[11];
      tag_v_r_10_sv2v_reg <= tag_mem_data_lo[10];
      tag_v_r_9_sv2v_reg <= tag_mem_data_lo[9];
      tag_v_r_8_sv2v_reg <= tag_mem_data_lo[8];
      tag_v_r_7_sv2v_reg <= tag_mem_data_lo[7];
      tag_v_r_6_sv2v_reg <= tag_mem_data_lo[6];
      tag_v_r_5_sv2v_reg <= tag_mem_data_lo[5];
      tag_v_r_4_sv2v_reg <= tag_mem_data_lo[4];
      tag_v_r_3_sv2v_reg <= tag_mem_data_lo[3];
      tag_v_r_2_sv2v_reg <= tag_mem_data_lo[2];
      tag_v_r_1_sv2v_reg <= tag_mem_data_lo[1];
      tag_v_r_0_sv2v_reg <= tag_mem_data_lo[0];
    end 
    if(reset_i) begin
      mask_v_r_1_sv2v_reg <= 1'b0;
      lock_v_r_3_sv2v_reg <= 1'b0;
      lock_v_r_2_sv2v_reg <= 1'b0;
      lock_v_r_1_sv2v_reg <= 1'b0;
      lock_v_r_0_sv2v_reg <= 1'b0;
      tag_v_r_71_sv2v_reg <= 1'b0;
      tag_v_r_70_sv2v_reg <= 1'b0;
      tag_v_r_69_sv2v_reg <= 1'b0;
      tag_v_r_68_sv2v_reg <= 1'b0;
      tag_v_r_67_sv2v_reg <= 1'b0;
      tag_v_r_66_sv2v_reg <= 1'b0;
      tag_v_r_65_sv2v_reg <= 1'b0;
      tag_v_r_64_sv2v_reg <= 1'b0;
      tag_v_r_63_sv2v_reg <= 1'b0;
      tag_v_r_62_sv2v_reg <= 1'b0;
      tag_v_r_61_sv2v_reg <= 1'b0;
      tag_v_r_60_sv2v_reg <= 1'b0;
      tag_v_r_59_sv2v_reg <= 1'b0;
      tag_v_r_58_sv2v_reg <= 1'b0;
      tag_v_r_57_sv2v_reg <= 1'b0;
      tag_v_r_56_sv2v_reg <= 1'b0;
      tag_v_r_55_sv2v_reg <= 1'b0;
      tag_v_r_54_sv2v_reg <= 1'b0;
      tag_v_r_53_sv2v_reg <= 1'b0;
      tag_v_r_52_sv2v_reg <= 1'b0;
      tag_v_r_51_sv2v_reg <= 1'b0;
      tag_v_r_50_sv2v_reg <= 1'b0;
      tag_v_r_49_sv2v_reg <= 1'b0;
      tag_v_r_48_sv2v_reg <= 1'b0;
      tag_v_r_47_sv2v_reg <= 1'b0;
      tag_v_r_46_sv2v_reg <= 1'b0;
      tag_v_r_45_sv2v_reg <= 1'b0;
      tag_v_r_44_sv2v_reg <= 1'b0;
      tag_v_r_43_sv2v_reg <= 1'b0;
      tag_v_r_42_sv2v_reg <= 1'b0;
      tag_v_r_41_sv2v_reg <= 1'b0;
      tag_v_r_40_sv2v_reg <= 1'b0;
      tag_v_r_39_sv2v_reg <= 1'b0;
      tag_v_r_38_sv2v_reg <= 1'b0;
      tag_v_r_37_sv2v_reg <= 1'b0;
      tag_v_r_36_sv2v_reg <= 1'b0;
      tag_v_r_35_sv2v_reg <= 1'b0;
      tag_v_r_34_sv2v_reg <= 1'b0;
      tag_v_r_33_sv2v_reg <= 1'b0;
      tag_v_r_32_sv2v_reg <= 1'b0;
      tag_v_r_31_sv2v_reg <= 1'b0;
      tag_v_r_30_sv2v_reg <= 1'b0;
      tag_v_r_29_sv2v_reg <= 1'b0;
      tag_v_r_28_sv2v_reg <= 1'b0;
      tag_v_r_27_sv2v_reg <= 1'b0;
      tag_v_r_26_sv2v_reg <= 1'b0;
      tag_v_r_25_sv2v_reg <= 1'b0;
      tag_v_r_24_sv2v_reg <= 1'b0;
      tag_v_r_23_sv2v_reg <= 1'b0;
      tag_v_r_22_sv2v_reg <= 1'b0;
    end else if(N79) begin
      mask_v_r_1_sv2v_reg <= mask_tl_r[1];
      lock_v_r_3_sv2v_reg <= tag_mem_data_lo[78];
      lock_v_r_2_sv2v_reg <= tag_mem_data_lo[58];
      lock_v_r_1_sv2v_reg <= tag_mem_data_lo[38];
      lock_v_r_0_sv2v_reg <= tag_mem_data_lo[18];
      tag_v_r_71_sv2v_reg <= tag_mem_data_lo[77];
      tag_v_r_70_sv2v_reg <= tag_mem_data_lo[76];
      tag_v_r_69_sv2v_reg <= tag_mem_data_lo[75];
      tag_v_r_68_sv2v_reg <= tag_mem_data_lo[74];
      tag_v_r_67_sv2v_reg <= tag_mem_data_lo[73];
      tag_v_r_66_sv2v_reg <= tag_mem_data_lo[72];
      tag_v_r_65_sv2v_reg <= tag_mem_data_lo[71];
      tag_v_r_64_sv2v_reg <= tag_mem_data_lo[70];
      tag_v_r_63_sv2v_reg <= tag_mem_data_lo[69];
      tag_v_r_62_sv2v_reg <= tag_mem_data_lo[68];
      tag_v_r_61_sv2v_reg <= tag_mem_data_lo[67];
      tag_v_r_60_sv2v_reg <= tag_mem_data_lo[66];
      tag_v_r_59_sv2v_reg <= tag_mem_data_lo[65];
      tag_v_r_58_sv2v_reg <= tag_mem_data_lo[64];
      tag_v_r_57_sv2v_reg <= tag_mem_data_lo[63];
      tag_v_r_56_sv2v_reg <= tag_mem_data_lo[62];
      tag_v_r_55_sv2v_reg <= tag_mem_data_lo[61];
      tag_v_r_54_sv2v_reg <= tag_mem_data_lo[60];
      tag_v_r_53_sv2v_reg <= tag_mem_data_lo[57];
      tag_v_r_52_sv2v_reg <= tag_mem_data_lo[56];
      tag_v_r_51_sv2v_reg <= tag_mem_data_lo[55];
      tag_v_r_50_sv2v_reg <= tag_mem_data_lo[54];
      tag_v_r_49_sv2v_reg <= tag_mem_data_lo[53];
      tag_v_r_48_sv2v_reg <= tag_mem_data_lo[52];
      tag_v_r_47_sv2v_reg <= tag_mem_data_lo[51];
      tag_v_r_46_sv2v_reg <= tag_mem_data_lo[50];
      tag_v_r_45_sv2v_reg <= tag_mem_data_lo[49];
      tag_v_r_44_sv2v_reg <= tag_mem_data_lo[48];
      tag_v_r_43_sv2v_reg <= tag_mem_data_lo[47];
      tag_v_r_42_sv2v_reg <= tag_mem_data_lo[46];
      tag_v_r_41_sv2v_reg <= tag_mem_data_lo[45];
      tag_v_r_40_sv2v_reg <= tag_mem_data_lo[44];
      tag_v_r_39_sv2v_reg <= tag_mem_data_lo[43];
      tag_v_r_38_sv2v_reg <= tag_mem_data_lo[42];
      tag_v_r_37_sv2v_reg <= tag_mem_data_lo[41];
      tag_v_r_36_sv2v_reg <= tag_mem_data_lo[40];
      tag_v_r_35_sv2v_reg <= tag_mem_data_lo[37];
      tag_v_r_34_sv2v_reg <= tag_mem_data_lo[36];
      tag_v_r_33_sv2v_reg <= tag_mem_data_lo[35];
      tag_v_r_32_sv2v_reg <= tag_mem_data_lo[34];
      tag_v_r_31_sv2v_reg <= tag_mem_data_lo[33];
      tag_v_r_30_sv2v_reg <= tag_mem_data_lo[32];
      tag_v_r_29_sv2v_reg <= tag_mem_data_lo[31];
      tag_v_r_28_sv2v_reg <= tag_mem_data_lo[30];
      tag_v_r_27_sv2v_reg <= tag_mem_data_lo[29];
      tag_v_r_26_sv2v_reg <= tag_mem_data_lo[28];
      tag_v_r_25_sv2v_reg <= tag_mem_data_lo[27];
      tag_v_r_24_sv2v_reg <= tag_mem_data_lo[26];
      tag_v_r_23_sv2v_reg <= tag_mem_data_lo[25];
      tag_v_r_22_sv2v_reg <= tag_mem_data_lo[24];
    end 
  end


endmodule

