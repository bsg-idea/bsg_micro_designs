

module top
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [1023:0] i;
  input [1023:0] sel_oi_one_hot_i;
  output [1023:0] o;

  bsg_crossbar_o_by_i
  wrapper
  (
    .i(i),
    .sel_oi_one_hot_i(sel_oi_one_hot_i),
    .o(o)
  );


endmodule



module bsg_mux_one_hot_width_p32_els_p32
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [1023:0] data_i;
  input [31:0] sel_one_hot_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959;
  wire [1023:0] data_masked;
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[1];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[1];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[1];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[1];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[1];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[1];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[1];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[1];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[1];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[1];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[1];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[1];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[1];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[1];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[1];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[1];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[1];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[1];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[1];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[1];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[1];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[1];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[1];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[1];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[1];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[1];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[1];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[1];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[1];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[2];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[2];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[2];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[2];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[2];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[2];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[2];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[2];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[2];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[2];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[2];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[2];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[2];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[2];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[2];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[2];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[2];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[2];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[2];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[2];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[2];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[2];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[2];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[2];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[2];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[2];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[2];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[2];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[2];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[2];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[2];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[2];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[3];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[3];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[3];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[3];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[3];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[3];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[3];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[3];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[3];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[3];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[3];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[3];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[3];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[3];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[3];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[3];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[3];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[3];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[3];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[3];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[3];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[3];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[3];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[3];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[3];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[3];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[3];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[3];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[3];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[3];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[3];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[3];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[4];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[4];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[4];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[4];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[4];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[4];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[4];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[4];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[4];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[4];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[4];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[4];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[4];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[4];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[4];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[4];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[4];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[4];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[4];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[4];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[4];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[4];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[4];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[4];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[4];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[4];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[4];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[4];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[4];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[4];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[4];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[4];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[5];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[5];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[5];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[5];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[5];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[5];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[5];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[5];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[5];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[5];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[5];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[5];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[5];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[5];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[5];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[5];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[5];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[5];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[5];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[5];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[5];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[5];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[5];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[5];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[5];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[5];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[5];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[5];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[5];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[5];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[5];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[5];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[6];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[6];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[6];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[6];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[6];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[6];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[6];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[6];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[6];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[6];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[6];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[6];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[6];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[6];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[6];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[6];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[6];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[6];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[6];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[6];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[6];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[6];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[6];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[6];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[6];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[6];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[6];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[6];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[6];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[6];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[6];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[6];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[7];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[7];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[7];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[7];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[7];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[7];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[7];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[7];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[7];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[7];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[7];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[7];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[7];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[7];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[7];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[7];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[7];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[7];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[7];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[7];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[7];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[7];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[7];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[7];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[7];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[7];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[7];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[7];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[7];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[7];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[7];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[7];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[8];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[8];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[8];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[8];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[8];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[8];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[8];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[8];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[8];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[8];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[8];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[8];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[8];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[8];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[8];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[8];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[8];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[8];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[8];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[8];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[8];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[8];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[8];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[8];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[8];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[8];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[8];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[8];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[8];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[8];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[8];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[8];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[9];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[9];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[9];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[9];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[9];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[9];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[9];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[9];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[9];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[9];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[9];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[9];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[9];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[9];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[9];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[9];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[9];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[9];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[9];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[9];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[9];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[9];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[9];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[9];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[9];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[9];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[9];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[9];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[9];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[9];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[9];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[9];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[10];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[10];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[10];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[10];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[10];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[10];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[10];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[10];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[10];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[10];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[10];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[10];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[10];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[10];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[10];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[10];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[10];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[10];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[10];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[10];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[10];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[10];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[10];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[10];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[10];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[10];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[10];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[10];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[10];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[10];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[10];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[10];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[11];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[11];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[11];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[11];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[11];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[11];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[11];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[11];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[11];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[11];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[11];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[11];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[11];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[11];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[11];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[11];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[11];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[11];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[11];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[11];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[11];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[11];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[11];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[11];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[11];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[11];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[11];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[11];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[11];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[11];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[11];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[11];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[12];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[12];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[12];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[12];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[12];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[12];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[12];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[12];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[12];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[12];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[12];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[12];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[12];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[12];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[12];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[12];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[12];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[12];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[12];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[12];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[12];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[12];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[12];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[12];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[12];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[12];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[12];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[12];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[12];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[12];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[12];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[12];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[13];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[13];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[13];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[13];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[13];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[13];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[13];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[13];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[13];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[13];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[13];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[13];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[13];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[13];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[13];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[13];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[13];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[13];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[13];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[13];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[13];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[13];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[13];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[13];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[13];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[13];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[13];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[13];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[13];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[13];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[13];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[13];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[14];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[14];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[14];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[14];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[14];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[14];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[14];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[14];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[14];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[14];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[14];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[14];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[14];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[14];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[14];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[14];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[14];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[14];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[14];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[14];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[14];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[14];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[14];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[14];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[14];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[14];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[14];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[14];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[14];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[14];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[14];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[14];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[15];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[15];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[15];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[15];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[15];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[15];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[15];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[15];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[15];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[15];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[15];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[15];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[15];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[15];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[15];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[15];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[15];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[15];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[15];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[15];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[15];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[15];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[15];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[15];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[15];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[15];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[15];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[15];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[15];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[15];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[15];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[15];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[16];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[16];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[16];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[16];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[16];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[16];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[16];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[16];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[16];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[16];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[16];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[16];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[16];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[16];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[16];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[16];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[16];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[16];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[16];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[16];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[16];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[16];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[16];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[16];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[16];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[16];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[16];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[16];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[16];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[16];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[16];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[16];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[17];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[17];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[17];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[17];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[17];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[17];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[17];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[17];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[17];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[17];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[17];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[17];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[17];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[17];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[17];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[17];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[17];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[17];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[17];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[17];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[17];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[17];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[17];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[17];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[17];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[17];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[17];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[17];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[17];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[17];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[17];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[17];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[18];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[18];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[18];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[18];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[18];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[18];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[18];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[18];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[18];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[18];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[18];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[18];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[18];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[18];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[18];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[18];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[18];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[18];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[18];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[18];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[18];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[18];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[18];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[18];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[18];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[18];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[18];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[18];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[18];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[18];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[18];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[18];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[19];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[19];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[19];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[19];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[19];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[19];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[19];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[19];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[19];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[19];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[19];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[19];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[19];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[19];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[19];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[19];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[19];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[19];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[19];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[19];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[19];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[19];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[19];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[19];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[19];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[19];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[19];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[19];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[19];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[19];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[19];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[19];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[20];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[20];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[20];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[20];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[20];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[20];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[20];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[20];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[20];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[20];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[20];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[20];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[20];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[20];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[20];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[20];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[20];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[20];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[20];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[20];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[20];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[20];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[20];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[20];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[20];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[20];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[20];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[20];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[20];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[20];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[20];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[20];
  assign data_masked[703] = data_i[703] & sel_one_hot_i[21];
  assign data_masked[702] = data_i[702] & sel_one_hot_i[21];
  assign data_masked[701] = data_i[701] & sel_one_hot_i[21];
  assign data_masked[700] = data_i[700] & sel_one_hot_i[21];
  assign data_masked[699] = data_i[699] & sel_one_hot_i[21];
  assign data_masked[698] = data_i[698] & sel_one_hot_i[21];
  assign data_masked[697] = data_i[697] & sel_one_hot_i[21];
  assign data_masked[696] = data_i[696] & sel_one_hot_i[21];
  assign data_masked[695] = data_i[695] & sel_one_hot_i[21];
  assign data_masked[694] = data_i[694] & sel_one_hot_i[21];
  assign data_masked[693] = data_i[693] & sel_one_hot_i[21];
  assign data_masked[692] = data_i[692] & sel_one_hot_i[21];
  assign data_masked[691] = data_i[691] & sel_one_hot_i[21];
  assign data_masked[690] = data_i[690] & sel_one_hot_i[21];
  assign data_masked[689] = data_i[689] & sel_one_hot_i[21];
  assign data_masked[688] = data_i[688] & sel_one_hot_i[21];
  assign data_masked[687] = data_i[687] & sel_one_hot_i[21];
  assign data_masked[686] = data_i[686] & sel_one_hot_i[21];
  assign data_masked[685] = data_i[685] & sel_one_hot_i[21];
  assign data_masked[684] = data_i[684] & sel_one_hot_i[21];
  assign data_masked[683] = data_i[683] & sel_one_hot_i[21];
  assign data_masked[682] = data_i[682] & sel_one_hot_i[21];
  assign data_masked[681] = data_i[681] & sel_one_hot_i[21];
  assign data_masked[680] = data_i[680] & sel_one_hot_i[21];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[21];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[21];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[21];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[21];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[21];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[21];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[21];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[21];
  assign data_masked[735] = data_i[735] & sel_one_hot_i[22];
  assign data_masked[734] = data_i[734] & sel_one_hot_i[22];
  assign data_masked[733] = data_i[733] & sel_one_hot_i[22];
  assign data_masked[732] = data_i[732] & sel_one_hot_i[22];
  assign data_masked[731] = data_i[731] & sel_one_hot_i[22];
  assign data_masked[730] = data_i[730] & sel_one_hot_i[22];
  assign data_masked[729] = data_i[729] & sel_one_hot_i[22];
  assign data_masked[728] = data_i[728] & sel_one_hot_i[22];
  assign data_masked[727] = data_i[727] & sel_one_hot_i[22];
  assign data_masked[726] = data_i[726] & sel_one_hot_i[22];
  assign data_masked[725] = data_i[725] & sel_one_hot_i[22];
  assign data_masked[724] = data_i[724] & sel_one_hot_i[22];
  assign data_masked[723] = data_i[723] & sel_one_hot_i[22];
  assign data_masked[722] = data_i[722] & sel_one_hot_i[22];
  assign data_masked[721] = data_i[721] & sel_one_hot_i[22];
  assign data_masked[720] = data_i[720] & sel_one_hot_i[22];
  assign data_masked[719] = data_i[719] & sel_one_hot_i[22];
  assign data_masked[718] = data_i[718] & sel_one_hot_i[22];
  assign data_masked[717] = data_i[717] & sel_one_hot_i[22];
  assign data_masked[716] = data_i[716] & sel_one_hot_i[22];
  assign data_masked[715] = data_i[715] & sel_one_hot_i[22];
  assign data_masked[714] = data_i[714] & sel_one_hot_i[22];
  assign data_masked[713] = data_i[713] & sel_one_hot_i[22];
  assign data_masked[712] = data_i[712] & sel_one_hot_i[22];
  assign data_masked[711] = data_i[711] & sel_one_hot_i[22];
  assign data_masked[710] = data_i[710] & sel_one_hot_i[22];
  assign data_masked[709] = data_i[709] & sel_one_hot_i[22];
  assign data_masked[708] = data_i[708] & sel_one_hot_i[22];
  assign data_masked[707] = data_i[707] & sel_one_hot_i[22];
  assign data_masked[706] = data_i[706] & sel_one_hot_i[22];
  assign data_masked[705] = data_i[705] & sel_one_hot_i[22];
  assign data_masked[704] = data_i[704] & sel_one_hot_i[22];
  assign data_masked[767] = data_i[767] & sel_one_hot_i[23];
  assign data_masked[766] = data_i[766] & sel_one_hot_i[23];
  assign data_masked[765] = data_i[765] & sel_one_hot_i[23];
  assign data_masked[764] = data_i[764] & sel_one_hot_i[23];
  assign data_masked[763] = data_i[763] & sel_one_hot_i[23];
  assign data_masked[762] = data_i[762] & sel_one_hot_i[23];
  assign data_masked[761] = data_i[761] & sel_one_hot_i[23];
  assign data_masked[760] = data_i[760] & sel_one_hot_i[23];
  assign data_masked[759] = data_i[759] & sel_one_hot_i[23];
  assign data_masked[758] = data_i[758] & sel_one_hot_i[23];
  assign data_masked[757] = data_i[757] & sel_one_hot_i[23];
  assign data_masked[756] = data_i[756] & sel_one_hot_i[23];
  assign data_masked[755] = data_i[755] & sel_one_hot_i[23];
  assign data_masked[754] = data_i[754] & sel_one_hot_i[23];
  assign data_masked[753] = data_i[753] & sel_one_hot_i[23];
  assign data_masked[752] = data_i[752] & sel_one_hot_i[23];
  assign data_masked[751] = data_i[751] & sel_one_hot_i[23];
  assign data_masked[750] = data_i[750] & sel_one_hot_i[23];
  assign data_masked[749] = data_i[749] & sel_one_hot_i[23];
  assign data_masked[748] = data_i[748] & sel_one_hot_i[23];
  assign data_masked[747] = data_i[747] & sel_one_hot_i[23];
  assign data_masked[746] = data_i[746] & sel_one_hot_i[23];
  assign data_masked[745] = data_i[745] & sel_one_hot_i[23];
  assign data_masked[744] = data_i[744] & sel_one_hot_i[23];
  assign data_masked[743] = data_i[743] & sel_one_hot_i[23];
  assign data_masked[742] = data_i[742] & sel_one_hot_i[23];
  assign data_masked[741] = data_i[741] & sel_one_hot_i[23];
  assign data_masked[740] = data_i[740] & sel_one_hot_i[23];
  assign data_masked[739] = data_i[739] & sel_one_hot_i[23];
  assign data_masked[738] = data_i[738] & sel_one_hot_i[23];
  assign data_masked[737] = data_i[737] & sel_one_hot_i[23];
  assign data_masked[736] = data_i[736] & sel_one_hot_i[23];
  assign data_masked[799] = data_i[799] & sel_one_hot_i[24];
  assign data_masked[798] = data_i[798] & sel_one_hot_i[24];
  assign data_masked[797] = data_i[797] & sel_one_hot_i[24];
  assign data_masked[796] = data_i[796] & sel_one_hot_i[24];
  assign data_masked[795] = data_i[795] & sel_one_hot_i[24];
  assign data_masked[794] = data_i[794] & sel_one_hot_i[24];
  assign data_masked[793] = data_i[793] & sel_one_hot_i[24];
  assign data_masked[792] = data_i[792] & sel_one_hot_i[24];
  assign data_masked[791] = data_i[791] & sel_one_hot_i[24];
  assign data_masked[790] = data_i[790] & sel_one_hot_i[24];
  assign data_masked[789] = data_i[789] & sel_one_hot_i[24];
  assign data_masked[788] = data_i[788] & sel_one_hot_i[24];
  assign data_masked[787] = data_i[787] & sel_one_hot_i[24];
  assign data_masked[786] = data_i[786] & sel_one_hot_i[24];
  assign data_masked[785] = data_i[785] & sel_one_hot_i[24];
  assign data_masked[784] = data_i[784] & sel_one_hot_i[24];
  assign data_masked[783] = data_i[783] & sel_one_hot_i[24];
  assign data_masked[782] = data_i[782] & sel_one_hot_i[24];
  assign data_masked[781] = data_i[781] & sel_one_hot_i[24];
  assign data_masked[780] = data_i[780] & sel_one_hot_i[24];
  assign data_masked[779] = data_i[779] & sel_one_hot_i[24];
  assign data_masked[778] = data_i[778] & sel_one_hot_i[24];
  assign data_masked[777] = data_i[777] & sel_one_hot_i[24];
  assign data_masked[776] = data_i[776] & sel_one_hot_i[24];
  assign data_masked[775] = data_i[775] & sel_one_hot_i[24];
  assign data_masked[774] = data_i[774] & sel_one_hot_i[24];
  assign data_masked[773] = data_i[773] & sel_one_hot_i[24];
  assign data_masked[772] = data_i[772] & sel_one_hot_i[24];
  assign data_masked[771] = data_i[771] & sel_one_hot_i[24];
  assign data_masked[770] = data_i[770] & sel_one_hot_i[24];
  assign data_masked[769] = data_i[769] & sel_one_hot_i[24];
  assign data_masked[768] = data_i[768] & sel_one_hot_i[24];
  assign data_masked[831] = data_i[831] & sel_one_hot_i[25];
  assign data_masked[830] = data_i[830] & sel_one_hot_i[25];
  assign data_masked[829] = data_i[829] & sel_one_hot_i[25];
  assign data_masked[828] = data_i[828] & sel_one_hot_i[25];
  assign data_masked[827] = data_i[827] & sel_one_hot_i[25];
  assign data_masked[826] = data_i[826] & sel_one_hot_i[25];
  assign data_masked[825] = data_i[825] & sel_one_hot_i[25];
  assign data_masked[824] = data_i[824] & sel_one_hot_i[25];
  assign data_masked[823] = data_i[823] & sel_one_hot_i[25];
  assign data_masked[822] = data_i[822] & sel_one_hot_i[25];
  assign data_masked[821] = data_i[821] & sel_one_hot_i[25];
  assign data_masked[820] = data_i[820] & sel_one_hot_i[25];
  assign data_masked[819] = data_i[819] & sel_one_hot_i[25];
  assign data_masked[818] = data_i[818] & sel_one_hot_i[25];
  assign data_masked[817] = data_i[817] & sel_one_hot_i[25];
  assign data_masked[816] = data_i[816] & sel_one_hot_i[25];
  assign data_masked[815] = data_i[815] & sel_one_hot_i[25];
  assign data_masked[814] = data_i[814] & sel_one_hot_i[25];
  assign data_masked[813] = data_i[813] & sel_one_hot_i[25];
  assign data_masked[812] = data_i[812] & sel_one_hot_i[25];
  assign data_masked[811] = data_i[811] & sel_one_hot_i[25];
  assign data_masked[810] = data_i[810] & sel_one_hot_i[25];
  assign data_masked[809] = data_i[809] & sel_one_hot_i[25];
  assign data_masked[808] = data_i[808] & sel_one_hot_i[25];
  assign data_masked[807] = data_i[807] & sel_one_hot_i[25];
  assign data_masked[806] = data_i[806] & sel_one_hot_i[25];
  assign data_masked[805] = data_i[805] & sel_one_hot_i[25];
  assign data_masked[804] = data_i[804] & sel_one_hot_i[25];
  assign data_masked[803] = data_i[803] & sel_one_hot_i[25];
  assign data_masked[802] = data_i[802] & sel_one_hot_i[25];
  assign data_masked[801] = data_i[801] & sel_one_hot_i[25];
  assign data_masked[800] = data_i[800] & sel_one_hot_i[25];
  assign data_masked[863] = data_i[863] & sel_one_hot_i[26];
  assign data_masked[862] = data_i[862] & sel_one_hot_i[26];
  assign data_masked[861] = data_i[861] & sel_one_hot_i[26];
  assign data_masked[860] = data_i[860] & sel_one_hot_i[26];
  assign data_masked[859] = data_i[859] & sel_one_hot_i[26];
  assign data_masked[858] = data_i[858] & sel_one_hot_i[26];
  assign data_masked[857] = data_i[857] & sel_one_hot_i[26];
  assign data_masked[856] = data_i[856] & sel_one_hot_i[26];
  assign data_masked[855] = data_i[855] & sel_one_hot_i[26];
  assign data_masked[854] = data_i[854] & sel_one_hot_i[26];
  assign data_masked[853] = data_i[853] & sel_one_hot_i[26];
  assign data_masked[852] = data_i[852] & sel_one_hot_i[26];
  assign data_masked[851] = data_i[851] & sel_one_hot_i[26];
  assign data_masked[850] = data_i[850] & sel_one_hot_i[26];
  assign data_masked[849] = data_i[849] & sel_one_hot_i[26];
  assign data_masked[848] = data_i[848] & sel_one_hot_i[26];
  assign data_masked[847] = data_i[847] & sel_one_hot_i[26];
  assign data_masked[846] = data_i[846] & sel_one_hot_i[26];
  assign data_masked[845] = data_i[845] & sel_one_hot_i[26];
  assign data_masked[844] = data_i[844] & sel_one_hot_i[26];
  assign data_masked[843] = data_i[843] & sel_one_hot_i[26];
  assign data_masked[842] = data_i[842] & sel_one_hot_i[26];
  assign data_masked[841] = data_i[841] & sel_one_hot_i[26];
  assign data_masked[840] = data_i[840] & sel_one_hot_i[26];
  assign data_masked[839] = data_i[839] & sel_one_hot_i[26];
  assign data_masked[838] = data_i[838] & sel_one_hot_i[26];
  assign data_masked[837] = data_i[837] & sel_one_hot_i[26];
  assign data_masked[836] = data_i[836] & sel_one_hot_i[26];
  assign data_masked[835] = data_i[835] & sel_one_hot_i[26];
  assign data_masked[834] = data_i[834] & sel_one_hot_i[26];
  assign data_masked[833] = data_i[833] & sel_one_hot_i[26];
  assign data_masked[832] = data_i[832] & sel_one_hot_i[26];
  assign data_masked[895] = data_i[895] & sel_one_hot_i[27];
  assign data_masked[894] = data_i[894] & sel_one_hot_i[27];
  assign data_masked[893] = data_i[893] & sel_one_hot_i[27];
  assign data_masked[892] = data_i[892] & sel_one_hot_i[27];
  assign data_masked[891] = data_i[891] & sel_one_hot_i[27];
  assign data_masked[890] = data_i[890] & sel_one_hot_i[27];
  assign data_masked[889] = data_i[889] & sel_one_hot_i[27];
  assign data_masked[888] = data_i[888] & sel_one_hot_i[27];
  assign data_masked[887] = data_i[887] & sel_one_hot_i[27];
  assign data_masked[886] = data_i[886] & sel_one_hot_i[27];
  assign data_masked[885] = data_i[885] & sel_one_hot_i[27];
  assign data_masked[884] = data_i[884] & sel_one_hot_i[27];
  assign data_masked[883] = data_i[883] & sel_one_hot_i[27];
  assign data_masked[882] = data_i[882] & sel_one_hot_i[27];
  assign data_masked[881] = data_i[881] & sel_one_hot_i[27];
  assign data_masked[880] = data_i[880] & sel_one_hot_i[27];
  assign data_masked[879] = data_i[879] & sel_one_hot_i[27];
  assign data_masked[878] = data_i[878] & sel_one_hot_i[27];
  assign data_masked[877] = data_i[877] & sel_one_hot_i[27];
  assign data_masked[876] = data_i[876] & sel_one_hot_i[27];
  assign data_masked[875] = data_i[875] & sel_one_hot_i[27];
  assign data_masked[874] = data_i[874] & sel_one_hot_i[27];
  assign data_masked[873] = data_i[873] & sel_one_hot_i[27];
  assign data_masked[872] = data_i[872] & sel_one_hot_i[27];
  assign data_masked[871] = data_i[871] & sel_one_hot_i[27];
  assign data_masked[870] = data_i[870] & sel_one_hot_i[27];
  assign data_masked[869] = data_i[869] & sel_one_hot_i[27];
  assign data_masked[868] = data_i[868] & sel_one_hot_i[27];
  assign data_masked[867] = data_i[867] & sel_one_hot_i[27];
  assign data_masked[866] = data_i[866] & sel_one_hot_i[27];
  assign data_masked[865] = data_i[865] & sel_one_hot_i[27];
  assign data_masked[864] = data_i[864] & sel_one_hot_i[27];
  assign data_masked[927] = data_i[927] & sel_one_hot_i[28];
  assign data_masked[926] = data_i[926] & sel_one_hot_i[28];
  assign data_masked[925] = data_i[925] & sel_one_hot_i[28];
  assign data_masked[924] = data_i[924] & sel_one_hot_i[28];
  assign data_masked[923] = data_i[923] & sel_one_hot_i[28];
  assign data_masked[922] = data_i[922] & sel_one_hot_i[28];
  assign data_masked[921] = data_i[921] & sel_one_hot_i[28];
  assign data_masked[920] = data_i[920] & sel_one_hot_i[28];
  assign data_masked[919] = data_i[919] & sel_one_hot_i[28];
  assign data_masked[918] = data_i[918] & sel_one_hot_i[28];
  assign data_masked[917] = data_i[917] & sel_one_hot_i[28];
  assign data_masked[916] = data_i[916] & sel_one_hot_i[28];
  assign data_masked[915] = data_i[915] & sel_one_hot_i[28];
  assign data_masked[914] = data_i[914] & sel_one_hot_i[28];
  assign data_masked[913] = data_i[913] & sel_one_hot_i[28];
  assign data_masked[912] = data_i[912] & sel_one_hot_i[28];
  assign data_masked[911] = data_i[911] & sel_one_hot_i[28];
  assign data_masked[910] = data_i[910] & sel_one_hot_i[28];
  assign data_masked[909] = data_i[909] & sel_one_hot_i[28];
  assign data_masked[908] = data_i[908] & sel_one_hot_i[28];
  assign data_masked[907] = data_i[907] & sel_one_hot_i[28];
  assign data_masked[906] = data_i[906] & sel_one_hot_i[28];
  assign data_masked[905] = data_i[905] & sel_one_hot_i[28];
  assign data_masked[904] = data_i[904] & sel_one_hot_i[28];
  assign data_masked[903] = data_i[903] & sel_one_hot_i[28];
  assign data_masked[902] = data_i[902] & sel_one_hot_i[28];
  assign data_masked[901] = data_i[901] & sel_one_hot_i[28];
  assign data_masked[900] = data_i[900] & sel_one_hot_i[28];
  assign data_masked[899] = data_i[899] & sel_one_hot_i[28];
  assign data_masked[898] = data_i[898] & sel_one_hot_i[28];
  assign data_masked[897] = data_i[897] & sel_one_hot_i[28];
  assign data_masked[896] = data_i[896] & sel_one_hot_i[28];
  assign data_masked[959] = data_i[959] & sel_one_hot_i[29];
  assign data_masked[958] = data_i[958] & sel_one_hot_i[29];
  assign data_masked[957] = data_i[957] & sel_one_hot_i[29];
  assign data_masked[956] = data_i[956] & sel_one_hot_i[29];
  assign data_masked[955] = data_i[955] & sel_one_hot_i[29];
  assign data_masked[954] = data_i[954] & sel_one_hot_i[29];
  assign data_masked[953] = data_i[953] & sel_one_hot_i[29];
  assign data_masked[952] = data_i[952] & sel_one_hot_i[29];
  assign data_masked[951] = data_i[951] & sel_one_hot_i[29];
  assign data_masked[950] = data_i[950] & sel_one_hot_i[29];
  assign data_masked[949] = data_i[949] & sel_one_hot_i[29];
  assign data_masked[948] = data_i[948] & sel_one_hot_i[29];
  assign data_masked[947] = data_i[947] & sel_one_hot_i[29];
  assign data_masked[946] = data_i[946] & sel_one_hot_i[29];
  assign data_masked[945] = data_i[945] & sel_one_hot_i[29];
  assign data_masked[944] = data_i[944] & sel_one_hot_i[29];
  assign data_masked[943] = data_i[943] & sel_one_hot_i[29];
  assign data_masked[942] = data_i[942] & sel_one_hot_i[29];
  assign data_masked[941] = data_i[941] & sel_one_hot_i[29];
  assign data_masked[940] = data_i[940] & sel_one_hot_i[29];
  assign data_masked[939] = data_i[939] & sel_one_hot_i[29];
  assign data_masked[938] = data_i[938] & sel_one_hot_i[29];
  assign data_masked[937] = data_i[937] & sel_one_hot_i[29];
  assign data_masked[936] = data_i[936] & sel_one_hot_i[29];
  assign data_masked[935] = data_i[935] & sel_one_hot_i[29];
  assign data_masked[934] = data_i[934] & sel_one_hot_i[29];
  assign data_masked[933] = data_i[933] & sel_one_hot_i[29];
  assign data_masked[932] = data_i[932] & sel_one_hot_i[29];
  assign data_masked[931] = data_i[931] & sel_one_hot_i[29];
  assign data_masked[930] = data_i[930] & sel_one_hot_i[29];
  assign data_masked[929] = data_i[929] & sel_one_hot_i[29];
  assign data_masked[928] = data_i[928] & sel_one_hot_i[29];
  assign data_masked[991] = data_i[991] & sel_one_hot_i[30];
  assign data_masked[990] = data_i[990] & sel_one_hot_i[30];
  assign data_masked[989] = data_i[989] & sel_one_hot_i[30];
  assign data_masked[988] = data_i[988] & sel_one_hot_i[30];
  assign data_masked[987] = data_i[987] & sel_one_hot_i[30];
  assign data_masked[986] = data_i[986] & sel_one_hot_i[30];
  assign data_masked[985] = data_i[985] & sel_one_hot_i[30];
  assign data_masked[984] = data_i[984] & sel_one_hot_i[30];
  assign data_masked[983] = data_i[983] & sel_one_hot_i[30];
  assign data_masked[982] = data_i[982] & sel_one_hot_i[30];
  assign data_masked[981] = data_i[981] & sel_one_hot_i[30];
  assign data_masked[980] = data_i[980] & sel_one_hot_i[30];
  assign data_masked[979] = data_i[979] & sel_one_hot_i[30];
  assign data_masked[978] = data_i[978] & sel_one_hot_i[30];
  assign data_masked[977] = data_i[977] & sel_one_hot_i[30];
  assign data_masked[976] = data_i[976] & sel_one_hot_i[30];
  assign data_masked[975] = data_i[975] & sel_one_hot_i[30];
  assign data_masked[974] = data_i[974] & sel_one_hot_i[30];
  assign data_masked[973] = data_i[973] & sel_one_hot_i[30];
  assign data_masked[972] = data_i[972] & sel_one_hot_i[30];
  assign data_masked[971] = data_i[971] & sel_one_hot_i[30];
  assign data_masked[970] = data_i[970] & sel_one_hot_i[30];
  assign data_masked[969] = data_i[969] & sel_one_hot_i[30];
  assign data_masked[968] = data_i[968] & sel_one_hot_i[30];
  assign data_masked[967] = data_i[967] & sel_one_hot_i[30];
  assign data_masked[966] = data_i[966] & sel_one_hot_i[30];
  assign data_masked[965] = data_i[965] & sel_one_hot_i[30];
  assign data_masked[964] = data_i[964] & sel_one_hot_i[30];
  assign data_masked[963] = data_i[963] & sel_one_hot_i[30];
  assign data_masked[962] = data_i[962] & sel_one_hot_i[30];
  assign data_masked[961] = data_i[961] & sel_one_hot_i[30];
  assign data_masked[960] = data_i[960] & sel_one_hot_i[30];
  assign data_masked[1023] = data_i[1023] & sel_one_hot_i[31];
  assign data_masked[1022] = data_i[1022] & sel_one_hot_i[31];
  assign data_masked[1021] = data_i[1021] & sel_one_hot_i[31];
  assign data_masked[1020] = data_i[1020] & sel_one_hot_i[31];
  assign data_masked[1019] = data_i[1019] & sel_one_hot_i[31];
  assign data_masked[1018] = data_i[1018] & sel_one_hot_i[31];
  assign data_masked[1017] = data_i[1017] & sel_one_hot_i[31];
  assign data_masked[1016] = data_i[1016] & sel_one_hot_i[31];
  assign data_masked[1015] = data_i[1015] & sel_one_hot_i[31];
  assign data_masked[1014] = data_i[1014] & sel_one_hot_i[31];
  assign data_masked[1013] = data_i[1013] & sel_one_hot_i[31];
  assign data_masked[1012] = data_i[1012] & sel_one_hot_i[31];
  assign data_masked[1011] = data_i[1011] & sel_one_hot_i[31];
  assign data_masked[1010] = data_i[1010] & sel_one_hot_i[31];
  assign data_masked[1009] = data_i[1009] & sel_one_hot_i[31];
  assign data_masked[1008] = data_i[1008] & sel_one_hot_i[31];
  assign data_masked[1007] = data_i[1007] & sel_one_hot_i[31];
  assign data_masked[1006] = data_i[1006] & sel_one_hot_i[31];
  assign data_masked[1005] = data_i[1005] & sel_one_hot_i[31];
  assign data_masked[1004] = data_i[1004] & sel_one_hot_i[31];
  assign data_masked[1003] = data_i[1003] & sel_one_hot_i[31];
  assign data_masked[1002] = data_i[1002] & sel_one_hot_i[31];
  assign data_masked[1001] = data_i[1001] & sel_one_hot_i[31];
  assign data_masked[1000] = data_i[1000] & sel_one_hot_i[31];
  assign data_masked[999] = data_i[999] & sel_one_hot_i[31];
  assign data_masked[998] = data_i[998] & sel_one_hot_i[31];
  assign data_masked[997] = data_i[997] & sel_one_hot_i[31];
  assign data_masked[996] = data_i[996] & sel_one_hot_i[31];
  assign data_masked[995] = data_i[995] & sel_one_hot_i[31];
  assign data_masked[994] = data_i[994] & sel_one_hot_i[31];
  assign data_masked[993] = data_i[993] & sel_one_hot_i[31];
  assign data_masked[992] = data_i[992] & sel_one_hot_i[31];
  assign data_o[0] = N29 | data_masked[0];
  assign N29 = N28 | data_masked[32];
  assign N28 = N27 | data_masked[64];
  assign N27 = N26 | data_masked[96];
  assign N26 = N25 | data_masked[128];
  assign N25 = N24 | data_masked[160];
  assign N24 = N23 | data_masked[192];
  assign N23 = N22 | data_masked[224];
  assign N22 = N21 | data_masked[256];
  assign N21 = N20 | data_masked[288];
  assign N20 = N19 | data_masked[320];
  assign N19 = N18 | data_masked[352];
  assign N18 = N17 | data_masked[384];
  assign N17 = N16 | data_masked[416];
  assign N16 = N15 | data_masked[448];
  assign N15 = N14 | data_masked[480];
  assign N14 = N13 | data_masked[512];
  assign N13 = N12 | data_masked[544];
  assign N12 = N11 | data_masked[576];
  assign N11 = N10 | data_masked[608];
  assign N10 = N9 | data_masked[640];
  assign N9 = N8 | data_masked[672];
  assign N8 = N7 | data_masked[704];
  assign N7 = N6 | data_masked[736];
  assign N6 = N5 | data_masked[768];
  assign N5 = N4 | data_masked[800];
  assign N4 = N3 | data_masked[832];
  assign N3 = N2 | data_masked[864];
  assign N2 = N1 | data_masked[896];
  assign N1 = N0 | data_masked[928];
  assign N0 = data_masked[992] | data_masked[960];
  assign data_o[1] = N59 | data_masked[1];
  assign N59 = N58 | data_masked[33];
  assign N58 = N57 | data_masked[65];
  assign N57 = N56 | data_masked[97];
  assign N56 = N55 | data_masked[129];
  assign N55 = N54 | data_masked[161];
  assign N54 = N53 | data_masked[193];
  assign N53 = N52 | data_masked[225];
  assign N52 = N51 | data_masked[257];
  assign N51 = N50 | data_masked[289];
  assign N50 = N49 | data_masked[321];
  assign N49 = N48 | data_masked[353];
  assign N48 = N47 | data_masked[385];
  assign N47 = N46 | data_masked[417];
  assign N46 = N45 | data_masked[449];
  assign N45 = N44 | data_masked[481];
  assign N44 = N43 | data_masked[513];
  assign N43 = N42 | data_masked[545];
  assign N42 = N41 | data_masked[577];
  assign N41 = N40 | data_masked[609];
  assign N40 = N39 | data_masked[641];
  assign N39 = N38 | data_masked[673];
  assign N38 = N37 | data_masked[705];
  assign N37 = N36 | data_masked[737];
  assign N36 = N35 | data_masked[769];
  assign N35 = N34 | data_masked[801];
  assign N34 = N33 | data_masked[833];
  assign N33 = N32 | data_masked[865];
  assign N32 = N31 | data_masked[897];
  assign N31 = N30 | data_masked[929];
  assign N30 = data_masked[993] | data_masked[961];
  assign data_o[2] = N89 | data_masked[2];
  assign N89 = N88 | data_masked[34];
  assign N88 = N87 | data_masked[66];
  assign N87 = N86 | data_masked[98];
  assign N86 = N85 | data_masked[130];
  assign N85 = N84 | data_masked[162];
  assign N84 = N83 | data_masked[194];
  assign N83 = N82 | data_masked[226];
  assign N82 = N81 | data_masked[258];
  assign N81 = N80 | data_masked[290];
  assign N80 = N79 | data_masked[322];
  assign N79 = N78 | data_masked[354];
  assign N78 = N77 | data_masked[386];
  assign N77 = N76 | data_masked[418];
  assign N76 = N75 | data_masked[450];
  assign N75 = N74 | data_masked[482];
  assign N74 = N73 | data_masked[514];
  assign N73 = N72 | data_masked[546];
  assign N72 = N71 | data_masked[578];
  assign N71 = N70 | data_masked[610];
  assign N70 = N69 | data_masked[642];
  assign N69 = N68 | data_masked[674];
  assign N68 = N67 | data_masked[706];
  assign N67 = N66 | data_masked[738];
  assign N66 = N65 | data_masked[770];
  assign N65 = N64 | data_masked[802];
  assign N64 = N63 | data_masked[834];
  assign N63 = N62 | data_masked[866];
  assign N62 = N61 | data_masked[898];
  assign N61 = N60 | data_masked[930];
  assign N60 = data_masked[994] | data_masked[962];
  assign data_o[3] = N119 | data_masked[3];
  assign N119 = N118 | data_masked[35];
  assign N118 = N117 | data_masked[67];
  assign N117 = N116 | data_masked[99];
  assign N116 = N115 | data_masked[131];
  assign N115 = N114 | data_masked[163];
  assign N114 = N113 | data_masked[195];
  assign N113 = N112 | data_masked[227];
  assign N112 = N111 | data_masked[259];
  assign N111 = N110 | data_masked[291];
  assign N110 = N109 | data_masked[323];
  assign N109 = N108 | data_masked[355];
  assign N108 = N107 | data_masked[387];
  assign N107 = N106 | data_masked[419];
  assign N106 = N105 | data_masked[451];
  assign N105 = N104 | data_masked[483];
  assign N104 = N103 | data_masked[515];
  assign N103 = N102 | data_masked[547];
  assign N102 = N101 | data_masked[579];
  assign N101 = N100 | data_masked[611];
  assign N100 = N99 | data_masked[643];
  assign N99 = N98 | data_masked[675];
  assign N98 = N97 | data_masked[707];
  assign N97 = N96 | data_masked[739];
  assign N96 = N95 | data_masked[771];
  assign N95 = N94 | data_masked[803];
  assign N94 = N93 | data_masked[835];
  assign N93 = N92 | data_masked[867];
  assign N92 = N91 | data_masked[899];
  assign N91 = N90 | data_masked[931];
  assign N90 = data_masked[995] | data_masked[963];
  assign data_o[4] = N149 | data_masked[4];
  assign N149 = N148 | data_masked[36];
  assign N148 = N147 | data_masked[68];
  assign N147 = N146 | data_masked[100];
  assign N146 = N145 | data_masked[132];
  assign N145 = N144 | data_masked[164];
  assign N144 = N143 | data_masked[196];
  assign N143 = N142 | data_masked[228];
  assign N142 = N141 | data_masked[260];
  assign N141 = N140 | data_masked[292];
  assign N140 = N139 | data_masked[324];
  assign N139 = N138 | data_masked[356];
  assign N138 = N137 | data_masked[388];
  assign N137 = N136 | data_masked[420];
  assign N136 = N135 | data_masked[452];
  assign N135 = N134 | data_masked[484];
  assign N134 = N133 | data_masked[516];
  assign N133 = N132 | data_masked[548];
  assign N132 = N131 | data_masked[580];
  assign N131 = N130 | data_masked[612];
  assign N130 = N129 | data_masked[644];
  assign N129 = N128 | data_masked[676];
  assign N128 = N127 | data_masked[708];
  assign N127 = N126 | data_masked[740];
  assign N126 = N125 | data_masked[772];
  assign N125 = N124 | data_masked[804];
  assign N124 = N123 | data_masked[836];
  assign N123 = N122 | data_masked[868];
  assign N122 = N121 | data_masked[900];
  assign N121 = N120 | data_masked[932];
  assign N120 = data_masked[996] | data_masked[964];
  assign data_o[5] = N179 | data_masked[5];
  assign N179 = N178 | data_masked[37];
  assign N178 = N177 | data_masked[69];
  assign N177 = N176 | data_masked[101];
  assign N176 = N175 | data_masked[133];
  assign N175 = N174 | data_masked[165];
  assign N174 = N173 | data_masked[197];
  assign N173 = N172 | data_masked[229];
  assign N172 = N171 | data_masked[261];
  assign N171 = N170 | data_masked[293];
  assign N170 = N169 | data_masked[325];
  assign N169 = N168 | data_masked[357];
  assign N168 = N167 | data_masked[389];
  assign N167 = N166 | data_masked[421];
  assign N166 = N165 | data_masked[453];
  assign N165 = N164 | data_masked[485];
  assign N164 = N163 | data_masked[517];
  assign N163 = N162 | data_masked[549];
  assign N162 = N161 | data_masked[581];
  assign N161 = N160 | data_masked[613];
  assign N160 = N159 | data_masked[645];
  assign N159 = N158 | data_masked[677];
  assign N158 = N157 | data_masked[709];
  assign N157 = N156 | data_masked[741];
  assign N156 = N155 | data_masked[773];
  assign N155 = N154 | data_masked[805];
  assign N154 = N153 | data_masked[837];
  assign N153 = N152 | data_masked[869];
  assign N152 = N151 | data_masked[901];
  assign N151 = N150 | data_masked[933];
  assign N150 = data_masked[997] | data_masked[965];
  assign data_o[6] = N209 | data_masked[6];
  assign N209 = N208 | data_masked[38];
  assign N208 = N207 | data_masked[70];
  assign N207 = N206 | data_masked[102];
  assign N206 = N205 | data_masked[134];
  assign N205 = N204 | data_masked[166];
  assign N204 = N203 | data_masked[198];
  assign N203 = N202 | data_masked[230];
  assign N202 = N201 | data_masked[262];
  assign N201 = N200 | data_masked[294];
  assign N200 = N199 | data_masked[326];
  assign N199 = N198 | data_masked[358];
  assign N198 = N197 | data_masked[390];
  assign N197 = N196 | data_masked[422];
  assign N196 = N195 | data_masked[454];
  assign N195 = N194 | data_masked[486];
  assign N194 = N193 | data_masked[518];
  assign N193 = N192 | data_masked[550];
  assign N192 = N191 | data_masked[582];
  assign N191 = N190 | data_masked[614];
  assign N190 = N189 | data_masked[646];
  assign N189 = N188 | data_masked[678];
  assign N188 = N187 | data_masked[710];
  assign N187 = N186 | data_masked[742];
  assign N186 = N185 | data_masked[774];
  assign N185 = N184 | data_masked[806];
  assign N184 = N183 | data_masked[838];
  assign N183 = N182 | data_masked[870];
  assign N182 = N181 | data_masked[902];
  assign N181 = N180 | data_masked[934];
  assign N180 = data_masked[998] | data_masked[966];
  assign data_o[7] = N239 | data_masked[7];
  assign N239 = N238 | data_masked[39];
  assign N238 = N237 | data_masked[71];
  assign N237 = N236 | data_masked[103];
  assign N236 = N235 | data_masked[135];
  assign N235 = N234 | data_masked[167];
  assign N234 = N233 | data_masked[199];
  assign N233 = N232 | data_masked[231];
  assign N232 = N231 | data_masked[263];
  assign N231 = N230 | data_masked[295];
  assign N230 = N229 | data_masked[327];
  assign N229 = N228 | data_masked[359];
  assign N228 = N227 | data_masked[391];
  assign N227 = N226 | data_masked[423];
  assign N226 = N225 | data_masked[455];
  assign N225 = N224 | data_masked[487];
  assign N224 = N223 | data_masked[519];
  assign N223 = N222 | data_masked[551];
  assign N222 = N221 | data_masked[583];
  assign N221 = N220 | data_masked[615];
  assign N220 = N219 | data_masked[647];
  assign N219 = N218 | data_masked[679];
  assign N218 = N217 | data_masked[711];
  assign N217 = N216 | data_masked[743];
  assign N216 = N215 | data_masked[775];
  assign N215 = N214 | data_masked[807];
  assign N214 = N213 | data_masked[839];
  assign N213 = N212 | data_masked[871];
  assign N212 = N211 | data_masked[903];
  assign N211 = N210 | data_masked[935];
  assign N210 = data_masked[999] | data_masked[967];
  assign data_o[8] = N269 | data_masked[8];
  assign N269 = N268 | data_masked[40];
  assign N268 = N267 | data_masked[72];
  assign N267 = N266 | data_masked[104];
  assign N266 = N265 | data_masked[136];
  assign N265 = N264 | data_masked[168];
  assign N264 = N263 | data_masked[200];
  assign N263 = N262 | data_masked[232];
  assign N262 = N261 | data_masked[264];
  assign N261 = N260 | data_masked[296];
  assign N260 = N259 | data_masked[328];
  assign N259 = N258 | data_masked[360];
  assign N258 = N257 | data_masked[392];
  assign N257 = N256 | data_masked[424];
  assign N256 = N255 | data_masked[456];
  assign N255 = N254 | data_masked[488];
  assign N254 = N253 | data_masked[520];
  assign N253 = N252 | data_masked[552];
  assign N252 = N251 | data_masked[584];
  assign N251 = N250 | data_masked[616];
  assign N250 = N249 | data_masked[648];
  assign N249 = N248 | data_masked[680];
  assign N248 = N247 | data_masked[712];
  assign N247 = N246 | data_masked[744];
  assign N246 = N245 | data_masked[776];
  assign N245 = N244 | data_masked[808];
  assign N244 = N243 | data_masked[840];
  assign N243 = N242 | data_masked[872];
  assign N242 = N241 | data_masked[904];
  assign N241 = N240 | data_masked[936];
  assign N240 = data_masked[1000] | data_masked[968];
  assign data_o[9] = N299 | data_masked[9];
  assign N299 = N298 | data_masked[41];
  assign N298 = N297 | data_masked[73];
  assign N297 = N296 | data_masked[105];
  assign N296 = N295 | data_masked[137];
  assign N295 = N294 | data_masked[169];
  assign N294 = N293 | data_masked[201];
  assign N293 = N292 | data_masked[233];
  assign N292 = N291 | data_masked[265];
  assign N291 = N290 | data_masked[297];
  assign N290 = N289 | data_masked[329];
  assign N289 = N288 | data_masked[361];
  assign N288 = N287 | data_masked[393];
  assign N287 = N286 | data_masked[425];
  assign N286 = N285 | data_masked[457];
  assign N285 = N284 | data_masked[489];
  assign N284 = N283 | data_masked[521];
  assign N283 = N282 | data_masked[553];
  assign N282 = N281 | data_masked[585];
  assign N281 = N280 | data_masked[617];
  assign N280 = N279 | data_masked[649];
  assign N279 = N278 | data_masked[681];
  assign N278 = N277 | data_masked[713];
  assign N277 = N276 | data_masked[745];
  assign N276 = N275 | data_masked[777];
  assign N275 = N274 | data_masked[809];
  assign N274 = N273 | data_masked[841];
  assign N273 = N272 | data_masked[873];
  assign N272 = N271 | data_masked[905];
  assign N271 = N270 | data_masked[937];
  assign N270 = data_masked[1001] | data_masked[969];
  assign data_o[10] = N329 | data_masked[10];
  assign N329 = N328 | data_masked[42];
  assign N328 = N327 | data_masked[74];
  assign N327 = N326 | data_masked[106];
  assign N326 = N325 | data_masked[138];
  assign N325 = N324 | data_masked[170];
  assign N324 = N323 | data_masked[202];
  assign N323 = N322 | data_masked[234];
  assign N322 = N321 | data_masked[266];
  assign N321 = N320 | data_masked[298];
  assign N320 = N319 | data_masked[330];
  assign N319 = N318 | data_masked[362];
  assign N318 = N317 | data_masked[394];
  assign N317 = N316 | data_masked[426];
  assign N316 = N315 | data_masked[458];
  assign N315 = N314 | data_masked[490];
  assign N314 = N313 | data_masked[522];
  assign N313 = N312 | data_masked[554];
  assign N312 = N311 | data_masked[586];
  assign N311 = N310 | data_masked[618];
  assign N310 = N309 | data_masked[650];
  assign N309 = N308 | data_masked[682];
  assign N308 = N307 | data_masked[714];
  assign N307 = N306 | data_masked[746];
  assign N306 = N305 | data_masked[778];
  assign N305 = N304 | data_masked[810];
  assign N304 = N303 | data_masked[842];
  assign N303 = N302 | data_masked[874];
  assign N302 = N301 | data_masked[906];
  assign N301 = N300 | data_masked[938];
  assign N300 = data_masked[1002] | data_masked[970];
  assign data_o[11] = N359 | data_masked[11];
  assign N359 = N358 | data_masked[43];
  assign N358 = N357 | data_masked[75];
  assign N357 = N356 | data_masked[107];
  assign N356 = N355 | data_masked[139];
  assign N355 = N354 | data_masked[171];
  assign N354 = N353 | data_masked[203];
  assign N353 = N352 | data_masked[235];
  assign N352 = N351 | data_masked[267];
  assign N351 = N350 | data_masked[299];
  assign N350 = N349 | data_masked[331];
  assign N349 = N348 | data_masked[363];
  assign N348 = N347 | data_masked[395];
  assign N347 = N346 | data_masked[427];
  assign N346 = N345 | data_masked[459];
  assign N345 = N344 | data_masked[491];
  assign N344 = N343 | data_masked[523];
  assign N343 = N342 | data_masked[555];
  assign N342 = N341 | data_masked[587];
  assign N341 = N340 | data_masked[619];
  assign N340 = N339 | data_masked[651];
  assign N339 = N338 | data_masked[683];
  assign N338 = N337 | data_masked[715];
  assign N337 = N336 | data_masked[747];
  assign N336 = N335 | data_masked[779];
  assign N335 = N334 | data_masked[811];
  assign N334 = N333 | data_masked[843];
  assign N333 = N332 | data_masked[875];
  assign N332 = N331 | data_masked[907];
  assign N331 = N330 | data_masked[939];
  assign N330 = data_masked[1003] | data_masked[971];
  assign data_o[12] = N389 | data_masked[12];
  assign N389 = N388 | data_masked[44];
  assign N388 = N387 | data_masked[76];
  assign N387 = N386 | data_masked[108];
  assign N386 = N385 | data_masked[140];
  assign N385 = N384 | data_masked[172];
  assign N384 = N383 | data_masked[204];
  assign N383 = N382 | data_masked[236];
  assign N382 = N381 | data_masked[268];
  assign N381 = N380 | data_masked[300];
  assign N380 = N379 | data_masked[332];
  assign N379 = N378 | data_masked[364];
  assign N378 = N377 | data_masked[396];
  assign N377 = N376 | data_masked[428];
  assign N376 = N375 | data_masked[460];
  assign N375 = N374 | data_masked[492];
  assign N374 = N373 | data_masked[524];
  assign N373 = N372 | data_masked[556];
  assign N372 = N371 | data_masked[588];
  assign N371 = N370 | data_masked[620];
  assign N370 = N369 | data_masked[652];
  assign N369 = N368 | data_masked[684];
  assign N368 = N367 | data_masked[716];
  assign N367 = N366 | data_masked[748];
  assign N366 = N365 | data_masked[780];
  assign N365 = N364 | data_masked[812];
  assign N364 = N363 | data_masked[844];
  assign N363 = N362 | data_masked[876];
  assign N362 = N361 | data_masked[908];
  assign N361 = N360 | data_masked[940];
  assign N360 = data_masked[1004] | data_masked[972];
  assign data_o[13] = N419 | data_masked[13];
  assign N419 = N418 | data_masked[45];
  assign N418 = N417 | data_masked[77];
  assign N417 = N416 | data_masked[109];
  assign N416 = N415 | data_masked[141];
  assign N415 = N414 | data_masked[173];
  assign N414 = N413 | data_masked[205];
  assign N413 = N412 | data_masked[237];
  assign N412 = N411 | data_masked[269];
  assign N411 = N410 | data_masked[301];
  assign N410 = N409 | data_masked[333];
  assign N409 = N408 | data_masked[365];
  assign N408 = N407 | data_masked[397];
  assign N407 = N406 | data_masked[429];
  assign N406 = N405 | data_masked[461];
  assign N405 = N404 | data_masked[493];
  assign N404 = N403 | data_masked[525];
  assign N403 = N402 | data_masked[557];
  assign N402 = N401 | data_masked[589];
  assign N401 = N400 | data_masked[621];
  assign N400 = N399 | data_masked[653];
  assign N399 = N398 | data_masked[685];
  assign N398 = N397 | data_masked[717];
  assign N397 = N396 | data_masked[749];
  assign N396 = N395 | data_masked[781];
  assign N395 = N394 | data_masked[813];
  assign N394 = N393 | data_masked[845];
  assign N393 = N392 | data_masked[877];
  assign N392 = N391 | data_masked[909];
  assign N391 = N390 | data_masked[941];
  assign N390 = data_masked[1005] | data_masked[973];
  assign data_o[14] = N449 | data_masked[14];
  assign N449 = N448 | data_masked[46];
  assign N448 = N447 | data_masked[78];
  assign N447 = N446 | data_masked[110];
  assign N446 = N445 | data_masked[142];
  assign N445 = N444 | data_masked[174];
  assign N444 = N443 | data_masked[206];
  assign N443 = N442 | data_masked[238];
  assign N442 = N441 | data_masked[270];
  assign N441 = N440 | data_masked[302];
  assign N440 = N439 | data_masked[334];
  assign N439 = N438 | data_masked[366];
  assign N438 = N437 | data_masked[398];
  assign N437 = N436 | data_masked[430];
  assign N436 = N435 | data_masked[462];
  assign N435 = N434 | data_masked[494];
  assign N434 = N433 | data_masked[526];
  assign N433 = N432 | data_masked[558];
  assign N432 = N431 | data_masked[590];
  assign N431 = N430 | data_masked[622];
  assign N430 = N429 | data_masked[654];
  assign N429 = N428 | data_masked[686];
  assign N428 = N427 | data_masked[718];
  assign N427 = N426 | data_masked[750];
  assign N426 = N425 | data_masked[782];
  assign N425 = N424 | data_masked[814];
  assign N424 = N423 | data_masked[846];
  assign N423 = N422 | data_masked[878];
  assign N422 = N421 | data_masked[910];
  assign N421 = N420 | data_masked[942];
  assign N420 = data_masked[1006] | data_masked[974];
  assign data_o[15] = N479 | data_masked[15];
  assign N479 = N478 | data_masked[47];
  assign N478 = N477 | data_masked[79];
  assign N477 = N476 | data_masked[111];
  assign N476 = N475 | data_masked[143];
  assign N475 = N474 | data_masked[175];
  assign N474 = N473 | data_masked[207];
  assign N473 = N472 | data_masked[239];
  assign N472 = N471 | data_masked[271];
  assign N471 = N470 | data_masked[303];
  assign N470 = N469 | data_masked[335];
  assign N469 = N468 | data_masked[367];
  assign N468 = N467 | data_masked[399];
  assign N467 = N466 | data_masked[431];
  assign N466 = N465 | data_masked[463];
  assign N465 = N464 | data_masked[495];
  assign N464 = N463 | data_masked[527];
  assign N463 = N462 | data_masked[559];
  assign N462 = N461 | data_masked[591];
  assign N461 = N460 | data_masked[623];
  assign N460 = N459 | data_masked[655];
  assign N459 = N458 | data_masked[687];
  assign N458 = N457 | data_masked[719];
  assign N457 = N456 | data_masked[751];
  assign N456 = N455 | data_masked[783];
  assign N455 = N454 | data_masked[815];
  assign N454 = N453 | data_masked[847];
  assign N453 = N452 | data_masked[879];
  assign N452 = N451 | data_masked[911];
  assign N451 = N450 | data_masked[943];
  assign N450 = data_masked[1007] | data_masked[975];
  assign data_o[16] = N509 | data_masked[16];
  assign N509 = N508 | data_masked[48];
  assign N508 = N507 | data_masked[80];
  assign N507 = N506 | data_masked[112];
  assign N506 = N505 | data_masked[144];
  assign N505 = N504 | data_masked[176];
  assign N504 = N503 | data_masked[208];
  assign N503 = N502 | data_masked[240];
  assign N502 = N501 | data_masked[272];
  assign N501 = N500 | data_masked[304];
  assign N500 = N499 | data_masked[336];
  assign N499 = N498 | data_masked[368];
  assign N498 = N497 | data_masked[400];
  assign N497 = N496 | data_masked[432];
  assign N496 = N495 | data_masked[464];
  assign N495 = N494 | data_masked[496];
  assign N494 = N493 | data_masked[528];
  assign N493 = N492 | data_masked[560];
  assign N492 = N491 | data_masked[592];
  assign N491 = N490 | data_masked[624];
  assign N490 = N489 | data_masked[656];
  assign N489 = N488 | data_masked[688];
  assign N488 = N487 | data_masked[720];
  assign N487 = N486 | data_masked[752];
  assign N486 = N485 | data_masked[784];
  assign N485 = N484 | data_masked[816];
  assign N484 = N483 | data_masked[848];
  assign N483 = N482 | data_masked[880];
  assign N482 = N481 | data_masked[912];
  assign N481 = N480 | data_masked[944];
  assign N480 = data_masked[1008] | data_masked[976];
  assign data_o[17] = N539 | data_masked[17];
  assign N539 = N538 | data_masked[49];
  assign N538 = N537 | data_masked[81];
  assign N537 = N536 | data_masked[113];
  assign N536 = N535 | data_masked[145];
  assign N535 = N534 | data_masked[177];
  assign N534 = N533 | data_masked[209];
  assign N533 = N532 | data_masked[241];
  assign N532 = N531 | data_masked[273];
  assign N531 = N530 | data_masked[305];
  assign N530 = N529 | data_masked[337];
  assign N529 = N528 | data_masked[369];
  assign N528 = N527 | data_masked[401];
  assign N527 = N526 | data_masked[433];
  assign N526 = N525 | data_masked[465];
  assign N525 = N524 | data_masked[497];
  assign N524 = N523 | data_masked[529];
  assign N523 = N522 | data_masked[561];
  assign N522 = N521 | data_masked[593];
  assign N521 = N520 | data_masked[625];
  assign N520 = N519 | data_masked[657];
  assign N519 = N518 | data_masked[689];
  assign N518 = N517 | data_masked[721];
  assign N517 = N516 | data_masked[753];
  assign N516 = N515 | data_masked[785];
  assign N515 = N514 | data_masked[817];
  assign N514 = N513 | data_masked[849];
  assign N513 = N512 | data_masked[881];
  assign N512 = N511 | data_masked[913];
  assign N511 = N510 | data_masked[945];
  assign N510 = data_masked[1009] | data_masked[977];
  assign data_o[18] = N569 | data_masked[18];
  assign N569 = N568 | data_masked[50];
  assign N568 = N567 | data_masked[82];
  assign N567 = N566 | data_masked[114];
  assign N566 = N565 | data_masked[146];
  assign N565 = N564 | data_masked[178];
  assign N564 = N563 | data_masked[210];
  assign N563 = N562 | data_masked[242];
  assign N562 = N561 | data_masked[274];
  assign N561 = N560 | data_masked[306];
  assign N560 = N559 | data_masked[338];
  assign N559 = N558 | data_masked[370];
  assign N558 = N557 | data_masked[402];
  assign N557 = N556 | data_masked[434];
  assign N556 = N555 | data_masked[466];
  assign N555 = N554 | data_masked[498];
  assign N554 = N553 | data_masked[530];
  assign N553 = N552 | data_masked[562];
  assign N552 = N551 | data_masked[594];
  assign N551 = N550 | data_masked[626];
  assign N550 = N549 | data_masked[658];
  assign N549 = N548 | data_masked[690];
  assign N548 = N547 | data_masked[722];
  assign N547 = N546 | data_masked[754];
  assign N546 = N545 | data_masked[786];
  assign N545 = N544 | data_masked[818];
  assign N544 = N543 | data_masked[850];
  assign N543 = N542 | data_masked[882];
  assign N542 = N541 | data_masked[914];
  assign N541 = N540 | data_masked[946];
  assign N540 = data_masked[1010] | data_masked[978];
  assign data_o[19] = N599 | data_masked[19];
  assign N599 = N598 | data_masked[51];
  assign N598 = N597 | data_masked[83];
  assign N597 = N596 | data_masked[115];
  assign N596 = N595 | data_masked[147];
  assign N595 = N594 | data_masked[179];
  assign N594 = N593 | data_masked[211];
  assign N593 = N592 | data_masked[243];
  assign N592 = N591 | data_masked[275];
  assign N591 = N590 | data_masked[307];
  assign N590 = N589 | data_masked[339];
  assign N589 = N588 | data_masked[371];
  assign N588 = N587 | data_masked[403];
  assign N587 = N586 | data_masked[435];
  assign N586 = N585 | data_masked[467];
  assign N585 = N584 | data_masked[499];
  assign N584 = N583 | data_masked[531];
  assign N583 = N582 | data_masked[563];
  assign N582 = N581 | data_masked[595];
  assign N581 = N580 | data_masked[627];
  assign N580 = N579 | data_masked[659];
  assign N579 = N578 | data_masked[691];
  assign N578 = N577 | data_masked[723];
  assign N577 = N576 | data_masked[755];
  assign N576 = N575 | data_masked[787];
  assign N575 = N574 | data_masked[819];
  assign N574 = N573 | data_masked[851];
  assign N573 = N572 | data_masked[883];
  assign N572 = N571 | data_masked[915];
  assign N571 = N570 | data_masked[947];
  assign N570 = data_masked[1011] | data_masked[979];
  assign data_o[20] = N629 | data_masked[20];
  assign N629 = N628 | data_masked[52];
  assign N628 = N627 | data_masked[84];
  assign N627 = N626 | data_masked[116];
  assign N626 = N625 | data_masked[148];
  assign N625 = N624 | data_masked[180];
  assign N624 = N623 | data_masked[212];
  assign N623 = N622 | data_masked[244];
  assign N622 = N621 | data_masked[276];
  assign N621 = N620 | data_masked[308];
  assign N620 = N619 | data_masked[340];
  assign N619 = N618 | data_masked[372];
  assign N618 = N617 | data_masked[404];
  assign N617 = N616 | data_masked[436];
  assign N616 = N615 | data_masked[468];
  assign N615 = N614 | data_masked[500];
  assign N614 = N613 | data_masked[532];
  assign N613 = N612 | data_masked[564];
  assign N612 = N611 | data_masked[596];
  assign N611 = N610 | data_masked[628];
  assign N610 = N609 | data_masked[660];
  assign N609 = N608 | data_masked[692];
  assign N608 = N607 | data_masked[724];
  assign N607 = N606 | data_masked[756];
  assign N606 = N605 | data_masked[788];
  assign N605 = N604 | data_masked[820];
  assign N604 = N603 | data_masked[852];
  assign N603 = N602 | data_masked[884];
  assign N602 = N601 | data_masked[916];
  assign N601 = N600 | data_masked[948];
  assign N600 = data_masked[1012] | data_masked[980];
  assign data_o[21] = N659 | data_masked[21];
  assign N659 = N658 | data_masked[53];
  assign N658 = N657 | data_masked[85];
  assign N657 = N656 | data_masked[117];
  assign N656 = N655 | data_masked[149];
  assign N655 = N654 | data_masked[181];
  assign N654 = N653 | data_masked[213];
  assign N653 = N652 | data_masked[245];
  assign N652 = N651 | data_masked[277];
  assign N651 = N650 | data_masked[309];
  assign N650 = N649 | data_masked[341];
  assign N649 = N648 | data_masked[373];
  assign N648 = N647 | data_masked[405];
  assign N647 = N646 | data_masked[437];
  assign N646 = N645 | data_masked[469];
  assign N645 = N644 | data_masked[501];
  assign N644 = N643 | data_masked[533];
  assign N643 = N642 | data_masked[565];
  assign N642 = N641 | data_masked[597];
  assign N641 = N640 | data_masked[629];
  assign N640 = N639 | data_masked[661];
  assign N639 = N638 | data_masked[693];
  assign N638 = N637 | data_masked[725];
  assign N637 = N636 | data_masked[757];
  assign N636 = N635 | data_masked[789];
  assign N635 = N634 | data_masked[821];
  assign N634 = N633 | data_masked[853];
  assign N633 = N632 | data_masked[885];
  assign N632 = N631 | data_masked[917];
  assign N631 = N630 | data_masked[949];
  assign N630 = data_masked[1013] | data_masked[981];
  assign data_o[22] = N689 | data_masked[22];
  assign N689 = N688 | data_masked[54];
  assign N688 = N687 | data_masked[86];
  assign N687 = N686 | data_masked[118];
  assign N686 = N685 | data_masked[150];
  assign N685 = N684 | data_masked[182];
  assign N684 = N683 | data_masked[214];
  assign N683 = N682 | data_masked[246];
  assign N682 = N681 | data_masked[278];
  assign N681 = N680 | data_masked[310];
  assign N680 = N679 | data_masked[342];
  assign N679 = N678 | data_masked[374];
  assign N678 = N677 | data_masked[406];
  assign N677 = N676 | data_masked[438];
  assign N676 = N675 | data_masked[470];
  assign N675 = N674 | data_masked[502];
  assign N674 = N673 | data_masked[534];
  assign N673 = N672 | data_masked[566];
  assign N672 = N671 | data_masked[598];
  assign N671 = N670 | data_masked[630];
  assign N670 = N669 | data_masked[662];
  assign N669 = N668 | data_masked[694];
  assign N668 = N667 | data_masked[726];
  assign N667 = N666 | data_masked[758];
  assign N666 = N665 | data_masked[790];
  assign N665 = N664 | data_masked[822];
  assign N664 = N663 | data_masked[854];
  assign N663 = N662 | data_masked[886];
  assign N662 = N661 | data_masked[918];
  assign N661 = N660 | data_masked[950];
  assign N660 = data_masked[1014] | data_masked[982];
  assign data_o[23] = N719 | data_masked[23];
  assign N719 = N718 | data_masked[55];
  assign N718 = N717 | data_masked[87];
  assign N717 = N716 | data_masked[119];
  assign N716 = N715 | data_masked[151];
  assign N715 = N714 | data_masked[183];
  assign N714 = N713 | data_masked[215];
  assign N713 = N712 | data_masked[247];
  assign N712 = N711 | data_masked[279];
  assign N711 = N710 | data_masked[311];
  assign N710 = N709 | data_masked[343];
  assign N709 = N708 | data_masked[375];
  assign N708 = N707 | data_masked[407];
  assign N707 = N706 | data_masked[439];
  assign N706 = N705 | data_masked[471];
  assign N705 = N704 | data_masked[503];
  assign N704 = N703 | data_masked[535];
  assign N703 = N702 | data_masked[567];
  assign N702 = N701 | data_masked[599];
  assign N701 = N700 | data_masked[631];
  assign N700 = N699 | data_masked[663];
  assign N699 = N698 | data_masked[695];
  assign N698 = N697 | data_masked[727];
  assign N697 = N696 | data_masked[759];
  assign N696 = N695 | data_masked[791];
  assign N695 = N694 | data_masked[823];
  assign N694 = N693 | data_masked[855];
  assign N693 = N692 | data_masked[887];
  assign N692 = N691 | data_masked[919];
  assign N691 = N690 | data_masked[951];
  assign N690 = data_masked[1015] | data_masked[983];
  assign data_o[24] = N749 | data_masked[24];
  assign N749 = N748 | data_masked[56];
  assign N748 = N747 | data_masked[88];
  assign N747 = N746 | data_masked[120];
  assign N746 = N745 | data_masked[152];
  assign N745 = N744 | data_masked[184];
  assign N744 = N743 | data_masked[216];
  assign N743 = N742 | data_masked[248];
  assign N742 = N741 | data_masked[280];
  assign N741 = N740 | data_masked[312];
  assign N740 = N739 | data_masked[344];
  assign N739 = N738 | data_masked[376];
  assign N738 = N737 | data_masked[408];
  assign N737 = N736 | data_masked[440];
  assign N736 = N735 | data_masked[472];
  assign N735 = N734 | data_masked[504];
  assign N734 = N733 | data_masked[536];
  assign N733 = N732 | data_masked[568];
  assign N732 = N731 | data_masked[600];
  assign N731 = N730 | data_masked[632];
  assign N730 = N729 | data_masked[664];
  assign N729 = N728 | data_masked[696];
  assign N728 = N727 | data_masked[728];
  assign N727 = N726 | data_masked[760];
  assign N726 = N725 | data_masked[792];
  assign N725 = N724 | data_masked[824];
  assign N724 = N723 | data_masked[856];
  assign N723 = N722 | data_masked[888];
  assign N722 = N721 | data_masked[920];
  assign N721 = N720 | data_masked[952];
  assign N720 = data_masked[1016] | data_masked[984];
  assign data_o[25] = N779 | data_masked[25];
  assign N779 = N778 | data_masked[57];
  assign N778 = N777 | data_masked[89];
  assign N777 = N776 | data_masked[121];
  assign N776 = N775 | data_masked[153];
  assign N775 = N774 | data_masked[185];
  assign N774 = N773 | data_masked[217];
  assign N773 = N772 | data_masked[249];
  assign N772 = N771 | data_masked[281];
  assign N771 = N770 | data_masked[313];
  assign N770 = N769 | data_masked[345];
  assign N769 = N768 | data_masked[377];
  assign N768 = N767 | data_masked[409];
  assign N767 = N766 | data_masked[441];
  assign N766 = N765 | data_masked[473];
  assign N765 = N764 | data_masked[505];
  assign N764 = N763 | data_masked[537];
  assign N763 = N762 | data_masked[569];
  assign N762 = N761 | data_masked[601];
  assign N761 = N760 | data_masked[633];
  assign N760 = N759 | data_masked[665];
  assign N759 = N758 | data_masked[697];
  assign N758 = N757 | data_masked[729];
  assign N757 = N756 | data_masked[761];
  assign N756 = N755 | data_masked[793];
  assign N755 = N754 | data_masked[825];
  assign N754 = N753 | data_masked[857];
  assign N753 = N752 | data_masked[889];
  assign N752 = N751 | data_masked[921];
  assign N751 = N750 | data_masked[953];
  assign N750 = data_masked[1017] | data_masked[985];
  assign data_o[26] = N809 | data_masked[26];
  assign N809 = N808 | data_masked[58];
  assign N808 = N807 | data_masked[90];
  assign N807 = N806 | data_masked[122];
  assign N806 = N805 | data_masked[154];
  assign N805 = N804 | data_masked[186];
  assign N804 = N803 | data_masked[218];
  assign N803 = N802 | data_masked[250];
  assign N802 = N801 | data_masked[282];
  assign N801 = N800 | data_masked[314];
  assign N800 = N799 | data_masked[346];
  assign N799 = N798 | data_masked[378];
  assign N798 = N797 | data_masked[410];
  assign N797 = N796 | data_masked[442];
  assign N796 = N795 | data_masked[474];
  assign N795 = N794 | data_masked[506];
  assign N794 = N793 | data_masked[538];
  assign N793 = N792 | data_masked[570];
  assign N792 = N791 | data_masked[602];
  assign N791 = N790 | data_masked[634];
  assign N790 = N789 | data_masked[666];
  assign N789 = N788 | data_masked[698];
  assign N788 = N787 | data_masked[730];
  assign N787 = N786 | data_masked[762];
  assign N786 = N785 | data_masked[794];
  assign N785 = N784 | data_masked[826];
  assign N784 = N783 | data_masked[858];
  assign N783 = N782 | data_masked[890];
  assign N782 = N781 | data_masked[922];
  assign N781 = N780 | data_masked[954];
  assign N780 = data_masked[1018] | data_masked[986];
  assign data_o[27] = N839 | data_masked[27];
  assign N839 = N838 | data_masked[59];
  assign N838 = N837 | data_masked[91];
  assign N837 = N836 | data_masked[123];
  assign N836 = N835 | data_masked[155];
  assign N835 = N834 | data_masked[187];
  assign N834 = N833 | data_masked[219];
  assign N833 = N832 | data_masked[251];
  assign N832 = N831 | data_masked[283];
  assign N831 = N830 | data_masked[315];
  assign N830 = N829 | data_masked[347];
  assign N829 = N828 | data_masked[379];
  assign N828 = N827 | data_masked[411];
  assign N827 = N826 | data_masked[443];
  assign N826 = N825 | data_masked[475];
  assign N825 = N824 | data_masked[507];
  assign N824 = N823 | data_masked[539];
  assign N823 = N822 | data_masked[571];
  assign N822 = N821 | data_masked[603];
  assign N821 = N820 | data_masked[635];
  assign N820 = N819 | data_masked[667];
  assign N819 = N818 | data_masked[699];
  assign N818 = N817 | data_masked[731];
  assign N817 = N816 | data_masked[763];
  assign N816 = N815 | data_masked[795];
  assign N815 = N814 | data_masked[827];
  assign N814 = N813 | data_masked[859];
  assign N813 = N812 | data_masked[891];
  assign N812 = N811 | data_masked[923];
  assign N811 = N810 | data_masked[955];
  assign N810 = data_masked[1019] | data_masked[987];
  assign data_o[28] = N869 | data_masked[28];
  assign N869 = N868 | data_masked[60];
  assign N868 = N867 | data_masked[92];
  assign N867 = N866 | data_masked[124];
  assign N866 = N865 | data_masked[156];
  assign N865 = N864 | data_masked[188];
  assign N864 = N863 | data_masked[220];
  assign N863 = N862 | data_masked[252];
  assign N862 = N861 | data_masked[284];
  assign N861 = N860 | data_masked[316];
  assign N860 = N859 | data_masked[348];
  assign N859 = N858 | data_masked[380];
  assign N858 = N857 | data_masked[412];
  assign N857 = N856 | data_masked[444];
  assign N856 = N855 | data_masked[476];
  assign N855 = N854 | data_masked[508];
  assign N854 = N853 | data_masked[540];
  assign N853 = N852 | data_masked[572];
  assign N852 = N851 | data_masked[604];
  assign N851 = N850 | data_masked[636];
  assign N850 = N849 | data_masked[668];
  assign N849 = N848 | data_masked[700];
  assign N848 = N847 | data_masked[732];
  assign N847 = N846 | data_masked[764];
  assign N846 = N845 | data_masked[796];
  assign N845 = N844 | data_masked[828];
  assign N844 = N843 | data_masked[860];
  assign N843 = N842 | data_masked[892];
  assign N842 = N841 | data_masked[924];
  assign N841 = N840 | data_masked[956];
  assign N840 = data_masked[1020] | data_masked[988];
  assign data_o[29] = N899 | data_masked[29];
  assign N899 = N898 | data_masked[61];
  assign N898 = N897 | data_masked[93];
  assign N897 = N896 | data_masked[125];
  assign N896 = N895 | data_masked[157];
  assign N895 = N894 | data_masked[189];
  assign N894 = N893 | data_masked[221];
  assign N893 = N892 | data_masked[253];
  assign N892 = N891 | data_masked[285];
  assign N891 = N890 | data_masked[317];
  assign N890 = N889 | data_masked[349];
  assign N889 = N888 | data_masked[381];
  assign N888 = N887 | data_masked[413];
  assign N887 = N886 | data_masked[445];
  assign N886 = N885 | data_masked[477];
  assign N885 = N884 | data_masked[509];
  assign N884 = N883 | data_masked[541];
  assign N883 = N882 | data_masked[573];
  assign N882 = N881 | data_masked[605];
  assign N881 = N880 | data_masked[637];
  assign N880 = N879 | data_masked[669];
  assign N879 = N878 | data_masked[701];
  assign N878 = N877 | data_masked[733];
  assign N877 = N876 | data_masked[765];
  assign N876 = N875 | data_masked[797];
  assign N875 = N874 | data_masked[829];
  assign N874 = N873 | data_masked[861];
  assign N873 = N872 | data_masked[893];
  assign N872 = N871 | data_masked[925];
  assign N871 = N870 | data_masked[957];
  assign N870 = data_masked[1021] | data_masked[989];
  assign data_o[30] = N929 | data_masked[30];
  assign N929 = N928 | data_masked[62];
  assign N928 = N927 | data_masked[94];
  assign N927 = N926 | data_masked[126];
  assign N926 = N925 | data_masked[158];
  assign N925 = N924 | data_masked[190];
  assign N924 = N923 | data_masked[222];
  assign N923 = N922 | data_masked[254];
  assign N922 = N921 | data_masked[286];
  assign N921 = N920 | data_masked[318];
  assign N920 = N919 | data_masked[350];
  assign N919 = N918 | data_masked[382];
  assign N918 = N917 | data_masked[414];
  assign N917 = N916 | data_masked[446];
  assign N916 = N915 | data_masked[478];
  assign N915 = N914 | data_masked[510];
  assign N914 = N913 | data_masked[542];
  assign N913 = N912 | data_masked[574];
  assign N912 = N911 | data_masked[606];
  assign N911 = N910 | data_masked[638];
  assign N910 = N909 | data_masked[670];
  assign N909 = N908 | data_masked[702];
  assign N908 = N907 | data_masked[734];
  assign N907 = N906 | data_masked[766];
  assign N906 = N905 | data_masked[798];
  assign N905 = N904 | data_masked[830];
  assign N904 = N903 | data_masked[862];
  assign N903 = N902 | data_masked[894];
  assign N902 = N901 | data_masked[926];
  assign N901 = N900 | data_masked[958];
  assign N900 = data_masked[1022] | data_masked[990];
  assign data_o[31] = N959 | data_masked[31];
  assign N959 = N958 | data_masked[63];
  assign N958 = N957 | data_masked[95];
  assign N957 = N956 | data_masked[127];
  assign N956 = N955 | data_masked[159];
  assign N955 = N954 | data_masked[191];
  assign N954 = N953 | data_masked[223];
  assign N953 = N952 | data_masked[255];
  assign N952 = N951 | data_masked[287];
  assign N951 = N950 | data_masked[319];
  assign N950 = N949 | data_masked[351];
  assign N949 = N948 | data_masked[383];
  assign N948 = N947 | data_masked[415];
  assign N947 = N946 | data_masked[447];
  assign N946 = N945 | data_masked[479];
  assign N945 = N944 | data_masked[511];
  assign N944 = N943 | data_masked[543];
  assign N943 = N942 | data_masked[575];
  assign N942 = N941 | data_masked[607];
  assign N941 = N940 | data_masked[639];
  assign N940 = N939 | data_masked[671];
  assign N939 = N938 | data_masked[703];
  assign N938 = N937 | data_masked[735];
  assign N937 = N936 | data_masked[767];
  assign N936 = N935 | data_masked[799];
  assign N935 = N934 | data_masked[831];
  assign N934 = N933 | data_masked[863];
  assign N933 = N932 | data_masked[895];
  assign N932 = N931 | data_masked[927];
  assign N931 = N930 | data_masked[959];
  assign N930 = data_masked[1023] | data_masked[991];

endmodule



module bsg_crossbar_o_by_i
(
  i,
  sel_oi_one_hot_i,
  o
);

  input [1023:0] i;
  input [1023:0] sel_oi_one_hot_i;
  output [1023:0] o;
  wire [1023:0] o;

  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_0_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[31:0]),
    .data_o(o[31:0])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_1_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[63:32]),
    .data_o(o[63:32])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_2_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[95:64]),
    .data_o(o[95:64])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_3_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[127:96]),
    .data_o(o[127:96])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_4_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[159:128]),
    .data_o(o[159:128])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_5_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[191:160]),
    .data_o(o[191:160])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_6_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[223:192]),
    .data_o(o[223:192])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_7_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[255:224]),
    .data_o(o[255:224])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_8_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[287:256]),
    .data_o(o[287:256])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_9_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[319:288]),
    .data_o(o[319:288])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_10_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[351:320]),
    .data_o(o[351:320])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_11_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[383:352]),
    .data_o(o[383:352])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_12_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[415:384]),
    .data_o(o[415:384])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_13_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[447:416]),
    .data_o(o[447:416])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_14_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[479:448]),
    .data_o(o[479:448])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_15_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[511:480]),
    .data_o(o[511:480])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_16_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[543:512]),
    .data_o(o[543:512])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_17_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[575:544]),
    .data_o(o[575:544])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_18_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[607:576]),
    .data_o(o[607:576])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_19_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[639:608]),
    .data_o(o[639:608])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_20_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[671:640]),
    .data_o(o[671:640])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_21_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[703:672]),
    .data_o(o[703:672])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_22_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[735:704]),
    .data_o(o[735:704])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_23_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[767:736]),
    .data_o(o[767:736])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_24_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[799:768]),
    .data_o(o[799:768])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_25_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[831:800]),
    .data_o(o[831:800])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_26_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[863:832]),
    .data_o(o[863:832])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_27_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[895:864]),
    .data_o(o[895:864])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_28_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[927:896]),
    .data_o(o[927:896])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_29_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[959:928]),
    .data_o(o[959:928])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_30_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[991:960]),
    .data_o(o[991:960])
  );


  bsg_mux_one_hot_width_p32_els_p32
  \genblk1_31_.mux_one_hot 
  (
    .data_i(i),
    .sel_one_hot_i(sel_oi_one_hot_i[1023:992]),
    .data_o(o[1023:992])
  );


endmodule

