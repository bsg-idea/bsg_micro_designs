

module top
(
  clk_i,
  reset_i,
  v_i,
  len_i,
  data_i,
  ready_o,
  v_o,
  len_v_o,
  data_o,
  yumi_i
);

  input [5:0] len_i;
  input [1599:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output len_v_o;

  bsg_parallel_in_serial_out_dynamic
  wrapper
  (
    .len_i(len_i),
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .v_o(v_o),
    .len_v_o(len_v_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p6_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [5:0] w_data_i;
  input [0:0] r_addr_i;
  output [5:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [5:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [11:0] mem;
  reg mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,
  mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,
  mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[11] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[10] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[9] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[8] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[7] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[6] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      mem_11_sv2v_reg <= w_data_i[5];
      mem_10_sv2v_reg <= w_data_i[4];
      mem_9_sv2v_reg <= w_data_i[3];
      mem_8_sv2v_reg <= w_data_i[2];
      mem_7_sv2v_reg <= w_data_i[1];
      mem_6_sv2v_reg <= w_data_i[0];
    end 
    if(N7) begin
      mem_5_sv2v_reg <= w_data_i[5];
      mem_4_sv2v_reg <= w_data_i[4];
      mem_3_sv2v_reg <= w_data_i[3];
      mem_2_sv2v_reg <= w_data_i[2];
      mem_1_sv2v_reg <= w_data_i[1];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p6_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [5:0] w_data_i;
  input [0:0] r_addr_i;
  output [5:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [5:0] r_data_o;

  bsg_mem_1r1w_synth_width_p6_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p6
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [5:0] data_i;
  output [5:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [5:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p6_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p1600_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [1599:0] w_data_i;
  input [0:0] r_addr_i;
  output [1599:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [1599:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38;
  wire [3199:0] mem;
  reg mem_3199_sv2v_reg,mem_3198_sv2v_reg,mem_3197_sv2v_reg,mem_3196_sv2v_reg,
  mem_3195_sv2v_reg,mem_3194_sv2v_reg,mem_3193_sv2v_reg,mem_3192_sv2v_reg,
  mem_3191_sv2v_reg,mem_3190_sv2v_reg,mem_3189_sv2v_reg,mem_3188_sv2v_reg,mem_3187_sv2v_reg,
  mem_3186_sv2v_reg,mem_3185_sv2v_reg,mem_3184_sv2v_reg,mem_3183_sv2v_reg,
  mem_3182_sv2v_reg,mem_3181_sv2v_reg,mem_3180_sv2v_reg,mem_3179_sv2v_reg,mem_3178_sv2v_reg,
  mem_3177_sv2v_reg,mem_3176_sv2v_reg,mem_3175_sv2v_reg,mem_3174_sv2v_reg,
  mem_3173_sv2v_reg,mem_3172_sv2v_reg,mem_3171_sv2v_reg,mem_3170_sv2v_reg,mem_3169_sv2v_reg,
  mem_3168_sv2v_reg,mem_3167_sv2v_reg,mem_3166_sv2v_reg,mem_3165_sv2v_reg,
  mem_3164_sv2v_reg,mem_3163_sv2v_reg,mem_3162_sv2v_reg,mem_3161_sv2v_reg,mem_3160_sv2v_reg,
  mem_3159_sv2v_reg,mem_3158_sv2v_reg,mem_3157_sv2v_reg,mem_3156_sv2v_reg,
  mem_3155_sv2v_reg,mem_3154_sv2v_reg,mem_3153_sv2v_reg,mem_3152_sv2v_reg,
  mem_3151_sv2v_reg,mem_3150_sv2v_reg,mem_3149_sv2v_reg,mem_3148_sv2v_reg,mem_3147_sv2v_reg,
  mem_3146_sv2v_reg,mem_3145_sv2v_reg,mem_3144_sv2v_reg,mem_3143_sv2v_reg,
  mem_3142_sv2v_reg,mem_3141_sv2v_reg,mem_3140_sv2v_reg,mem_3139_sv2v_reg,mem_3138_sv2v_reg,
  mem_3137_sv2v_reg,mem_3136_sv2v_reg,mem_3135_sv2v_reg,mem_3134_sv2v_reg,
  mem_3133_sv2v_reg,mem_3132_sv2v_reg,mem_3131_sv2v_reg,mem_3130_sv2v_reg,mem_3129_sv2v_reg,
  mem_3128_sv2v_reg,mem_3127_sv2v_reg,mem_3126_sv2v_reg,mem_3125_sv2v_reg,
  mem_3124_sv2v_reg,mem_3123_sv2v_reg,mem_3122_sv2v_reg,mem_3121_sv2v_reg,mem_3120_sv2v_reg,
  mem_3119_sv2v_reg,mem_3118_sv2v_reg,mem_3117_sv2v_reg,mem_3116_sv2v_reg,
  mem_3115_sv2v_reg,mem_3114_sv2v_reg,mem_3113_sv2v_reg,mem_3112_sv2v_reg,
  mem_3111_sv2v_reg,mem_3110_sv2v_reg,mem_3109_sv2v_reg,mem_3108_sv2v_reg,mem_3107_sv2v_reg,
  mem_3106_sv2v_reg,mem_3105_sv2v_reg,mem_3104_sv2v_reg,mem_3103_sv2v_reg,
  mem_3102_sv2v_reg,mem_3101_sv2v_reg,mem_3100_sv2v_reg,mem_3099_sv2v_reg,mem_3098_sv2v_reg,
  mem_3097_sv2v_reg,mem_3096_sv2v_reg,mem_3095_sv2v_reg,mem_3094_sv2v_reg,
  mem_3093_sv2v_reg,mem_3092_sv2v_reg,mem_3091_sv2v_reg,mem_3090_sv2v_reg,mem_3089_sv2v_reg,
  mem_3088_sv2v_reg,mem_3087_sv2v_reg,mem_3086_sv2v_reg,mem_3085_sv2v_reg,
  mem_3084_sv2v_reg,mem_3083_sv2v_reg,mem_3082_sv2v_reg,mem_3081_sv2v_reg,mem_3080_sv2v_reg,
  mem_3079_sv2v_reg,mem_3078_sv2v_reg,mem_3077_sv2v_reg,mem_3076_sv2v_reg,
  mem_3075_sv2v_reg,mem_3074_sv2v_reg,mem_3073_sv2v_reg,mem_3072_sv2v_reg,
  mem_3071_sv2v_reg,mem_3070_sv2v_reg,mem_3069_sv2v_reg,mem_3068_sv2v_reg,mem_3067_sv2v_reg,
  mem_3066_sv2v_reg,mem_3065_sv2v_reg,mem_3064_sv2v_reg,mem_3063_sv2v_reg,
  mem_3062_sv2v_reg,mem_3061_sv2v_reg,mem_3060_sv2v_reg,mem_3059_sv2v_reg,mem_3058_sv2v_reg,
  mem_3057_sv2v_reg,mem_3056_sv2v_reg,mem_3055_sv2v_reg,mem_3054_sv2v_reg,
  mem_3053_sv2v_reg,mem_3052_sv2v_reg,mem_3051_sv2v_reg,mem_3050_sv2v_reg,mem_3049_sv2v_reg,
  mem_3048_sv2v_reg,mem_3047_sv2v_reg,mem_3046_sv2v_reg,mem_3045_sv2v_reg,
  mem_3044_sv2v_reg,mem_3043_sv2v_reg,mem_3042_sv2v_reg,mem_3041_sv2v_reg,mem_3040_sv2v_reg,
  mem_3039_sv2v_reg,mem_3038_sv2v_reg,mem_3037_sv2v_reg,mem_3036_sv2v_reg,
  mem_3035_sv2v_reg,mem_3034_sv2v_reg,mem_3033_sv2v_reg,mem_3032_sv2v_reg,
  mem_3031_sv2v_reg,mem_3030_sv2v_reg,mem_3029_sv2v_reg,mem_3028_sv2v_reg,mem_3027_sv2v_reg,
  mem_3026_sv2v_reg,mem_3025_sv2v_reg,mem_3024_sv2v_reg,mem_3023_sv2v_reg,
  mem_3022_sv2v_reg,mem_3021_sv2v_reg,mem_3020_sv2v_reg,mem_3019_sv2v_reg,mem_3018_sv2v_reg,
  mem_3017_sv2v_reg,mem_3016_sv2v_reg,mem_3015_sv2v_reg,mem_3014_sv2v_reg,
  mem_3013_sv2v_reg,mem_3012_sv2v_reg,mem_3011_sv2v_reg,mem_3010_sv2v_reg,mem_3009_sv2v_reg,
  mem_3008_sv2v_reg,mem_3007_sv2v_reg,mem_3006_sv2v_reg,mem_3005_sv2v_reg,
  mem_3004_sv2v_reg,mem_3003_sv2v_reg,mem_3002_sv2v_reg,mem_3001_sv2v_reg,mem_3000_sv2v_reg,
  mem_2999_sv2v_reg,mem_2998_sv2v_reg,mem_2997_sv2v_reg,mem_2996_sv2v_reg,
  mem_2995_sv2v_reg,mem_2994_sv2v_reg,mem_2993_sv2v_reg,mem_2992_sv2v_reg,
  mem_2991_sv2v_reg,mem_2990_sv2v_reg,mem_2989_sv2v_reg,mem_2988_sv2v_reg,mem_2987_sv2v_reg,
  mem_2986_sv2v_reg,mem_2985_sv2v_reg,mem_2984_sv2v_reg,mem_2983_sv2v_reg,
  mem_2982_sv2v_reg,mem_2981_sv2v_reg,mem_2980_sv2v_reg,mem_2979_sv2v_reg,mem_2978_sv2v_reg,
  mem_2977_sv2v_reg,mem_2976_sv2v_reg,mem_2975_sv2v_reg,mem_2974_sv2v_reg,
  mem_2973_sv2v_reg,mem_2972_sv2v_reg,mem_2971_sv2v_reg,mem_2970_sv2v_reg,mem_2969_sv2v_reg,
  mem_2968_sv2v_reg,mem_2967_sv2v_reg,mem_2966_sv2v_reg,mem_2965_sv2v_reg,
  mem_2964_sv2v_reg,mem_2963_sv2v_reg,mem_2962_sv2v_reg,mem_2961_sv2v_reg,mem_2960_sv2v_reg,
  mem_2959_sv2v_reg,mem_2958_sv2v_reg,mem_2957_sv2v_reg,mem_2956_sv2v_reg,
  mem_2955_sv2v_reg,mem_2954_sv2v_reg,mem_2953_sv2v_reg,mem_2952_sv2v_reg,
  mem_2951_sv2v_reg,mem_2950_sv2v_reg,mem_2949_sv2v_reg,mem_2948_sv2v_reg,mem_2947_sv2v_reg,
  mem_2946_sv2v_reg,mem_2945_sv2v_reg,mem_2944_sv2v_reg,mem_2943_sv2v_reg,
  mem_2942_sv2v_reg,mem_2941_sv2v_reg,mem_2940_sv2v_reg,mem_2939_sv2v_reg,mem_2938_sv2v_reg,
  mem_2937_sv2v_reg,mem_2936_sv2v_reg,mem_2935_sv2v_reg,mem_2934_sv2v_reg,
  mem_2933_sv2v_reg,mem_2932_sv2v_reg,mem_2931_sv2v_reg,mem_2930_sv2v_reg,mem_2929_sv2v_reg,
  mem_2928_sv2v_reg,mem_2927_sv2v_reg,mem_2926_sv2v_reg,mem_2925_sv2v_reg,
  mem_2924_sv2v_reg,mem_2923_sv2v_reg,mem_2922_sv2v_reg,mem_2921_sv2v_reg,mem_2920_sv2v_reg,
  mem_2919_sv2v_reg,mem_2918_sv2v_reg,mem_2917_sv2v_reg,mem_2916_sv2v_reg,
  mem_2915_sv2v_reg,mem_2914_sv2v_reg,mem_2913_sv2v_reg,mem_2912_sv2v_reg,
  mem_2911_sv2v_reg,mem_2910_sv2v_reg,mem_2909_sv2v_reg,mem_2908_sv2v_reg,mem_2907_sv2v_reg,
  mem_2906_sv2v_reg,mem_2905_sv2v_reg,mem_2904_sv2v_reg,mem_2903_sv2v_reg,
  mem_2902_sv2v_reg,mem_2901_sv2v_reg,mem_2900_sv2v_reg,mem_2899_sv2v_reg,mem_2898_sv2v_reg,
  mem_2897_sv2v_reg,mem_2896_sv2v_reg,mem_2895_sv2v_reg,mem_2894_sv2v_reg,
  mem_2893_sv2v_reg,mem_2892_sv2v_reg,mem_2891_sv2v_reg,mem_2890_sv2v_reg,mem_2889_sv2v_reg,
  mem_2888_sv2v_reg,mem_2887_sv2v_reg,mem_2886_sv2v_reg,mem_2885_sv2v_reg,
  mem_2884_sv2v_reg,mem_2883_sv2v_reg,mem_2882_sv2v_reg,mem_2881_sv2v_reg,mem_2880_sv2v_reg,
  mem_2879_sv2v_reg,mem_2878_sv2v_reg,mem_2877_sv2v_reg,mem_2876_sv2v_reg,
  mem_2875_sv2v_reg,mem_2874_sv2v_reg,mem_2873_sv2v_reg,mem_2872_sv2v_reg,
  mem_2871_sv2v_reg,mem_2870_sv2v_reg,mem_2869_sv2v_reg,mem_2868_sv2v_reg,mem_2867_sv2v_reg,
  mem_2866_sv2v_reg,mem_2865_sv2v_reg,mem_2864_sv2v_reg,mem_2863_sv2v_reg,
  mem_2862_sv2v_reg,mem_2861_sv2v_reg,mem_2860_sv2v_reg,mem_2859_sv2v_reg,mem_2858_sv2v_reg,
  mem_2857_sv2v_reg,mem_2856_sv2v_reg,mem_2855_sv2v_reg,mem_2854_sv2v_reg,
  mem_2853_sv2v_reg,mem_2852_sv2v_reg,mem_2851_sv2v_reg,mem_2850_sv2v_reg,mem_2849_sv2v_reg,
  mem_2848_sv2v_reg,mem_2847_sv2v_reg,mem_2846_sv2v_reg,mem_2845_sv2v_reg,
  mem_2844_sv2v_reg,mem_2843_sv2v_reg,mem_2842_sv2v_reg,mem_2841_sv2v_reg,mem_2840_sv2v_reg,
  mem_2839_sv2v_reg,mem_2838_sv2v_reg,mem_2837_sv2v_reg,mem_2836_sv2v_reg,
  mem_2835_sv2v_reg,mem_2834_sv2v_reg,mem_2833_sv2v_reg,mem_2832_sv2v_reg,
  mem_2831_sv2v_reg,mem_2830_sv2v_reg,mem_2829_sv2v_reg,mem_2828_sv2v_reg,mem_2827_sv2v_reg,
  mem_2826_sv2v_reg,mem_2825_sv2v_reg,mem_2824_sv2v_reg,mem_2823_sv2v_reg,
  mem_2822_sv2v_reg,mem_2821_sv2v_reg,mem_2820_sv2v_reg,mem_2819_sv2v_reg,mem_2818_sv2v_reg,
  mem_2817_sv2v_reg,mem_2816_sv2v_reg,mem_2815_sv2v_reg,mem_2814_sv2v_reg,
  mem_2813_sv2v_reg,mem_2812_sv2v_reg,mem_2811_sv2v_reg,mem_2810_sv2v_reg,mem_2809_sv2v_reg,
  mem_2808_sv2v_reg,mem_2807_sv2v_reg,mem_2806_sv2v_reg,mem_2805_sv2v_reg,
  mem_2804_sv2v_reg,mem_2803_sv2v_reg,mem_2802_sv2v_reg,mem_2801_sv2v_reg,mem_2800_sv2v_reg,
  mem_2799_sv2v_reg,mem_2798_sv2v_reg,mem_2797_sv2v_reg,mem_2796_sv2v_reg,
  mem_2795_sv2v_reg,mem_2794_sv2v_reg,mem_2793_sv2v_reg,mem_2792_sv2v_reg,
  mem_2791_sv2v_reg,mem_2790_sv2v_reg,mem_2789_sv2v_reg,mem_2788_sv2v_reg,mem_2787_sv2v_reg,
  mem_2786_sv2v_reg,mem_2785_sv2v_reg,mem_2784_sv2v_reg,mem_2783_sv2v_reg,
  mem_2782_sv2v_reg,mem_2781_sv2v_reg,mem_2780_sv2v_reg,mem_2779_sv2v_reg,mem_2778_sv2v_reg,
  mem_2777_sv2v_reg,mem_2776_sv2v_reg,mem_2775_sv2v_reg,mem_2774_sv2v_reg,
  mem_2773_sv2v_reg,mem_2772_sv2v_reg,mem_2771_sv2v_reg,mem_2770_sv2v_reg,mem_2769_sv2v_reg,
  mem_2768_sv2v_reg,mem_2767_sv2v_reg,mem_2766_sv2v_reg,mem_2765_sv2v_reg,
  mem_2764_sv2v_reg,mem_2763_sv2v_reg,mem_2762_sv2v_reg,mem_2761_sv2v_reg,mem_2760_sv2v_reg,
  mem_2759_sv2v_reg,mem_2758_sv2v_reg,mem_2757_sv2v_reg,mem_2756_sv2v_reg,
  mem_2755_sv2v_reg,mem_2754_sv2v_reg,mem_2753_sv2v_reg,mem_2752_sv2v_reg,
  mem_2751_sv2v_reg,mem_2750_sv2v_reg,mem_2749_sv2v_reg,mem_2748_sv2v_reg,mem_2747_sv2v_reg,
  mem_2746_sv2v_reg,mem_2745_sv2v_reg,mem_2744_sv2v_reg,mem_2743_sv2v_reg,
  mem_2742_sv2v_reg,mem_2741_sv2v_reg,mem_2740_sv2v_reg,mem_2739_sv2v_reg,mem_2738_sv2v_reg,
  mem_2737_sv2v_reg,mem_2736_sv2v_reg,mem_2735_sv2v_reg,mem_2734_sv2v_reg,
  mem_2733_sv2v_reg,mem_2732_sv2v_reg,mem_2731_sv2v_reg,mem_2730_sv2v_reg,mem_2729_sv2v_reg,
  mem_2728_sv2v_reg,mem_2727_sv2v_reg,mem_2726_sv2v_reg,mem_2725_sv2v_reg,
  mem_2724_sv2v_reg,mem_2723_sv2v_reg,mem_2722_sv2v_reg,mem_2721_sv2v_reg,mem_2720_sv2v_reg,
  mem_2719_sv2v_reg,mem_2718_sv2v_reg,mem_2717_sv2v_reg,mem_2716_sv2v_reg,
  mem_2715_sv2v_reg,mem_2714_sv2v_reg,mem_2713_sv2v_reg,mem_2712_sv2v_reg,
  mem_2711_sv2v_reg,mem_2710_sv2v_reg,mem_2709_sv2v_reg,mem_2708_sv2v_reg,mem_2707_sv2v_reg,
  mem_2706_sv2v_reg,mem_2705_sv2v_reg,mem_2704_sv2v_reg,mem_2703_sv2v_reg,
  mem_2702_sv2v_reg,mem_2701_sv2v_reg,mem_2700_sv2v_reg,mem_2699_sv2v_reg,mem_2698_sv2v_reg,
  mem_2697_sv2v_reg,mem_2696_sv2v_reg,mem_2695_sv2v_reg,mem_2694_sv2v_reg,
  mem_2693_sv2v_reg,mem_2692_sv2v_reg,mem_2691_sv2v_reg,mem_2690_sv2v_reg,mem_2689_sv2v_reg,
  mem_2688_sv2v_reg,mem_2687_sv2v_reg,mem_2686_sv2v_reg,mem_2685_sv2v_reg,
  mem_2684_sv2v_reg,mem_2683_sv2v_reg,mem_2682_sv2v_reg,mem_2681_sv2v_reg,mem_2680_sv2v_reg,
  mem_2679_sv2v_reg,mem_2678_sv2v_reg,mem_2677_sv2v_reg,mem_2676_sv2v_reg,
  mem_2675_sv2v_reg,mem_2674_sv2v_reg,mem_2673_sv2v_reg,mem_2672_sv2v_reg,
  mem_2671_sv2v_reg,mem_2670_sv2v_reg,mem_2669_sv2v_reg,mem_2668_sv2v_reg,mem_2667_sv2v_reg,
  mem_2666_sv2v_reg,mem_2665_sv2v_reg,mem_2664_sv2v_reg,mem_2663_sv2v_reg,
  mem_2662_sv2v_reg,mem_2661_sv2v_reg,mem_2660_sv2v_reg,mem_2659_sv2v_reg,mem_2658_sv2v_reg,
  mem_2657_sv2v_reg,mem_2656_sv2v_reg,mem_2655_sv2v_reg,mem_2654_sv2v_reg,
  mem_2653_sv2v_reg,mem_2652_sv2v_reg,mem_2651_sv2v_reg,mem_2650_sv2v_reg,mem_2649_sv2v_reg,
  mem_2648_sv2v_reg,mem_2647_sv2v_reg,mem_2646_sv2v_reg,mem_2645_sv2v_reg,
  mem_2644_sv2v_reg,mem_2643_sv2v_reg,mem_2642_sv2v_reg,mem_2641_sv2v_reg,mem_2640_sv2v_reg,
  mem_2639_sv2v_reg,mem_2638_sv2v_reg,mem_2637_sv2v_reg,mem_2636_sv2v_reg,
  mem_2635_sv2v_reg,mem_2634_sv2v_reg,mem_2633_sv2v_reg,mem_2632_sv2v_reg,
  mem_2631_sv2v_reg,mem_2630_sv2v_reg,mem_2629_sv2v_reg,mem_2628_sv2v_reg,mem_2627_sv2v_reg,
  mem_2626_sv2v_reg,mem_2625_sv2v_reg,mem_2624_sv2v_reg,mem_2623_sv2v_reg,
  mem_2622_sv2v_reg,mem_2621_sv2v_reg,mem_2620_sv2v_reg,mem_2619_sv2v_reg,mem_2618_sv2v_reg,
  mem_2617_sv2v_reg,mem_2616_sv2v_reg,mem_2615_sv2v_reg,mem_2614_sv2v_reg,
  mem_2613_sv2v_reg,mem_2612_sv2v_reg,mem_2611_sv2v_reg,mem_2610_sv2v_reg,mem_2609_sv2v_reg,
  mem_2608_sv2v_reg,mem_2607_sv2v_reg,mem_2606_sv2v_reg,mem_2605_sv2v_reg,
  mem_2604_sv2v_reg,mem_2603_sv2v_reg,mem_2602_sv2v_reg,mem_2601_sv2v_reg,mem_2600_sv2v_reg,
  mem_2599_sv2v_reg,mem_2598_sv2v_reg,mem_2597_sv2v_reg,mem_2596_sv2v_reg,
  mem_2595_sv2v_reg,mem_2594_sv2v_reg,mem_2593_sv2v_reg,mem_2592_sv2v_reg,
  mem_2591_sv2v_reg,mem_2590_sv2v_reg,mem_2589_sv2v_reg,mem_2588_sv2v_reg,mem_2587_sv2v_reg,
  mem_2586_sv2v_reg,mem_2585_sv2v_reg,mem_2584_sv2v_reg,mem_2583_sv2v_reg,
  mem_2582_sv2v_reg,mem_2581_sv2v_reg,mem_2580_sv2v_reg,mem_2579_sv2v_reg,mem_2578_sv2v_reg,
  mem_2577_sv2v_reg,mem_2576_sv2v_reg,mem_2575_sv2v_reg,mem_2574_sv2v_reg,
  mem_2573_sv2v_reg,mem_2572_sv2v_reg,mem_2571_sv2v_reg,mem_2570_sv2v_reg,mem_2569_sv2v_reg,
  mem_2568_sv2v_reg,mem_2567_sv2v_reg,mem_2566_sv2v_reg,mem_2565_sv2v_reg,
  mem_2564_sv2v_reg,mem_2563_sv2v_reg,mem_2562_sv2v_reg,mem_2561_sv2v_reg,mem_2560_sv2v_reg,
  mem_2559_sv2v_reg,mem_2558_sv2v_reg,mem_2557_sv2v_reg,mem_2556_sv2v_reg,
  mem_2555_sv2v_reg,mem_2554_sv2v_reg,mem_2553_sv2v_reg,mem_2552_sv2v_reg,
  mem_2551_sv2v_reg,mem_2550_sv2v_reg,mem_2549_sv2v_reg,mem_2548_sv2v_reg,mem_2547_sv2v_reg,
  mem_2546_sv2v_reg,mem_2545_sv2v_reg,mem_2544_sv2v_reg,mem_2543_sv2v_reg,
  mem_2542_sv2v_reg,mem_2541_sv2v_reg,mem_2540_sv2v_reg,mem_2539_sv2v_reg,mem_2538_sv2v_reg,
  mem_2537_sv2v_reg,mem_2536_sv2v_reg,mem_2535_sv2v_reg,mem_2534_sv2v_reg,
  mem_2533_sv2v_reg,mem_2532_sv2v_reg,mem_2531_sv2v_reg,mem_2530_sv2v_reg,mem_2529_sv2v_reg,
  mem_2528_sv2v_reg,mem_2527_sv2v_reg,mem_2526_sv2v_reg,mem_2525_sv2v_reg,
  mem_2524_sv2v_reg,mem_2523_sv2v_reg,mem_2522_sv2v_reg,mem_2521_sv2v_reg,mem_2520_sv2v_reg,
  mem_2519_sv2v_reg,mem_2518_sv2v_reg,mem_2517_sv2v_reg,mem_2516_sv2v_reg,
  mem_2515_sv2v_reg,mem_2514_sv2v_reg,mem_2513_sv2v_reg,mem_2512_sv2v_reg,
  mem_2511_sv2v_reg,mem_2510_sv2v_reg,mem_2509_sv2v_reg,mem_2508_sv2v_reg,mem_2507_sv2v_reg,
  mem_2506_sv2v_reg,mem_2505_sv2v_reg,mem_2504_sv2v_reg,mem_2503_sv2v_reg,
  mem_2502_sv2v_reg,mem_2501_sv2v_reg,mem_2500_sv2v_reg,mem_2499_sv2v_reg,mem_2498_sv2v_reg,
  mem_2497_sv2v_reg,mem_2496_sv2v_reg,mem_2495_sv2v_reg,mem_2494_sv2v_reg,
  mem_2493_sv2v_reg,mem_2492_sv2v_reg,mem_2491_sv2v_reg,mem_2490_sv2v_reg,mem_2489_sv2v_reg,
  mem_2488_sv2v_reg,mem_2487_sv2v_reg,mem_2486_sv2v_reg,mem_2485_sv2v_reg,
  mem_2484_sv2v_reg,mem_2483_sv2v_reg,mem_2482_sv2v_reg,mem_2481_sv2v_reg,mem_2480_sv2v_reg,
  mem_2479_sv2v_reg,mem_2478_sv2v_reg,mem_2477_sv2v_reg,mem_2476_sv2v_reg,
  mem_2475_sv2v_reg,mem_2474_sv2v_reg,mem_2473_sv2v_reg,mem_2472_sv2v_reg,
  mem_2471_sv2v_reg,mem_2470_sv2v_reg,mem_2469_sv2v_reg,mem_2468_sv2v_reg,mem_2467_sv2v_reg,
  mem_2466_sv2v_reg,mem_2465_sv2v_reg,mem_2464_sv2v_reg,mem_2463_sv2v_reg,
  mem_2462_sv2v_reg,mem_2461_sv2v_reg,mem_2460_sv2v_reg,mem_2459_sv2v_reg,mem_2458_sv2v_reg,
  mem_2457_sv2v_reg,mem_2456_sv2v_reg,mem_2455_sv2v_reg,mem_2454_sv2v_reg,
  mem_2453_sv2v_reg,mem_2452_sv2v_reg,mem_2451_sv2v_reg,mem_2450_sv2v_reg,mem_2449_sv2v_reg,
  mem_2448_sv2v_reg,mem_2447_sv2v_reg,mem_2446_sv2v_reg,mem_2445_sv2v_reg,
  mem_2444_sv2v_reg,mem_2443_sv2v_reg,mem_2442_sv2v_reg,mem_2441_sv2v_reg,mem_2440_sv2v_reg,
  mem_2439_sv2v_reg,mem_2438_sv2v_reg,mem_2437_sv2v_reg,mem_2436_sv2v_reg,
  mem_2435_sv2v_reg,mem_2434_sv2v_reg,mem_2433_sv2v_reg,mem_2432_sv2v_reg,
  mem_2431_sv2v_reg,mem_2430_sv2v_reg,mem_2429_sv2v_reg,mem_2428_sv2v_reg,mem_2427_sv2v_reg,
  mem_2426_sv2v_reg,mem_2425_sv2v_reg,mem_2424_sv2v_reg,mem_2423_sv2v_reg,
  mem_2422_sv2v_reg,mem_2421_sv2v_reg,mem_2420_sv2v_reg,mem_2419_sv2v_reg,mem_2418_sv2v_reg,
  mem_2417_sv2v_reg,mem_2416_sv2v_reg,mem_2415_sv2v_reg,mem_2414_sv2v_reg,
  mem_2413_sv2v_reg,mem_2412_sv2v_reg,mem_2411_sv2v_reg,mem_2410_sv2v_reg,mem_2409_sv2v_reg,
  mem_2408_sv2v_reg,mem_2407_sv2v_reg,mem_2406_sv2v_reg,mem_2405_sv2v_reg,
  mem_2404_sv2v_reg,mem_2403_sv2v_reg,mem_2402_sv2v_reg,mem_2401_sv2v_reg,mem_2400_sv2v_reg,
  mem_2399_sv2v_reg,mem_2398_sv2v_reg,mem_2397_sv2v_reg,mem_2396_sv2v_reg,
  mem_2395_sv2v_reg,mem_2394_sv2v_reg,mem_2393_sv2v_reg,mem_2392_sv2v_reg,
  mem_2391_sv2v_reg,mem_2390_sv2v_reg,mem_2389_sv2v_reg,mem_2388_sv2v_reg,mem_2387_sv2v_reg,
  mem_2386_sv2v_reg,mem_2385_sv2v_reg,mem_2384_sv2v_reg,mem_2383_sv2v_reg,
  mem_2382_sv2v_reg,mem_2381_sv2v_reg,mem_2380_sv2v_reg,mem_2379_sv2v_reg,mem_2378_sv2v_reg,
  mem_2377_sv2v_reg,mem_2376_sv2v_reg,mem_2375_sv2v_reg,mem_2374_sv2v_reg,
  mem_2373_sv2v_reg,mem_2372_sv2v_reg,mem_2371_sv2v_reg,mem_2370_sv2v_reg,mem_2369_sv2v_reg,
  mem_2368_sv2v_reg,mem_2367_sv2v_reg,mem_2366_sv2v_reg,mem_2365_sv2v_reg,
  mem_2364_sv2v_reg,mem_2363_sv2v_reg,mem_2362_sv2v_reg,mem_2361_sv2v_reg,mem_2360_sv2v_reg,
  mem_2359_sv2v_reg,mem_2358_sv2v_reg,mem_2357_sv2v_reg,mem_2356_sv2v_reg,
  mem_2355_sv2v_reg,mem_2354_sv2v_reg,mem_2353_sv2v_reg,mem_2352_sv2v_reg,
  mem_2351_sv2v_reg,mem_2350_sv2v_reg,mem_2349_sv2v_reg,mem_2348_sv2v_reg,mem_2347_sv2v_reg,
  mem_2346_sv2v_reg,mem_2345_sv2v_reg,mem_2344_sv2v_reg,mem_2343_sv2v_reg,
  mem_2342_sv2v_reg,mem_2341_sv2v_reg,mem_2340_sv2v_reg,mem_2339_sv2v_reg,mem_2338_sv2v_reg,
  mem_2337_sv2v_reg,mem_2336_sv2v_reg,mem_2335_sv2v_reg,mem_2334_sv2v_reg,
  mem_2333_sv2v_reg,mem_2332_sv2v_reg,mem_2331_sv2v_reg,mem_2330_sv2v_reg,mem_2329_sv2v_reg,
  mem_2328_sv2v_reg,mem_2327_sv2v_reg,mem_2326_sv2v_reg,mem_2325_sv2v_reg,
  mem_2324_sv2v_reg,mem_2323_sv2v_reg,mem_2322_sv2v_reg,mem_2321_sv2v_reg,mem_2320_sv2v_reg,
  mem_2319_sv2v_reg,mem_2318_sv2v_reg,mem_2317_sv2v_reg,mem_2316_sv2v_reg,
  mem_2315_sv2v_reg,mem_2314_sv2v_reg,mem_2313_sv2v_reg,mem_2312_sv2v_reg,
  mem_2311_sv2v_reg,mem_2310_sv2v_reg,mem_2309_sv2v_reg,mem_2308_sv2v_reg,mem_2307_sv2v_reg,
  mem_2306_sv2v_reg,mem_2305_sv2v_reg,mem_2304_sv2v_reg,mem_2303_sv2v_reg,
  mem_2302_sv2v_reg,mem_2301_sv2v_reg,mem_2300_sv2v_reg,mem_2299_sv2v_reg,mem_2298_sv2v_reg,
  mem_2297_sv2v_reg,mem_2296_sv2v_reg,mem_2295_sv2v_reg,mem_2294_sv2v_reg,
  mem_2293_sv2v_reg,mem_2292_sv2v_reg,mem_2291_sv2v_reg,mem_2290_sv2v_reg,mem_2289_sv2v_reg,
  mem_2288_sv2v_reg,mem_2287_sv2v_reg,mem_2286_sv2v_reg,mem_2285_sv2v_reg,
  mem_2284_sv2v_reg,mem_2283_sv2v_reg,mem_2282_sv2v_reg,mem_2281_sv2v_reg,mem_2280_sv2v_reg,
  mem_2279_sv2v_reg,mem_2278_sv2v_reg,mem_2277_sv2v_reg,mem_2276_sv2v_reg,
  mem_2275_sv2v_reg,mem_2274_sv2v_reg,mem_2273_sv2v_reg,mem_2272_sv2v_reg,
  mem_2271_sv2v_reg,mem_2270_sv2v_reg,mem_2269_sv2v_reg,mem_2268_sv2v_reg,mem_2267_sv2v_reg,
  mem_2266_sv2v_reg,mem_2265_sv2v_reg,mem_2264_sv2v_reg,mem_2263_sv2v_reg,
  mem_2262_sv2v_reg,mem_2261_sv2v_reg,mem_2260_sv2v_reg,mem_2259_sv2v_reg,mem_2258_sv2v_reg,
  mem_2257_sv2v_reg,mem_2256_sv2v_reg,mem_2255_sv2v_reg,mem_2254_sv2v_reg,
  mem_2253_sv2v_reg,mem_2252_sv2v_reg,mem_2251_sv2v_reg,mem_2250_sv2v_reg,mem_2249_sv2v_reg,
  mem_2248_sv2v_reg,mem_2247_sv2v_reg,mem_2246_sv2v_reg,mem_2245_sv2v_reg,
  mem_2244_sv2v_reg,mem_2243_sv2v_reg,mem_2242_sv2v_reg,mem_2241_sv2v_reg,mem_2240_sv2v_reg,
  mem_2239_sv2v_reg,mem_2238_sv2v_reg,mem_2237_sv2v_reg,mem_2236_sv2v_reg,
  mem_2235_sv2v_reg,mem_2234_sv2v_reg,mem_2233_sv2v_reg,mem_2232_sv2v_reg,
  mem_2231_sv2v_reg,mem_2230_sv2v_reg,mem_2229_sv2v_reg,mem_2228_sv2v_reg,mem_2227_sv2v_reg,
  mem_2226_sv2v_reg,mem_2225_sv2v_reg,mem_2224_sv2v_reg,mem_2223_sv2v_reg,
  mem_2222_sv2v_reg,mem_2221_sv2v_reg,mem_2220_sv2v_reg,mem_2219_sv2v_reg,mem_2218_sv2v_reg,
  mem_2217_sv2v_reg,mem_2216_sv2v_reg,mem_2215_sv2v_reg,mem_2214_sv2v_reg,
  mem_2213_sv2v_reg,mem_2212_sv2v_reg,mem_2211_sv2v_reg,mem_2210_sv2v_reg,mem_2209_sv2v_reg,
  mem_2208_sv2v_reg,mem_2207_sv2v_reg,mem_2206_sv2v_reg,mem_2205_sv2v_reg,
  mem_2204_sv2v_reg,mem_2203_sv2v_reg,mem_2202_sv2v_reg,mem_2201_sv2v_reg,mem_2200_sv2v_reg,
  mem_2199_sv2v_reg,mem_2198_sv2v_reg,mem_2197_sv2v_reg,mem_2196_sv2v_reg,
  mem_2195_sv2v_reg,mem_2194_sv2v_reg,mem_2193_sv2v_reg,mem_2192_sv2v_reg,
  mem_2191_sv2v_reg,mem_2190_sv2v_reg,mem_2189_sv2v_reg,mem_2188_sv2v_reg,mem_2187_sv2v_reg,
  mem_2186_sv2v_reg,mem_2185_sv2v_reg,mem_2184_sv2v_reg,mem_2183_sv2v_reg,
  mem_2182_sv2v_reg,mem_2181_sv2v_reg,mem_2180_sv2v_reg,mem_2179_sv2v_reg,mem_2178_sv2v_reg,
  mem_2177_sv2v_reg,mem_2176_sv2v_reg,mem_2175_sv2v_reg,mem_2174_sv2v_reg,
  mem_2173_sv2v_reg,mem_2172_sv2v_reg,mem_2171_sv2v_reg,mem_2170_sv2v_reg,mem_2169_sv2v_reg,
  mem_2168_sv2v_reg,mem_2167_sv2v_reg,mem_2166_sv2v_reg,mem_2165_sv2v_reg,
  mem_2164_sv2v_reg,mem_2163_sv2v_reg,mem_2162_sv2v_reg,mem_2161_sv2v_reg,mem_2160_sv2v_reg,
  mem_2159_sv2v_reg,mem_2158_sv2v_reg,mem_2157_sv2v_reg,mem_2156_sv2v_reg,
  mem_2155_sv2v_reg,mem_2154_sv2v_reg,mem_2153_sv2v_reg,mem_2152_sv2v_reg,
  mem_2151_sv2v_reg,mem_2150_sv2v_reg,mem_2149_sv2v_reg,mem_2148_sv2v_reg,mem_2147_sv2v_reg,
  mem_2146_sv2v_reg,mem_2145_sv2v_reg,mem_2144_sv2v_reg,mem_2143_sv2v_reg,
  mem_2142_sv2v_reg,mem_2141_sv2v_reg,mem_2140_sv2v_reg,mem_2139_sv2v_reg,mem_2138_sv2v_reg,
  mem_2137_sv2v_reg,mem_2136_sv2v_reg,mem_2135_sv2v_reg,mem_2134_sv2v_reg,
  mem_2133_sv2v_reg,mem_2132_sv2v_reg,mem_2131_sv2v_reg,mem_2130_sv2v_reg,mem_2129_sv2v_reg,
  mem_2128_sv2v_reg,mem_2127_sv2v_reg,mem_2126_sv2v_reg,mem_2125_sv2v_reg,
  mem_2124_sv2v_reg,mem_2123_sv2v_reg,mem_2122_sv2v_reg,mem_2121_sv2v_reg,mem_2120_sv2v_reg,
  mem_2119_sv2v_reg,mem_2118_sv2v_reg,mem_2117_sv2v_reg,mem_2116_sv2v_reg,
  mem_2115_sv2v_reg,mem_2114_sv2v_reg,mem_2113_sv2v_reg,mem_2112_sv2v_reg,
  mem_2111_sv2v_reg,mem_2110_sv2v_reg,mem_2109_sv2v_reg,mem_2108_sv2v_reg,mem_2107_sv2v_reg,
  mem_2106_sv2v_reg,mem_2105_sv2v_reg,mem_2104_sv2v_reg,mem_2103_sv2v_reg,
  mem_2102_sv2v_reg,mem_2101_sv2v_reg,mem_2100_sv2v_reg,mem_2099_sv2v_reg,mem_2098_sv2v_reg,
  mem_2097_sv2v_reg,mem_2096_sv2v_reg,mem_2095_sv2v_reg,mem_2094_sv2v_reg,
  mem_2093_sv2v_reg,mem_2092_sv2v_reg,mem_2091_sv2v_reg,mem_2090_sv2v_reg,mem_2089_sv2v_reg,
  mem_2088_sv2v_reg,mem_2087_sv2v_reg,mem_2086_sv2v_reg,mem_2085_sv2v_reg,
  mem_2084_sv2v_reg,mem_2083_sv2v_reg,mem_2082_sv2v_reg,mem_2081_sv2v_reg,mem_2080_sv2v_reg,
  mem_2079_sv2v_reg,mem_2078_sv2v_reg,mem_2077_sv2v_reg,mem_2076_sv2v_reg,
  mem_2075_sv2v_reg,mem_2074_sv2v_reg,mem_2073_sv2v_reg,mem_2072_sv2v_reg,
  mem_2071_sv2v_reg,mem_2070_sv2v_reg,mem_2069_sv2v_reg,mem_2068_sv2v_reg,mem_2067_sv2v_reg,
  mem_2066_sv2v_reg,mem_2065_sv2v_reg,mem_2064_sv2v_reg,mem_2063_sv2v_reg,
  mem_2062_sv2v_reg,mem_2061_sv2v_reg,mem_2060_sv2v_reg,mem_2059_sv2v_reg,mem_2058_sv2v_reg,
  mem_2057_sv2v_reg,mem_2056_sv2v_reg,mem_2055_sv2v_reg,mem_2054_sv2v_reg,
  mem_2053_sv2v_reg,mem_2052_sv2v_reg,mem_2051_sv2v_reg,mem_2050_sv2v_reg,mem_2049_sv2v_reg,
  mem_2048_sv2v_reg,mem_2047_sv2v_reg,mem_2046_sv2v_reg,mem_2045_sv2v_reg,
  mem_2044_sv2v_reg,mem_2043_sv2v_reg,mem_2042_sv2v_reg,mem_2041_sv2v_reg,mem_2040_sv2v_reg,
  mem_2039_sv2v_reg,mem_2038_sv2v_reg,mem_2037_sv2v_reg,mem_2036_sv2v_reg,
  mem_2035_sv2v_reg,mem_2034_sv2v_reg,mem_2033_sv2v_reg,mem_2032_sv2v_reg,
  mem_2031_sv2v_reg,mem_2030_sv2v_reg,mem_2029_sv2v_reg,mem_2028_sv2v_reg,mem_2027_sv2v_reg,
  mem_2026_sv2v_reg,mem_2025_sv2v_reg,mem_2024_sv2v_reg,mem_2023_sv2v_reg,
  mem_2022_sv2v_reg,mem_2021_sv2v_reg,mem_2020_sv2v_reg,mem_2019_sv2v_reg,mem_2018_sv2v_reg,
  mem_2017_sv2v_reg,mem_2016_sv2v_reg,mem_2015_sv2v_reg,mem_2014_sv2v_reg,
  mem_2013_sv2v_reg,mem_2012_sv2v_reg,mem_2011_sv2v_reg,mem_2010_sv2v_reg,mem_2009_sv2v_reg,
  mem_2008_sv2v_reg,mem_2007_sv2v_reg,mem_2006_sv2v_reg,mem_2005_sv2v_reg,
  mem_2004_sv2v_reg,mem_2003_sv2v_reg,mem_2002_sv2v_reg,mem_2001_sv2v_reg,mem_2000_sv2v_reg,
  mem_1999_sv2v_reg,mem_1998_sv2v_reg,mem_1997_sv2v_reg,mem_1996_sv2v_reg,
  mem_1995_sv2v_reg,mem_1994_sv2v_reg,mem_1993_sv2v_reg,mem_1992_sv2v_reg,
  mem_1991_sv2v_reg,mem_1990_sv2v_reg,mem_1989_sv2v_reg,mem_1988_sv2v_reg,mem_1987_sv2v_reg,
  mem_1986_sv2v_reg,mem_1985_sv2v_reg,mem_1984_sv2v_reg,mem_1983_sv2v_reg,
  mem_1982_sv2v_reg,mem_1981_sv2v_reg,mem_1980_sv2v_reg,mem_1979_sv2v_reg,mem_1978_sv2v_reg,
  mem_1977_sv2v_reg,mem_1976_sv2v_reg,mem_1975_sv2v_reg,mem_1974_sv2v_reg,
  mem_1973_sv2v_reg,mem_1972_sv2v_reg,mem_1971_sv2v_reg,mem_1970_sv2v_reg,mem_1969_sv2v_reg,
  mem_1968_sv2v_reg,mem_1967_sv2v_reg,mem_1966_sv2v_reg,mem_1965_sv2v_reg,
  mem_1964_sv2v_reg,mem_1963_sv2v_reg,mem_1962_sv2v_reg,mem_1961_sv2v_reg,mem_1960_sv2v_reg,
  mem_1959_sv2v_reg,mem_1958_sv2v_reg,mem_1957_sv2v_reg,mem_1956_sv2v_reg,
  mem_1955_sv2v_reg,mem_1954_sv2v_reg,mem_1953_sv2v_reg,mem_1952_sv2v_reg,
  mem_1951_sv2v_reg,mem_1950_sv2v_reg,mem_1949_sv2v_reg,mem_1948_sv2v_reg,mem_1947_sv2v_reg,
  mem_1946_sv2v_reg,mem_1945_sv2v_reg,mem_1944_sv2v_reg,mem_1943_sv2v_reg,
  mem_1942_sv2v_reg,mem_1941_sv2v_reg,mem_1940_sv2v_reg,mem_1939_sv2v_reg,mem_1938_sv2v_reg,
  mem_1937_sv2v_reg,mem_1936_sv2v_reg,mem_1935_sv2v_reg,mem_1934_sv2v_reg,
  mem_1933_sv2v_reg,mem_1932_sv2v_reg,mem_1931_sv2v_reg,mem_1930_sv2v_reg,mem_1929_sv2v_reg,
  mem_1928_sv2v_reg,mem_1927_sv2v_reg,mem_1926_sv2v_reg,mem_1925_sv2v_reg,
  mem_1924_sv2v_reg,mem_1923_sv2v_reg,mem_1922_sv2v_reg,mem_1921_sv2v_reg,mem_1920_sv2v_reg,
  mem_1919_sv2v_reg,mem_1918_sv2v_reg,mem_1917_sv2v_reg,mem_1916_sv2v_reg,
  mem_1915_sv2v_reg,mem_1914_sv2v_reg,mem_1913_sv2v_reg,mem_1912_sv2v_reg,
  mem_1911_sv2v_reg,mem_1910_sv2v_reg,mem_1909_sv2v_reg,mem_1908_sv2v_reg,mem_1907_sv2v_reg,
  mem_1906_sv2v_reg,mem_1905_sv2v_reg,mem_1904_sv2v_reg,mem_1903_sv2v_reg,
  mem_1902_sv2v_reg,mem_1901_sv2v_reg,mem_1900_sv2v_reg,mem_1899_sv2v_reg,mem_1898_sv2v_reg,
  mem_1897_sv2v_reg,mem_1896_sv2v_reg,mem_1895_sv2v_reg,mem_1894_sv2v_reg,
  mem_1893_sv2v_reg,mem_1892_sv2v_reg,mem_1891_sv2v_reg,mem_1890_sv2v_reg,mem_1889_sv2v_reg,
  mem_1888_sv2v_reg,mem_1887_sv2v_reg,mem_1886_sv2v_reg,mem_1885_sv2v_reg,
  mem_1884_sv2v_reg,mem_1883_sv2v_reg,mem_1882_sv2v_reg,mem_1881_sv2v_reg,mem_1880_sv2v_reg,
  mem_1879_sv2v_reg,mem_1878_sv2v_reg,mem_1877_sv2v_reg,mem_1876_sv2v_reg,
  mem_1875_sv2v_reg,mem_1874_sv2v_reg,mem_1873_sv2v_reg,mem_1872_sv2v_reg,
  mem_1871_sv2v_reg,mem_1870_sv2v_reg,mem_1869_sv2v_reg,mem_1868_sv2v_reg,mem_1867_sv2v_reg,
  mem_1866_sv2v_reg,mem_1865_sv2v_reg,mem_1864_sv2v_reg,mem_1863_sv2v_reg,
  mem_1862_sv2v_reg,mem_1861_sv2v_reg,mem_1860_sv2v_reg,mem_1859_sv2v_reg,mem_1858_sv2v_reg,
  mem_1857_sv2v_reg,mem_1856_sv2v_reg,mem_1855_sv2v_reg,mem_1854_sv2v_reg,
  mem_1853_sv2v_reg,mem_1852_sv2v_reg,mem_1851_sv2v_reg,mem_1850_sv2v_reg,mem_1849_sv2v_reg,
  mem_1848_sv2v_reg,mem_1847_sv2v_reg,mem_1846_sv2v_reg,mem_1845_sv2v_reg,
  mem_1844_sv2v_reg,mem_1843_sv2v_reg,mem_1842_sv2v_reg,mem_1841_sv2v_reg,mem_1840_sv2v_reg,
  mem_1839_sv2v_reg,mem_1838_sv2v_reg,mem_1837_sv2v_reg,mem_1836_sv2v_reg,
  mem_1835_sv2v_reg,mem_1834_sv2v_reg,mem_1833_sv2v_reg,mem_1832_sv2v_reg,
  mem_1831_sv2v_reg,mem_1830_sv2v_reg,mem_1829_sv2v_reg,mem_1828_sv2v_reg,mem_1827_sv2v_reg,
  mem_1826_sv2v_reg,mem_1825_sv2v_reg,mem_1824_sv2v_reg,mem_1823_sv2v_reg,
  mem_1822_sv2v_reg,mem_1821_sv2v_reg,mem_1820_sv2v_reg,mem_1819_sv2v_reg,mem_1818_sv2v_reg,
  mem_1817_sv2v_reg,mem_1816_sv2v_reg,mem_1815_sv2v_reg,mem_1814_sv2v_reg,
  mem_1813_sv2v_reg,mem_1812_sv2v_reg,mem_1811_sv2v_reg,mem_1810_sv2v_reg,mem_1809_sv2v_reg,
  mem_1808_sv2v_reg,mem_1807_sv2v_reg,mem_1806_sv2v_reg,mem_1805_sv2v_reg,
  mem_1804_sv2v_reg,mem_1803_sv2v_reg,mem_1802_sv2v_reg,mem_1801_sv2v_reg,mem_1800_sv2v_reg,
  mem_1799_sv2v_reg,mem_1798_sv2v_reg,mem_1797_sv2v_reg,mem_1796_sv2v_reg,
  mem_1795_sv2v_reg,mem_1794_sv2v_reg,mem_1793_sv2v_reg,mem_1792_sv2v_reg,
  mem_1791_sv2v_reg,mem_1790_sv2v_reg,mem_1789_sv2v_reg,mem_1788_sv2v_reg,mem_1787_sv2v_reg,
  mem_1786_sv2v_reg,mem_1785_sv2v_reg,mem_1784_sv2v_reg,mem_1783_sv2v_reg,
  mem_1782_sv2v_reg,mem_1781_sv2v_reg,mem_1780_sv2v_reg,mem_1779_sv2v_reg,mem_1778_sv2v_reg,
  mem_1777_sv2v_reg,mem_1776_sv2v_reg,mem_1775_sv2v_reg,mem_1774_sv2v_reg,
  mem_1773_sv2v_reg,mem_1772_sv2v_reg,mem_1771_sv2v_reg,mem_1770_sv2v_reg,mem_1769_sv2v_reg,
  mem_1768_sv2v_reg,mem_1767_sv2v_reg,mem_1766_sv2v_reg,mem_1765_sv2v_reg,
  mem_1764_sv2v_reg,mem_1763_sv2v_reg,mem_1762_sv2v_reg,mem_1761_sv2v_reg,mem_1760_sv2v_reg,
  mem_1759_sv2v_reg,mem_1758_sv2v_reg,mem_1757_sv2v_reg,mem_1756_sv2v_reg,
  mem_1755_sv2v_reg,mem_1754_sv2v_reg,mem_1753_sv2v_reg,mem_1752_sv2v_reg,
  mem_1751_sv2v_reg,mem_1750_sv2v_reg,mem_1749_sv2v_reg,mem_1748_sv2v_reg,mem_1747_sv2v_reg,
  mem_1746_sv2v_reg,mem_1745_sv2v_reg,mem_1744_sv2v_reg,mem_1743_sv2v_reg,
  mem_1742_sv2v_reg,mem_1741_sv2v_reg,mem_1740_sv2v_reg,mem_1739_sv2v_reg,mem_1738_sv2v_reg,
  mem_1737_sv2v_reg,mem_1736_sv2v_reg,mem_1735_sv2v_reg,mem_1734_sv2v_reg,
  mem_1733_sv2v_reg,mem_1732_sv2v_reg,mem_1731_sv2v_reg,mem_1730_sv2v_reg,mem_1729_sv2v_reg,
  mem_1728_sv2v_reg,mem_1727_sv2v_reg,mem_1726_sv2v_reg,mem_1725_sv2v_reg,
  mem_1724_sv2v_reg,mem_1723_sv2v_reg,mem_1722_sv2v_reg,mem_1721_sv2v_reg,mem_1720_sv2v_reg,
  mem_1719_sv2v_reg,mem_1718_sv2v_reg,mem_1717_sv2v_reg,mem_1716_sv2v_reg,
  mem_1715_sv2v_reg,mem_1714_sv2v_reg,mem_1713_sv2v_reg,mem_1712_sv2v_reg,
  mem_1711_sv2v_reg,mem_1710_sv2v_reg,mem_1709_sv2v_reg,mem_1708_sv2v_reg,mem_1707_sv2v_reg,
  mem_1706_sv2v_reg,mem_1705_sv2v_reg,mem_1704_sv2v_reg,mem_1703_sv2v_reg,
  mem_1702_sv2v_reg,mem_1701_sv2v_reg,mem_1700_sv2v_reg,mem_1699_sv2v_reg,mem_1698_sv2v_reg,
  mem_1697_sv2v_reg,mem_1696_sv2v_reg,mem_1695_sv2v_reg,mem_1694_sv2v_reg,
  mem_1693_sv2v_reg,mem_1692_sv2v_reg,mem_1691_sv2v_reg,mem_1690_sv2v_reg,mem_1689_sv2v_reg,
  mem_1688_sv2v_reg,mem_1687_sv2v_reg,mem_1686_sv2v_reg,mem_1685_sv2v_reg,
  mem_1684_sv2v_reg,mem_1683_sv2v_reg,mem_1682_sv2v_reg,mem_1681_sv2v_reg,mem_1680_sv2v_reg,
  mem_1679_sv2v_reg,mem_1678_sv2v_reg,mem_1677_sv2v_reg,mem_1676_sv2v_reg,
  mem_1675_sv2v_reg,mem_1674_sv2v_reg,mem_1673_sv2v_reg,mem_1672_sv2v_reg,
  mem_1671_sv2v_reg,mem_1670_sv2v_reg,mem_1669_sv2v_reg,mem_1668_sv2v_reg,mem_1667_sv2v_reg,
  mem_1666_sv2v_reg,mem_1665_sv2v_reg,mem_1664_sv2v_reg,mem_1663_sv2v_reg,
  mem_1662_sv2v_reg,mem_1661_sv2v_reg,mem_1660_sv2v_reg,mem_1659_sv2v_reg,mem_1658_sv2v_reg,
  mem_1657_sv2v_reg,mem_1656_sv2v_reg,mem_1655_sv2v_reg,mem_1654_sv2v_reg,
  mem_1653_sv2v_reg,mem_1652_sv2v_reg,mem_1651_sv2v_reg,mem_1650_sv2v_reg,mem_1649_sv2v_reg,
  mem_1648_sv2v_reg,mem_1647_sv2v_reg,mem_1646_sv2v_reg,mem_1645_sv2v_reg,
  mem_1644_sv2v_reg,mem_1643_sv2v_reg,mem_1642_sv2v_reg,mem_1641_sv2v_reg,mem_1640_sv2v_reg,
  mem_1639_sv2v_reg,mem_1638_sv2v_reg,mem_1637_sv2v_reg,mem_1636_sv2v_reg,
  mem_1635_sv2v_reg,mem_1634_sv2v_reg,mem_1633_sv2v_reg,mem_1632_sv2v_reg,
  mem_1631_sv2v_reg,mem_1630_sv2v_reg,mem_1629_sv2v_reg,mem_1628_sv2v_reg,mem_1627_sv2v_reg,
  mem_1626_sv2v_reg,mem_1625_sv2v_reg,mem_1624_sv2v_reg,mem_1623_sv2v_reg,
  mem_1622_sv2v_reg,mem_1621_sv2v_reg,mem_1620_sv2v_reg,mem_1619_sv2v_reg,mem_1618_sv2v_reg,
  mem_1617_sv2v_reg,mem_1616_sv2v_reg,mem_1615_sv2v_reg,mem_1614_sv2v_reg,
  mem_1613_sv2v_reg,mem_1612_sv2v_reg,mem_1611_sv2v_reg,mem_1610_sv2v_reg,mem_1609_sv2v_reg,
  mem_1608_sv2v_reg,mem_1607_sv2v_reg,mem_1606_sv2v_reg,mem_1605_sv2v_reg,
  mem_1604_sv2v_reg,mem_1603_sv2v_reg,mem_1602_sv2v_reg,mem_1601_sv2v_reg,mem_1600_sv2v_reg,
  mem_1599_sv2v_reg,mem_1598_sv2v_reg,mem_1597_sv2v_reg,mem_1596_sv2v_reg,
  mem_1595_sv2v_reg,mem_1594_sv2v_reg,mem_1593_sv2v_reg,mem_1592_sv2v_reg,
  mem_1591_sv2v_reg,mem_1590_sv2v_reg,mem_1589_sv2v_reg,mem_1588_sv2v_reg,mem_1587_sv2v_reg,
  mem_1586_sv2v_reg,mem_1585_sv2v_reg,mem_1584_sv2v_reg,mem_1583_sv2v_reg,
  mem_1582_sv2v_reg,mem_1581_sv2v_reg,mem_1580_sv2v_reg,mem_1579_sv2v_reg,mem_1578_sv2v_reg,
  mem_1577_sv2v_reg,mem_1576_sv2v_reg,mem_1575_sv2v_reg,mem_1574_sv2v_reg,
  mem_1573_sv2v_reg,mem_1572_sv2v_reg,mem_1571_sv2v_reg,mem_1570_sv2v_reg,mem_1569_sv2v_reg,
  mem_1568_sv2v_reg,mem_1567_sv2v_reg,mem_1566_sv2v_reg,mem_1565_sv2v_reg,
  mem_1564_sv2v_reg,mem_1563_sv2v_reg,mem_1562_sv2v_reg,mem_1561_sv2v_reg,mem_1560_sv2v_reg,
  mem_1559_sv2v_reg,mem_1558_sv2v_reg,mem_1557_sv2v_reg,mem_1556_sv2v_reg,
  mem_1555_sv2v_reg,mem_1554_sv2v_reg,mem_1553_sv2v_reg,mem_1552_sv2v_reg,
  mem_1551_sv2v_reg,mem_1550_sv2v_reg,mem_1549_sv2v_reg,mem_1548_sv2v_reg,mem_1547_sv2v_reg,
  mem_1546_sv2v_reg,mem_1545_sv2v_reg,mem_1544_sv2v_reg,mem_1543_sv2v_reg,
  mem_1542_sv2v_reg,mem_1541_sv2v_reg,mem_1540_sv2v_reg,mem_1539_sv2v_reg,mem_1538_sv2v_reg,
  mem_1537_sv2v_reg,mem_1536_sv2v_reg,mem_1535_sv2v_reg,mem_1534_sv2v_reg,
  mem_1533_sv2v_reg,mem_1532_sv2v_reg,mem_1531_sv2v_reg,mem_1530_sv2v_reg,mem_1529_sv2v_reg,
  mem_1528_sv2v_reg,mem_1527_sv2v_reg,mem_1526_sv2v_reg,mem_1525_sv2v_reg,
  mem_1524_sv2v_reg,mem_1523_sv2v_reg,mem_1522_sv2v_reg,mem_1521_sv2v_reg,mem_1520_sv2v_reg,
  mem_1519_sv2v_reg,mem_1518_sv2v_reg,mem_1517_sv2v_reg,mem_1516_sv2v_reg,
  mem_1515_sv2v_reg,mem_1514_sv2v_reg,mem_1513_sv2v_reg,mem_1512_sv2v_reg,
  mem_1511_sv2v_reg,mem_1510_sv2v_reg,mem_1509_sv2v_reg,mem_1508_sv2v_reg,mem_1507_sv2v_reg,
  mem_1506_sv2v_reg,mem_1505_sv2v_reg,mem_1504_sv2v_reg,mem_1503_sv2v_reg,
  mem_1502_sv2v_reg,mem_1501_sv2v_reg,mem_1500_sv2v_reg,mem_1499_sv2v_reg,mem_1498_sv2v_reg,
  mem_1497_sv2v_reg,mem_1496_sv2v_reg,mem_1495_sv2v_reg,mem_1494_sv2v_reg,
  mem_1493_sv2v_reg,mem_1492_sv2v_reg,mem_1491_sv2v_reg,mem_1490_sv2v_reg,mem_1489_sv2v_reg,
  mem_1488_sv2v_reg,mem_1487_sv2v_reg,mem_1486_sv2v_reg,mem_1485_sv2v_reg,
  mem_1484_sv2v_reg,mem_1483_sv2v_reg,mem_1482_sv2v_reg,mem_1481_sv2v_reg,mem_1480_sv2v_reg,
  mem_1479_sv2v_reg,mem_1478_sv2v_reg,mem_1477_sv2v_reg,mem_1476_sv2v_reg,
  mem_1475_sv2v_reg,mem_1474_sv2v_reg,mem_1473_sv2v_reg,mem_1472_sv2v_reg,
  mem_1471_sv2v_reg,mem_1470_sv2v_reg,mem_1469_sv2v_reg,mem_1468_sv2v_reg,mem_1467_sv2v_reg,
  mem_1466_sv2v_reg,mem_1465_sv2v_reg,mem_1464_sv2v_reg,mem_1463_sv2v_reg,
  mem_1462_sv2v_reg,mem_1461_sv2v_reg,mem_1460_sv2v_reg,mem_1459_sv2v_reg,mem_1458_sv2v_reg,
  mem_1457_sv2v_reg,mem_1456_sv2v_reg,mem_1455_sv2v_reg,mem_1454_sv2v_reg,
  mem_1453_sv2v_reg,mem_1452_sv2v_reg,mem_1451_sv2v_reg,mem_1450_sv2v_reg,mem_1449_sv2v_reg,
  mem_1448_sv2v_reg,mem_1447_sv2v_reg,mem_1446_sv2v_reg,mem_1445_sv2v_reg,
  mem_1444_sv2v_reg,mem_1443_sv2v_reg,mem_1442_sv2v_reg,mem_1441_sv2v_reg,mem_1440_sv2v_reg,
  mem_1439_sv2v_reg,mem_1438_sv2v_reg,mem_1437_sv2v_reg,mem_1436_sv2v_reg,
  mem_1435_sv2v_reg,mem_1434_sv2v_reg,mem_1433_sv2v_reg,mem_1432_sv2v_reg,
  mem_1431_sv2v_reg,mem_1430_sv2v_reg,mem_1429_sv2v_reg,mem_1428_sv2v_reg,mem_1427_sv2v_reg,
  mem_1426_sv2v_reg,mem_1425_sv2v_reg,mem_1424_sv2v_reg,mem_1423_sv2v_reg,
  mem_1422_sv2v_reg,mem_1421_sv2v_reg,mem_1420_sv2v_reg,mem_1419_sv2v_reg,mem_1418_sv2v_reg,
  mem_1417_sv2v_reg,mem_1416_sv2v_reg,mem_1415_sv2v_reg,mem_1414_sv2v_reg,
  mem_1413_sv2v_reg,mem_1412_sv2v_reg,mem_1411_sv2v_reg,mem_1410_sv2v_reg,mem_1409_sv2v_reg,
  mem_1408_sv2v_reg,mem_1407_sv2v_reg,mem_1406_sv2v_reg,mem_1405_sv2v_reg,
  mem_1404_sv2v_reg,mem_1403_sv2v_reg,mem_1402_sv2v_reg,mem_1401_sv2v_reg,mem_1400_sv2v_reg,
  mem_1399_sv2v_reg,mem_1398_sv2v_reg,mem_1397_sv2v_reg,mem_1396_sv2v_reg,
  mem_1395_sv2v_reg,mem_1394_sv2v_reg,mem_1393_sv2v_reg,mem_1392_sv2v_reg,
  mem_1391_sv2v_reg,mem_1390_sv2v_reg,mem_1389_sv2v_reg,mem_1388_sv2v_reg,mem_1387_sv2v_reg,
  mem_1386_sv2v_reg,mem_1385_sv2v_reg,mem_1384_sv2v_reg,mem_1383_sv2v_reg,
  mem_1382_sv2v_reg,mem_1381_sv2v_reg,mem_1380_sv2v_reg,mem_1379_sv2v_reg,mem_1378_sv2v_reg,
  mem_1377_sv2v_reg,mem_1376_sv2v_reg,mem_1375_sv2v_reg,mem_1374_sv2v_reg,
  mem_1373_sv2v_reg,mem_1372_sv2v_reg,mem_1371_sv2v_reg,mem_1370_sv2v_reg,mem_1369_sv2v_reg,
  mem_1368_sv2v_reg,mem_1367_sv2v_reg,mem_1366_sv2v_reg,mem_1365_sv2v_reg,
  mem_1364_sv2v_reg,mem_1363_sv2v_reg,mem_1362_sv2v_reg,mem_1361_sv2v_reg,mem_1360_sv2v_reg,
  mem_1359_sv2v_reg,mem_1358_sv2v_reg,mem_1357_sv2v_reg,mem_1356_sv2v_reg,
  mem_1355_sv2v_reg,mem_1354_sv2v_reg,mem_1353_sv2v_reg,mem_1352_sv2v_reg,
  mem_1351_sv2v_reg,mem_1350_sv2v_reg,mem_1349_sv2v_reg,mem_1348_sv2v_reg,mem_1347_sv2v_reg,
  mem_1346_sv2v_reg,mem_1345_sv2v_reg,mem_1344_sv2v_reg,mem_1343_sv2v_reg,
  mem_1342_sv2v_reg,mem_1341_sv2v_reg,mem_1340_sv2v_reg,mem_1339_sv2v_reg,mem_1338_sv2v_reg,
  mem_1337_sv2v_reg,mem_1336_sv2v_reg,mem_1335_sv2v_reg,mem_1334_sv2v_reg,
  mem_1333_sv2v_reg,mem_1332_sv2v_reg,mem_1331_sv2v_reg,mem_1330_sv2v_reg,mem_1329_sv2v_reg,
  mem_1328_sv2v_reg,mem_1327_sv2v_reg,mem_1326_sv2v_reg,mem_1325_sv2v_reg,
  mem_1324_sv2v_reg,mem_1323_sv2v_reg,mem_1322_sv2v_reg,mem_1321_sv2v_reg,mem_1320_sv2v_reg,
  mem_1319_sv2v_reg,mem_1318_sv2v_reg,mem_1317_sv2v_reg,mem_1316_sv2v_reg,
  mem_1315_sv2v_reg,mem_1314_sv2v_reg,mem_1313_sv2v_reg,mem_1312_sv2v_reg,
  mem_1311_sv2v_reg,mem_1310_sv2v_reg,mem_1309_sv2v_reg,mem_1308_sv2v_reg,mem_1307_sv2v_reg,
  mem_1306_sv2v_reg,mem_1305_sv2v_reg,mem_1304_sv2v_reg,mem_1303_sv2v_reg,
  mem_1302_sv2v_reg,mem_1301_sv2v_reg,mem_1300_sv2v_reg,mem_1299_sv2v_reg,mem_1298_sv2v_reg,
  mem_1297_sv2v_reg,mem_1296_sv2v_reg,mem_1295_sv2v_reg,mem_1294_sv2v_reg,
  mem_1293_sv2v_reg,mem_1292_sv2v_reg,mem_1291_sv2v_reg,mem_1290_sv2v_reg,mem_1289_sv2v_reg,
  mem_1288_sv2v_reg,mem_1287_sv2v_reg,mem_1286_sv2v_reg,mem_1285_sv2v_reg,
  mem_1284_sv2v_reg,mem_1283_sv2v_reg,mem_1282_sv2v_reg,mem_1281_sv2v_reg,mem_1280_sv2v_reg,
  mem_1279_sv2v_reg,mem_1278_sv2v_reg,mem_1277_sv2v_reg,mem_1276_sv2v_reg,
  mem_1275_sv2v_reg,mem_1274_sv2v_reg,mem_1273_sv2v_reg,mem_1272_sv2v_reg,
  mem_1271_sv2v_reg,mem_1270_sv2v_reg,mem_1269_sv2v_reg,mem_1268_sv2v_reg,mem_1267_sv2v_reg,
  mem_1266_sv2v_reg,mem_1265_sv2v_reg,mem_1264_sv2v_reg,mem_1263_sv2v_reg,
  mem_1262_sv2v_reg,mem_1261_sv2v_reg,mem_1260_sv2v_reg,mem_1259_sv2v_reg,mem_1258_sv2v_reg,
  mem_1257_sv2v_reg,mem_1256_sv2v_reg,mem_1255_sv2v_reg,mem_1254_sv2v_reg,
  mem_1253_sv2v_reg,mem_1252_sv2v_reg,mem_1251_sv2v_reg,mem_1250_sv2v_reg,mem_1249_sv2v_reg,
  mem_1248_sv2v_reg,mem_1247_sv2v_reg,mem_1246_sv2v_reg,mem_1245_sv2v_reg,
  mem_1244_sv2v_reg,mem_1243_sv2v_reg,mem_1242_sv2v_reg,mem_1241_sv2v_reg,mem_1240_sv2v_reg,
  mem_1239_sv2v_reg,mem_1238_sv2v_reg,mem_1237_sv2v_reg,mem_1236_sv2v_reg,
  mem_1235_sv2v_reg,mem_1234_sv2v_reg,mem_1233_sv2v_reg,mem_1232_sv2v_reg,
  mem_1231_sv2v_reg,mem_1230_sv2v_reg,mem_1229_sv2v_reg,mem_1228_sv2v_reg,mem_1227_sv2v_reg,
  mem_1226_sv2v_reg,mem_1225_sv2v_reg,mem_1224_sv2v_reg,mem_1223_sv2v_reg,
  mem_1222_sv2v_reg,mem_1221_sv2v_reg,mem_1220_sv2v_reg,mem_1219_sv2v_reg,mem_1218_sv2v_reg,
  mem_1217_sv2v_reg,mem_1216_sv2v_reg,mem_1215_sv2v_reg,mem_1214_sv2v_reg,
  mem_1213_sv2v_reg,mem_1212_sv2v_reg,mem_1211_sv2v_reg,mem_1210_sv2v_reg,mem_1209_sv2v_reg,
  mem_1208_sv2v_reg,mem_1207_sv2v_reg,mem_1206_sv2v_reg,mem_1205_sv2v_reg,
  mem_1204_sv2v_reg,mem_1203_sv2v_reg,mem_1202_sv2v_reg,mem_1201_sv2v_reg,mem_1200_sv2v_reg,
  mem_1199_sv2v_reg,mem_1198_sv2v_reg,mem_1197_sv2v_reg,mem_1196_sv2v_reg,
  mem_1195_sv2v_reg,mem_1194_sv2v_reg,mem_1193_sv2v_reg,mem_1192_sv2v_reg,
  mem_1191_sv2v_reg,mem_1190_sv2v_reg,mem_1189_sv2v_reg,mem_1188_sv2v_reg,mem_1187_sv2v_reg,
  mem_1186_sv2v_reg,mem_1185_sv2v_reg,mem_1184_sv2v_reg,mem_1183_sv2v_reg,
  mem_1182_sv2v_reg,mem_1181_sv2v_reg,mem_1180_sv2v_reg,mem_1179_sv2v_reg,mem_1178_sv2v_reg,
  mem_1177_sv2v_reg,mem_1176_sv2v_reg,mem_1175_sv2v_reg,mem_1174_sv2v_reg,
  mem_1173_sv2v_reg,mem_1172_sv2v_reg,mem_1171_sv2v_reg,mem_1170_sv2v_reg,mem_1169_sv2v_reg,
  mem_1168_sv2v_reg,mem_1167_sv2v_reg,mem_1166_sv2v_reg,mem_1165_sv2v_reg,
  mem_1164_sv2v_reg,mem_1163_sv2v_reg,mem_1162_sv2v_reg,mem_1161_sv2v_reg,mem_1160_sv2v_reg,
  mem_1159_sv2v_reg,mem_1158_sv2v_reg,mem_1157_sv2v_reg,mem_1156_sv2v_reg,
  mem_1155_sv2v_reg,mem_1154_sv2v_reg,mem_1153_sv2v_reg,mem_1152_sv2v_reg,
  mem_1151_sv2v_reg,mem_1150_sv2v_reg,mem_1149_sv2v_reg,mem_1148_sv2v_reg,mem_1147_sv2v_reg,
  mem_1146_sv2v_reg,mem_1145_sv2v_reg,mem_1144_sv2v_reg,mem_1143_sv2v_reg,
  mem_1142_sv2v_reg,mem_1141_sv2v_reg,mem_1140_sv2v_reg,mem_1139_sv2v_reg,mem_1138_sv2v_reg,
  mem_1137_sv2v_reg,mem_1136_sv2v_reg,mem_1135_sv2v_reg,mem_1134_sv2v_reg,
  mem_1133_sv2v_reg,mem_1132_sv2v_reg,mem_1131_sv2v_reg,mem_1130_sv2v_reg,mem_1129_sv2v_reg,
  mem_1128_sv2v_reg,mem_1127_sv2v_reg,mem_1126_sv2v_reg,mem_1125_sv2v_reg,
  mem_1124_sv2v_reg,mem_1123_sv2v_reg,mem_1122_sv2v_reg,mem_1121_sv2v_reg,mem_1120_sv2v_reg,
  mem_1119_sv2v_reg,mem_1118_sv2v_reg,mem_1117_sv2v_reg,mem_1116_sv2v_reg,
  mem_1115_sv2v_reg,mem_1114_sv2v_reg,mem_1113_sv2v_reg,mem_1112_sv2v_reg,
  mem_1111_sv2v_reg,mem_1110_sv2v_reg,mem_1109_sv2v_reg,mem_1108_sv2v_reg,mem_1107_sv2v_reg,
  mem_1106_sv2v_reg,mem_1105_sv2v_reg,mem_1104_sv2v_reg,mem_1103_sv2v_reg,
  mem_1102_sv2v_reg,mem_1101_sv2v_reg,mem_1100_sv2v_reg,mem_1099_sv2v_reg,mem_1098_sv2v_reg,
  mem_1097_sv2v_reg,mem_1096_sv2v_reg,mem_1095_sv2v_reg,mem_1094_sv2v_reg,
  mem_1093_sv2v_reg,mem_1092_sv2v_reg,mem_1091_sv2v_reg,mem_1090_sv2v_reg,mem_1089_sv2v_reg,
  mem_1088_sv2v_reg,mem_1087_sv2v_reg,mem_1086_sv2v_reg,mem_1085_sv2v_reg,
  mem_1084_sv2v_reg,mem_1083_sv2v_reg,mem_1082_sv2v_reg,mem_1081_sv2v_reg,mem_1080_sv2v_reg,
  mem_1079_sv2v_reg,mem_1078_sv2v_reg,mem_1077_sv2v_reg,mem_1076_sv2v_reg,
  mem_1075_sv2v_reg,mem_1074_sv2v_reg,mem_1073_sv2v_reg,mem_1072_sv2v_reg,
  mem_1071_sv2v_reg,mem_1070_sv2v_reg,mem_1069_sv2v_reg,mem_1068_sv2v_reg,mem_1067_sv2v_reg,
  mem_1066_sv2v_reg,mem_1065_sv2v_reg,mem_1064_sv2v_reg,mem_1063_sv2v_reg,
  mem_1062_sv2v_reg,mem_1061_sv2v_reg,mem_1060_sv2v_reg,mem_1059_sv2v_reg,mem_1058_sv2v_reg,
  mem_1057_sv2v_reg,mem_1056_sv2v_reg,mem_1055_sv2v_reg,mem_1054_sv2v_reg,
  mem_1053_sv2v_reg,mem_1052_sv2v_reg,mem_1051_sv2v_reg,mem_1050_sv2v_reg,mem_1049_sv2v_reg,
  mem_1048_sv2v_reg,mem_1047_sv2v_reg,mem_1046_sv2v_reg,mem_1045_sv2v_reg,
  mem_1044_sv2v_reg,mem_1043_sv2v_reg,mem_1042_sv2v_reg,mem_1041_sv2v_reg,mem_1040_sv2v_reg,
  mem_1039_sv2v_reg,mem_1038_sv2v_reg,mem_1037_sv2v_reg,mem_1036_sv2v_reg,
  mem_1035_sv2v_reg,mem_1034_sv2v_reg,mem_1033_sv2v_reg,mem_1032_sv2v_reg,
  mem_1031_sv2v_reg,mem_1030_sv2v_reg,mem_1029_sv2v_reg,mem_1028_sv2v_reg,mem_1027_sv2v_reg,
  mem_1026_sv2v_reg,mem_1025_sv2v_reg,mem_1024_sv2v_reg,mem_1023_sv2v_reg,
  mem_1022_sv2v_reg,mem_1021_sv2v_reg,mem_1020_sv2v_reg,mem_1019_sv2v_reg,mem_1018_sv2v_reg,
  mem_1017_sv2v_reg,mem_1016_sv2v_reg,mem_1015_sv2v_reg,mem_1014_sv2v_reg,
  mem_1013_sv2v_reg,mem_1012_sv2v_reg,mem_1011_sv2v_reg,mem_1010_sv2v_reg,mem_1009_sv2v_reg,
  mem_1008_sv2v_reg,mem_1007_sv2v_reg,mem_1006_sv2v_reg,mem_1005_sv2v_reg,
  mem_1004_sv2v_reg,mem_1003_sv2v_reg,mem_1002_sv2v_reg,mem_1001_sv2v_reg,mem_1000_sv2v_reg,
  mem_999_sv2v_reg,mem_998_sv2v_reg,mem_997_sv2v_reg,mem_996_sv2v_reg,
  mem_995_sv2v_reg,mem_994_sv2v_reg,mem_993_sv2v_reg,mem_992_sv2v_reg,mem_991_sv2v_reg,
  mem_990_sv2v_reg,mem_989_sv2v_reg,mem_988_sv2v_reg,mem_987_sv2v_reg,mem_986_sv2v_reg,
  mem_985_sv2v_reg,mem_984_sv2v_reg,mem_983_sv2v_reg,mem_982_sv2v_reg,
  mem_981_sv2v_reg,mem_980_sv2v_reg,mem_979_sv2v_reg,mem_978_sv2v_reg,mem_977_sv2v_reg,
  mem_976_sv2v_reg,mem_975_sv2v_reg,mem_974_sv2v_reg,mem_973_sv2v_reg,mem_972_sv2v_reg,
  mem_971_sv2v_reg,mem_970_sv2v_reg,mem_969_sv2v_reg,mem_968_sv2v_reg,
  mem_967_sv2v_reg,mem_966_sv2v_reg,mem_965_sv2v_reg,mem_964_sv2v_reg,mem_963_sv2v_reg,
  mem_962_sv2v_reg,mem_961_sv2v_reg,mem_960_sv2v_reg,mem_959_sv2v_reg,mem_958_sv2v_reg,
  mem_957_sv2v_reg,mem_956_sv2v_reg,mem_955_sv2v_reg,mem_954_sv2v_reg,mem_953_sv2v_reg,
  mem_952_sv2v_reg,mem_951_sv2v_reg,mem_950_sv2v_reg,mem_949_sv2v_reg,
  mem_948_sv2v_reg,mem_947_sv2v_reg,mem_946_sv2v_reg,mem_945_sv2v_reg,mem_944_sv2v_reg,
  mem_943_sv2v_reg,mem_942_sv2v_reg,mem_941_sv2v_reg,mem_940_sv2v_reg,mem_939_sv2v_reg,
  mem_938_sv2v_reg,mem_937_sv2v_reg,mem_936_sv2v_reg,mem_935_sv2v_reg,
  mem_934_sv2v_reg,mem_933_sv2v_reg,mem_932_sv2v_reg,mem_931_sv2v_reg,mem_930_sv2v_reg,
  mem_929_sv2v_reg,mem_928_sv2v_reg,mem_927_sv2v_reg,mem_926_sv2v_reg,mem_925_sv2v_reg,
  mem_924_sv2v_reg,mem_923_sv2v_reg,mem_922_sv2v_reg,mem_921_sv2v_reg,mem_920_sv2v_reg,
  mem_919_sv2v_reg,mem_918_sv2v_reg,mem_917_sv2v_reg,mem_916_sv2v_reg,
  mem_915_sv2v_reg,mem_914_sv2v_reg,mem_913_sv2v_reg,mem_912_sv2v_reg,mem_911_sv2v_reg,
  mem_910_sv2v_reg,mem_909_sv2v_reg,mem_908_sv2v_reg,mem_907_sv2v_reg,mem_906_sv2v_reg,
  mem_905_sv2v_reg,mem_904_sv2v_reg,mem_903_sv2v_reg,mem_902_sv2v_reg,
  mem_901_sv2v_reg,mem_900_sv2v_reg,mem_899_sv2v_reg,mem_898_sv2v_reg,mem_897_sv2v_reg,
  mem_896_sv2v_reg,mem_895_sv2v_reg,mem_894_sv2v_reg,mem_893_sv2v_reg,mem_892_sv2v_reg,
  mem_891_sv2v_reg,mem_890_sv2v_reg,mem_889_sv2v_reg,mem_888_sv2v_reg,
  mem_887_sv2v_reg,mem_886_sv2v_reg,mem_885_sv2v_reg,mem_884_sv2v_reg,mem_883_sv2v_reg,
  mem_882_sv2v_reg,mem_881_sv2v_reg,mem_880_sv2v_reg,mem_879_sv2v_reg,mem_878_sv2v_reg,
  mem_877_sv2v_reg,mem_876_sv2v_reg,mem_875_sv2v_reg,mem_874_sv2v_reg,mem_873_sv2v_reg,
  mem_872_sv2v_reg,mem_871_sv2v_reg,mem_870_sv2v_reg,mem_869_sv2v_reg,
  mem_868_sv2v_reg,mem_867_sv2v_reg,mem_866_sv2v_reg,mem_865_sv2v_reg,mem_864_sv2v_reg,
  mem_863_sv2v_reg,mem_862_sv2v_reg,mem_861_sv2v_reg,mem_860_sv2v_reg,mem_859_sv2v_reg,
  mem_858_sv2v_reg,mem_857_sv2v_reg,mem_856_sv2v_reg,mem_855_sv2v_reg,
  mem_854_sv2v_reg,mem_853_sv2v_reg,mem_852_sv2v_reg,mem_851_sv2v_reg,mem_850_sv2v_reg,
  mem_849_sv2v_reg,mem_848_sv2v_reg,mem_847_sv2v_reg,mem_846_sv2v_reg,mem_845_sv2v_reg,
  mem_844_sv2v_reg,mem_843_sv2v_reg,mem_842_sv2v_reg,mem_841_sv2v_reg,mem_840_sv2v_reg,
  mem_839_sv2v_reg,mem_838_sv2v_reg,mem_837_sv2v_reg,mem_836_sv2v_reg,
  mem_835_sv2v_reg,mem_834_sv2v_reg,mem_833_sv2v_reg,mem_832_sv2v_reg,mem_831_sv2v_reg,
  mem_830_sv2v_reg,mem_829_sv2v_reg,mem_828_sv2v_reg,mem_827_sv2v_reg,mem_826_sv2v_reg,
  mem_825_sv2v_reg,mem_824_sv2v_reg,mem_823_sv2v_reg,mem_822_sv2v_reg,
  mem_821_sv2v_reg,mem_820_sv2v_reg,mem_819_sv2v_reg,mem_818_sv2v_reg,mem_817_sv2v_reg,
  mem_816_sv2v_reg,mem_815_sv2v_reg,mem_814_sv2v_reg,mem_813_sv2v_reg,mem_812_sv2v_reg,
  mem_811_sv2v_reg,mem_810_sv2v_reg,mem_809_sv2v_reg,mem_808_sv2v_reg,
  mem_807_sv2v_reg,mem_806_sv2v_reg,mem_805_sv2v_reg,mem_804_sv2v_reg,mem_803_sv2v_reg,
  mem_802_sv2v_reg,mem_801_sv2v_reg,mem_800_sv2v_reg,mem_799_sv2v_reg,mem_798_sv2v_reg,
  mem_797_sv2v_reg,mem_796_sv2v_reg,mem_795_sv2v_reg,mem_794_sv2v_reg,mem_793_sv2v_reg,
  mem_792_sv2v_reg,mem_791_sv2v_reg,mem_790_sv2v_reg,mem_789_sv2v_reg,
  mem_788_sv2v_reg,mem_787_sv2v_reg,mem_786_sv2v_reg,mem_785_sv2v_reg,mem_784_sv2v_reg,
  mem_783_sv2v_reg,mem_782_sv2v_reg,mem_781_sv2v_reg,mem_780_sv2v_reg,mem_779_sv2v_reg,
  mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,mem_775_sv2v_reg,
  mem_774_sv2v_reg,mem_773_sv2v_reg,mem_772_sv2v_reg,mem_771_sv2v_reg,mem_770_sv2v_reg,
  mem_769_sv2v_reg,mem_768_sv2v_reg,mem_767_sv2v_reg,mem_766_sv2v_reg,mem_765_sv2v_reg,
  mem_764_sv2v_reg,mem_763_sv2v_reg,mem_762_sv2v_reg,mem_761_sv2v_reg,mem_760_sv2v_reg,
  mem_759_sv2v_reg,mem_758_sv2v_reg,mem_757_sv2v_reg,mem_756_sv2v_reg,
  mem_755_sv2v_reg,mem_754_sv2v_reg,mem_753_sv2v_reg,mem_752_sv2v_reg,mem_751_sv2v_reg,
  mem_750_sv2v_reg,mem_749_sv2v_reg,mem_748_sv2v_reg,mem_747_sv2v_reg,mem_746_sv2v_reg,
  mem_745_sv2v_reg,mem_744_sv2v_reg,mem_743_sv2v_reg,mem_742_sv2v_reg,
  mem_741_sv2v_reg,mem_740_sv2v_reg,mem_739_sv2v_reg,mem_738_sv2v_reg,mem_737_sv2v_reg,
  mem_736_sv2v_reg,mem_735_sv2v_reg,mem_734_sv2v_reg,mem_733_sv2v_reg,mem_732_sv2v_reg,
  mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,mem_728_sv2v_reg,
  mem_727_sv2v_reg,mem_726_sv2v_reg,mem_725_sv2v_reg,mem_724_sv2v_reg,mem_723_sv2v_reg,
  mem_722_sv2v_reg,mem_721_sv2v_reg,mem_720_sv2v_reg,mem_719_sv2v_reg,mem_718_sv2v_reg,
  mem_717_sv2v_reg,mem_716_sv2v_reg,mem_715_sv2v_reg,mem_714_sv2v_reg,mem_713_sv2v_reg,
  mem_712_sv2v_reg,mem_711_sv2v_reg,mem_710_sv2v_reg,mem_709_sv2v_reg,
  mem_708_sv2v_reg,mem_707_sv2v_reg,mem_706_sv2v_reg,mem_705_sv2v_reg,mem_704_sv2v_reg,
  mem_703_sv2v_reg,mem_702_sv2v_reg,mem_701_sv2v_reg,mem_700_sv2v_reg,mem_699_sv2v_reg,
  mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,mem_695_sv2v_reg,
  mem_694_sv2v_reg,mem_693_sv2v_reg,mem_692_sv2v_reg,mem_691_sv2v_reg,mem_690_sv2v_reg,
  mem_689_sv2v_reg,mem_688_sv2v_reg,mem_687_sv2v_reg,mem_686_sv2v_reg,mem_685_sv2v_reg,
  mem_684_sv2v_reg,mem_683_sv2v_reg,mem_682_sv2v_reg,mem_681_sv2v_reg,mem_680_sv2v_reg,
  mem_679_sv2v_reg,mem_678_sv2v_reg,mem_677_sv2v_reg,mem_676_sv2v_reg,
  mem_675_sv2v_reg,mem_674_sv2v_reg,mem_673_sv2v_reg,mem_672_sv2v_reg,mem_671_sv2v_reg,
  mem_670_sv2v_reg,mem_669_sv2v_reg,mem_668_sv2v_reg,mem_667_sv2v_reg,mem_666_sv2v_reg,
  mem_665_sv2v_reg,mem_664_sv2v_reg,mem_663_sv2v_reg,mem_662_sv2v_reg,
  mem_661_sv2v_reg,mem_660_sv2v_reg,mem_659_sv2v_reg,mem_658_sv2v_reg,mem_657_sv2v_reg,
  mem_656_sv2v_reg,mem_655_sv2v_reg,mem_654_sv2v_reg,mem_653_sv2v_reg,mem_652_sv2v_reg,
  mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,mem_648_sv2v_reg,
  mem_647_sv2v_reg,mem_646_sv2v_reg,mem_645_sv2v_reg,mem_644_sv2v_reg,mem_643_sv2v_reg,
  mem_642_sv2v_reg,mem_641_sv2v_reg,mem_640_sv2v_reg,mem_639_sv2v_reg,mem_638_sv2v_reg,
  mem_637_sv2v_reg,mem_636_sv2v_reg,mem_635_sv2v_reg,mem_634_sv2v_reg,mem_633_sv2v_reg,
  mem_632_sv2v_reg,mem_631_sv2v_reg,mem_630_sv2v_reg,mem_629_sv2v_reg,
  mem_628_sv2v_reg,mem_627_sv2v_reg,mem_626_sv2v_reg,mem_625_sv2v_reg,mem_624_sv2v_reg,
  mem_623_sv2v_reg,mem_622_sv2v_reg,mem_621_sv2v_reg,mem_620_sv2v_reg,mem_619_sv2v_reg,
  mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,mem_615_sv2v_reg,
  mem_614_sv2v_reg,mem_613_sv2v_reg,mem_612_sv2v_reg,mem_611_sv2v_reg,mem_610_sv2v_reg,
  mem_609_sv2v_reg,mem_608_sv2v_reg,mem_607_sv2v_reg,mem_606_sv2v_reg,mem_605_sv2v_reg,
  mem_604_sv2v_reg,mem_603_sv2v_reg,mem_602_sv2v_reg,mem_601_sv2v_reg,mem_600_sv2v_reg,
  mem_599_sv2v_reg,mem_598_sv2v_reg,mem_597_sv2v_reg,mem_596_sv2v_reg,
  mem_595_sv2v_reg,mem_594_sv2v_reg,mem_593_sv2v_reg,mem_592_sv2v_reg,mem_591_sv2v_reg,
  mem_590_sv2v_reg,mem_589_sv2v_reg,mem_588_sv2v_reg,mem_587_sv2v_reg,mem_586_sv2v_reg,
  mem_585_sv2v_reg,mem_584_sv2v_reg,mem_583_sv2v_reg,mem_582_sv2v_reg,
  mem_581_sv2v_reg,mem_580_sv2v_reg,mem_579_sv2v_reg,mem_578_sv2v_reg,mem_577_sv2v_reg,
  mem_576_sv2v_reg,mem_575_sv2v_reg,mem_574_sv2v_reg,mem_573_sv2v_reg,mem_572_sv2v_reg,
  mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,mem_568_sv2v_reg,
  mem_567_sv2v_reg,mem_566_sv2v_reg,mem_565_sv2v_reg,mem_564_sv2v_reg,mem_563_sv2v_reg,
  mem_562_sv2v_reg,mem_561_sv2v_reg,mem_560_sv2v_reg,mem_559_sv2v_reg,mem_558_sv2v_reg,
  mem_557_sv2v_reg,mem_556_sv2v_reg,mem_555_sv2v_reg,mem_554_sv2v_reg,mem_553_sv2v_reg,
  mem_552_sv2v_reg,mem_551_sv2v_reg,mem_550_sv2v_reg,mem_549_sv2v_reg,
  mem_548_sv2v_reg,mem_547_sv2v_reg,mem_546_sv2v_reg,mem_545_sv2v_reg,mem_544_sv2v_reg,
  mem_543_sv2v_reg,mem_542_sv2v_reg,mem_541_sv2v_reg,mem_540_sv2v_reg,mem_539_sv2v_reg,
  mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,mem_535_sv2v_reg,
  mem_534_sv2v_reg,mem_533_sv2v_reg,mem_532_sv2v_reg,mem_531_sv2v_reg,mem_530_sv2v_reg,
  mem_529_sv2v_reg,mem_528_sv2v_reg,mem_527_sv2v_reg,mem_526_sv2v_reg,mem_525_sv2v_reg,
  mem_524_sv2v_reg,mem_523_sv2v_reg,mem_522_sv2v_reg,mem_521_sv2v_reg,mem_520_sv2v_reg,
  mem_519_sv2v_reg,mem_518_sv2v_reg,mem_517_sv2v_reg,mem_516_sv2v_reg,
  mem_515_sv2v_reg,mem_514_sv2v_reg,mem_513_sv2v_reg,mem_512_sv2v_reg,mem_511_sv2v_reg,
  mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,mem_507_sv2v_reg,mem_506_sv2v_reg,
  mem_505_sv2v_reg,mem_504_sv2v_reg,mem_503_sv2v_reg,mem_502_sv2v_reg,
  mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,mem_497_sv2v_reg,
  mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,mem_493_sv2v_reg,mem_492_sv2v_reg,
  mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,mem_488_sv2v_reg,
  mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,mem_483_sv2v_reg,
  mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,mem_479_sv2v_reg,mem_478_sv2v_reg,
  mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,mem_474_sv2v_reg,mem_473_sv2v_reg,
  mem_472_sv2v_reg,mem_471_sv2v_reg,mem_470_sv2v_reg,mem_469_sv2v_reg,
  mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,mem_464_sv2v_reg,
  mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,mem_460_sv2v_reg,mem_459_sv2v_reg,
  mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,mem_455_sv2v_reg,
  mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,mem_450_sv2v_reg,
  mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,mem_446_sv2v_reg,mem_445_sv2v_reg,
  mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,mem_441_sv2v_reg,mem_440_sv2v_reg,
  mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,mem_436_sv2v_reg,
  mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,mem_431_sv2v_reg,
  mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,mem_427_sv2v_reg,mem_426_sv2v_reg,
  mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,mem_422_sv2v_reg,
  mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,mem_417_sv2v_reg,
  mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,mem_413_sv2v_reg,mem_412_sv2v_reg,
  mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,mem_408_sv2v_reg,
  mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,mem_403_sv2v_reg,
  mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,mem_399_sv2v_reg,mem_398_sv2v_reg,
  mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,mem_394_sv2v_reg,mem_393_sv2v_reg,
  mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,mem_389_sv2v_reg,
  mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,mem_384_sv2v_reg,
  mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,mem_380_sv2v_reg,mem_379_sv2v_reg,
  mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,mem_375_sv2v_reg,
  mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,mem_370_sv2v_reg,
  mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,mem_366_sv2v_reg,mem_365_sv2v_reg,
  mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,mem_361_sv2v_reg,mem_360_sv2v_reg,
  mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,mem_356_sv2v_reg,
  mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,mem_351_sv2v_reg,
  mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,mem_347_sv2v_reg,mem_346_sv2v_reg,
  mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,mem_342_sv2v_reg,
  mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,mem_337_sv2v_reg,
  mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,mem_333_sv2v_reg,mem_332_sv2v_reg,
  mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,mem_328_sv2v_reg,
  mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,mem_323_sv2v_reg,
  mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,mem_319_sv2v_reg,mem_318_sv2v_reg,
  mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,mem_314_sv2v_reg,mem_313_sv2v_reg,
  mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,mem_309_sv2v_reg,
  mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,mem_304_sv2v_reg,
  mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,mem_300_sv2v_reg,mem_299_sv2v_reg,
  mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,mem_295_sv2v_reg,
  mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,mem_290_sv2v_reg,
  mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,mem_286_sv2v_reg,mem_285_sv2v_reg,
  mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,mem_281_sv2v_reg,mem_280_sv2v_reg,
  mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,mem_276_sv2v_reg,
  mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,mem_271_sv2v_reg,
  mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,mem_267_sv2v_reg,mem_266_sv2v_reg,
  mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,mem_262_sv2v_reg,
  mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,mem_257_sv2v_reg,
  mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,
  mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,
  mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,
  mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,
  mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,mem_233_sv2v_reg,
  mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,mem_229_sv2v_reg,
  mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,
  mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,mem_219_sv2v_reg,
  mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,mem_215_sv2v_reg,
  mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,
  mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,
  mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,mem_200_sv2v_reg,
  mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,mem_196_sv2v_reg,
  mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,
  mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,mem_186_sv2v_reg,
  mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,mem_182_sv2v_reg,
  mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,
  mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,
  mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,
  mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,
  mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,
  mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,mem_153_sv2v_reg,
  mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,mem_149_sv2v_reg,
  mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,
  mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,mem_139_sv2v_reg,
  mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,mem_135_sv2v_reg,
  mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,
  mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,
  mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,mem_120_sv2v_reg,
  mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,mem_116_sv2v_reg,
  mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,
  mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,mem_106_sv2v_reg,
  mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,mem_102_sv2v_reg,
  mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,
  mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,
  mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,
  mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,
  mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,
  mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,
  mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,
  mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,
  mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,
  mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,
  mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,
  mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,
  mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,
  mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,
  mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,
  mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,
  mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,
  mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,
  mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,
  mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,
  mem_0_sv2v_reg;
  assign mem[3199] = mem_3199_sv2v_reg;
  assign mem[3198] = mem_3198_sv2v_reg;
  assign mem[3197] = mem_3197_sv2v_reg;
  assign mem[3196] = mem_3196_sv2v_reg;
  assign mem[3195] = mem_3195_sv2v_reg;
  assign mem[3194] = mem_3194_sv2v_reg;
  assign mem[3193] = mem_3193_sv2v_reg;
  assign mem[3192] = mem_3192_sv2v_reg;
  assign mem[3191] = mem_3191_sv2v_reg;
  assign mem[3190] = mem_3190_sv2v_reg;
  assign mem[3189] = mem_3189_sv2v_reg;
  assign mem[3188] = mem_3188_sv2v_reg;
  assign mem[3187] = mem_3187_sv2v_reg;
  assign mem[3186] = mem_3186_sv2v_reg;
  assign mem[3185] = mem_3185_sv2v_reg;
  assign mem[3184] = mem_3184_sv2v_reg;
  assign mem[3183] = mem_3183_sv2v_reg;
  assign mem[3182] = mem_3182_sv2v_reg;
  assign mem[3181] = mem_3181_sv2v_reg;
  assign mem[3180] = mem_3180_sv2v_reg;
  assign mem[3179] = mem_3179_sv2v_reg;
  assign mem[3178] = mem_3178_sv2v_reg;
  assign mem[3177] = mem_3177_sv2v_reg;
  assign mem[3176] = mem_3176_sv2v_reg;
  assign mem[3175] = mem_3175_sv2v_reg;
  assign mem[3174] = mem_3174_sv2v_reg;
  assign mem[3173] = mem_3173_sv2v_reg;
  assign mem[3172] = mem_3172_sv2v_reg;
  assign mem[3171] = mem_3171_sv2v_reg;
  assign mem[3170] = mem_3170_sv2v_reg;
  assign mem[3169] = mem_3169_sv2v_reg;
  assign mem[3168] = mem_3168_sv2v_reg;
  assign mem[3167] = mem_3167_sv2v_reg;
  assign mem[3166] = mem_3166_sv2v_reg;
  assign mem[3165] = mem_3165_sv2v_reg;
  assign mem[3164] = mem_3164_sv2v_reg;
  assign mem[3163] = mem_3163_sv2v_reg;
  assign mem[3162] = mem_3162_sv2v_reg;
  assign mem[3161] = mem_3161_sv2v_reg;
  assign mem[3160] = mem_3160_sv2v_reg;
  assign mem[3159] = mem_3159_sv2v_reg;
  assign mem[3158] = mem_3158_sv2v_reg;
  assign mem[3157] = mem_3157_sv2v_reg;
  assign mem[3156] = mem_3156_sv2v_reg;
  assign mem[3155] = mem_3155_sv2v_reg;
  assign mem[3154] = mem_3154_sv2v_reg;
  assign mem[3153] = mem_3153_sv2v_reg;
  assign mem[3152] = mem_3152_sv2v_reg;
  assign mem[3151] = mem_3151_sv2v_reg;
  assign mem[3150] = mem_3150_sv2v_reg;
  assign mem[3149] = mem_3149_sv2v_reg;
  assign mem[3148] = mem_3148_sv2v_reg;
  assign mem[3147] = mem_3147_sv2v_reg;
  assign mem[3146] = mem_3146_sv2v_reg;
  assign mem[3145] = mem_3145_sv2v_reg;
  assign mem[3144] = mem_3144_sv2v_reg;
  assign mem[3143] = mem_3143_sv2v_reg;
  assign mem[3142] = mem_3142_sv2v_reg;
  assign mem[3141] = mem_3141_sv2v_reg;
  assign mem[3140] = mem_3140_sv2v_reg;
  assign mem[3139] = mem_3139_sv2v_reg;
  assign mem[3138] = mem_3138_sv2v_reg;
  assign mem[3137] = mem_3137_sv2v_reg;
  assign mem[3136] = mem_3136_sv2v_reg;
  assign mem[3135] = mem_3135_sv2v_reg;
  assign mem[3134] = mem_3134_sv2v_reg;
  assign mem[3133] = mem_3133_sv2v_reg;
  assign mem[3132] = mem_3132_sv2v_reg;
  assign mem[3131] = mem_3131_sv2v_reg;
  assign mem[3130] = mem_3130_sv2v_reg;
  assign mem[3129] = mem_3129_sv2v_reg;
  assign mem[3128] = mem_3128_sv2v_reg;
  assign mem[3127] = mem_3127_sv2v_reg;
  assign mem[3126] = mem_3126_sv2v_reg;
  assign mem[3125] = mem_3125_sv2v_reg;
  assign mem[3124] = mem_3124_sv2v_reg;
  assign mem[3123] = mem_3123_sv2v_reg;
  assign mem[3122] = mem_3122_sv2v_reg;
  assign mem[3121] = mem_3121_sv2v_reg;
  assign mem[3120] = mem_3120_sv2v_reg;
  assign mem[3119] = mem_3119_sv2v_reg;
  assign mem[3118] = mem_3118_sv2v_reg;
  assign mem[3117] = mem_3117_sv2v_reg;
  assign mem[3116] = mem_3116_sv2v_reg;
  assign mem[3115] = mem_3115_sv2v_reg;
  assign mem[3114] = mem_3114_sv2v_reg;
  assign mem[3113] = mem_3113_sv2v_reg;
  assign mem[3112] = mem_3112_sv2v_reg;
  assign mem[3111] = mem_3111_sv2v_reg;
  assign mem[3110] = mem_3110_sv2v_reg;
  assign mem[3109] = mem_3109_sv2v_reg;
  assign mem[3108] = mem_3108_sv2v_reg;
  assign mem[3107] = mem_3107_sv2v_reg;
  assign mem[3106] = mem_3106_sv2v_reg;
  assign mem[3105] = mem_3105_sv2v_reg;
  assign mem[3104] = mem_3104_sv2v_reg;
  assign mem[3103] = mem_3103_sv2v_reg;
  assign mem[3102] = mem_3102_sv2v_reg;
  assign mem[3101] = mem_3101_sv2v_reg;
  assign mem[3100] = mem_3100_sv2v_reg;
  assign mem[3099] = mem_3099_sv2v_reg;
  assign mem[3098] = mem_3098_sv2v_reg;
  assign mem[3097] = mem_3097_sv2v_reg;
  assign mem[3096] = mem_3096_sv2v_reg;
  assign mem[3095] = mem_3095_sv2v_reg;
  assign mem[3094] = mem_3094_sv2v_reg;
  assign mem[3093] = mem_3093_sv2v_reg;
  assign mem[3092] = mem_3092_sv2v_reg;
  assign mem[3091] = mem_3091_sv2v_reg;
  assign mem[3090] = mem_3090_sv2v_reg;
  assign mem[3089] = mem_3089_sv2v_reg;
  assign mem[3088] = mem_3088_sv2v_reg;
  assign mem[3087] = mem_3087_sv2v_reg;
  assign mem[3086] = mem_3086_sv2v_reg;
  assign mem[3085] = mem_3085_sv2v_reg;
  assign mem[3084] = mem_3084_sv2v_reg;
  assign mem[3083] = mem_3083_sv2v_reg;
  assign mem[3082] = mem_3082_sv2v_reg;
  assign mem[3081] = mem_3081_sv2v_reg;
  assign mem[3080] = mem_3080_sv2v_reg;
  assign mem[3079] = mem_3079_sv2v_reg;
  assign mem[3078] = mem_3078_sv2v_reg;
  assign mem[3077] = mem_3077_sv2v_reg;
  assign mem[3076] = mem_3076_sv2v_reg;
  assign mem[3075] = mem_3075_sv2v_reg;
  assign mem[3074] = mem_3074_sv2v_reg;
  assign mem[3073] = mem_3073_sv2v_reg;
  assign mem[3072] = mem_3072_sv2v_reg;
  assign mem[3071] = mem_3071_sv2v_reg;
  assign mem[3070] = mem_3070_sv2v_reg;
  assign mem[3069] = mem_3069_sv2v_reg;
  assign mem[3068] = mem_3068_sv2v_reg;
  assign mem[3067] = mem_3067_sv2v_reg;
  assign mem[3066] = mem_3066_sv2v_reg;
  assign mem[3065] = mem_3065_sv2v_reg;
  assign mem[3064] = mem_3064_sv2v_reg;
  assign mem[3063] = mem_3063_sv2v_reg;
  assign mem[3062] = mem_3062_sv2v_reg;
  assign mem[3061] = mem_3061_sv2v_reg;
  assign mem[3060] = mem_3060_sv2v_reg;
  assign mem[3059] = mem_3059_sv2v_reg;
  assign mem[3058] = mem_3058_sv2v_reg;
  assign mem[3057] = mem_3057_sv2v_reg;
  assign mem[3056] = mem_3056_sv2v_reg;
  assign mem[3055] = mem_3055_sv2v_reg;
  assign mem[3054] = mem_3054_sv2v_reg;
  assign mem[3053] = mem_3053_sv2v_reg;
  assign mem[3052] = mem_3052_sv2v_reg;
  assign mem[3051] = mem_3051_sv2v_reg;
  assign mem[3050] = mem_3050_sv2v_reg;
  assign mem[3049] = mem_3049_sv2v_reg;
  assign mem[3048] = mem_3048_sv2v_reg;
  assign mem[3047] = mem_3047_sv2v_reg;
  assign mem[3046] = mem_3046_sv2v_reg;
  assign mem[3045] = mem_3045_sv2v_reg;
  assign mem[3044] = mem_3044_sv2v_reg;
  assign mem[3043] = mem_3043_sv2v_reg;
  assign mem[3042] = mem_3042_sv2v_reg;
  assign mem[3041] = mem_3041_sv2v_reg;
  assign mem[3040] = mem_3040_sv2v_reg;
  assign mem[3039] = mem_3039_sv2v_reg;
  assign mem[3038] = mem_3038_sv2v_reg;
  assign mem[3037] = mem_3037_sv2v_reg;
  assign mem[3036] = mem_3036_sv2v_reg;
  assign mem[3035] = mem_3035_sv2v_reg;
  assign mem[3034] = mem_3034_sv2v_reg;
  assign mem[3033] = mem_3033_sv2v_reg;
  assign mem[3032] = mem_3032_sv2v_reg;
  assign mem[3031] = mem_3031_sv2v_reg;
  assign mem[3030] = mem_3030_sv2v_reg;
  assign mem[3029] = mem_3029_sv2v_reg;
  assign mem[3028] = mem_3028_sv2v_reg;
  assign mem[3027] = mem_3027_sv2v_reg;
  assign mem[3026] = mem_3026_sv2v_reg;
  assign mem[3025] = mem_3025_sv2v_reg;
  assign mem[3024] = mem_3024_sv2v_reg;
  assign mem[3023] = mem_3023_sv2v_reg;
  assign mem[3022] = mem_3022_sv2v_reg;
  assign mem[3021] = mem_3021_sv2v_reg;
  assign mem[3020] = mem_3020_sv2v_reg;
  assign mem[3019] = mem_3019_sv2v_reg;
  assign mem[3018] = mem_3018_sv2v_reg;
  assign mem[3017] = mem_3017_sv2v_reg;
  assign mem[3016] = mem_3016_sv2v_reg;
  assign mem[3015] = mem_3015_sv2v_reg;
  assign mem[3014] = mem_3014_sv2v_reg;
  assign mem[3013] = mem_3013_sv2v_reg;
  assign mem[3012] = mem_3012_sv2v_reg;
  assign mem[3011] = mem_3011_sv2v_reg;
  assign mem[3010] = mem_3010_sv2v_reg;
  assign mem[3009] = mem_3009_sv2v_reg;
  assign mem[3008] = mem_3008_sv2v_reg;
  assign mem[3007] = mem_3007_sv2v_reg;
  assign mem[3006] = mem_3006_sv2v_reg;
  assign mem[3005] = mem_3005_sv2v_reg;
  assign mem[3004] = mem_3004_sv2v_reg;
  assign mem[3003] = mem_3003_sv2v_reg;
  assign mem[3002] = mem_3002_sv2v_reg;
  assign mem[3001] = mem_3001_sv2v_reg;
  assign mem[3000] = mem_3000_sv2v_reg;
  assign mem[2999] = mem_2999_sv2v_reg;
  assign mem[2998] = mem_2998_sv2v_reg;
  assign mem[2997] = mem_2997_sv2v_reg;
  assign mem[2996] = mem_2996_sv2v_reg;
  assign mem[2995] = mem_2995_sv2v_reg;
  assign mem[2994] = mem_2994_sv2v_reg;
  assign mem[2993] = mem_2993_sv2v_reg;
  assign mem[2992] = mem_2992_sv2v_reg;
  assign mem[2991] = mem_2991_sv2v_reg;
  assign mem[2990] = mem_2990_sv2v_reg;
  assign mem[2989] = mem_2989_sv2v_reg;
  assign mem[2988] = mem_2988_sv2v_reg;
  assign mem[2987] = mem_2987_sv2v_reg;
  assign mem[2986] = mem_2986_sv2v_reg;
  assign mem[2985] = mem_2985_sv2v_reg;
  assign mem[2984] = mem_2984_sv2v_reg;
  assign mem[2983] = mem_2983_sv2v_reg;
  assign mem[2982] = mem_2982_sv2v_reg;
  assign mem[2981] = mem_2981_sv2v_reg;
  assign mem[2980] = mem_2980_sv2v_reg;
  assign mem[2979] = mem_2979_sv2v_reg;
  assign mem[2978] = mem_2978_sv2v_reg;
  assign mem[2977] = mem_2977_sv2v_reg;
  assign mem[2976] = mem_2976_sv2v_reg;
  assign mem[2975] = mem_2975_sv2v_reg;
  assign mem[2974] = mem_2974_sv2v_reg;
  assign mem[2973] = mem_2973_sv2v_reg;
  assign mem[2972] = mem_2972_sv2v_reg;
  assign mem[2971] = mem_2971_sv2v_reg;
  assign mem[2970] = mem_2970_sv2v_reg;
  assign mem[2969] = mem_2969_sv2v_reg;
  assign mem[2968] = mem_2968_sv2v_reg;
  assign mem[2967] = mem_2967_sv2v_reg;
  assign mem[2966] = mem_2966_sv2v_reg;
  assign mem[2965] = mem_2965_sv2v_reg;
  assign mem[2964] = mem_2964_sv2v_reg;
  assign mem[2963] = mem_2963_sv2v_reg;
  assign mem[2962] = mem_2962_sv2v_reg;
  assign mem[2961] = mem_2961_sv2v_reg;
  assign mem[2960] = mem_2960_sv2v_reg;
  assign mem[2959] = mem_2959_sv2v_reg;
  assign mem[2958] = mem_2958_sv2v_reg;
  assign mem[2957] = mem_2957_sv2v_reg;
  assign mem[2956] = mem_2956_sv2v_reg;
  assign mem[2955] = mem_2955_sv2v_reg;
  assign mem[2954] = mem_2954_sv2v_reg;
  assign mem[2953] = mem_2953_sv2v_reg;
  assign mem[2952] = mem_2952_sv2v_reg;
  assign mem[2951] = mem_2951_sv2v_reg;
  assign mem[2950] = mem_2950_sv2v_reg;
  assign mem[2949] = mem_2949_sv2v_reg;
  assign mem[2948] = mem_2948_sv2v_reg;
  assign mem[2947] = mem_2947_sv2v_reg;
  assign mem[2946] = mem_2946_sv2v_reg;
  assign mem[2945] = mem_2945_sv2v_reg;
  assign mem[2944] = mem_2944_sv2v_reg;
  assign mem[2943] = mem_2943_sv2v_reg;
  assign mem[2942] = mem_2942_sv2v_reg;
  assign mem[2941] = mem_2941_sv2v_reg;
  assign mem[2940] = mem_2940_sv2v_reg;
  assign mem[2939] = mem_2939_sv2v_reg;
  assign mem[2938] = mem_2938_sv2v_reg;
  assign mem[2937] = mem_2937_sv2v_reg;
  assign mem[2936] = mem_2936_sv2v_reg;
  assign mem[2935] = mem_2935_sv2v_reg;
  assign mem[2934] = mem_2934_sv2v_reg;
  assign mem[2933] = mem_2933_sv2v_reg;
  assign mem[2932] = mem_2932_sv2v_reg;
  assign mem[2931] = mem_2931_sv2v_reg;
  assign mem[2930] = mem_2930_sv2v_reg;
  assign mem[2929] = mem_2929_sv2v_reg;
  assign mem[2928] = mem_2928_sv2v_reg;
  assign mem[2927] = mem_2927_sv2v_reg;
  assign mem[2926] = mem_2926_sv2v_reg;
  assign mem[2925] = mem_2925_sv2v_reg;
  assign mem[2924] = mem_2924_sv2v_reg;
  assign mem[2923] = mem_2923_sv2v_reg;
  assign mem[2922] = mem_2922_sv2v_reg;
  assign mem[2921] = mem_2921_sv2v_reg;
  assign mem[2920] = mem_2920_sv2v_reg;
  assign mem[2919] = mem_2919_sv2v_reg;
  assign mem[2918] = mem_2918_sv2v_reg;
  assign mem[2917] = mem_2917_sv2v_reg;
  assign mem[2916] = mem_2916_sv2v_reg;
  assign mem[2915] = mem_2915_sv2v_reg;
  assign mem[2914] = mem_2914_sv2v_reg;
  assign mem[2913] = mem_2913_sv2v_reg;
  assign mem[2912] = mem_2912_sv2v_reg;
  assign mem[2911] = mem_2911_sv2v_reg;
  assign mem[2910] = mem_2910_sv2v_reg;
  assign mem[2909] = mem_2909_sv2v_reg;
  assign mem[2908] = mem_2908_sv2v_reg;
  assign mem[2907] = mem_2907_sv2v_reg;
  assign mem[2906] = mem_2906_sv2v_reg;
  assign mem[2905] = mem_2905_sv2v_reg;
  assign mem[2904] = mem_2904_sv2v_reg;
  assign mem[2903] = mem_2903_sv2v_reg;
  assign mem[2902] = mem_2902_sv2v_reg;
  assign mem[2901] = mem_2901_sv2v_reg;
  assign mem[2900] = mem_2900_sv2v_reg;
  assign mem[2899] = mem_2899_sv2v_reg;
  assign mem[2898] = mem_2898_sv2v_reg;
  assign mem[2897] = mem_2897_sv2v_reg;
  assign mem[2896] = mem_2896_sv2v_reg;
  assign mem[2895] = mem_2895_sv2v_reg;
  assign mem[2894] = mem_2894_sv2v_reg;
  assign mem[2893] = mem_2893_sv2v_reg;
  assign mem[2892] = mem_2892_sv2v_reg;
  assign mem[2891] = mem_2891_sv2v_reg;
  assign mem[2890] = mem_2890_sv2v_reg;
  assign mem[2889] = mem_2889_sv2v_reg;
  assign mem[2888] = mem_2888_sv2v_reg;
  assign mem[2887] = mem_2887_sv2v_reg;
  assign mem[2886] = mem_2886_sv2v_reg;
  assign mem[2885] = mem_2885_sv2v_reg;
  assign mem[2884] = mem_2884_sv2v_reg;
  assign mem[2883] = mem_2883_sv2v_reg;
  assign mem[2882] = mem_2882_sv2v_reg;
  assign mem[2881] = mem_2881_sv2v_reg;
  assign mem[2880] = mem_2880_sv2v_reg;
  assign mem[2879] = mem_2879_sv2v_reg;
  assign mem[2878] = mem_2878_sv2v_reg;
  assign mem[2877] = mem_2877_sv2v_reg;
  assign mem[2876] = mem_2876_sv2v_reg;
  assign mem[2875] = mem_2875_sv2v_reg;
  assign mem[2874] = mem_2874_sv2v_reg;
  assign mem[2873] = mem_2873_sv2v_reg;
  assign mem[2872] = mem_2872_sv2v_reg;
  assign mem[2871] = mem_2871_sv2v_reg;
  assign mem[2870] = mem_2870_sv2v_reg;
  assign mem[2869] = mem_2869_sv2v_reg;
  assign mem[2868] = mem_2868_sv2v_reg;
  assign mem[2867] = mem_2867_sv2v_reg;
  assign mem[2866] = mem_2866_sv2v_reg;
  assign mem[2865] = mem_2865_sv2v_reg;
  assign mem[2864] = mem_2864_sv2v_reg;
  assign mem[2863] = mem_2863_sv2v_reg;
  assign mem[2862] = mem_2862_sv2v_reg;
  assign mem[2861] = mem_2861_sv2v_reg;
  assign mem[2860] = mem_2860_sv2v_reg;
  assign mem[2859] = mem_2859_sv2v_reg;
  assign mem[2858] = mem_2858_sv2v_reg;
  assign mem[2857] = mem_2857_sv2v_reg;
  assign mem[2856] = mem_2856_sv2v_reg;
  assign mem[2855] = mem_2855_sv2v_reg;
  assign mem[2854] = mem_2854_sv2v_reg;
  assign mem[2853] = mem_2853_sv2v_reg;
  assign mem[2852] = mem_2852_sv2v_reg;
  assign mem[2851] = mem_2851_sv2v_reg;
  assign mem[2850] = mem_2850_sv2v_reg;
  assign mem[2849] = mem_2849_sv2v_reg;
  assign mem[2848] = mem_2848_sv2v_reg;
  assign mem[2847] = mem_2847_sv2v_reg;
  assign mem[2846] = mem_2846_sv2v_reg;
  assign mem[2845] = mem_2845_sv2v_reg;
  assign mem[2844] = mem_2844_sv2v_reg;
  assign mem[2843] = mem_2843_sv2v_reg;
  assign mem[2842] = mem_2842_sv2v_reg;
  assign mem[2841] = mem_2841_sv2v_reg;
  assign mem[2840] = mem_2840_sv2v_reg;
  assign mem[2839] = mem_2839_sv2v_reg;
  assign mem[2838] = mem_2838_sv2v_reg;
  assign mem[2837] = mem_2837_sv2v_reg;
  assign mem[2836] = mem_2836_sv2v_reg;
  assign mem[2835] = mem_2835_sv2v_reg;
  assign mem[2834] = mem_2834_sv2v_reg;
  assign mem[2833] = mem_2833_sv2v_reg;
  assign mem[2832] = mem_2832_sv2v_reg;
  assign mem[2831] = mem_2831_sv2v_reg;
  assign mem[2830] = mem_2830_sv2v_reg;
  assign mem[2829] = mem_2829_sv2v_reg;
  assign mem[2828] = mem_2828_sv2v_reg;
  assign mem[2827] = mem_2827_sv2v_reg;
  assign mem[2826] = mem_2826_sv2v_reg;
  assign mem[2825] = mem_2825_sv2v_reg;
  assign mem[2824] = mem_2824_sv2v_reg;
  assign mem[2823] = mem_2823_sv2v_reg;
  assign mem[2822] = mem_2822_sv2v_reg;
  assign mem[2821] = mem_2821_sv2v_reg;
  assign mem[2820] = mem_2820_sv2v_reg;
  assign mem[2819] = mem_2819_sv2v_reg;
  assign mem[2818] = mem_2818_sv2v_reg;
  assign mem[2817] = mem_2817_sv2v_reg;
  assign mem[2816] = mem_2816_sv2v_reg;
  assign mem[2815] = mem_2815_sv2v_reg;
  assign mem[2814] = mem_2814_sv2v_reg;
  assign mem[2813] = mem_2813_sv2v_reg;
  assign mem[2812] = mem_2812_sv2v_reg;
  assign mem[2811] = mem_2811_sv2v_reg;
  assign mem[2810] = mem_2810_sv2v_reg;
  assign mem[2809] = mem_2809_sv2v_reg;
  assign mem[2808] = mem_2808_sv2v_reg;
  assign mem[2807] = mem_2807_sv2v_reg;
  assign mem[2806] = mem_2806_sv2v_reg;
  assign mem[2805] = mem_2805_sv2v_reg;
  assign mem[2804] = mem_2804_sv2v_reg;
  assign mem[2803] = mem_2803_sv2v_reg;
  assign mem[2802] = mem_2802_sv2v_reg;
  assign mem[2801] = mem_2801_sv2v_reg;
  assign mem[2800] = mem_2800_sv2v_reg;
  assign mem[2799] = mem_2799_sv2v_reg;
  assign mem[2798] = mem_2798_sv2v_reg;
  assign mem[2797] = mem_2797_sv2v_reg;
  assign mem[2796] = mem_2796_sv2v_reg;
  assign mem[2795] = mem_2795_sv2v_reg;
  assign mem[2794] = mem_2794_sv2v_reg;
  assign mem[2793] = mem_2793_sv2v_reg;
  assign mem[2792] = mem_2792_sv2v_reg;
  assign mem[2791] = mem_2791_sv2v_reg;
  assign mem[2790] = mem_2790_sv2v_reg;
  assign mem[2789] = mem_2789_sv2v_reg;
  assign mem[2788] = mem_2788_sv2v_reg;
  assign mem[2787] = mem_2787_sv2v_reg;
  assign mem[2786] = mem_2786_sv2v_reg;
  assign mem[2785] = mem_2785_sv2v_reg;
  assign mem[2784] = mem_2784_sv2v_reg;
  assign mem[2783] = mem_2783_sv2v_reg;
  assign mem[2782] = mem_2782_sv2v_reg;
  assign mem[2781] = mem_2781_sv2v_reg;
  assign mem[2780] = mem_2780_sv2v_reg;
  assign mem[2779] = mem_2779_sv2v_reg;
  assign mem[2778] = mem_2778_sv2v_reg;
  assign mem[2777] = mem_2777_sv2v_reg;
  assign mem[2776] = mem_2776_sv2v_reg;
  assign mem[2775] = mem_2775_sv2v_reg;
  assign mem[2774] = mem_2774_sv2v_reg;
  assign mem[2773] = mem_2773_sv2v_reg;
  assign mem[2772] = mem_2772_sv2v_reg;
  assign mem[2771] = mem_2771_sv2v_reg;
  assign mem[2770] = mem_2770_sv2v_reg;
  assign mem[2769] = mem_2769_sv2v_reg;
  assign mem[2768] = mem_2768_sv2v_reg;
  assign mem[2767] = mem_2767_sv2v_reg;
  assign mem[2766] = mem_2766_sv2v_reg;
  assign mem[2765] = mem_2765_sv2v_reg;
  assign mem[2764] = mem_2764_sv2v_reg;
  assign mem[2763] = mem_2763_sv2v_reg;
  assign mem[2762] = mem_2762_sv2v_reg;
  assign mem[2761] = mem_2761_sv2v_reg;
  assign mem[2760] = mem_2760_sv2v_reg;
  assign mem[2759] = mem_2759_sv2v_reg;
  assign mem[2758] = mem_2758_sv2v_reg;
  assign mem[2757] = mem_2757_sv2v_reg;
  assign mem[2756] = mem_2756_sv2v_reg;
  assign mem[2755] = mem_2755_sv2v_reg;
  assign mem[2754] = mem_2754_sv2v_reg;
  assign mem[2753] = mem_2753_sv2v_reg;
  assign mem[2752] = mem_2752_sv2v_reg;
  assign mem[2751] = mem_2751_sv2v_reg;
  assign mem[2750] = mem_2750_sv2v_reg;
  assign mem[2749] = mem_2749_sv2v_reg;
  assign mem[2748] = mem_2748_sv2v_reg;
  assign mem[2747] = mem_2747_sv2v_reg;
  assign mem[2746] = mem_2746_sv2v_reg;
  assign mem[2745] = mem_2745_sv2v_reg;
  assign mem[2744] = mem_2744_sv2v_reg;
  assign mem[2743] = mem_2743_sv2v_reg;
  assign mem[2742] = mem_2742_sv2v_reg;
  assign mem[2741] = mem_2741_sv2v_reg;
  assign mem[2740] = mem_2740_sv2v_reg;
  assign mem[2739] = mem_2739_sv2v_reg;
  assign mem[2738] = mem_2738_sv2v_reg;
  assign mem[2737] = mem_2737_sv2v_reg;
  assign mem[2736] = mem_2736_sv2v_reg;
  assign mem[2735] = mem_2735_sv2v_reg;
  assign mem[2734] = mem_2734_sv2v_reg;
  assign mem[2733] = mem_2733_sv2v_reg;
  assign mem[2732] = mem_2732_sv2v_reg;
  assign mem[2731] = mem_2731_sv2v_reg;
  assign mem[2730] = mem_2730_sv2v_reg;
  assign mem[2729] = mem_2729_sv2v_reg;
  assign mem[2728] = mem_2728_sv2v_reg;
  assign mem[2727] = mem_2727_sv2v_reg;
  assign mem[2726] = mem_2726_sv2v_reg;
  assign mem[2725] = mem_2725_sv2v_reg;
  assign mem[2724] = mem_2724_sv2v_reg;
  assign mem[2723] = mem_2723_sv2v_reg;
  assign mem[2722] = mem_2722_sv2v_reg;
  assign mem[2721] = mem_2721_sv2v_reg;
  assign mem[2720] = mem_2720_sv2v_reg;
  assign mem[2719] = mem_2719_sv2v_reg;
  assign mem[2718] = mem_2718_sv2v_reg;
  assign mem[2717] = mem_2717_sv2v_reg;
  assign mem[2716] = mem_2716_sv2v_reg;
  assign mem[2715] = mem_2715_sv2v_reg;
  assign mem[2714] = mem_2714_sv2v_reg;
  assign mem[2713] = mem_2713_sv2v_reg;
  assign mem[2712] = mem_2712_sv2v_reg;
  assign mem[2711] = mem_2711_sv2v_reg;
  assign mem[2710] = mem_2710_sv2v_reg;
  assign mem[2709] = mem_2709_sv2v_reg;
  assign mem[2708] = mem_2708_sv2v_reg;
  assign mem[2707] = mem_2707_sv2v_reg;
  assign mem[2706] = mem_2706_sv2v_reg;
  assign mem[2705] = mem_2705_sv2v_reg;
  assign mem[2704] = mem_2704_sv2v_reg;
  assign mem[2703] = mem_2703_sv2v_reg;
  assign mem[2702] = mem_2702_sv2v_reg;
  assign mem[2701] = mem_2701_sv2v_reg;
  assign mem[2700] = mem_2700_sv2v_reg;
  assign mem[2699] = mem_2699_sv2v_reg;
  assign mem[2698] = mem_2698_sv2v_reg;
  assign mem[2697] = mem_2697_sv2v_reg;
  assign mem[2696] = mem_2696_sv2v_reg;
  assign mem[2695] = mem_2695_sv2v_reg;
  assign mem[2694] = mem_2694_sv2v_reg;
  assign mem[2693] = mem_2693_sv2v_reg;
  assign mem[2692] = mem_2692_sv2v_reg;
  assign mem[2691] = mem_2691_sv2v_reg;
  assign mem[2690] = mem_2690_sv2v_reg;
  assign mem[2689] = mem_2689_sv2v_reg;
  assign mem[2688] = mem_2688_sv2v_reg;
  assign mem[2687] = mem_2687_sv2v_reg;
  assign mem[2686] = mem_2686_sv2v_reg;
  assign mem[2685] = mem_2685_sv2v_reg;
  assign mem[2684] = mem_2684_sv2v_reg;
  assign mem[2683] = mem_2683_sv2v_reg;
  assign mem[2682] = mem_2682_sv2v_reg;
  assign mem[2681] = mem_2681_sv2v_reg;
  assign mem[2680] = mem_2680_sv2v_reg;
  assign mem[2679] = mem_2679_sv2v_reg;
  assign mem[2678] = mem_2678_sv2v_reg;
  assign mem[2677] = mem_2677_sv2v_reg;
  assign mem[2676] = mem_2676_sv2v_reg;
  assign mem[2675] = mem_2675_sv2v_reg;
  assign mem[2674] = mem_2674_sv2v_reg;
  assign mem[2673] = mem_2673_sv2v_reg;
  assign mem[2672] = mem_2672_sv2v_reg;
  assign mem[2671] = mem_2671_sv2v_reg;
  assign mem[2670] = mem_2670_sv2v_reg;
  assign mem[2669] = mem_2669_sv2v_reg;
  assign mem[2668] = mem_2668_sv2v_reg;
  assign mem[2667] = mem_2667_sv2v_reg;
  assign mem[2666] = mem_2666_sv2v_reg;
  assign mem[2665] = mem_2665_sv2v_reg;
  assign mem[2664] = mem_2664_sv2v_reg;
  assign mem[2663] = mem_2663_sv2v_reg;
  assign mem[2662] = mem_2662_sv2v_reg;
  assign mem[2661] = mem_2661_sv2v_reg;
  assign mem[2660] = mem_2660_sv2v_reg;
  assign mem[2659] = mem_2659_sv2v_reg;
  assign mem[2658] = mem_2658_sv2v_reg;
  assign mem[2657] = mem_2657_sv2v_reg;
  assign mem[2656] = mem_2656_sv2v_reg;
  assign mem[2655] = mem_2655_sv2v_reg;
  assign mem[2654] = mem_2654_sv2v_reg;
  assign mem[2653] = mem_2653_sv2v_reg;
  assign mem[2652] = mem_2652_sv2v_reg;
  assign mem[2651] = mem_2651_sv2v_reg;
  assign mem[2650] = mem_2650_sv2v_reg;
  assign mem[2649] = mem_2649_sv2v_reg;
  assign mem[2648] = mem_2648_sv2v_reg;
  assign mem[2647] = mem_2647_sv2v_reg;
  assign mem[2646] = mem_2646_sv2v_reg;
  assign mem[2645] = mem_2645_sv2v_reg;
  assign mem[2644] = mem_2644_sv2v_reg;
  assign mem[2643] = mem_2643_sv2v_reg;
  assign mem[2642] = mem_2642_sv2v_reg;
  assign mem[2641] = mem_2641_sv2v_reg;
  assign mem[2640] = mem_2640_sv2v_reg;
  assign mem[2639] = mem_2639_sv2v_reg;
  assign mem[2638] = mem_2638_sv2v_reg;
  assign mem[2637] = mem_2637_sv2v_reg;
  assign mem[2636] = mem_2636_sv2v_reg;
  assign mem[2635] = mem_2635_sv2v_reg;
  assign mem[2634] = mem_2634_sv2v_reg;
  assign mem[2633] = mem_2633_sv2v_reg;
  assign mem[2632] = mem_2632_sv2v_reg;
  assign mem[2631] = mem_2631_sv2v_reg;
  assign mem[2630] = mem_2630_sv2v_reg;
  assign mem[2629] = mem_2629_sv2v_reg;
  assign mem[2628] = mem_2628_sv2v_reg;
  assign mem[2627] = mem_2627_sv2v_reg;
  assign mem[2626] = mem_2626_sv2v_reg;
  assign mem[2625] = mem_2625_sv2v_reg;
  assign mem[2624] = mem_2624_sv2v_reg;
  assign mem[2623] = mem_2623_sv2v_reg;
  assign mem[2622] = mem_2622_sv2v_reg;
  assign mem[2621] = mem_2621_sv2v_reg;
  assign mem[2620] = mem_2620_sv2v_reg;
  assign mem[2619] = mem_2619_sv2v_reg;
  assign mem[2618] = mem_2618_sv2v_reg;
  assign mem[2617] = mem_2617_sv2v_reg;
  assign mem[2616] = mem_2616_sv2v_reg;
  assign mem[2615] = mem_2615_sv2v_reg;
  assign mem[2614] = mem_2614_sv2v_reg;
  assign mem[2613] = mem_2613_sv2v_reg;
  assign mem[2612] = mem_2612_sv2v_reg;
  assign mem[2611] = mem_2611_sv2v_reg;
  assign mem[2610] = mem_2610_sv2v_reg;
  assign mem[2609] = mem_2609_sv2v_reg;
  assign mem[2608] = mem_2608_sv2v_reg;
  assign mem[2607] = mem_2607_sv2v_reg;
  assign mem[2606] = mem_2606_sv2v_reg;
  assign mem[2605] = mem_2605_sv2v_reg;
  assign mem[2604] = mem_2604_sv2v_reg;
  assign mem[2603] = mem_2603_sv2v_reg;
  assign mem[2602] = mem_2602_sv2v_reg;
  assign mem[2601] = mem_2601_sv2v_reg;
  assign mem[2600] = mem_2600_sv2v_reg;
  assign mem[2599] = mem_2599_sv2v_reg;
  assign mem[2598] = mem_2598_sv2v_reg;
  assign mem[2597] = mem_2597_sv2v_reg;
  assign mem[2596] = mem_2596_sv2v_reg;
  assign mem[2595] = mem_2595_sv2v_reg;
  assign mem[2594] = mem_2594_sv2v_reg;
  assign mem[2593] = mem_2593_sv2v_reg;
  assign mem[2592] = mem_2592_sv2v_reg;
  assign mem[2591] = mem_2591_sv2v_reg;
  assign mem[2590] = mem_2590_sv2v_reg;
  assign mem[2589] = mem_2589_sv2v_reg;
  assign mem[2588] = mem_2588_sv2v_reg;
  assign mem[2587] = mem_2587_sv2v_reg;
  assign mem[2586] = mem_2586_sv2v_reg;
  assign mem[2585] = mem_2585_sv2v_reg;
  assign mem[2584] = mem_2584_sv2v_reg;
  assign mem[2583] = mem_2583_sv2v_reg;
  assign mem[2582] = mem_2582_sv2v_reg;
  assign mem[2581] = mem_2581_sv2v_reg;
  assign mem[2580] = mem_2580_sv2v_reg;
  assign mem[2579] = mem_2579_sv2v_reg;
  assign mem[2578] = mem_2578_sv2v_reg;
  assign mem[2577] = mem_2577_sv2v_reg;
  assign mem[2576] = mem_2576_sv2v_reg;
  assign mem[2575] = mem_2575_sv2v_reg;
  assign mem[2574] = mem_2574_sv2v_reg;
  assign mem[2573] = mem_2573_sv2v_reg;
  assign mem[2572] = mem_2572_sv2v_reg;
  assign mem[2571] = mem_2571_sv2v_reg;
  assign mem[2570] = mem_2570_sv2v_reg;
  assign mem[2569] = mem_2569_sv2v_reg;
  assign mem[2568] = mem_2568_sv2v_reg;
  assign mem[2567] = mem_2567_sv2v_reg;
  assign mem[2566] = mem_2566_sv2v_reg;
  assign mem[2565] = mem_2565_sv2v_reg;
  assign mem[2564] = mem_2564_sv2v_reg;
  assign mem[2563] = mem_2563_sv2v_reg;
  assign mem[2562] = mem_2562_sv2v_reg;
  assign mem[2561] = mem_2561_sv2v_reg;
  assign mem[2560] = mem_2560_sv2v_reg;
  assign mem[2559] = mem_2559_sv2v_reg;
  assign mem[2558] = mem_2558_sv2v_reg;
  assign mem[2557] = mem_2557_sv2v_reg;
  assign mem[2556] = mem_2556_sv2v_reg;
  assign mem[2555] = mem_2555_sv2v_reg;
  assign mem[2554] = mem_2554_sv2v_reg;
  assign mem[2553] = mem_2553_sv2v_reg;
  assign mem[2552] = mem_2552_sv2v_reg;
  assign mem[2551] = mem_2551_sv2v_reg;
  assign mem[2550] = mem_2550_sv2v_reg;
  assign mem[2549] = mem_2549_sv2v_reg;
  assign mem[2548] = mem_2548_sv2v_reg;
  assign mem[2547] = mem_2547_sv2v_reg;
  assign mem[2546] = mem_2546_sv2v_reg;
  assign mem[2545] = mem_2545_sv2v_reg;
  assign mem[2544] = mem_2544_sv2v_reg;
  assign mem[2543] = mem_2543_sv2v_reg;
  assign mem[2542] = mem_2542_sv2v_reg;
  assign mem[2541] = mem_2541_sv2v_reg;
  assign mem[2540] = mem_2540_sv2v_reg;
  assign mem[2539] = mem_2539_sv2v_reg;
  assign mem[2538] = mem_2538_sv2v_reg;
  assign mem[2537] = mem_2537_sv2v_reg;
  assign mem[2536] = mem_2536_sv2v_reg;
  assign mem[2535] = mem_2535_sv2v_reg;
  assign mem[2534] = mem_2534_sv2v_reg;
  assign mem[2533] = mem_2533_sv2v_reg;
  assign mem[2532] = mem_2532_sv2v_reg;
  assign mem[2531] = mem_2531_sv2v_reg;
  assign mem[2530] = mem_2530_sv2v_reg;
  assign mem[2529] = mem_2529_sv2v_reg;
  assign mem[2528] = mem_2528_sv2v_reg;
  assign mem[2527] = mem_2527_sv2v_reg;
  assign mem[2526] = mem_2526_sv2v_reg;
  assign mem[2525] = mem_2525_sv2v_reg;
  assign mem[2524] = mem_2524_sv2v_reg;
  assign mem[2523] = mem_2523_sv2v_reg;
  assign mem[2522] = mem_2522_sv2v_reg;
  assign mem[2521] = mem_2521_sv2v_reg;
  assign mem[2520] = mem_2520_sv2v_reg;
  assign mem[2519] = mem_2519_sv2v_reg;
  assign mem[2518] = mem_2518_sv2v_reg;
  assign mem[2517] = mem_2517_sv2v_reg;
  assign mem[2516] = mem_2516_sv2v_reg;
  assign mem[2515] = mem_2515_sv2v_reg;
  assign mem[2514] = mem_2514_sv2v_reg;
  assign mem[2513] = mem_2513_sv2v_reg;
  assign mem[2512] = mem_2512_sv2v_reg;
  assign mem[2511] = mem_2511_sv2v_reg;
  assign mem[2510] = mem_2510_sv2v_reg;
  assign mem[2509] = mem_2509_sv2v_reg;
  assign mem[2508] = mem_2508_sv2v_reg;
  assign mem[2507] = mem_2507_sv2v_reg;
  assign mem[2506] = mem_2506_sv2v_reg;
  assign mem[2505] = mem_2505_sv2v_reg;
  assign mem[2504] = mem_2504_sv2v_reg;
  assign mem[2503] = mem_2503_sv2v_reg;
  assign mem[2502] = mem_2502_sv2v_reg;
  assign mem[2501] = mem_2501_sv2v_reg;
  assign mem[2500] = mem_2500_sv2v_reg;
  assign mem[2499] = mem_2499_sv2v_reg;
  assign mem[2498] = mem_2498_sv2v_reg;
  assign mem[2497] = mem_2497_sv2v_reg;
  assign mem[2496] = mem_2496_sv2v_reg;
  assign mem[2495] = mem_2495_sv2v_reg;
  assign mem[2494] = mem_2494_sv2v_reg;
  assign mem[2493] = mem_2493_sv2v_reg;
  assign mem[2492] = mem_2492_sv2v_reg;
  assign mem[2491] = mem_2491_sv2v_reg;
  assign mem[2490] = mem_2490_sv2v_reg;
  assign mem[2489] = mem_2489_sv2v_reg;
  assign mem[2488] = mem_2488_sv2v_reg;
  assign mem[2487] = mem_2487_sv2v_reg;
  assign mem[2486] = mem_2486_sv2v_reg;
  assign mem[2485] = mem_2485_sv2v_reg;
  assign mem[2484] = mem_2484_sv2v_reg;
  assign mem[2483] = mem_2483_sv2v_reg;
  assign mem[2482] = mem_2482_sv2v_reg;
  assign mem[2481] = mem_2481_sv2v_reg;
  assign mem[2480] = mem_2480_sv2v_reg;
  assign mem[2479] = mem_2479_sv2v_reg;
  assign mem[2478] = mem_2478_sv2v_reg;
  assign mem[2477] = mem_2477_sv2v_reg;
  assign mem[2476] = mem_2476_sv2v_reg;
  assign mem[2475] = mem_2475_sv2v_reg;
  assign mem[2474] = mem_2474_sv2v_reg;
  assign mem[2473] = mem_2473_sv2v_reg;
  assign mem[2472] = mem_2472_sv2v_reg;
  assign mem[2471] = mem_2471_sv2v_reg;
  assign mem[2470] = mem_2470_sv2v_reg;
  assign mem[2469] = mem_2469_sv2v_reg;
  assign mem[2468] = mem_2468_sv2v_reg;
  assign mem[2467] = mem_2467_sv2v_reg;
  assign mem[2466] = mem_2466_sv2v_reg;
  assign mem[2465] = mem_2465_sv2v_reg;
  assign mem[2464] = mem_2464_sv2v_reg;
  assign mem[2463] = mem_2463_sv2v_reg;
  assign mem[2462] = mem_2462_sv2v_reg;
  assign mem[2461] = mem_2461_sv2v_reg;
  assign mem[2460] = mem_2460_sv2v_reg;
  assign mem[2459] = mem_2459_sv2v_reg;
  assign mem[2458] = mem_2458_sv2v_reg;
  assign mem[2457] = mem_2457_sv2v_reg;
  assign mem[2456] = mem_2456_sv2v_reg;
  assign mem[2455] = mem_2455_sv2v_reg;
  assign mem[2454] = mem_2454_sv2v_reg;
  assign mem[2453] = mem_2453_sv2v_reg;
  assign mem[2452] = mem_2452_sv2v_reg;
  assign mem[2451] = mem_2451_sv2v_reg;
  assign mem[2450] = mem_2450_sv2v_reg;
  assign mem[2449] = mem_2449_sv2v_reg;
  assign mem[2448] = mem_2448_sv2v_reg;
  assign mem[2447] = mem_2447_sv2v_reg;
  assign mem[2446] = mem_2446_sv2v_reg;
  assign mem[2445] = mem_2445_sv2v_reg;
  assign mem[2444] = mem_2444_sv2v_reg;
  assign mem[2443] = mem_2443_sv2v_reg;
  assign mem[2442] = mem_2442_sv2v_reg;
  assign mem[2441] = mem_2441_sv2v_reg;
  assign mem[2440] = mem_2440_sv2v_reg;
  assign mem[2439] = mem_2439_sv2v_reg;
  assign mem[2438] = mem_2438_sv2v_reg;
  assign mem[2437] = mem_2437_sv2v_reg;
  assign mem[2436] = mem_2436_sv2v_reg;
  assign mem[2435] = mem_2435_sv2v_reg;
  assign mem[2434] = mem_2434_sv2v_reg;
  assign mem[2433] = mem_2433_sv2v_reg;
  assign mem[2432] = mem_2432_sv2v_reg;
  assign mem[2431] = mem_2431_sv2v_reg;
  assign mem[2430] = mem_2430_sv2v_reg;
  assign mem[2429] = mem_2429_sv2v_reg;
  assign mem[2428] = mem_2428_sv2v_reg;
  assign mem[2427] = mem_2427_sv2v_reg;
  assign mem[2426] = mem_2426_sv2v_reg;
  assign mem[2425] = mem_2425_sv2v_reg;
  assign mem[2424] = mem_2424_sv2v_reg;
  assign mem[2423] = mem_2423_sv2v_reg;
  assign mem[2422] = mem_2422_sv2v_reg;
  assign mem[2421] = mem_2421_sv2v_reg;
  assign mem[2420] = mem_2420_sv2v_reg;
  assign mem[2419] = mem_2419_sv2v_reg;
  assign mem[2418] = mem_2418_sv2v_reg;
  assign mem[2417] = mem_2417_sv2v_reg;
  assign mem[2416] = mem_2416_sv2v_reg;
  assign mem[2415] = mem_2415_sv2v_reg;
  assign mem[2414] = mem_2414_sv2v_reg;
  assign mem[2413] = mem_2413_sv2v_reg;
  assign mem[2412] = mem_2412_sv2v_reg;
  assign mem[2411] = mem_2411_sv2v_reg;
  assign mem[2410] = mem_2410_sv2v_reg;
  assign mem[2409] = mem_2409_sv2v_reg;
  assign mem[2408] = mem_2408_sv2v_reg;
  assign mem[2407] = mem_2407_sv2v_reg;
  assign mem[2406] = mem_2406_sv2v_reg;
  assign mem[2405] = mem_2405_sv2v_reg;
  assign mem[2404] = mem_2404_sv2v_reg;
  assign mem[2403] = mem_2403_sv2v_reg;
  assign mem[2402] = mem_2402_sv2v_reg;
  assign mem[2401] = mem_2401_sv2v_reg;
  assign mem[2400] = mem_2400_sv2v_reg;
  assign mem[2399] = mem_2399_sv2v_reg;
  assign mem[2398] = mem_2398_sv2v_reg;
  assign mem[2397] = mem_2397_sv2v_reg;
  assign mem[2396] = mem_2396_sv2v_reg;
  assign mem[2395] = mem_2395_sv2v_reg;
  assign mem[2394] = mem_2394_sv2v_reg;
  assign mem[2393] = mem_2393_sv2v_reg;
  assign mem[2392] = mem_2392_sv2v_reg;
  assign mem[2391] = mem_2391_sv2v_reg;
  assign mem[2390] = mem_2390_sv2v_reg;
  assign mem[2389] = mem_2389_sv2v_reg;
  assign mem[2388] = mem_2388_sv2v_reg;
  assign mem[2387] = mem_2387_sv2v_reg;
  assign mem[2386] = mem_2386_sv2v_reg;
  assign mem[2385] = mem_2385_sv2v_reg;
  assign mem[2384] = mem_2384_sv2v_reg;
  assign mem[2383] = mem_2383_sv2v_reg;
  assign mem[2382] = mem_2382_sv2v_reg;
  assign mem[2381] = mem_2381_sv2v_reg;
  assign mem[2380] = mem_2380_sv2v_reg;
  assign mem[2379] = mem_2379_sv2v_reg;
  assign mem[2378] = mem_2378_sv2v_reg;
  assign mem[2377] = mem_2377_sv2v_reg;
  assign mem[2376] = mem_2376_sv2v_reg;
  assign mem[2375] = mem_2375_sv2v_reg;
  assign mem[2374] = mem_2374_sv2v_reg;
  assign mem[2373] = mem_2373_sv2v_reg;
  assign mem[2372] = mem_2372_sv2v_reg;
  assign mem[2371] = mem_2371_sv2v_reg;
  assign mem[2370] = mem_2370_sv2v_reg;
  assign mem[2369] = mem_2369_sv2v_reg;
  assign mem[2368] = mem_2368_sv2v_reg;
  assign mem[2367] = mem_2367_sv2v_reg;
  assign mem[2366] = mem_2366_sv2v_reg;
  assign mem[2365] = mem_2365_sv2v_reg;
  assign mem[2364] = mem_2364_sv2v_reg;
  assign mem[2363] = mem_2363_sv2v_reg;
  assign mem[2362] = mem_2362_sv2v_reg;
  assign mem[2361] = mem_2361_sv2v_reg;
  assign mem[2360] = mem_2360_sv2v_reg;
  assign mem[2359] = mem_2359_sv2v_reg;
  assign mem[2358] = mem_2358_sv2v_reg;
  assign mem[2357] = mem_2357_sv2v_reg;
  assign mem[2356] = mem_2356_sv2v_reg;
  assign mem[2355] = mem_2355_sv2v_reg;
  assign mem[2354] = mem_2354_sv2v_reg;
  assign mem[2353] = mem_2353_sv2v_reg;
  assign mem[2352] = mem_2352_sv2v_reg;
  assign mem[2351] = mem_2351_sv2v_reg;
  assign mem[2350] = mem_2350_sv2v_reg;
  assign mem[2349] = mem_2349_sv2v_reg;
  assign mem[2348] = mem_2348_sv2v_reg;
  assign mem[2347] = mem_2347_sv2v_reg;
  assign mem[2346] = mem_2346_sv2v_reg;
  assign mem[2345] = mem_2345_sv2v_reg;
  assign mem[2344] = mem_2344_sv2v_reg;
  assign mem[2343] = mem_2343_sv2v_reg;
  assign mem[2342] = mem_2342_sv2v_reg;
  assign mem[2341] = mem_2341_sv2v_reg;
  assign mem[2340] = mem_2340_sv2v_reg;
  assign mem[2339] = mem_2339_sv2v_reg;
  assign mem[2338] = mem_2338_sv2v_reg;
  assign mem[2337] = mem_2337_sv2v_reg;
  assign mem[2336] = mem_2336_sv2v_reg;
  assign mem[2335] = mem_2335_sv2v_reg;
  assign mem[2334] = mem_2334_sv2v_reg;
  assign mem[2333] = mem_2333_sv2v_reg;
  assign mem[2332] = mem_2332_sv2v_reg;
  assign mem[2331] = mem_2331_sv2v_reg;
  assign mem[2330] = mem_2330_sv2v_reg;
  assign mem[2329] = mem_2329_sv2v_reg;
  assign mem[2328] = mem_2328_sv2v_reg;
  assign mem[2327] = mem_2327_sv2v_reg;
  assign mem[2326] = mem_2326_sv2v_reg;
  assign mem[2325] = mem_2325_sv2v_reg;
  assign mem[2324] = mem_2324_sv2v_reg;
  assign mem[2323] = mem_2323_sv2v_reg;
  assign mem[2322] = mem_2322_sv2v_reg;
  assign mem[2321] = mem_2321_sv2v_reg;
  assign mem[2320] = mem_2320_sv2v_reg;
  assign mem[2319] = mem_2319_sv2v_reg;
  assign mem[2318] = mem_2318_sv2v_reg;
  assign mem[2317] = mem_2317_sv2v_reg;
  assign mem[2316] = mem_2316_sv2v_reg;
  assign mem[2315] = mem_2315_sv2v_reg;
  assign mem[2314] = mem_2314_sv2v_reg;
  assign mem[2313] = mem_2313_sv2v_reg;
  assign mem[2312] = mem_2312_sv2v_reg;
  assign mem[2311] = mem_2311_sv2v_reg;
  assign mem[2310] = mem_2310_sv2v_reg;
  assign mem[2309] = mem_2309_sv2v_reg;
  assign mem[2308] = mem_2308_sv2v_reg;
  assign mem[2307] = mem_2307_sv2v_reg;
  assign mem[2306] = mem_2306_sv2v_reg;
  assign mem[2305] = mem_2305_sv2v_reg;
  assign mem[2304] = mem_2304_sv2v_reg;
  assign mem[2303] = mem_2303_sv2v_reg;
  assign mem[2302] = mem_2302_sv2v_reg;
  assign mem[2301] = mem_2301_sv2v_reg;
  assign mem[2300] = mem_2300_sv2v_reg;
  assign mem[2299] = mem_2299_sv2v_reg;
  assign mem[2298] = mem_2298_sv2v_reg;
  assign mem[2297] = mem_2297_sv2v_reg;
  assign mem[2296] = mem_2296_sv2v_reg;
  assign mem[2295] = mem_2295_sv2v_reg;
  assign mem[2294] = mem_2294_sv2v_reg;
  assign mem[2293] = mem_2293_sv2v_reg;
  assign mem[2292] = mem_2292_sv2v_reg;
  assign mem[2291] = mem_2291_sv2v_reg;
  assign mem[2290] = mem_2290_sv2v_reg;
  assign mem[2289] = mem_2289_sv2v_reg;
  assign mem[2288] = mem_2288_sv2v_reg;
  assign mem[2287] = mem_2287_sv2v_reg;
  assign mem[2286] = mem_2286_sv2v_reg;
  assign mem[2285] = mem_2285_sv2v_reg;
  assign mem[2284] = mem_2284_sv2v_reg;
  assign mem[2283] = mem_2283_sv2v_reg;
  assign mem[2282] = mem_2282_sv2v_reg;
  assign mem[2281] = mem_2281_sv2v_reg;
  assign mem[2280] = mem_2280_sv2v_reg;
  assign mem[2279] = mem_2279_sv2v_reg;
  assign mem[2278] = mem_2278_sv2v_reg;
  assign mem[2277] = mem_2277_sv2v_reg;
  assign mem[2276] = mem_2276_sv2v_reg;
  assign mem[2275] = mem_2275_sv2v_reg;
  assign mem[2274] = mem_2274_sv2v_reg;
  assign mem[2273] = mem_2273_sv2v_reg;
  assign mem[2272] = mem_2272_sv2v_reg;
  assign mem[2271] = mem_2271_sv2v_reg;
  assign mem[2270] = mem_2270_sv2v_reg;
  assign mem[2269] = mem_2269_sv2v_reg;
  assign mem[2268] = mem_2268_sv2v_reg;
  assign mem[2267] = mem_2267_sv2v_reg;
  assign mem[2266] = mem_2266_sv2v_reg;
  assign mem[2265] = mem_2265_sv2v_reg;
  assign mem[2264] = mem_2264_sv2v_reg;
  assign mem[2263] = mem_2263_sv2v_reg;
  assign mem[2262] = mem_2262_sv2v_reg;
  assign mem[2261] = mem_2261_sv2v_reg;
  assign mem[2260] = mem_2260_sv2v_reg;
  assign mem[2259] = mem_2259_sv2v_reg;
  assign mem[2258] = mem_2258_sv2v_reg;
  assign mem[2257] = mem_2257_sv2v_reg;
  assign mem[2256] = mem_2256_sv2v_reg;
  assign mem[2255] = mem_2255_sv2v_reg;
  assign mem[2254] = mem_2254_sv2v_reg;
  assign mem[2253] = mem_2253_sv2v_reg;
  assign mem[2252] = mem_2252_sv2v_reg;
  assign mem[2251] = mem_2251_sv2v_reg;
  assign mem[2250] = mem_2250_sv2v_reg;
  assign mem[2249] = mem_2249_sv2v_reg;
  assign mem[2248] = mem_2248_sv2v_reg;
  assign mem[2247] = mem_2247_sv2v_reg;
  assign mem[2246] = mem_2246_sv2v_reg;
  assign mem[2245] = mem_2245_sv2v_reg;
  assign mem[2244] = mem_2244_sv2v_reg;
  assign mem[2243] = mem_2243_sv2v_reg;
  assign mem[2242] = mem_2242_sv2v_reg;
  assign mem[2241] = mem_2241_sv2v_reg;
  assign mem[2240] = mem_2240_sv2v_reg;
  assign mem[2239] = mem_2239_sv2v_reg;
  assign mem[2238] = mem_2238_sv2v_reg;
  assign mem[2237] = mem_2237_sv2v_reg;
  assign mem[2236] = mem_2236_sv2v_reg;
  assign mem[2235] = mem_2235_sv2v_reg;
  assign mem[2234] = mem_2234_sv2v_reg;
  assign mem[2233] = mem_2233_sv2v_reg;
  assign mem[2232] = mem_2232_sv2v_reg;
  assign mem[2231] = mem_2231_sv2v_reg;
  assign mem[2230] = mem_2230_sv2v_reg;
  assign mem[2229] = mem_2229_sv2v_reg;
  assign mem[2228] = mem_2228_sv2v_reg;
  assign mem[2227] = mem_2227_sv2v_reg;
  assign mem[2226] = mem_2226_sv2v_reg;
  assign mem[2225] = mem_2225_sv2v_reg;
  assign mem[2224] = mem_2224_sv2v_reg;
  assign mem[2223] = mem_2223_sv2v_reg;
  assign mem[2222] = mem_2222_sv2v_reg;
  assign mem[2221] = mem_2221_sv2v_reg;
  assign mem[2220] = mem_2220_sv2v_reg;
  assign mem[2219] = mem_2219_sv2v_reg;
  assign mem[2218] = mem_2218_sv2v_reg;
  assign mem[2217] = mem_2217_sv2v_reg;
  assign mem[2216] = mem_2216_sv2v_reg;
  assign mem[2215] = mem_2215_sv2v_reg;
  assign mem[2214] = mem_2214_sv2v_reg;
  assign mem[2213] = mem_2213_sv2v_reg;
  assign mem[2212] = mem_2212_sv2v_reg;
  assign mem[2211] = mem_2211_sv2v_reg;
  assign mem[2210] = mem_2210_sv2v_reg;
  assign mem[2209] = mem_2209_sv2v_reg;
  assign mem[2208] = mem_2208_sv2v_reg;
  assign mem[2207] = mem_2207_sv2v_reg;
  assign mem[2206] = mem_2206_sv2v_reg;
  assign mem[2205] = mem_2205_sv2v_reg;
  assign mem[2204] = mem_2204_sv2v_reg;
  assign mem[2203] = mem_2203_sv2v_reg;
  assign mem[2202] = mem_2202_sv2v_reg;
  assign mem[2201] = mem_2201_sv2v_reg;
  assign mem[2200] = mem_2200_sv2v_reg;
  assign mem[2199] = mem_2199_sv2v_reg;
  assign mem[2198] = mem_2198_sv2v_reg;
  assign mem[2197] = mem_2197_sv2v_reg;
  assign mem[2196] = mem_2196_sv2v_reg;
  assign mem[2195] = mem_2195_sv2v_reg;
  assign mem[2194] = mem_2194_sv2v_reg;
  assign mem[2193] = mem_2193_sv2v_reg;
  assign mem[2192] = mem_2192_sv2v_reg;
  assign mem[2191] = mem_2191_sv2v_reg;
  assign mem[2190] = mem_2190_sv2v_reg;
  assign mem[2189] = mem_2189_sv2v_reg;
  assign mem[2188] = mem_2188_sv2v_reg;
  assign mem[2187] = mem_2187_sv2v_reg;
  assign mem[2186] = mem_2186_sv2v_reg;
  assign mem[2185] = mem_2185_sv2v_reg;
  assign mem[2184] = mem_2184_sv2v_reg;
  assign mem[2183] = mem_2183_sv2v_reg;
  assign mem[2182] = mem_2182_sv2v_reg;
  assign mem[2181] = mem_2181_sv2v_reg;
  assign mem[2180] = mem_2180_sv2v_reg;
  assign mem[2179] = mem_2179_sv2v_reg;
  assign mem[2178] = mem_2178_sv2v_reg;
  assign mem[2177] = mem_2177_sv2v_reg;
  assign mem[2176] = mem_2176_sv2v_reg;
  assign mem[2175] = mem_2175_sv2v_reg;
  assign mem[2174] = mem_2174_sv2v_reg;
  assign mem[2173] = mem_2173_sv2v_reg;
  assign mem[2172] = mem_2172_sv2v_reg;
  assign mem[2171] = mem_2171_sv2v_reg;
  assign mem[2170] = mem_2170_sv2v_reg;
  assign mem[2169] = mem_2169_sv2v_reg;
  assign mem[2168] = mem_2168_sv2v_reg;
  assign mem[2167] = mem_2167_sv2v_reg;
  assign mem[2166] = mem_2166_sv2v_reg;
  assign mem[2165] = mem_2165_sv2v_reg;
  assign mem[2164] = mem_2164_sv2v_reg;
  assign mem[2163] = mem_2163_sv2v_reg;
  assign mem[2162] = mem_2162_sv2v_reg;
  assign mem[2161] = mem_2161_sv2v_reg;
  assign mem[2160] = mem_2160_sv2v_reg;
  assign mem[2159] = mem_2159_sv2v_reg;
  assign mem[2158] = mem_2158_sv2v_reg;
  assign mem[2157] = mem_2157_sv2v_reg;
  assign mem[2156] = mem_2156_sv2v_reg;
  assign mem[2155] = mem_2155_sv2v_reg;
  assign mem[2154] = mem_2154_sv2v_reg;
  assign mem[2153] = mem_2153_sv2v_reg;
  assign mem[2152] = mem_2152_sv2v_reg;
  assign mem[2151] = mem_2151_sv2v_reg;
  assign mem[2150] = mem_2150_sv2v_reg;
  assign mem[2149] = mem_2149_sv2v_reg;
  assign mem[2148] = mem_2148_sv2v_reg;
  assign mem[2147] = mem_2147_sv2v_reg;
  assign mem[2146] = mem_2146_sv2v_reg;
  assign mem[2145] = mem_2145_sv2v_reg;
  assign mem[2144] = mem_2144_sv2v_reg;
  assign mem[2143] = mem_2143_sv2v_reg;
  assign mem[2142] = mem_2142_sv2v_reg;
  assign mem[2141] = mem_2141_sv2v_reg;
  assign mem[2140] = mem_2140_sv2v_reg;
  assign mem[2139] = mem_2139_sv2v_reg;
  assign mem[2138] = mem_2138_sv2v_reg;
  assign mem[2137] = mem_2137_sv2v_reg;
  assign mem[2136] = mem_2136_sv2v_reg;
  assign mem[2135] = mem_2135_sv2v_reg;
  assign mem[2134] = mem_2134_sv2v_reg;
  assign mem[2133] = mem_2133_sv2v_reg;
  assign mem[2132] = mem_2132_sv2v_reg;
  assign mem[2131] = mem_2131_sv2v_reg;
  assign mem[2130] = mem_2130_sv2v_reg;
  assign mem[2129] = mem_2129_sv2v_reg;
  assign mem[2128] = mem_2128_sv2v_reg;
  assign mem[2127] = mem_2127_sv2v_reg;
  assign mem[2126] = mem_2126_sv2v_reg;
  assign mem[2125] = mem_2125_sv2v_reg;
  assign mem[2124] = mem_2124_sv2v_reg;
  assign mem[2123] = mem_2123_sv2v_reg;
  assign mem[2122] = mem_2122_sv2v_reg;
  assign mem[2121] = mem_2121_sv2v_reg;
  assign mem[2120] = mem_2120_sv2v_reg;
  assign mem[2119] = mem_2119_sv2v_reg;
  assign mem[2118] = mem_2118_sv2v_reg;
  assign mem[2117] = mem_2117_sv2v_reg;
  assign mem[2116] = mem_2116_sv2v_reg;
  assign mem[2115] = mem_2115_sv2v_reg;
  assign mem[2114] = mem_2114_sv2v_reg;
  assign mem[2113] = mem_2113_sv2v_reg;
  assign mem[2112] = mem_2112_sv2v_reg;
  assign mem[2111] = mem_2111_sv2v_reg;
  assign mem[2110] = mem_2110_sv2v_reg;
  assign mem[2109] = mem_2109_sv2v_reg;
  assign mem[2108] = mem_2108_sv2v_reg;
  assign mem[2107] = mem_2107_sv2v_reg;
  assign mem[2106] = mem_2106_sv2v_reg;
  assign mem[2105] = mem_2105_sv2v_reg;
  assign mem[2104] = mem_2104_sv2v_reg;
  assign mem[2103] = mem_2103_sv2v_reg;
  assign mem[2102] = mem_2102_sv2v_reg;
  assign mem[2101] = mem_2101_sv2v_reg;
  assign mem[2100] = mem_2100_sv2v_reg;
  assign mem[2099] = mem_2099_sv2v_reg;
  assign mem[2098] = mem_2098_sv2v_reg;
  assign mem[2097] = mem_2097_sv2v_reg;
  assign mem[2096] = mem_2096_sv2v_reg;
  assign mem[2095] = mem_2095_sv2v_reg;
  assign mem[2094] = mem_2094_sv2v_reg;
  assign mem[2093] = mem_2093_sv2v_reg;
  assign mem[2092] = mem_2092_sv2v_reg;
  assign mem[2091] = mem_2091_sv2v_reg;
  assign mem[2090] = mem_2090_sv2v_reg;
  assign mem[2089] = mem_2089_sv2v_reg;
  assign mem[2088] = mem_2088_sv2v_reg;
  assign mem[2087] = mem_2087_sv2v_reg;
  assign mem[2086] = mem_2086_sv2v_reg;
  assign mem[2085] = mem_2085_sv2v_reg;
  assign mem[2084] = mem_2084_sv2v_reg;
  assign mem[2083] = mem_2083_sv2v_reg;
  assign mem[2082] = mem_2082_sv2v_reg;
  assign mem[2081] = mem_2081_sv2v_reg;
  assign mem[2080] = mem_2080_sv2v_reg;
  assign mem[2079] = mem_2079_sv2v_reg;
  assign mem[2078] = mem_2078_sv2v_reg;
  assign mem[2077] = mem_2077_sv2v_reg;
  assign mem[2076] = mem_2076_sv2v_reg;
  assign mem[2075] = mem_2075_sv2v_reg;
  assign mem[2074] = mem_2074_sv2v_reg;
  assign mem[2073] = mem_2073_sv2v_reg;
  assign mem[2072] = mem_2072_sv2v_reg;
  assign mem[2071] = mem_2071_sv2v_reg;
  assign mem[2070] = mem_2070_sv2v_reg;
  assign mem[2069] = mem_2069_sv2v_reg;
  assign mem[2068] = mem_2068_sv2v_reg;
  assign mem[2067] = mem_2067_sv2v_reg;
  assign mem[2066] = mem_2066_sv2v_reg;
  assign mem[2065] = mem_2065_sv2v_reg;
  assign mem[2064] = mem_2064_sv2v_reg;
  assign mem[2063] = mem_2063_sv2v_reg;
  assign mem[2062] = mem_2062_sv2v_reg;
  assign mem[2061] = mem_2061_sv2v_reg;
  assign mem[2060] = mem_2060_sv2v_reg;
  assign mem[2059] = mem_2059_sv2v_reg;
  assign mem[2058] = mem_2058_sv2v_reg;
  assign mem[2057] = mem_2057_sv2v_reg;
  assign mem[2056] = mem_2056_sv2v_reg;
  assign mem[2055] = mem_2055_sv2v_reg;
  assign mem[2054] = mem_2054_sv2v_reg;
  assign mem[2053] = mem_2053_sv2v_reg;
  assign mem[2052] = mem_2052_sv2v_reg;
  assign mem[2051] = mem_2051_sv2v_reg;
  assign mem[2050] = mem_2050_sv2v_reg;
  assign mem[2049] = mem_2049_sv2v_reg;
  assign mem[2048] = mem_2048_sv2v_reg;
  assign mem[2047] = mem_2047_sv2v_reg;
  assign mem[2046] = mem_2046_sv2v_reg;
  assign mem[2045] = mem_2045_sv2v_reg;
  assign mem[2044] = mem_2044_sv2v_reg;
  assign mem[2043] = mem_2043_sv2v_reg;
  assign mem[2042] = mem_2042_sv2v_reg;
  assign mem[2041] = mem_2041_sv2v_reg;
  assign mem[2040] = mem_2040_sv2v_reg;
  assign mem[2039] = mem_2039_sv2v_reg;
  assign mem[2038] = mem_2038_sv2v_reg;
  assign mem[2037] = mem_2037_sv2v_reg;
  assign mem[2036] = mem_2036_sv2v_reg;
  assign mem[2035] = mem_2035_sv2v_reg;
  assign mem[2034] = mem_2034_sv2v_reg;
  assign mem[2033] = mem_2033_sv2v_reg;
  assign mem[2032] = mem_2032_sv2v_reg;
  assign mem[2031] = mem_2031_sv2v_reg;
  assign mem[2030] = mem_2030_sv2v_reg;
  assign mem[2029] = mem_2029_sv2v_reg;
  assign mem[2028] = mem_2028_sv2v_reg;
  assign mem[2027] = mem_2027_sv2v_reg;
  assign mem[2026] = mem_2026_sv2v_reg;
  assign mem[2025] = mem_2025_sv2v_reg;
  assign mem[2024] = mem_2024_sv2v_reg;
  assign mem[2023] = mem_2023_sv2v_reg;
  assign mem[2022] = mem_2022_sv2v_reg;
  assign mem[2021] = mem_2021_sv2v_reg;
  assign mem[2020] = mem_2020_sv2v_reg;
  assign mem[2019] = mem_2019_sv2v_reg;
  assign mem[2018] = mem_2018_sv2v_reg;
  assign mem[2017] = mem_2017_sv2v_reg;
  assign mem[2016] = mem_2016_sv2v_reg;
  assign mem[2015] = mem_2015_sv2v_reg;
  assign mem[2014] = mem_2014_sv2v_reg;
  assign mem[2013] = mem_2013_sv2v_reg;
  assign mem[2012] = mem_2012_sv2v_reg;
  assign mem[2011] = mem_2011_sv2v_reg;
  assign mem[2010] = mem_2010_sv2v_reg;
  assign mem[2009] = mem_2009_sv2v_reg;
  assign mem[2008] = mem_2008_sv2v_reg;
  assign mem[2007] = mem_2007_sv2v_reg;
  assign mem[2006] = mem_2006_sv2v_reg;
  assign mem[2005] = mem_2005_sv2v_reg;
  assign mem[2004] = mem_2004_sv2v_reg;
  assign mem[2003] = mem_2003_sv2v_reg;
  assign mem[2002] = mem_2002_sv2v_reg;
  assign mem[2001] = mem_2001_sv2v_reg;
  assign mem[2000] = mem_2000_sv2v_reg;
  assign mem[1999] = mem_1999_sv2v_reg;
  assign mem[1998] = mem_1998_sv2v_reg;
  assign mem[1997] = mem_1997_sv2v_reg;
  assign mem[1996] = mem_1996_sv2v_reg;
  assign mem[1995] = mem_1995_sv2v_reg;
  assign mem[1994] = mem_1994_sv2v_reg;
  assign mem[1993] = mem_1993_sv2v_reg;
  assign mem[1992] = mem_1992_sv2v_reg;
  assign mem[1991] = mem_1991_sv2v_reg;
  assign mem[1990] = mem_1990_sv2v_reg;
  assign mem[1989] = mem_1989_sv2v_reg;
  assign mem[1988] = mem_1988_sv2v_reg;
  assign mem[1987] = mem_1987_sv2v_reg;
  assign mem[1986] = mem_1986_sv2v_reg;
  assign mem[1985] = mem_1985_sv2v_reg;
  assign mem[1984] = mem_1984_sv2v_reg;
  assign mem[1983] = mem_1983_sv2v_reg;
  assign mem[1982] = mem_1982_sv2v_reg;
  assign mem[1981] = mem_1981_sv2v_reg;
  assign mem[1980] = mem_1980_sv2v_reg;
  assign mem[1979] = mem_1979_sv2v_reg;
  assign mem[1978] = mem_1978_sv2v_reg;
  assign mem[1977] = mem_1977_sv2v_reg;
  assign mem[1976] = mem_1976_sv2v_reg;
  assign mem[1975] = mem_1975_sv2v_reg;
  assign mem[1974] = mem_1974_sv2v_reg;
  assign mem[1973] = mem_1973_sv2v_reg;
  assign mem[1972] = mem_1972_sv2v_reg;
  assign mem[1971] = mem_1971_sv2v_reg;
  assign mem[1970] = mem_1970_sv2v_reg;
  assign mem[1969] = mem_1969_sv2v_reg;
  assign mem[1968] = mem_1968_sv2v_reg;
  assign mem[1967] = mem_1967_sv2v_reg;
  assign mem[1966] = mem_1966_sv2v_reg;
  assign mem[1965] = mem_1965_sv2v_reg;
  assign mem[1964] = mem_1964_sv2v_reg;
  assign mem[1963] = mem_1963_sv2v_reg;
  assign mem[1962] = mem_1962_sv2v_reg;
  assign mem[1961] = mem_1961_sv2v_reg;
  assign mem[1960] = mem_1960_sv2v_reg;
  assign mem[1959] = mem_1959_sv2v_reg;
  assign mem[1958] = mem_1958_sv2v_reg;
  assign mem[1957] = mem_1957_sv2v_reg;
  assign mem[1956] = mem_1956_sv2v_reg;
  assign mem[1955] = mem_1955_sv2v_reg;
  assign mem[1954] = mem_1954_sv2v_reg;
  assign mem[1953] = mem_1953_sv2v_reg;
  assign mem[1952] = mem_1952_sv2v_reg;
  assign mem[1951] = mem_1951_sv2v_reg;
  assign mem[1950] = mem_1950_sv2v_reg;
  assign mem[1949] = mem_1949_sv2v_reg;
  assign mem[1948] = mem_1948_sv2v_reg;
  assign mem[1947] = mem_1947_sv2v_reg;
  assign mem[1946] = mem_1946_sv2v_reg;
  assign mem[1945] = mem_1945_sv2v_reg;
  assign mem[1944] = mem_1944_sv2v_reg;
  assign mem[1943] = mem_1943_sv2v_reg;
  assign mem[1942] = mem_1942_sv2v_reg;
  assign mem[1941] = mem_1941_sv2v_reg;
  assign mem[1940] = mem_1940_sv2v_reg;
  assign mem[1939] = mem_1939_sv2v_reg;
  assign mem[1938] = mem_1938_sv2v_reg;
  assign mem[1937] = mem_1937_sv2v_reg;
  assign mem[1936] = mem_1936_sv2v_reg;
  assign mem[1935] = mem_1935_sv2v_reg;
  assign mem[1934] = mem_1934_sv2v_reg;
  assign mem[1933] = mem_1933_sv2v_reg;
  assign mem[1932] = mem_1932_sv2v_reg;
  assign mem[1931] = mem_1931_sv2v_reg;
  assign mem[1930] = mem_1930_sv2v_reg;
  assign mem[1929] = mem_1929_sv2v_reg;
  assign mem[1928] = mem_1928_sv2v_reg;
  assign mem[1927] = mem_1927_sv2v_reg;
  assign mem[1926] = mem_1926_sv2v_reg;
  assign mem[1925] = mem_1925_sv2v_reg;
  assign mem[1924] = mem_1924_sv2v_reg;
  assign mem[1923] = mem_1923_sv2v_reg;
  assign mem[1922] = mem_1922_sv2v_reg;
  assign mem[1921] = mem_1921_sv2v_reg;
  assign mem[1920] = mem_1920_sv2v_reg;
  assign mem[1919] = mem_1919_sv2v_reg;
  assign mem[1918] = mem_1918_sv2v_reg;
  assign mem[1917] = mem_1917_sv2v_reg;
  assign mem[1916] = mem_1916_sv2v_reg;
  assign mem[1915] = mem_1915_sv2v_reg;
  assign mem[1914] = mem_1914_sv2v_reg;
  assign mem[1913] = mem_1913_sv2v_reg;
  assign mem[1912] = mem_1912_sv2v_reg;
  assign mem[1911] = mem_1911_sv2v_reg;
  assign mem[1910] = mem_1910_sv2v_reg;
  assign mem[1909] = mem_1909_sv2v_reg;
  assign mem[1908] = mem_1908_sv2v_reg;
  assign mem[1907] = mem_1907_sv2v_reg;
  assign mem[1906] = mem_1906_sv2v_reg;
  assign mem[1905] = mem_1905_sv2v_reg;
  assign mem[1904] = mem_1904_sv2v_reg;
  assign mem[1903] = mem_1903_sv2v_reg;
  assign mem[1902] = mem_1902_sv2v_reg;
  assign mem[1901] = mem_1901_sv2v_reg;
  assign mem[1900] = mem_1900_sv2v_reg;
  assign mem[1899] = mem_1899_sv2v_reg;
  assign mem[1898] = mem_1898_sv2v_reg;
  assign mem[1897] = mem_1897_sv2v_reg;
  assign mem[1896] = mem_1896_sv2v_reg;
  assign mem[1895] = mem_1895_sv2v_reg;
  assign mem[1894] = mem_1894_sv2v_reg;
  assign mem[1893] = mem_1893_sv2v_reg;
  assign mem[1892] = mem_1892_sv2v_reg;
  assign mem[1891] = mem_1891_sv2v_reg;
  assign mem[1890] = mem_1890_sv2v_reg;
  assign mem[1889] = mem_1889_sv2v_reg;
  assign mem[1888] = mem_1888_sv2v_reg;
  assign mem[1887] = mem_1887_sv2v_reg;
  assign mem[1886] = mem_1886_sv2v_reg;
  assign mem[1885] = mem_1885_sv2v_reg;
  assign mem[1884] = mem_1884_sv2v_reg;
  assign mem[1883] = mem_1883_sv2v_reg;
  assign mem[1882] = mem_1882_sv2v_reg;
  assign mem[1881] = mem_1881_sv2v_reg;
  assign mem[1880] = mem_1880_sv2v_reg;
  assign mem[1879] = mem_1879_sv2v_reg;
  assign mem[1878] = mem_1878_sv2v_reg;
  assign mem[1877] = mem_1877_sv2v_reg;
  assign mem[1876] = mem_1876_sv2v_reg;
  assign mem[1875] = mem_1875_sv2v_reg;
  assign mem[1874] = mem_1874_sv2v_reg;
  assign mem[1873] = mem_1873_sv2v_reg;
  assign mem[1872] = mem_1872_sv2v_reg;
  assign mem[1871] = mem_1871_sv2v_reg;
  assign mem[1870] = mem_1870_sv2v_reg;
  assign mem[1869] = mem_1869_sv2v_reg;
  assign mem[1868] = mem_1868_sv2v_reg;
  assign mem[1867] = mem_1867_sv2v_reg;
  assign mem[1866] = mem_1866_sv2v_reg;
  assign mem[1865] = mem_1865_sv2v_reg;
  assign mem[1864] = mem_1864_sv2v_reg;
  assign mem[1863] = mem_1863_sv2v_reg;
  assign mem[1862] = mem_1862_sv2v_reg;
  assign mem[1861] = mem_1861_sv2v_reg;
  assign mem[1860] = mem_1860_sv2v_reg;
  assign mem[1859] = mem_1859_sv2v_reg;
  assign mem[1858] = mem_1858_sv2v_reg;
  assign mem[1857] = mem_1857_sv2v_reg;
  assign mem[1856] = mem_1856_sv2v_reg;
  assign mem[1855] = mem_1855_sv2v_reg;
  assign mem[1854] = mem_1854_sv2v_reg;
  assign mem[1853] = mem_1853_sv2v_reg;
  assign mem[1852] = mem_1852_sv2v_reg;
  assign mem[1851] = mem_1851_sv2v_reg;
  assign mem[1850] = mem_1850_sv2v_reg;
  assign mem[1849] = mem_1849_sv2v_reg;
  assign mem[1848] = mem_1848_sv2v_reg;
  assign mem[1847] = mem_1847_sv2v_reg;
  assign mem[1846] = mem_1846_sv2v_reg;
  assign mem[1845] = mem_1845_sv2v_reg;
  assign mem[1844] = mem_1844_sv2v_reg;
  assign mem[1843] = mem_1843_sv2v_reg;
  assign mem[1842] = mem_1842_sv2v_reg;
  assign mem[1841] = mem_1841_sv2v_reg;
  assign mem[1840] = mem_1840_sv2v_reg;
  assign mem[1839] = mem_1839_sv2v_reg;
  assign mem[1838] = mem_1838_sv2v_reg;
  assign mem[1837] = mem_1837_sv2v_reg;
  assign mem[1836] = mem_1836_sv2v_reg;
  assign mem[1835] = mem_1835_sv2v_reg;
  assign mem[1834] = mem_1834_sv2v_reg;
  assign mem[1833] = mem_1833_sv2v_reg;
  assign mem[1832] = mem_1832_sv2v_reg;
  assign mem[1831] = mem_1831_sv2v_reg;
  assign mem[1830] = mem_1830_sv2v_reg;
  assign mem[1829] = mem_1829_sv2v_reg;
  assign mem[1828] = mem_1828_sv2v_reg;
  assign mem[1827] = mem_1827_sv2v_reg;
  assign mem[1826] = mem_1826_sv2v_reg;
  assign mem[1825] = mem_1825_sv2v_reg;
  assign mem[1824] = mem_1824_sv2v_reg;
  assign mem[1823] = mem_1823_sv2v_reg;
  assign mem[1822] = mem_1822_sv2v_reg;
  assign mem[1821] = mem_1821_sv2v_reg;
  assign mem[1820] = mem_1820_sv2v_reg;
  assign mem[1819] = mem_1819_sv2v_reg;
  assign mem[1818] = mem_1818_sv2v_reg;
  assign mem[1817] = mem_1817_sv2v_reg;
  assign mem[1816] = mem_1816_sv2v_reg;
  assign mem[1815] = mem_1815_sv2v_reg;
  assign mem[1814] = mem_1814_sv2v_reg;
  assign mem[1813] = mem_1813_sv2v_reg;
  assign mem[1812] = mem_1812_sv2v_reg;
  assign mem[1811] = mem_1811_sv2v_reg;
  assign mem[1810] = mem_1810_sv2v_reg;
  assign mem[1809] = mem_1809_sv2v_reg;
  assign mem[1808] = mem_1808_sv2v_reg;
  assign mem[1807] = mem_1807_sv2v_reg;
  assign mem[1806] = mem_1806_sv2v_reg;
  assign mem[1805] = mem_1805_sv2v_reg;
  assign mem[1804] = mem_1804_sv2v_reg;
  assign mem[1803] = mem_1803_sv2v_reg;
  assign mem[1802] = mem_1802_sv2v_reg;
  assign mem[1801] = mem_1801_sv2v_reg;
  assign mem[1800] = mem_1800_sv2v_reg;
  assign mem[1799] = mem_1799_sv2v_reg;
  assign mem[1798] = mem_1798_sv2v_reg;
  assign mem[1797] = mem_1797_sv2v_reg;
  assign mem[1796] = mem_1796_sv2v_reg;
  assign mem[1795] = mem_1795_sv2v_reg;
  assign mem[1794] = mem_1794_sv2v_reg;
  assign mem[1793] = mem_1793_sv2v_reg;
  assign mem[1792] = mem_1792_sv2v_reg;
  assign mem[1791] = mem_1791_sv2v_reg;
  assign mem[1790] = mem_1790_sv2v_reg;
  assign mem[1789] = mem_1789_sv2v_reg;
  assign mem[1788] = mem_1788_sv2v_reg;
  assign mem[1787] = mem_1787_sv2v_reg;
  assign mem[1786] = mem_1786_sv2v_reg;
  assign mem[1785] = mem_1785_sv2v_reg;
  assign mem[1784] = mem_1784_sv2v_reg;
  assign mem[1783] = mem_1783_sv2v_reg;
  assign mem[1782] = mem_1782_sv2v_reg;
  assign mem[1781] = mem_1781_sv2v_reg;
  assign mem[1780] = mem_1780_sv2v_reg;
  assign mem[1779] = mem_1779_sv2v_reg;
  assign mem[1778] = mem_1778_sv2v_reg;
  assign mem[1777] = mem_1777_sv2v_reg;
  assign mem[1776] = mem_1776_sv2v_reg;
  assign mem[1775] = mem_1775_sv2v_reg;
  assign mem[1774] = mem_1774_sv2v_reg;
  assign mem[1773] = mem_1773_sv2v_reg;
  assign mem[1772] = mem_1772_sv2v_reg;
  assign mem[1771] = mem_1771_sv2v_reg;
  assign mem[1770] = mem_1770_sv2v_reg;
  assign mem[1769] = mem_1769_sv2v_reg;
  assign mem[1768] = mem_1768_sv2v_reg;
  assign mem[1767] = mem_1767_sv2v_reg;
  assign mem[1766] = mem_1766_sv2v_reg;
  assign mem[1765] = mem_1765_sv2v_reg;
  assign mem[1764] = mem_1764_sv2v_reg;
  assign mem[1763] = mem_1763_sv2v_reg;
  assign mem[1762] = mem_1762_sv2v_reg;
  assign mem[1761] = mem_1761_sv2v_reg;
  assign mem[1760] = mem_1760_sv2v_reg;
  assign mem[1759] = mem_1759_sv2v_reg;
  assign mem[1758] = mem_1758_sv2v_reg;
  assign mem[1757] = mem_1757_sv2v_reg;
  assign mem[1756] = mem_1756_sv2v_reg;
  assign mem[1755] = mem_1755_sv2v_reg;
  assign mem[1754] = mem_1754_sv2v_reg;
  assign mem[1753] = mem_1753_sv2v_reg;
  assign mem[1752] = mem_1752_sv2v_reg;
  assign mem[1751] = mem_1751_sv2v_reg;
  assign mem[1750] = mem_1750_sv2v_reg;
  assign mem[1749] = mem_1749_sv2v_reg;
  assign mem[1748] = mem_1748_sv2v_reg;
  assign mem[1747] = mem_1747_sv2v_reg;
  assign mem[1746] = mem_1746_sv2v_reg;
  assign mem[1745] = mem_1745_sv2v_reg;
  assign mem[1744] = mem_1744_sv2v_reg;
  assign mem[1743] = mem_1743_sv2v_reg;
  assign mem[1742] = mem_1742_sv2v_reg;
  assign mem[1741] = mem_1741_sv2v_reg;
  assign mem[1740] = mem_1740_sv2v_reg;
  assign mem[1739] = mem_1739_sv2v_reg;
  assign mem[1738] = mem_1738_sv2v_reg;
  assign mem[1737] = mem_1737_sv2v_reg;
  assign mem[1736] = mem_1736_sv2v_reg;
  assign mem[1735] = mem_1735_sv2v_reg;
  assign mem[1734] = mem_1734_sv2v_reg;
  assign mem[1733] = mem_1733_sv2v_reg;
  assign mem[1732] = mem_1732_sv2v_reg;
  assign mem[1731] = mem_1731_sv2v_reg;
  assign mem[1730] = mem_1730_sv2v_reg;
  assign mem[1729] = mem_1729_sv2v_reg;
  assign mem[1728] = mem_1728_sv2v_reg;
  assign mem[1727] = mem_1727_sv2v_reg;
  assign mem[1726] = mem_1726_sv2v_reg;
  assign mem[1725] = mem_1725_sv2v_reg;
  assign mem[1724] = mem_1724_sv2v_reg;
  assign mem[1723] = mem_1723_sv2v_reg;
  assign mem[1722] = mem_1722_sv2v_reg;
  assign mem[1721] = mem_1721_sv2v_reg;
  assign mem[1720] = mem_1720_sv2v_reg;
  assign mem[1719] = mem_1719_sv2v_reg;
  assign mem[1718] = mem_1718_sv2v_reg;
  assign mem[1717] = mem_1717_sv2v_reg;
  assign mem[1716] = mem_1716_sv2v_reg;
  assign mem[1715] = mem_1715_sv2v_reg;
  assign mem[1714] = mem_1714_sv2v_reg;
  assign mem[1713] = mem_1713_sv2v_reg;
  assign mem[1712] = mem_1712_sv2v_reg;
  assign mem[1711] = mem_1711_sv2v_reg;
  assign mem[1710] = mem_1710_sv2v_reg;
  assign mem[1709] = mem_1709_sv2v_reg;
  assign mem[1708] = mem_1708_sv2v_reg;
  assign mem[1707] = mem_1707_sv2v_reg;
  assign mem[1706] = mem_1706_sv2v_reg;
  assign mem[1705] = mem_1705_sv2v_reg;
  assign mem[1704] = mem_1704_sv2v_reg;
  assign mem[1703] = mem_1703_sv2v_reg;
  assign mem[1702] = mem_1702_sv2v_reg;
  assign mem[1701] = mem_1701_sv2v_reg;
  assign mem[1700] = mem_1700_sv2v_reg;
  assign mem[1699] = mem_1699_sv2v_reg;
  assign mem[1698] = mem_1698_sv2v_reg;
  assign mem[1697] = mem_1697_sv2v_reg;
  assign mem[1696] = mem_1696_sv2v_reg;
  assign mem[1695] = mem_1695_sv2v_reg;
  assign mem[1694] = mem_1694_sv2v_reg;
  assign mem[1693] = mem_1693_sv2v_reg;
  assign mem[1692] = mem_1692_sv2v_reg;
  assign mem[1691] = mem_1691_sv2v_reg;
  assign mem[1690] = mem_1690_sv2v_reg;
  assign mem[1689] = mem_1689_sv2v_reg;
  assign mem[1688] = mem_1688_sv2v_reg;
  assign mem[1687] = mem_1687_sv2v_reg;
  assign mem[1686] = mem_1686_sv2v_reg;
  assign mem[1685] = mem_1685_sv2v_reg;
  assign mem[1684] = mem_1684_sv2v_reg;
  assign mem[1683] = mem_1683_sv2v_reg;
  assign mem[1682] = mem_1682_sv2v_reg;
  assign mem[1681] = mem_1681_sv2v_reg;
  assign mem[1680] = mem_1680_sv2v_reg;
  assign mem[1679] = mem_1679_sv2v_reg;
  assign mem[1678] = mem_1678_sv2v_reg;
  assign mem[1677] = mem_1677_sv2v_reg;
  assign mem[1676] = mem_1676_sv2v_reg;
  assign mem[1675] = mem_1675_sv2v_reg;
  assign mem[1674] = mem_1674_sv2v_reg;
  assign mem[1673] = mem_1673_sv2v_reg;
  assign mem[1672] = mem_1672_sv2v_reg;
  assign mem[1671] = mem_1671_sv2v_reg;
  assign mem[1670] = mem_1670_sv2v_reg;
  assign mem[1669] = mem_1669_sv2v_reg;
  assign mem[1668] = mem_1668_sv2v_reg;
  assign mem[1667] = mem_1667_sv2v_reg;
  assign mem[1666] = mem_1666_sv2v_reg;
  assign mem[1665] = mem_1665_sv2v_reg;
  assign mem[1664] = mem_1664_sv2v_reg;
  assign mem[1663] = mem_1663_sv2v_reg;
  assign mem[1662] = mem_1662_sv2v_reg;
  assign mem[1661] = mem_1661_sv2v_reg;
  assign mem[1660] = mem_1660_sv2v_reg;
  assign mem[1659] = mem_1659_sv2v_reg;
  assign mem[1658] = mem_1658_sv2v_reg;
  assign mem[1657] = mem_1657_sv2v_reg;
  assign mem[1656] = mem_1656_sv2v_reg;
  assign mem[1655] = mem_1655_sv2v_reg;
  assign mem[1654] = mem_1654_sv2v_reg;
  assign mem[1653] = mem_1653_sv2v_reg;
  assign mem[1652] = mem_1652_sv2v_reg;
  assign mem[1651] = mem_1651_sv2v_reg;
  assign mem[1650] = mem_1650_sv2v_reg;
  assign mem[1649] = mem_1649_sv2v_reg;
  assign mem[1648] = mem_1648_sv2v_reg;
  assign mem[1647] = mem_1647_sv2v_reg;
  assign mem[1646] = mem_1646_sv2v_reg;
  assign mem[1645] = mem_1645_sv2v_reg;
  assign mem[1644] = mem_1644_sv2v_reg;
  assign mem[1643] = mem_1643_sv2v_reg;
  assign mem[1642] = mem_1642_sv2v_reg;
  assign mem[1641] = mem_1641_sv2v_reg;
  assign mem[1640] = mem_1640_sv2v_reg;
  assign mem[1639] = mem_1639_sv2v_reg;
  assign mem[1638] = mem_1638_sv2v_reg;
  assign mem[1637] = mem_1637_sv2v_reg;
  assign mem[1636] = mem_1636_sv2v_reg;
  assign mem[1635] = mem_1635_sv2v_reg;
  assign mem[1634] = mem_1634_sv2v_reg;
  assign mem[1633] = mem_1633_sv2v_reg;
  assign mem[1632] = mem_1632_sv2v_reg;
  assign mem[1631] = mem_1631_sv2v_reg;
  assign mem[1630] = mem_1630_sv2v_reg;
  assign mem[1629] = mem_1629_sv2v_reg;
  assign mem[1628] = mem_1628_sv2v_reg;
  assign mem[1627] = mem_1627_sv2v_reg;
  assign mem[1626] = mem_1626_sv2v_reg;
  assign mem[1625] = mem_1625_sv2v_reg;
  assign mem[1624] = mem_1624_sv2v_reg;
  assign mem[1623] = mem_1623_sv2v_reg;
  assign mem[1622] = mem_1622_sv2v_reg;
  assign mem[1621] = mem_1621_sv2v_reg;
  assign mem[1620] = mem_1620_sv2v_reg;
  assign mem[1619] = mem_1619_sv2v_reg;
  assign mem[1618] = mem_1618_sv2v_reg;
  assign mem[1617] = mem_1617_sv2v_reg;
  assign mem[1616] = mem_1616_sv2v_reg;
  assign mem[1615] = mem_1615_sv2v_reg;
  assign mem[1614] = mem_1614_sv2v_reg;
  assign mem[1613] = mem_1613_sv2v_reg;
  assign mem[1612] = mem_1612_sv2v_reg;
  assign mem[1611] = mem_1611_sv2v_reg;
  assign mem[1610] = mem_1610_sv2v_reg;
  assign mem[1609] = mem_1609_sv2v_reg;
  assign mem[1608] = mem_1608_sv2v_reg;
  assign mem[1607] = mem_1607_sv2v_reg;
  assign mem[1606] = mem_1606_sv2v_reg;
  assign mem[1605] = mem_1605_sv2v_reg;
  assign mem[1604] = mem_1604_sv2v_reg;
  assign mem[1603] = mem_1603_sv2v_reg;
  assign mem[1602] = mem_1602_sv2v_reg;
  assign mem[1601] = mem_1601_sv2v_reg;
  assign mem[1600] = mem_1600_sv2v_reg;
  assign mem[1599] = mem_1599_sv2v_reg;
  assign mem[1598] = mem_1598_sv2v_reg;
  assign mem[1597] = mem_1597_sv2v_reg;
  assign mem[1596] = mem_1596_sv2v_reg;
  assign mem[1595] = mem_1595_sv2v_reg;
  assign mem[1594] = mem_1594_sv2v_reg;
  assign mem[1593] = mem_1593_sv2v_reg;
  assign mem[1592] = mem_1592_sv2v_reg;
  assign mem[1591] = mem_1591_sv2v_reg;
  assign mem[1590] = mem_1590_sv2v_reg;
  assign mem[1589] = mem_1589_sv2v_reg;
  assign mem[1588] = mem_1588_sv2v_reg;
  assign mem[1587] = mem_1587_sv2v_reg;
  assign mem[1586] = mem_1586_sv2v_reg;
  assign mem[1585] = mem_1585_sv2v_reg;
  assign mem[1584] = mem_1584_sv2v_reg;
  assign mem[1583] = mem_1583_sv2v_reg;
  assign mem[1582] = mem_1582_sv2v_reg;
  assign mem[1581] = mem_1581_sv2v_reg;
  assign mem[1580] = mem_1580_sv2v_reg;
  assign mem[1579] = mem_1579_sv2v_reg;
  assign mem[1578] = mem_1578_sv2v_reg;
  assign mem[1577] = mem_1577_sv2v_reg;
  assign mem[1576] = mem_1576_sv2v_reg;
  assign mem[1575] = mem_1575_sv2v_reg;
  assign mem[1574] = mem_1574_sv2v_reg;
  assign mem[1573] = mem_1573_sv2v_reg;
  assign mem[1572] = mem_1572_sv2v_reg;
  assign mem[1571] = mem_1571_sv2v_reg;
  assign mem[1570] = mem_1570_sv2v_reg;
  assign mem[1569] = mem_1569_sv2v_reg;
  assign mem[1568] = mem_1568_sv2v_reg;
  assign mem[1567] = mem_1567_sv2v_reg;
  assign mem[1566] = mem_1566_sv2v_reg;
  assign mem[1565] = mem_1565_sv2v_reg;
  assign mem[1564] = mem_1564_sv2v_reg;
  assign mem[1563] = mem_1563_sv2v_reg;
  assign mem[1562] = mem_1562_sv2v_reg;
  assign mem[1561] = mem_1561_sv2v_reg;
  assign mem[1560] = mem_1560_sv2v_reg;
  assign mem[1559] = mem_1559_sv2v_reg;
  assign mem[1558] = mem_1558_sv2v_reg;
  assign mem[1557] = mem_1557_sv2v_reg;
  assign mem[1556] = mem_1556_sv2v_reg;
  assign mem[1555] = mem_1555_sv2v_reg;
  assign mem[1554] = mem_1554_sv2v_reg;
  assign mem[1553] = mem_1553_sv2v_reg;
  assign mem[1552] = mem_1552_sv2v_reg;
  assign mem[1551] = mem_1551_sv2v_reg;
  assign mem[1550] = mem_1550_sv2v_reg;
  assign mem[1549] = mem_1549_sv2v_reg;
  assign mem[1548] = mem_1548_sv2v_reg;
  assign mem[1547] = mem_1547_sv2v_reg;
  assign mem[1546] = mem_1546_sv2v_reg;
  assign mem[1545] = mem_1545_sv2v_reg;
  assign mem[1544] = mem_1544_sv2v_reg;
  assign mem[1543] = mem_1543_sv2v_reg;
  assign mem[1542] = mem_1542_sv2v_reg;
  assign mem[1541] = mem_1541_sv2v_reg;
  assign mem[1540] = mem_1540_sv2v_reg;
  assign mem[1539] = mem_1539_sv2v_reg;
  assign mem[1538] = mem_1538_sv2v_reg;
  assign mem[1537] = mem_1537_sv2v_reg;
  assign mem[1536] = mem_1536_sv2v_reg;
  assign mem[1535] = mem_1535_sv2v_reg;
  assign mem[1534] = mem_1534_sv2v_reg;
  assign mem[1533] = mem_1533_sv2v_reg;
  assign mem[1532] = mem_1532_sv2v_reg;
  assign mem[1531] = mem_1531_sv2v_reg;
  assign mem[1530] = mem_1530_sv2v_reg;
  assign mem[1529] = mem_1529_sv2v_reg;
  assign mem[1528] = mem_1528_sv2v_reg;
  assign mem[1527] = mem_1527_sv2v_reg;
  assign mem[1526] = mem_1526_sv2v_reg;
  assign mem[1525] = mem_1525_sv2v_reg;
  assign mem[1524] = mem_1524_sv2v_reg;
  assign mem[1523] = mem_1523_sv2v_reg;
  assign mem[1522] = mem_1522_sv2v_reg;
  assign mem[1521] = mem_1521_sv2v_reg;
  assign mem[1520] = mem_1520_sv2v_reg;
  assign mem[1519] = mem_1519_sv2v_reg;
  assign mem[1518] = mem_1518_sv2v_reg;
  assign mem[1517] = mem_1517_sv2v_reg;
  assign mem[1516] = mem_1516_sv2v_reg;
  assign mem[1515] = mem_1515_sv2v_reg;
  assign mem[1514] = mem_1514_sv2v_reg;
  assign mem[1513] = mem_1513_sv2v_reg;
  assign mem[1512] = mem_1512_sv2v_reg;
  assign mem[1511] = mem_1511_sv2v_reg;
  assign mem[1510] = mem_1510_sv2v_reg;
  assign mem[1509] = mem_1509_sv2v_reg;
  assign mem[1508] = mem_1508_sv2v_reg;
  assign mem[1507] = mem_1507_sv2v_reg;
  assign mem[1506] = mem_1506_sv2v_reg;
  assign mem[1505] = mem_1505_sv2v_reg;
  assign mem[1504] = mem_1504_sv2v_reg;
  assign mem[1503] = mem_1503_sv2v_reg;
  assign mem[1502] = mem_1502_sv2v_reg;
  assign mem[1501] = mem_1501_sv2v_reg;
  assign mem[1500] = mem_1500_sv2v_reg;
  assign mem[1499] = mem_1499_sv2v_reg;
  assign mem[1498] = mem_1498_sv2v_reg;
  assign mem[1497] = mem_1497_sv2v_reg;
  assign mem[1496] = mem_1496_sv2v_reg;
  assign mem[1495] = mem_1495_sv2v_reg;
  assign mem[1494] = mem_1494_sv2v_reg;
  assign mem[1493] = mem_1493_sv2v_reg;
  assign mem[1492] = mem_1492_sv2v_reg;
  assign mem[1491] = mem_1491_sv2v_reg;
  assign mem[1490] = mem_1490_sv2v_reg;
  assign mem[1489] = mem_1489_sv2v_reg;
  assign mem[1488] = mem_1488_sv2v_reg;
  assign mem[1487] = mem_1487_sv2v_reg;
  assign mem[1486] = mem_1486_sv2v_reg;
  assign mem[1485] = mem_1485_sv2v_reg;
  assign mem[1484] = mem_1484_sv2v_reg;
  assign mem[1483] = mem_1483_sv2v_reg;
  assign mem[1482] = mem_1482_sv2v_reg;
  assign mem[1481] = mem_1481_sv2v_reg;
  assign mem[1480] = mem_1480_sv2v_reg;
  assign mem[1479] = mem_1479_sv2v_reg;
  assign mem[1478] = mem_1478_sv2v_reg;
  assign mem[1477] = mem_1477_sv2v_reg;
  assign mem[1476] = mem_1476_sv2v_reg;
  assign mem[1475] = mem_1475_sv2v_reg;
  assign mem[1474] = mem_1474_sv2v_reg;
  assign mem[1473] = mem_1473_sv2v_reg;
  assign mem[1472] = mem_1472_sv2v_reg;
  assign mem[1471] = mem_1471_sv2v_reg;
  assign mem[1470] = mem_1470_sv2v_reg;
  assign mem[1469] = mem_1469_sv2v_reg;
  assign mem[1468] = mem_1468_sv2v_reg;
  assign mem[1467] = mem_1467_sv2v_reg;
  assign mem[1466] = mem_1466_sv2v_reg;
  assign mem[1465] = mem_1465_sv2v_reg;
  assign mem[1464] = mem_1464_sv2v_reg;
  assign mem[1463] = mem_1463_sv2v_reg;
  assign mem[1462] = mem_1462_sv2v_reg;
  assign mem[1461] = mem_1461_sv2v_reg;
  assign mem[1460] = mem_1460_sv2v_reg;
  assign mem[1459] = mem_1459_sv2v_reg;
  assign mem[1458] = mem_1458_sv2v_reg;
  assign mem[1457] = mem_1457_sv2v_reg;
  assign mem[1456] = mem_1456_sv2v_reg;
  assign mem[1455] = mem_1455_sv2v_reg;
  assign mem[1454] = mem_1454_sv2v_reg;
  assign mem[1453] = mem_1453_sv2v_reg;
  assign mem[1452] = mem_1452_sv2v_reg;
  assign mem[1451] = mem_1451_sv2v_reg;
  assign mem[1450] = mem_1450_sv2v_reg;
  assign mem[1449] = mem_1449_sv2v_reg;
  assign mem[1448] = mem_1448_sv2v_reg;
  assign mem[1447] = mem_1447_sv2v_reg;
  assign mem[1446] = mem_1446_sv2v_reg;
  assign mem[1445] = mem_1445_sv2v_reg;
  assign mem[1444] = mem_1444_sv2v_reg;
  assign mem[1443] = mem_1443_sv2v_reg;
  assign mem[1442] = mem_1442_sv2v_reg;
  assign mem[1441] = mem_1441_sv2v_reg;
  assign mem[1440] = mem_1440_sv2v_reg;
  assign mem[1439] = mem_1439_sv2v_reg;
  assign mem[1438] = mem_1438_sv2v_reg;
  assign mem[1437] = mem_1437_sv2v_reg;
  assign mem[1436] = mem_1436_sv2v_reg;
  assign mem[1435] = mem_1435_sv2v_reg;
  assign mem[1434] = mem_1434_sv2v_reg;
  assign mem[1433] = mem_1433_sv2v_reg;
  assign mem[1432] = mem_1432_sv2v_reg;
  assign mem[1431] = mem_1431_sv2v_reg;
  assign mem[1430] = mem_1430_sv2v_reg;
  assign mem[1429] = mem_1429_sv2v_reg;
  assign mem[1428] = mem_1428_sv2v_reg;
  assign mem[1427] = mem_1427_sv2v_reg;
  assign mem[1426] = mem_1426_sv2v_reg;
  assign mem[1425] = mem_1425_sv2v_reg;
  assign mem[1424] = mem_1424_sv2v_reg;
  assign mem[1423] = mem_1423_sv2v_reg;
  assign mem[1422] = mem_1422_sv2v_reg;
  assign mem[1421] = mem_1421_sv2v_reg;
  assign mem[1420] = mem_1420_sv2v_reg;
  assign mem[1419] = mem_1419_sv2v_reg;
  assign mem[1418] = mem_1418_sv2v_reg;
  assign mem[1417] = mem_1417_sv2v_reg;
  assign mem[1416] = mem_1416_sv2v_reg;
  assign mem[1415] = mem_1415_sv2v_reg;
  assign mem[1414] = mem_1414_sv2v_reg;
  assign mem[1413] = mem_1413_sv2v_reg;
  assign mem[1412] = mem_1412_sv2v_reg;
  assign mem[1411] = mem_1411_sv2v_reg;
  assign mem[1410] = mem_1410_sv2v_reg;
  assign mem[1409] = mem_1409_sv2v_reg;
  assign mem[1408] = mem_1408_sv2v_reg;
  assign mem[1407] = mem_1407_sv2v_reg;
  assign mem[1406] = mem_1406_sv2v_reg;
  assign mem[1405] = mem_1405_sv2v_reg;
  assign mem[1404] = mem_1404_sv2v_reg;
  assign mem[1403] = mem_1403_sv2v_reg;
  assign mem[1402] = mem_1402_sv2v_reg;
  assign mem[1401] = mem_1401_sv2v_reg;
  assign mem[1400] = mem_1400_sv2v_reg;
  assign mem[1399] = mem_1399_sv2v_reg;
  assign mem[1398] = mem_1398_sv2v_reg;
  assign mem[1397] = mem_1397_sv2v_reg;
  assign mem[1396] = mem_1396_sv2v_reg;
  assign mem[1395] = mem_1395_sv2v_reg;
  assign mem[1394] = mem_1394_sv2v_reg;
  assign mem[1393] = mem_1393_sv2v_reg;
  assign mem[1392] = mem_1392_sv2v_reg;
  assign mem[1391] = mem_1391_sv2v_reg;
  assign mem[1390] = mem_1390_sv2v_reg;
  assign mem[1389] = mem_1389_sv2v_reg;
  assign mem[1388] = mem_1388_sv2v_reg;
  assign mem[1387] = mem_1387_sv2v_reg;
  assign mem[1386] = mem_1386_sv2v_reg;
  assign mem[1385] = mem_1385_sv2v_reg;
  assign mem[1384] = mem_1384_sv2v_reg;
  assign mem[1383] = mem_1383_sv2v_reg;
  assign mem[1382] = mem_1382_sv2v_reg;
  assign mem[1381] = mem_1381_sv2v_reg;
  assign mem[1380] = mem_1380_sv2v_reg;
  assign mem[1379] = mem_1379_sv2v_reg;
  assign mem[1378] = mem_1378_sv2v_reg;
  assign mem[1377] = mem_1377_sv2v_reg;
  assign mem[1376] = mem_1376_sv2v_reg;
  assign mem[1375] = mem_1375_sv2v_reg;
  assign mem[1374] = mem_1374_sv2v_reg;
  assign mem[1373] = mem_1373_sv2v_reg;
  assign mem[1372] = mem_1372_sv2v_reg;
  assign mem[1371] = mem_1371_sv2v_reg;
  assign mem[1370] = mem_1370_sv2v_reg;
  assign mem[1369] = mem_1369_sv2v_reg;
  assign mem[1368] = mem_1368_sv2v_reg;
  assign mem[1367] = mem_1367_sv2v_reg;
  assign mem[1366] = mem_1366_sv2v_reg;
  assign mem[1365] = mem_1365_sv2v_reg;
  assign mem[1364] = mem_1364_sv2v_reg;
  assign mem[1363] = mem_1363_sv2v_reg;
  assign mem[1362] = mem_1362_sv2v_reg;
  assign mem[1361] = mem_1361_sv2v_reg;
  assign mem[1360] = mem_1360_sv2v_reg;
  assign mem[1359] = mem_1359_sv2v_reg;
  assign mem[1358] = mem_1358_sv2v_reg;
  assign mem[1357] = mem_1357_sv2v_reg;
  assign mem[1356] = mem_1356_sv2v_reg;
  assign mem[1355] = mem_1355_sv2v_reg;
  assign mem[1354] = mem_1354_sv2v_reg;
  assign mem[1353] = mem_1353_sv2v_reg;
  assign mem[1352] = mem_1352_sv2v_reg;
  assign mem[1351] = mem_1351_sv2v_reg;
  assign mem[1350] = mem_1350_sv2v_reg;
  assign mem[1349] = mem_1349_sv2v_reg;
  assign mem[1348] = mem_1348_sv2v_reg;
  assign mem[1347] = mem_1347_sv2v_reg;
  assign mem[1346] = mem_1346_sv2v_reg;
  assign mem[1345] = mem_1345_sv2v_reg;
  assign mem[1344] = mem_1344_sv2v_reg;
  assign mem[1343] = mem_1343_sv2v_reg;
  assign mem[1342] = mem_1342_sv2v_reg;
  assign mem[1341] = mem_1341_sv2v_reg;
  assign mem[1340] = mem_1340_sv2v_reg;
  assign mem[1339] = mem_1339_sv2v_reg;
  assign mem[1338] = mem_1338_sv2v_reg;
  assign mem[1337] = mem_1337_sv2v_reg;
  assign mem[1336] = mem_1336_sv2v_reg;
  assign mem[1335] = mem_1335_sv2v_reg;
  assign mem[1334] = mem_1334_sv2v_reg;
  assign mem[1333] = mem_1333_sv2v_reg;
  assign mem[1332] = mem_1332_sv2v_reg;
  assign mem[1331] = mem_1331_sv2v_reg;
  assign mem[1330] = mem_1330_sv2v_reg;
  assign mem[1329] = mem_1329_sv2v_reg;
  assign mem[1328] = mem_1328_sv2v_reg;
  assign mem[1327] = mem_1327_sv2v_reg;
  assign mem[1326] = mem_1326_sv2v_reg;
  assign mem[1325] = mem_1325_sv2v_reg;
  assign mem[1324] = mem_1324_sv2v_reg;
  assign mem[1323] = mem_1323_sv2v_reg;
  assign mem[1322] = mem_1322_sv2v_reg;
  assign mem[1321] = mem_1321_sv2v_reg;
  assign mem[1320] = mem_1320_sv2v_reg;
  assign mem[1319] = mem_1319_sv2v_reg;
  assign mem[1318] = mem_1318_sv2v_reg;
  assign mem[1317] = mem_1317_sv2v_reg;
  assign mem[1316] = mem_1316_sv2v_reg;
  assign mem[1315] = mem_1315_sv2v_reg;
  assign mem[1314] = mem_1314_sv2v_reg;
  assign mem[1313] = mem_1313_sv2v_reg;
  assign mem[1312] = mem_1312_sv2v_reg;
  assign mem[1311] = mem_1311_sv2v_reg;
  assign mem[1310] = mem_1310_sv2v_reg;
  assign mem[1309] = mem_1309_sv2v_reg;
  assign mem[1308] = mem_1308_sv2v_reg;
  assign mem[1307] = mem_1307_sv2v_reg;
  assign mem[1306] = mem_1306_sv2v_reg;
  assign mem[1305] = mem_1305_sv2v_reg;
  assign mem[1304] = mem_1304_sv2v_reg;
  assign mem[1303] = mem_1303_sv2v_reg;
  assign mem[1302] = mem_1302_sv2v_reg;
  assign mem[1301] = mem_1301_sv2v_reg;
  assign mem[1300] = mem_1300_sv2v_reg;
  assign mem[1299] = mem_1299_sv2v_reg;
  assign mem[1298] = mem_1298_sv2v_reg;
  assign mem[1297] = mem_1297_sv2v_reg;
  assign mem[1296] = mem_1296_sv2v_reg;
  assign mem[1295] = mem_1295_sv2v_reg;
  assign mem[1294] = mem_1294_sv2v_reg;
  assign mem[1293] = mem_1293_sv2v_reg;
  assign mem[1292] = mem_1292_sv2v_reg;
  assign mem[1291] = mem_1291_sv2v_reg;
  assign mem[1290] = mem_1290_sv2v_reg;
  assign mem[1289] = mem_1289_sv2v_reg;
  assign mem[1288] = mem_1288_sv2v_reg;
  assign mem[1287] = mem_1287_sv2v_reg;
  assign mem[1286] = mem_1286_sv2v_reg;
  assign mem[1285] = mem_1285_sv2v_reg;
  assign mem[1284] = mem_1284_sv2v_reg;
  assign mem[1283] = mem_1283_sv2v_reg;
  assign mem[1282] = mem_1282_sv2v_reg;
  assign mem[1281] = mem_1281_sv2v_reg;
  assign mem[1280] = mem_1280_sv2v_reg;
  assign mem[1279] = mem_1279_sv2v_reg;
  assign mem[1278] = mem_1278_sv2v_reg;
  assign mem[1277] = mem_1277_sv2v_reg;
  assign mem[1276] = mem_1276_sv2v_reg;
  assign mem[1275] = mem_1275_sv2v_reg;
  assign mem[1274] = mem_1274_sv2v_reg;
  assign mem[1273] = mem_1273_sv2v_reg;
  assign mem[1272] = mem_1272_sv2v_reg;
  assign mem[1271] = mem_1271_sv2v_reg;
  assign mem[1270] = mem_1270_sv2v_reg;
  assign mem[1269] = mem_1269_sv2v_reg;
  assign mem[1268] = mem_1268_sv2v_reg;
  assign mem[1267] = mem_1267_sv2v_reg;
  assign mem[1266] = mem_1266_sv2v_reg;
  assign mem[1265] = mem_1265_sv2v_reg;
  assign mem[1264] = mem_1264_sv2v_reg;
  assign mem[1263] = mem_1263_sv2v_reg;
  assign mem[1262] = mem_1262_sv2v_reg;
  assign mem[1261] = mem_1261_sv2v_reg;
  assign mem[1260] = mem_1260_sv2v_reg;
  assign mem[1259] = mem_1259_sv2v_reg;
  assign mem[1258] = mem_1258_sv2v_reg;
  assign mem[1257] = mem_1257_sv2v_reg;
  assign mem[1256] = mem_1256_sv2v_reg;
  assign mem[1255] = mem_1255_sv2v_reg;
  assign mem[1254] = mem_1254_sv2v_reg;
  assign mem[1253] = mem_1253_sv2v_reg;
  assign mem[1252] = mem_1252_sv2v_reg;
  assign mem[1251] = mem_1251_sv2v_reg;
  assign mem[1250] = mem_1250_sv2v_reg;
  assign mem[1249] = mem_1249_sv2v_reg;
  assign mem[1248] = mem_1248_sv2v_reg;
  assign mem[1247] = mem_1247_sv2v_reg;
  assign mem[1246] = mem_1246_sv2v_reg;
  assign mem[1245] = mem_1245_sv2v_reg;
  assign mem[1244] = mem_1244_sv2v_reg;
  assign mem[1243] = mem_1243_sv2v_reg;
  assign mem[1242] = mem_1242_sv2v_reg;
  assign mem[1241] = mem_1241_sv2v_reg;
  assign mem[1240] = mem_1240_sv2v_reg;
  assign mem[1239] = mem_1239_sv2v_reg;
  assign mem[1238] = mem_1238_sv2v_reg;
  assign mem[1237] = mem_1237_sv2v_reg;
  assign mem[1236] = mem_1236_sv2v_reg;
  assign mem[1235] = mem_1235_sv2v_reg;
  assign mem[1234] = mem_1234_sv2v_reg;
  assign mem[1233] = mem_1233_sv2v_reg;
  assign mem[1232] = mem_1232_sv2v_reg;
  assign mem[1231] = mem_1231_sv2v_reg;
  assign mem[1230] = mem_1230_sv2v_reg;
  assign mem[1229] = mem_1229_sv2v_reg;
  assign mem[1228] = mem_1228_sv2v_reg;
  assign mem[1227] = mem_1227_sv2v_reg;
  assign mem[1226] = mem_1226_sv2v_reg;
  assign mem[1225] = mem_1225_sv2v_reg;
  assign mem[1224] = mem_1224_sv2v_reg;
  assign mem[1223] = mem_1223_sv2v_reg;
  assign mem[1222] = mem_1222_sv2v_reg;
  assign mem[1221] = mem_1221_sv2v_reg;
  assign mem[1220] = mem_1220_sv2v_reg;
  assign mem[1219] = mem_1219_sv2v_reg;
  assign mem[1218] = mem_1218_sv2v_reg;
  assign mem[1217] = mem_1217_sv2v_reg;
  assign mem[1216] = mem_1216_sv2v_reg;
  assign mem[1215] = mem_1215_sv2v_reg;
  assign mem[1214] = mem_1214_sv2v_reg;
  assign mem[1213] = mem_1213_sv2v_reg;
  assign mem[1212] = mem_1212_sv2v_reg;
  assign mem[1211] = mem_1211_sv2v_reg;
  assign mem[1210] = mem_1210_sv2v_reg;
  assign mem[1209] = mem_1209_sv2v_reg;
  assign mem[1208] = mem_1208_sv2v_reg;
  assign mem[1207] = mem_1207_sv2v_reg;
  assign mem[1206] = mem_1206_sv2v_reg;
  assign mem[1205] = mem_1205_sv2v_reg;
  assign mem[1204] = mem_1204_sv2v_reg;
  assign mem[1203] = mem_1203_sv2v_reg;
  assign mem[1202] = mem_1202_sv2v_reg;
  assign mem[1201] = mem_1201_sv2v_reg;
  assign mem[1200] = mem_1200_sv2v_reg;
  assign mem[1199] = mem_1199_sv2v_reg;
  assign mem[1198] = mem_1198_sv2v_reg;
  assign mem[1197] = mem_1197_sv2v_reg;
  assign mem[1196] = mem_1196_sv2v_reg;
  assign mem[1195] = mem_1195_sv2v_reg;
  assign mem[1194] = mem_1194_sv2v_reg;
  assign mem[1193] = mem_1193_sv2v_reg;
  assign mem[1192] = mem_1192_sv2v_reg;
  assign mem[1191] = mem_1191_sv2v_reg;
  assign mem[1190] = mem_1190_sv2v_reg;
  assign mem[1189] = mem_1189_sv2v_reg;
  assign mem[1188] = mem_1188_sv2v_reg;
  assign mem[1187] = mem_1187_sv2v_reg;
  assign mem[1186] = mem_1186_sv2v_reg;
  assign mem[1185] = mem_1185_sv2v_reg;
  assign mem[1184] = mem_1184_sv2v_reg;
  assign mem[1183] = mem_1183_sv2v_reg;
  assign mem[1182] = mem_1182_sv2v_reg;
  assign mem[1181] = mem_1181_sv2v_reg;
  assign mem[1180] = mem_1180_sv2v_reg;
  assign mem[1179] = mem_1179_sv2v_reg;
  assign mem[1178] = mem_1178_sv2v_reg;
  assign mem[1177] = mem_1177_sv2v_reg;
  assign mem[1176] = mem_1176_sv2v_reg;
  assign mem[1175] = mem_1175_sv2v_reg;
  assign mem[1174] = mem_1174_sv2v_reg;
  assign mem[1173] = mem_1173_sv2v_reg;
  assign mem[1172] = mem_1172_sv2v_reg;
  assign mem[1171] = mem_1171_sv2v_reg;
  assign mem[1170] = mem_1170_sv2v_reg;
  assign mem[1169] = mem_1169_sv2v_reg;
  assign mem[1168] = mem_1168_sv2v_reg;
  assign mem[1167] = mem_1167_sv2v_reg;
  assign mem[1166] = mem_1166_sv2v_reg;
  assign mem[1165] = mem_1165_sv2v_reg;
  assign mem[1164] = mem_1164_sv2v_reg;
  assign mem[1163] = mem_1163_sv2v_reg;
  assign mem[1162] = mem_1162_sv2v_reg;
  assign mem[1161] = mem_1161_sv2v_reg;
  assign mem[1160] = mem_1160_sv2v_reg;
  assign mem[1159] = mem_1159_sv2v_reg;
  assign mem[1158] = mem_1158_sv2v_reg;
  assign mem[1157] = mem_1157_sv2v_reg;
  assign mem[1156] = mem_1156_sv2v_reg;
  assign mem[1155] = mem_1155_sv2v_reg;
  assign mem[1154] = mem_1154_sv2v_reg;
  assign mem[1153] = mem_1153_sv2v_reg;
  assign mem[1152] = mem_1152_sv2v_reg;
  assign mem[1151] = mem_1151_sv2v_reg;
  assign mem[1150] = mem_1150_sv2v_reg;
  assign mem[1149] = mem_1149_sv2v_reg;
  assign mem[1148] = mem_1148_sv2v_reg;
  assign mem[1147] = mem_1147_sv2v_reg;
  assign mem[1146] = mem_1146_sv2v_reg;
  assign mem[1145] = mem_1145_sv2v_reg;
  assign mem[1144] = mem_1144_sv2v_reg;
  assign mem[1143] = mem_1143_sv2v_reg;
  assign mem[1142] = mem_1142_sv2v_reg;
  assign mem[1141] = mem_1141_sv2v_reg;
  assign mem[1140] = mem_1140_sv2v_reg;
  assign mem[1139] = mem_1139_sv2v_reg;
  assign mem[1138] = mem_1138_sv2v_reg;
  assign mem[1137] = mem_1137_sv2v_reg;
  assign mem[1136] = mem_1136_sv2v_reg;
  assign mem[1135] = mem_1135_sv2v_reg;
  assign mem[1134] = mem_1134_sv2v_reg;
  assign mem[1133] = mem_1133_sv2v_reg;
  assign mem[1132] = mem_1132_sv2v_reg;
  assign mem[1131] = mem_1131_sv2v_reg;
  assign mem[1130] = mem_1130_sv2v_reg;
  assign mem[1129] = mem_1129_sv2v_reg;
  assign mem[1128] = mem_1128_sv2v_reg;
  assign mem[1127] = mem_1127_sv2v_reg;
  assign mem[1126] = mem_1126_sv2v_reg;
  assign mem[1125] = mem_1125_sv2v_reg;
  assign mem[1124] = mem_1124_sv2v_reg;
  assign mem[1123] = mem_1123_sv2v_reg;
  assign mem[1122] = mem_1122_sv2v_reg;
  assign mem[1121] = mem_1121_sv2v_reg;
  assign mem[1120] = mem_1120_sv2v_reg;
  assign mem[1119] = mem_1119_sv2v_reg;
  assign mem[1118] = mem_1118_sv2v_reg;
  assign mem[1117] = mem_1117_sv2v_reg;
  assign mem[1116] = mem_1116_sv2v_reg;
  assign mem[1115] = mem_1115_sv2v_reg;
  assign mem[1114] = mem_1114_sv2v_reg;
  assign mem[1113] = mem_1113_sv2v_reg;
  assign mem[1112] = mem_1112_sv2v_reg;
  assign mem[1111] = mem_1111_sv2v_reg;
  assign mem[1110] = mem_1110_sv2v_reg;
  assign mem[1109] = mem_1109_sv2v_reg;
  assign mem[1108] = mem_1108_sv2v_reg;
  assign mem[1107] = mem_1107_sv2v_reg;
  assign mem[1106] = mem_1106_sv2v_reg;
  assign mem[1105] = mem_1105_sv2v_reg;
  assign mem[1104] = mem_1104_sv2v_reg;
  assign mem[1103] = mem_1103_sv2v_reg;
  assign mem[1102] = mem_1102_sv2v_reg;
  assign mem[1101] = mem_1101_sv2v_reg;
  assign mem[1100] = mem_1100_sv2v_reg;
  assign mem[1099] = mem_1099_sv2v_reg;
  assign mem[1098] = mem_1098_sv2v_reg;
  assign mem[1097] = mem_1097_sv2v_reg;
  assign mem[1096] = mem_1096_sv2v_reg;
  assign mem[1095] = mem_1095_sv2v_reg;
  assign mem[1094] = mem_1094_sv2v_reg;
  assign mem[1093] = mem_1093_sv2v_reg;
  assign mem[1092] = mem_1092_sv2v_reg;
  assign mem[1091] = mem_1091_sv2v_reg;
  assign mem[1090] = mem_1090_sv2v_reg;
  assign mem[1089] = mem_1089_sv2v_reg;
  assign mem[1088] = mem_1088_sv2v_reg;
  assign mem[1087] = mem_1087_sv2v_reg;
  assign mem[1086] = mem_1086_sv2v_reg;
  assign mem[1085] = mem_1085_sv2v_reg;
  assign mem[1084] = mem_1084_sv2v_reg;
  assign mem[1083] = mem_1083_sv2v_reg;
  assign mem[1082] = mem_1082_sv2v_reg;
  assign mem[1081] = mem_1081_sv2v_reg;
  assign mem[1080] = mem_1080_sv2v_reg;
  assign mem[1079] = mem_1079_sv2v_reg;
  assign mem[1078] = mem_1078_sv2v_reg;
  assign mem[1077] = mem_1077_sv2v_reg;
  assign mem[1076] = mem_1076_sv2v_reg;
  assign mem[1075] = mem_1075_sv2v_reg;
  assign mem[1074] = mem_1074_sv2v_reg;
  assign mem[1073] = mem_1073_sv2v_reg;
  assign mem[1072] = mem_1072_sv2v_reg;
  assign mem[1071] = mem_1071_sv2v_reg;
  assign mem[1070] = mem_1070_sv2v_reg;
  assign mem[1069] = mem_1069_sv2v_reg;
  assign mem[1068] = mem_1068_sv2v_reg;
  assign mem[1067] = mem_1067_sv2v_reg;
  assign mem[1066] = mem_1066_sv2v_reg;
  assign mem[1065] = mem_1065_sv2v_reg;
  assign mem[1064] = mem_1064_sv2v_reg;
  assign mem[1063] = mem_1063_sv2v_reg;
  assign mem[1062] = mem_1062_sv2v_reg;
  assign mem[1061] = mem_1061_sv2v_reg;
  assign mem[1060] = mem_1060_sv2v_reg;
  assign mem[1059] = mem_1059_sv2v_reg;
  assign mem[1058] = mem_1058_sv2v_reg;
  assign mem[1057] = mem_1057_sv2v_reg;
  assign mem[1056] = mem_1056_sv2v_reg;
  assign mem[1055] = mem_1055_sv2v_reg;
  assign mem[1054] = mem_1054_sv2v_reg;
  assign mem[1053] = mem_1053_sv2v_reg;
  assign mem[1052] = mem_1052_sv2v_reg;
  assign mem[1051] = mem_1051_sv2v_reg;
  assign mem[1050] = mem_1050_sv2v_reg;
  assign mem[1049] = mem_1049_sv2v_reg;
  assign mem[1048] = mem_1048_sv2v_reg;
  assign mem[1047] = mem_1047_sv2v_reg;
  assign mem[1046] = mem_1046_sv2v_reg;
  assign mem[1045] = mem_1045_sv2v_reg;
  assign mem[1044] = mem_1044_sv2v_reg;
  assign mem[1043] = mem_1043_sv2v_reg;
  assign mem[1042] = mem_1042_sv2v_reg;
  assign mem[1041] = mem_1041_sv2v_reg;
  assign mem[1040] = mem_1040_sv2v_reg;
  assign mem[1039] = mem_1039_sv2v_reg;
  assign mem[1038] = mem_1038_sv2v_reg;
  assign mem[1037] = mem_1037_sv2v_reg;
  assign mem[1036] = mem_1036_sv2v_reg;
  assign mem[1035] = mem_1035_sv2v_reg;
  assign mem[1034] = mem_1034_sv2v_reg;
  assign mem[1033] = mem_1033_sv2v_reg;
  assign mem[1032] = mem_1032_sv2v_reg;
  assign mem[1031] = mem_1031_sv2v_reg;
  assign mem[1030] = mem_1030_sv2v_reg;
  assign mem[1029] = mem_1029_sv2v_reg;
  assign mem[1028] = mem_1028_sv2v_reg;
  assign mem[1027] = mem_1027_sv2v_reg;
  assign mem[1026] = mem_1026_sv2v_reg;
  assign mem[1025] = mem_1025_sv2v_reg;
  assign mem[1024] = mem_1024_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[1599] = (N3)? mem[1599] : 
                          (N0)? mem[3199] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[1598] = (N3)? mem[1598] : 
                          (N0)? mem[3198] : 1'b0;
  assign r_data_o[1597] = (N3)? mem[1597] : 
                          (N0)? mem[3197] : 1'b0;
  assign r_data_o[1596] = (N3)? mem[1596] : 
                          (N0)? mem[3196] : 1'b0;
  assign r_data_o[1595] = (N3)? mem[1595] : 
                          (N0)? mem[3195] : 1'b0;
  assign r_data_o[1594] = (N3)? mem[1594] : 
                          (N0)? mem[3194] : 1'b0;
  assign r_data_o[1593] = (N3)? mem[1593] : 
                          (N0)? mem[3193] : 1'b0;
  assign r_data_o[1592] = (N3)? mem[1592] : 
                          (N0)? mem[3192] : 1'b0;
  assign r_data_o[1591] = (N3)? mem[1591] : 
                          (N0)? mem[3191] : 1'b0;
  assign r_data_o[1590] = (N3)? mem[1590] : 
                          (N0)? mem[3190] : 1'b0;
  assign r_data_o[1589] = (N3)? mem[1589] : 
                          (N0)? mem[3189] : 1'b0;
  assign r_data_o[1588] = (N3)? mem[1588] : 
                          (N0)? mem[3188] : 1'b0;
  assign r_data_o[1587] = (N3)? mem[1587] : 
                          (N0)? mem[3187] : 1'b0;
  assign r_data_o[1586] = (N3)? mem[1586] : 
                          (N0)? mem[3186] : 1'b0;
  assign r_data_o[1585] = (N3)? mem[1585] : 
                          (N0)? mem[3185] : 1'b0;
  assign r_data_o[1584] = (N3)? mem[1584] : 
                          (N0)? mem[3184] : 1'b0;
  assign r_data_o[1583] = (N3)? mem[1583] : 
                          (N0)? mem[3183] : 1'b0;
  assign r_data_o[1582] = (N3)? mem[1582] : 
                          (N0)? mem[3182] : 1'b0;
  assign r_data_o[1581] = (N3)? mem[1581] : 
                          (N0)? mem[3181] : 1'b0;
  assign r_data_o[1580] = (N3)? mem[1580] : 
                          (N0)? mem[3180] : 1'b0;
  assign r_data_o[1579] = (N3)? mem[1579] : 
                          (N0)? mem[3179] : 1'b0;
  assign r_data_o[1578] = (N3)? mem[1578] : 
                          (N0)? mem[3178] : 1'b0;
  assign r_data_o[1577] = (N3)? mem[1577] : 
                          (N0)? mem[3177] : 1'b0;
  assign r_data_o[1576] = (N3)? mem[1576] : 
                          (N0)? mem[3176] : 1'b0;
  assign r_data_o[1575] = (N3)? mem[1575] : 
                          (N0)? mem[3175] : 1'b0;
  assign r_data_o[1574] = (N3)? mem[1574] : 
                          (N0)? mem[3174] : 1'b0;
  assign r_data_o[1573] = (N3)? mem[1573] : 
                          (N0)? mem[3173] : 1'b0;
  assign r_data_o[1572] = (N3)? mem[1572] : 
                          (N0)? mem[3172] : 1'b0;
  assign r_data_o[1571] = (N3)? mem[1571] : 
                          (N0)? mem[3171] : 1'b0;
  assign r_data_o[1570] = (N3)? mem[1570] : 
                          (N0)? mem[3170] : 1'b0;
  assign r_data_o[1569] = (N3)? mem[1569] : 
                          (N0)? mem[3169] : 1'b0;
  assign r_data_o[1568] = (N3)? mem[1568] : 
                          (N0)? mem[3168] : 1'b0;
  assign r_data_o[1567] = (N3)? mem[1567] : 
                          (N0)? mem[3167] : 1'b0;
  assign r_data_o[1566] = (N3)? mem[1566] : 
                          (N0)? mem[3166] : 1'b0;
  assign r_data_o[1565] = (N3)? mem[1565] : 
                          (N0)? mem[3165] : 1'b0;
  assign r_data_o[1564] = (N3)? mem[1564] : 
                          (N0)? mem[3164] : 1'b0;
  assign r_data_o[1563] = (N3)? mem[1563] : 
                          (N0)? mem[3163] : 1'b0;
  assign r_data_o[1562] = (N3)? mem[1562] : 
                          (N0)? mem[3162] : 1'b0;
  assign r_data_o[1561] = (N3)? mem[1561] : 
                          (N0)? mem[3161] : 1'b0;
  assign r_data_o[1560] = (N3)? mem[1560] : 
                          (N0)? mem[3160] : 1'b0;
  assign r_data_o[1559] = (N3)? mem[1559] : 
                          (N0)? mem[3159] : 1'b0;
  assign r_data_o[1558] = (N3)? mem[1558] : 
                          (N0)? mem[3158] : 1'b0;
  assign r_data_o[1557] = (N3)? mem[1557] : 
                          (N0)? mem[3157] : 1'b0;
  assign r_data_o[1556] = (N3)? mem[1556] : 
                          (N0)? mem[3156] : 1'b0;
  assign r_data_o[1555] = (N3)? mem[1555] : 
                          (N0)? mem[3155] : 1'b0;
  assign r_data_o[1554] = (N3)? mem[1554] : 
                          (N0)? mem[3154] : 1'b0;
  assign r_data_o[1553] = (N3)? mem[1553] : 
                          (N0)? mem[3153] : 1'b0;
  assign r_data_o[1552] = (N3)? mem[1552] : 
                          (N0)? mem[3152] : 1'b0;
  assign r_data_o[1551] = (N3)? mem[1551] : 
                          (N0)? mem[3151] : 1'b0;
  assign r_data_o[1550] = (N3)? mem[1550] : 
                          (N0)? mem[3150] : 1'b0;
  assign r_data_o[1549] = (N3)? mem[1549] : 
                          (N0)? mem[3149] : 1'b0;
  assign r_data_o[1548] = (N3)? mem[1548] : 
                          (N0)? mem[3148] : 1'b0;
  assign r_data_o[1547] = (N3)? mem[1547] : 
                          (N0)? mem[3147] : 1'b0;
  assign r_data_o[1546] = (N3)? mem[1546] : 
                          (N0)? mem[3146] : 1'b0;
  assign r_data_o[1545] = (N3)? mem[1545] : 
                          (N0)? mem[3145] : 1'b0;
  assign r_data_o[1544] = (N3)? mem[1544] : 
                          (N0)? mem[3144] : 1'b0;
  assign r_data_o[1543] = (N3)? mem[1543] : 
                          (N0)? mem[3143] : 1'b0;
  assign r_data_o[1542] = (N3)? mem[1542] : 
                          (N0)? mem[3142] : 1'b0;
  assign r_data_o[1541] = (N3)? mem[1541] : 
                          (N0)? mem[3141] : 1'b0;
  assign r_data_o[1540] = (N3)? mem[1540] : 
                          (N0)? mem[3140] : 1'b0;
  assign r_data_o[1539] = (N3)? mem[1539] : 
                          (N0)? mem[3139] : 1'b0;
  assign r_data_o[1538] = (N3)? mem[1538] : 
                          (N0)? mem[3138] : 1'b0;
  assign r_data_o[1537] = (N3)? mem[1537] : 
                          (N0)? mem[3137] : 1'b0;
  assign r_data_o[1536] = (N3)? mem[1536] : 
                          (N0)? mem[3136] : 1'b0;
  assign r_data_o[1535] = (N3)? mem[1535] : 
                          (N0)? mem[3135] : 1'b0;
  assign r_data_o[1534] = (N3)? mem[1534] : 
                          (N0)? mem[3134] : 1'b0;
  assign r_data_o[1533] = (N3)? mem[1533] : 
                          (N0)? mem[3133] : 1'b0;
  assign r_data_o[1532] = (N3)? mem[1532] : 
                          (N0)? mem[3132] : 1'b0;
  assign r_data_o[1531] = (N3)? mem[1531] : 
                          (N0)? mem[3131] : 1'b0;
  assign r_data_o[1530] = (N3)? mem[1530] : 
                          (N0)? mem[3130] : 1'b0;
  assign r_data_o[1529] = (N3)? mem[1529] : 
                          (N0)? mem[3129] : 1'b0;
  assign r_data_o[1528] = (N3)? mem[1528] : 
                          (N0)? mem[3128] : 1'b0;
  assign r_data_o[1527] = (N3)? mem[1527] : 
                          (N0)? mem[3127] : 1'b0;
  assign r_data_o[1526] = (N3)? mem[1526] : 
                          (N0)? mem[3126] : 1'b0;
  assign r_data_o[1525] = (N3)? mem[1525] : 
                          (N0)? mem[3125] : 1'b0;
  assign r_data_o[1524] = (N3)? mem[1524] : 
                          (N0)? mem[3124] : 1'b0;
  assign r_data_o[1523] = (N3)? mem[1523] : 
                          (N0)? mem[3123] : 1'b0;
  assign r_data_o[1522] = (N3)? mem[1522] : 
                          (N0)? mem[3122] : 1'b0;
  assign r_data_o[1521] = (N3)? mem[1521] : 
                          (N0)? mem[3121] : 1'b0;
  assign r_data_o[1520] = (N3)? mem[1520] : 
                          (N0)? mem[3120] : 1'b0;
  assign r_data_o[1519] = (N3)? mem[1519] : 
                          (N0)? mem[3119] : 1'b0;
  assign r_data_o[1518] = (N3)? mem[1518] : 
                          (N0)? mem[3118] : 1'b0;
  assign r_data_o[1517] = (N3)? mem[1517] : 
                          (N0)? mem[3117] : 1'b0;
  assign r_data_o[1516] = (N3)? mem[1516] : 
                          (N0)? mem[3116] : 1'b0;
  assign r_data_o[1515] = (N3)? mem[1515] : 
                          (N0)? mem[3115] : 1'b0;
  assign r_data_o[1514] = (N3)? mem[1514] : 
                          (N0)? mem[3114] : 1'b0;
  assign r_data_o[1513] = (N3)? mem[1513] : 
                          (N0)? mem[3113] : 1'b0;
  assign r_data_o[1512] = (N3)? mem[1512] : 
                          (N0)? mem[3112] : 1'b0;
  assign r_data_o[1511] = (N3)? mem[1511] : 
                          (N0)? mem[3111] : 1'b0;
  assign r_data_o[1510] = (N3)? mem[1510] : 
                          (N0)? mem[3110] : 1'b0;
  assign r_data_o[1509] = (N3)? mem[1509] : 
                          (N0)? mem[3109] : 1'b0;
  assign r_data_o[1508] = (N3)? mem[1508] : 
                          (N0)? mem[3108] : 1'b0;
  assign r_data_o[1507] = (N3)? mem[1507] : 
                          (N0)? mem[3107] : 1'b0;
  assign r_data_o[1506] = (N3)? mem[1506] : 
                          (N0)? mem[3106] : 1'b0;
  assign r_data_o[1505] = (N3)? mem[1505] : 
                          (N0)? mem[3105] : 1'b0;
  assign r_data_o[1504] = (N3)? mem[1504] : 
                          (N0)? mem[3104] : 1'b0;
  assign r_data_o[1503] = (N3)? mem[1503] : 
                          (N0)? mem[3103] : 1'b0;
  assign r_data_o[1502] = (N3)? mem[1502] : 
                          (N0)? mem[3102] : 1'b0;
  assign r_data_o[1501] = (N3)? mem[1501] : 
                          (N0)? mem[3101] : 1'b0;
  assign r_data_o[1500] = (N3)? mem[1500] : 
                          (N0)? mem[3100] : 1'b0;
  assign r_data_o[1499] = (N3)? mem[1499] : 
                          (N0)? mem[3099] : 1'b0;
  assign r_data_o[1498] = (N3)? mem[1498] : 
                          (N0)? mem[3098] : 1'b0;
  assign r_data_o[1497] = (N3)? mem[1497] : 
                          (N0)? mem[3097] : 1'b0;
  assign r_data_o[1496] = (N3)? mem[1496] : 
                          (N0)? mem[3096] : 1'b0;
  assign r_data_o[1495] = (N3)? mem[1495] : 
                          (N0)? mem[3095] : 1'b0;
  assign r_data_o[1494] = (N3)? mem[1494] : 
                          (N0)? mem[3094] : 1'b0;
  assign r_data_o[1493] = (N3)? mem[1493] : 
                          (N0)? mem[3093] : 1'b0;
  assign r_data_o[1492] = (N3)? mem[1492] : 
                          (N0)? mem[3092] : 1'b0;
  assign r_data_o[1491] = (N3)? mem[1491] : 
                          (N0)? mem[3091] : 1'b0;
  assign r_data_o[1490] = (N3)? mem[1490] : 
                          (N0)? mem[3090] : 1'b0;
  assign r_data_o[1489] = (N3)? mem[1489] : 
                          (N0)? mem[3089] : 1'b0;
  assign r_data_o[1488] = (N3)? mem[1488] : 
                          (N0)? mem[3088] : 1'b0;
  assign r_data_o[1487] = (N3)? mem[1487] : 
                          (N0)? mem[3087] : 1'b0;
  assign r_data_o[1486] = (N3)? mem[1486] : 
                          (N0)? mem[3086] : 1'b0;
  assign r_data_o[1485] = (N3)? mem[1485] : 
                          (N0)? mem[3085] : 1'b0;
  assign r_data_o[1484] = (N3)? mem[1484] : 
                          (N0)? mem[3084] : 1'b0;
  assign r_data_o[1483] = (N3)? mem[1483] : 
                          (N0)? mem[3083] : 1'b0;
  assign r_data_o[1482] = (N3)? mem[1482] : 
                          (N0)? mem[3082] : 1'b0;
  assign r_data_o[1481] = (N3)? mem[1481] : 
                          (N0)? mem[3081] : 1'b0;
  assign r_data_o[1480] = (N3)? mem[1480] : 
                          (N0)? mem[3080] : 1'b0;
  assign r_data_o[1479] = (N3)? mem[1479] : 
                          (N0)? mem[3079] : 1'b0;
  assign r_data_o[1478] = (N3)? mem[1478] : 
                          (N0)? mem[3078] : 1'b0;
  assign r_data_o[1477] = (N3)? mem[1477] : 
                          (N0)? mem[3077] : 1'b0;
  assign r_data_o[1476] = (N3)? mem[1476] : 
                          (N0)? mem[3076] : 1'b0;
  assign r_data_o[1475] = (N3)? mem[1475] : 
                          (N0)? mem[3075] : 1'b0;
  assign r_data_o[1474] = (N3)? mem[1474] : 
                          (N0)? mem[3074] : 1'b0;
  assign r_data_o[1473] = (N3)? mem[1473] : 
                          (N0)? mem[3073] : 1'b0;
  assign r_data_o[1472] = (N3)? mem[1472] : 
                          (N0)? mem[3072] : 1'b0;
  assign r_data_o[1471] = (N3)? mem[1471] : 
                          (N0)? mem[3071] : 1'b0;
  assign r_data_o[1470] = (N3)? mem[1470] : 
                          (N0)? mem[3070] : 1'b0;
  assign r_data_o[1469] = (N3)? mem[1469] : 
                          (N0)? mem[3069] : 1'b0;
  assign r_data_o[1468] = (N3)? mem[1468] : 
                          (N0)? mem[3068] : 1'b0;
  assign r_data_o[1467] = (N3)? mem[1467] : 
                          (N0)? mem[3067] : 1'b0;
  assign r_data_o[1466] = (N3)? mem[1466] : 
                          (N0)? mem[3066] : 1'b0;
  assign r_data_o[1465] = (N3)? mem[1465] : 
                          (N0)? mem[3065] : 1'b0;
  assign r_data_o[1464] = (N3)? mem[1464] : 
                          (N0)? mem[3064] : 1'b0;
  assign r_data_o[1463] = (N3)? mem[1463] : 
                          (N0)? mem[3063] : 1'b0;
  assign r_data_o[1462] = (N3)? mem[1462] : 
                          (N0)? mem[3062] : 1'b0;
  assign r_data_o[1461] = (N3)? mem[1461] : 
                          (N0)? mem[3061] : 1'b0;
  assign r_data_o[1460] = (N3)? mem[1460] : 
                          (N0)? mem[3060] : 1'b0;
  assign r_data_o[1459] = (N3)? mem[1459] : 
                          (N0)? mem[3059] : 1'b0;
  assign r_data_o[1458] = (N3)? mem[1458] : 
                          (N0)? mem[3058] : 1'b0;
  assign r_data_o[1457] = (N3)? mem[1457] : 
                          (N0)? mem[3057] : 1'b0;
  assign r_data_o[1456] = (N3)? mem[1456] : 
                          (N0)? mem[3056] : 1'b0;
  assign r_data_o[1455] = (N3)? mem[1455] : 
                          (N0)? mem[3055] : 1'b0;
  assign r_data_o[1454] = (N3)? mem[1454] : 
                          (N0)? mem[3054] : 1'b0;
  assign r_data_o[1453] = (N3)? mem[1453] : 
                          (N0)? mem[3053] : 1'b0;
  assign r_data_o[1452] = (N3)? mem[1452] : 
                          (N0)? mem[3052] : 1'b0;
  assign r_data_o[1451] = (N3)? mem[1451] : 
                          (N0)? mem[3051] : 1'b0;
  assign r_data_o[1450] = (N3)? mem[1450] : 
                          (N0)? mem[3050] : 1'b0;
  assign r_data_o[1449] = (N3)? mem[1449] : 
                          (N0)? mem[3049] : 1'b0;
  assign r_data_o[1448] = (N3)? mem[1448] : 
                          (N0)? mem[3048] : 1'b0;
  assign r_data_o[1447] = (N3)? mem[1447] : 
                          (N0)? mem[3047] : 1'b0;
  assign r_data_o[1446] = (N3)? mem[1446] : 
                          (N0)? mem[3046] : 1'b0;
  assign r_data_o[1445] = (N3)? mem[1445] : 
                          (N0)? mem[3045] : 1'b0;
  assign r_data_o[1444] = (N3)? mem[1444] : 
                          (N0)? mem[3044] : 1'b0;
  assign r_data_o[1443] = (N3)? mem[1443] : 
                          (N0)? mem[3043] : 1'b0;
  assign r_data_o[1442] = (N3)? mem[1442] : 
                          (N0)? mem[3042] : 1'b0;
  assign r_data_o[1441] = (N3)? mem[1441] : 
                          (N0)? mem[3041] : 1'b0;
  assign r_data_o[1440] = (N3)? mem[1440] : 
                          (N0)? mem[3040] : 1'b0;
  assign r_data_o[1439] = (N3)? mem[1439] : 
                          (N0)? mem[3039] : 1'b0;
  assign r_data_o[1438] = (N3)? mem[1438] : 
                          (N0)? mem[3038] : 1'b0;
  assign r_data_o[1437] = (N3)? mem[1437] : 
                          (N0)? mem[3037] : 1'b0;
  assign r_data_o[1436] = (N3)? mem[1436] : 
                          (N0)? mem[3036] : 1'b0;
  assign r_data_o[1435] = (N3)? mem[1435] : 
                          (N0)? mem[3035] : 1'b0;
  assign r_data_o[1434] = (N3)? mem[1434] : 
                          (N0)? mem[3034] : 1'b0;
  assign r_data_o[1433] = (N3)? mem[1433] : 
                          (N0)? mem[3033] : 1'b0;
  assign r_data_o[1432] = (N3)? mem[1432] : 
                          (N0)? mem[3032] : 1'b0;
  assign r_data_o[1431] = (N3)? mem[1431] : 
                          (N0)? mem[3031] : 1'b0;
  assign r_data_o[1430] = (N3)? mem[1430] : 
                          (N0)? mem[3030] : 1'b0;
  assign r_data_o[1429] = (N3)? mem[1429] : 
                          (N0)? mem[3029] : 1'b0;
  assign r_data_o[1428] = (N3)? mem[1428] : 
                          (N0)? mem[3028] : 1'b0;
  assign r_data_o[1427] = (N3)? mem[1427] : 
                          (N0)? mem[3027] : 1'b0;
  assign r_data_o[1426] = (N3)? mem[1426] : 
                          (N0)? mem[3026] : 1'b0;
  assign r_data_o[1425] = (N3)? mem[1425] : 
                          (N0)? mem[3025] : 1'b0;
  assign r_data_o[1424] = (N3)? mem[1424] : 
                          (N0)? mem[3024] : 1'b0;
  assign r_data_o[1423] = (N3)? mem[1423] : 
                          (N0)? mem[3023] : 1'b0;
  assign r_data_o[1422] = (N3)? mem[1422] : 
                          (N0)? mem[3022] : 1'b0;
  assign r_data_o[1421] = (N3)? mem[1421] : 
                          (N0)? mem[3021] : 1'b0;
  assign r_data_o[1420] = (N3)? mem[1420] : 
                          (N0)? mem[3020] : 1'b0;
  assign r_data_o[1419] = (N3)? mem[1419] : 
                          (N0)? mem[3019] : 1'b0;
  assign r_data_o[1418] = (N3)? mem[1418] : 
                          (N0)? mem[3018] : 1'b0;
  assign r_data_o[1417] = (N3)? mem[1417] : 
                          (N0)? mem[3017] : 1'b0;
  assign r_data_o[1416] = (N3)? mem[1416] : 
                          (N0)? mem[3016] : 1'b0;
  assign r_data_o[1415] = (N3)? mem[1415] : 
                          (N0)? mem[3015] : 1'b0;
  assign r_data_o[1414] = (N3)? mem[1414] : 
                          (N0)? mem[3014] : 1'b0;
  assign r_data_o[1413] = (N3)? mem[1413] : 
                          (N0)? mem[3013] : 1'b0;
  assign r_data_o[1412] = (N3)? mem[1412] : 
                          (N0)? mem[3012] : 1'b0;
  assign r_data_o[1411] = (N3)? mem[1411] : 
                          (N0)? mem[3011] : 1'b0;
  assign r_data_o[1410] = (N3)? mem[1410] : 
                          (N0)? mem[3010] : 1'b0;
  assign r_data_o[1409] = (N3)? mem[1409] : 
                          (N0)? mem[3009] : 1'b0;
  assign r_data_o[1408] = (N3)? mem[1408] : 
                          (N0)? mem[3008] : 1'b0;
  assign r_data_o[1407] = (N3)? mem[1407] : 
                          (N0)? mem[3007] : 1'b0;
  assign r_data_o[1406] = (N3)? mem[1406] : 
                          (N0)? mem[3006] : 1'b0;
  assign r_data_o[1405] = (N3)? mem[1405] : 
                          (N0)? mem[3005] : 1'b0;
  assign r_data_o[1404] = (N3)? mem[1404] : 
                          (N0)? mem[3004] : 1'b0;
  assign r_data_o[1403] = (N3)? mem[1403] : 
                          (N0)? mem[3003] : 1'b0;
  assign r_data_o[1402] = (N3)? mem[1402] : 
                          (N0)? mem[3002] : 1'b0;
  assign r_data_o[1401] = (N3)? mem[1401] : 
                          (N0)? mem[3001] : 1'b0;
  assign r_data_o[1400] = (N3)? mem[1400] : 
                          (N0)? mem[3000] : 1'b0;
  assign r_data_o[1399] = (N3)? mem[1399] : 
                          (N0)? mem[2999] : 1'b0;
  assign r_data_o[1398] = (N3)? mem[1398] : 
                          (N0)? mem[2998] : 1'b0;
  assign r_data_o[1397] = (N3)? mem[1397] : 
                          (N0)? mem[2997] : 1'b0;
  assign r_data_o[1396] = (N3)? mem[1396] : 
                          (N0)? mem[2996] : 1'b0;
  assign r_data_o[1395] = (N3)? mem[1395] : 
                          (N0)? mem[2995] : 1'b0;
  assign r_data_o[1394] = (N3)? mem[1394] : 
                          (N0)? mem[2994] : 1'b0;
  assign r_data_o[1393] = (N3)? mem[1393] : 
                          (N0)? mem[2993] : 1'b0;
  assign r_data_o[1392] = (N3)? mem[1392] : 
                          (N0)? mem[2992] : 1'b0;
  assign r_data_o[1391] = (N3)? mem[1391] : 
                          (N0)? mem[2991] : 1'b0;
  assign r_data_o[1390] = (N3)? mem[1390] : 
                          (N0)? mem[2990] : 1'b0;
  assign r_data_o[1389] = (N3)? mem[1389] : 
                          (N0)? mem[2989] : 1'b0;
  assign r_data_o[1388] = (N3)? mem[1388] : 
                          (N0)? mem[2988] : 1'b0;
  assign r_data_o[1387] = (N3)? mem[1387] : 
                          (N0)? mem[2987] : 1'b0;
  assign r_data_o[1386] = (N3)? mem[1386] : 
                          (N0)? mem[2986] : 1'b0;
  assign r_data_o[1385] = (N3)? mem[1385] : 
                          (N0)? mem[2985] : 1'b0;
  assign r_data_o[1384] = (N3)? mem[1384] : 
                          (N0)? mem[2984] : 1'b0;
  assign r_data_o[1383] = (N3)? mem[1383] : 
                          (N0)? mem[2983] : 1'b0;
  assign r_data_o[1382] = (N3)? mem[1382] : 
                          (N0)? mem[2982] : 1'b0;
  assign r_data_o[1381] = (N3)? mem[1381] : 
                          (N0)? mem[2981] : 1'b0;
  assign r_data_o[1380] = (N3)? mem[1380] : 
                          (N0)? mem[2980] : 1'b0;
  assign r_data_o[1379] = (N3)? mem[1379] : 
                          (N0)? mem[2979] : 1'b0;
  assign r_data_o[1378] = (N3)? mem[1378] : 
                          (N0)? mem[2978] : 1'b0;
  assign r_data_o[1377] = (N3)? mem[1377] : 
                          (N0)? mem[2977] : 1'b0;
  assign r_data_o[1376] = (N3)? mem[1376] : 
                          (N0)? mem[2976] : 1'b0;
  assign r_data_o[1375] = (N3)? mem[1375] : 
                          (N0)? mem[2975] : 1'b0;
  assign r_data_o[1374] = (N3)? mem[1374] : 
                          (N0)? mem[2974] : 1'b0;
  assign r_data_o[1373] = (N3)? mem[1373] : 
                          (N0)? mem[2973] : 1'b0;
  assign r_data_o[1372] = (N3)? mem[1372] : 
                          (N0)? mem[2972] : 1'b0;
  assign r_data_o[1371] = (N3)? mem[1371] : 
                          (N0)? mem[2971] : 1'b0;
  assign r_data_o[1370] = (N3)? mem[1370] : 
                          (N0)? mem[2970] : 1'b0;
  assign r_data_o[1369] = (N3)? mem[1369] : 
                          (N0)? mem[2969] : 1'b0;
  assign r_data_o[1368] = (N3)? mem[1368] : 
                          (N0)? mem[2968] : 1'b0;
  assign r_data_o[1367] = (N3)? mem[1367] : 
                          (N0)? mem[2967] : 1'b0;
  assign r_data_o[1366] = (N3)? mem[1366] : 
                          (N0)? mem[2966] : 1'b0;
  assign r_data_o[1365] = (N3)? mem[1365] : 
                          (N0)? mem[2965] : 1'b0;
  assign r_data_o[1364] = (N3)? mem[1364] : 
                          (N0)? mem[2964] : 1'b0;
  assign r_data_o[1363] = (N3)? mem[1363] : 
                          (N0)? mem[2963] : 1'b0;
  assign r_data_o[1362] = (N3)? mem[1362] : 
                          (N0)? mem[2962] : 1'b0;
  assign r_data_o[1361] = (N3)? mem[1361] : 
                          (N0)? mem[2961] : 1'b0;
  assign r_data_o[1360] = (N3)? mem[1360] : 
                          (N0)? mem[2960] : 1'b0;
  assign r_data_o[1359] = (N3)? mem[1359] : 
                          (N0)? mem[2959] : 1'b0;
  assign r_data_o[1358] = (N3)? mem[1358] : 
                          (N0)? mem[2958] : 1'b0;
  assign r_data_o[1357] = (N3)? mem[1357] : 
                          (N0)? mem[2957] : 1'b0;
  assign r_data_o[1356] = (N3)? mem[1356] : 
                          (N0)? mem[2956] : 1'b0;
  assign r_data_o[1355] = (N3)? mem[1355] : 
                          (N0)? mem[2955] : 1'b0;
  assign r_data_o[1354] = (N3)? mem[1354] : 
                          (N0)? mem[2954] : 1'b0;
  assign r_data_o[1353] = (N3)? mem[1353] : 
                          (N0)? mem[2953] : 1'b0;
  assign r_data_o[1352] = (N3)? mem[1352] : 
                          (N0)? mem[2952] : 1'b0;
  assign r_data_o[1351] = (N3)? mem[1351] : 
                          (N0)? mem[2951] : 1'b0;
  assign r_data_o[1350] = (N3)? mem[1350] : 
                          (N0)? mem[2950] : 1'b0;
  assign r_data_o[1349] = (N3)? mem[1349] : 
                          (N0)? mem[2949] : 1'b0;
  assign r_data_o[1348] = (N3)? mem[1348] : 
                          (N0)? mem[2948] : 1'b0;
  assign r_data_o[1347] = (N3)? mem[1347] : 
                          (N0)? mem[2947] : 1'b0;
  assign r_data_o[1346] = (N3)? mem[1346] : 
                          (N0)? mem[2946] : 1'b0;
  assign r_data_o[1345] = (N3)? mem[1345] : 
                          (N0)? mem[2945] : 1'b0;
  assign r_data_o[1344] = (N3)? mem[1344] : 
                          (N0)? mem[2944] : 1'b0;
  assign r_data_o[1343] = (N3)? mem[1343] : 
                          (N0)? mem[2943] : 1'b0;
  assign r_data_o[1342] = (N3)? mem[1342] : 
                          (N0)? mem[2942] : 1'b0;
  assign r_data_o[1341] = (N3)? mem[1341] : 
                          (N0)? mem[2941] : 1'b0;
  assign r_data_o[1340] = (N3)? mem[1340] : 
                          (N0)? mem[2940] : 1'b0;
  assign r_data_o[1339] = (N3)? mem[1339] : 
                          (N0)? mem[2939] : 1'b0;
  assign r_data_o[1338] = (N3)? mem[1338] : 
                          (N0)? mem[2938] : 1'b0;
  assign r_data_o[1337] = (N3)? mem[1337] : 
                          (N0)? mem[2937] : 1'b0;
  assign r_data_o[1336] = (N3)? mem[1336] : 
                          (N0)? mem[2936] : 1'b0;
  assign r_data_o[1335] = (N3)? mem[1335] : 
                          (N0)? mem[2935] : 1'b0;
  assign r_data_o[1334] = (N3)? mem[1334] : 
                          (N0)? mem[2934] : 1'b0;
  assign r_data_o[1333] = (N3)? mem[1333] : 
                          (N0)? mem[2933] : 1'b0;
  assign r_data_o[1332] = (N3)? mem[1332] : 
                          (N0)? mem[2932] : 1'b0;
  assign r_data_o[1331] = (N3)? mem[1331] : 
                          (N0)? mem[2931] : 1'b0;
  assign r_data_o[1330] = (N3)? mem[1330] : 
                          (N0)? mem[2930] : 1'b0;
  assign r_data_o[1329] = (N3)? mem[1329] : 
                          (N0)? mem[2929] : 1'b0;
  assign r_data_o[1328] = (N3)? mem[1328] : 
                          (N0)? mem[2928] : 1'b0;
  assign r_data_o[1327] = (N3)? mem[1327] : 
                          (N0)? mem[2927] : 1'b0;
  assign r_data_o[1326] = (N3)? mem[1326] : 
                          (N0)? mem[2926] : 1'b0;
  assign r_data_o[1325] = (N3)? mem[1325] : 
                          (N0)? mem[2925] : 1'b0;
  assign r_data_o[1324] = (N3)? mem[1324] : 
                          (N0)? mem[2924] : 1'b0;
  assign r_data_o[1323] = (N3)? mem[1323] : 
                          (N0)? mem[2923] : 1'b0;
  assign r_data_o[1322] = (N3)? mem[1322] : 
                          (N0)? mem[2922] : 1'b0;
  assign r_data_o[1321] = (N3)? mem[1321] : 
                          (N0)? mem[2921] : 1'b0;
  assign r_data_o[1320] = (N3)? mem[1320] : 
                          (N0)? mem[2920] : 1'b0;
  assign r_data_o[1319] = (N3)? mem[1319] : 
                          (N0)? mem[2919] : 1'b0;
  assign r_data_o[1318] = (N3)? mem[1318] : 
                          (N0)? mem[2918] : 1'b0;
  assign r_data_o[1317] = (N3)? mem[1317] : 
                          (N0)? mem[2917] : 1'b0;
  assign r_data_o[1316] = (N3)? mem[1316] : 
                          (N0)? mem[2916] : 1'b0;
  assign r_data_o[1315] = (N3)? mem[1315] : 
                          (N0)? mem[2915] : 1'b0;
  assign r_data_o[1314] = (N3)? mem[1314] : 
                          (N0)? mem[2914] : 1'b0;
  assign r_data_o[1313] = (N3)? mem[1313] : 
                          (N0)? mem[2913] : 1'b0;
  assign r_data_o[1312] = (N3)? mem[1312] : 
                          (N0)? mem[2912] : 1'b0;
  assign r_data_o[1311] = (N3)? mem[1311] : 
                          (N0)? mem[2911] : 1'b0;
  assign r_data_o[1310] = (N3)? mem[1310] : 
                          (N0)? mem[2910] : 1'b0;
  assign r_data_o[1309] = (N3)? mem[1309] : 
                          (N0)? mem[2909] : 1'b0;
  assign r_data_o[1308] = (N3)? mem[1308] : 
                          (N0)? mem[2908] : 1'b0;
  assign r_data_o[1307] = (N3)? mem[1307] : 
                          (N0)? mem[2907] : 1'b0;
  assign r_data_o[1306] = (N3)? mem[1306] : 
                          (N0)? mem[2906] : 1'b0;
  assign r_data_o[1305] = (N3)? mem[1305] : 
                          (N0)? mem[2905] : 1'b0;
  assign r_data_o[1304] = (N3)? mem[1304] : 
                          (N0)? mem[2904] : 1'b0;
  assign r_data_o[1303] = (N3)? mem[1303] : 
                          (N0)? mem[2903] : 1'b0;
  assign r_data_o[1302] = (N3)? mem[1302] : 
                          (N0)? mem[2902] : 1'b0;
  assign r_data_o[1301] = (N3)? mem[1301] : 
                          (N0)? mem[2901] : 1'b0;
  assign r_data_o[1300] = (N3)? mem[1300] : 
                          (N0)? mem[2900] : 1'b0;
  assign r_data_o[1299] = (N3)? mem[1299] : 
                          (N0)? mem[2899] : 1'b0;
  assign r_data_o[1298] = (N3)? mem[1298] : 
                          (N0)? mem[2898] : 1'b0;
  assign r_data_o[1297] = (N3)? mem[1297] : 
                          (N0)? mem[2897] : 1'b0;
  assign r_data_o[1296] = (N3)? mem[1296] : 
                          (N0)? mem[2896] : 1'b0;
  assign r_data_o[1295] = (N3)? mem[1295] : 
                          (N0)? mem[2895] : 1'b0;
  assign r_data_o[1294] = (N3)? mem[1294] : 
                          (N0)? mem[2894] : 1'b0;
  assign r_data_o[1293] = (N3)? mem[1293] : 
                          (N0)? mem[2893] : 1'b0;
  assign r_data_o[1292] = (N3)? mem[1292] : 
                          (N0)? mem[2892] : 1'b0;
  assign r_data_o[1291] = (N3)? mem[1291] : 
                          (N0)? mem[2891] : 1'b0;
  assign r_data_o[1290] = (N3)? mem[1290] : 
                          (N0)? mem[2890] : 1'b0;
  assign r_data_o[1289] = (N3)? mem[1289] : 
                          (N0)? mem[2889] : 1'b0;
  assign r_data_o[1288] = (N3)? mem[1288] : 
                          (N0)? mem[2888] : 1'b0;
  assign r_data_o[1287] = (N3)? mem[1287] : 
                          (N0)? mem[2887] : 1'b0;
  assign r_data_o[1286] = (N3)? mem[1286] : 
                          (N0)? mem[2886] : 1'b0;
  assign r_data_o[1285] = (N3)? mem[1285] : 
                          (N0)? mem[2885] : 1'b0;
  assign r_data_o[1284] = (N3)? mem[1284] : 
                          (N0)? mem[2884] : 1'b0;
  assign r_data_o[1283] = (N3)? mem[1283] : 
                          (N0)? mem[2883] : 1'b0;
  assign r_data_o[1282] = (N3)? mem[1282] : 
                          (N0)? mem[2882] : 1'b0;
  assign r_data_o[1281] = (N3)? mem[1281] : 
                          (N0)? mem[2881] : 1'b0;
  assign r_data_o[1280] = (N3)? mem[1280] : 
                          (N0)? mem[2880] : 1'b0;
  assign r_data_o[1279] = (N3)? mem[1279] : 
                          (N0)? mem[2879] : 1'b0;
  assign r_data_o[1278] = (N3)? mem[1278] : 
                          (N0)? mem[2878] : 1'b0;
  assign r_data_o[1277] = (N3)? mem[1277] : 
                          (N0)? mem[2877] : 1'b0;
  assign r_data_o[1276] = (N3)? mem[1276] : 
                          (N0)? mem[2876] : 1'b0;
  assign r_data_o[1275] = (N3)? mem[1275] : 
                          (N0)? mem[2875] : 1'b0;
  assign r_data_o[1274] = (N3)? mem[1274] : 
                          (N0)? mem[2874] : 1'b0;
  assign r_data_o[1273] = (N3)? mem[1273] : 
                          (N0)? mem[2873] : 1'b0;
  assign r_data_o[1272] = (N3)? mem[1272] : 
                          (N0)? mem[2872] : 1'b0;
  assign r_data_o[1271] = (N3)? mem[1271] : 
                          (N0)? mem[2871] : 1'b0;
  assign r_data_o[1270] = (N3)? mem[1270] : 
                          (N0)? mem[2870] : 1'b0;
  assign r_data_o[1269] = (N3)? mem[1269] : 
                          (N0)? mem[2869] : 1'b0;
  assign r_data_o[1268] = (N3)? mem[1268] : 
                          (N0)? mem[2868] : 1'b0;
  assign r_data_o[1267] = (N3)? mem[1267] : 
                          (N0)? mem[2867] : 1'b0;
  assign r_data_o[1266] = (N3)? mem[1266] : 
                          (N0)? mem[2866] : 1'b0;
  assign r_data_o[1265] = (N3)? mem[1265] : 
                          (N0)? mem[2865] : 1'b0;
  assign r_data_o[1264] = (N3)? mem[1264] : 
                          (N0)? mem[2864] : 1'b0;
  assign r_data_o[1263] = (N3)? mem[1263] : 
                          (N0)? mem[2863] : 1'b0;
  assign r_data_o[1262] = (N3)? mem[1262] : 
                          (N0)? mem[2862] : 1'b0;
  assign r_data_o[1261] = (N3)? mem[1261] : 
                          (N0)? mem[2861] : 1'b0;
  assign r_data_o[1260] = (N3)? mem[1260] : 
                          (N0)? mem[2860] : 1'b0;
  assign r_data_o[1259] = (N3)? mem[1259] : 
                          (N0)? mem[2859] : 1'b0;
  assign r_data_o[1258] = (N3)? mem[1258] : 
                          (N0)? mem[2858] : 1'b0;
  assign r_data_o[1257] = (N3)? mem[1257] : 
                          (N0)? mem[2857] : 1'b0;
  assign r_data_o[1256] = (N3)? mem[1256] : 
                          (N0)? mem[2856] : 1'b0;
  assign r_data_o[1255] = (N3)? mem[1255] : 
                          (N0)? mem[2855] : 1'b0;
  assign r_data_o[1254] = (N3)? mem[1254] : 
                          (N0)? mem[2854] : 1'b0;
  assign r_data_o[1253] = (N3)? mem[1253] : 
                          (N0)? mem[2853] : 1'b0;
  assign r_data_o[1252] = (N3)? mem[1252] : 
                          (N0)? mem[2852] : 1'b0;
  assign r_data_o[1251] = (N3)? mem[1251] : 
                          (N0)? mem[2851] : 1'b0;
  assign r_data_o[1250] = (N3)? mem[1250] : 
                          (N0)? mem[2850] : 1'b0;
  assign r_data_o[1249] = (N3)? mem[1249] : 
                          (N0)? mem[2849] : 1'b0;
  assign r_data_o[1248] = (N3)? mem[1248] : 
                          (N0)? mem[2848] : 1'b0;
  assign r_data_o[1247] = (N3)? mem[1247] : 
                          (N0)? mem[2847] : 1'b0;
  assign r_data_o[1246] = (N3)? mem[1246] : 
                          (N0)? mem[2846] : 1'b0;
  assign r_data_o[1245] = (N3)? mem[1245] : 
                          (N0)? mem[2845] : 1'b0;
  assign r_data_o[1244] = (N3)? mem[1244] : 
                          (N0)? mem[2844] : 1'b0;
  assign r_data_o[1243] = (N3)? mem[1243] : 
                          (N0)? mem[2843] : 1'b0;
  assign r_data_o[1242] = (N3)? mem[1242] : 
                          (N0)? mem[2842] : 1'b0;
  assign r_data_o[1241] = (N3)? mem[1241] : 
                          (N0)? mem[2841] : 1'b0;
  assign r_data_o[1240] = (N3)? mem[1240] : 
                          (N0)? mem[2840] : 1'b0;
  assign r_data_o[1239] = (N3)? mem[1239] : 
                          (N0)? mem[2839] : 1'b0;
  assign r_data_o[1238] = (N3)? mem[1238] : 
                          (N0)? mem[2838] : 1'b0;
  assign r_data_o[1237] = (N3)? mem[1237] : 
                          (N0)? mem[2837] : 1'b0;
  assign r_data_o[1236] = (N3)? mem[1236] : 
                          (N0)? mem[2836] : 1'b0;
  assign r_data_o[1235] = (N3)? mem[1235] : 
                          (N0)? mem[2835] : 1'b0;
  assign r_data_o[1234] = (N3)? mem[1234] : 
                          (N0)? mem[2834] : 1'b0;
  assign r_data_o[1233] = (N3)? mem[1233] : 
                          (N0)? mem[2833] : 1'b0;
  assign r_data_o[1232] = (N3)? mem[1232] : 
                          (N0)? mem[2832] : 1'b0;
  assign r_data_o[1231] = (N3)? mem[1231] : 
                          (N0)? mem[2831] : 1'b0;
  assign r_data_o[1230] = (N3)? mem[1230] : 
                          (N0)? mem[2830] : 1'b0;
  assign r_data_o[1229] = (N3)? mem[1229] : 
                          (N0)? mem[2829] : 1'b0;
  assign r_data_o[1228] = (N3)? mem[1228] : 
                          (N0)? mem[2828] : 1'b0;
  assign r_data_o[1227] = (N3)? mem[1227] : 
                          (N0)? mem[2827] : 1'b0;
  assign r_data_o[1226] = (N3)? mem[1226] : 
                          (N0)? mem[2826] : 1'b0;
  assign r_data_o[1225] = (N3)? mem[1225] : 
                          (N0)? mem[2825] : 1'b0;
  assign r_data_o[1224] = (N3)? mem[1224] : 
                          (N0)? mem[2824] : 1'b0;
  assign r_data_o[1223] = (N3)? mem[1223] : 
                          (N0)? mem[2823] : 1'b0;
  assign r_data_o[1222] = (N3)? mem[1222] : 
                          (N0)? mem[2822] : 1'b0;
  assign r_data_o[1221] = (N3)? mem[1221] : 
                          (N0)? mem[2821] : 1'b0;
  assign r_data_o[1220] = (N3)? mem[1220] : 
                          (N0)? mem[2820] : 1'b0;
  assign r_data_o[1219] = (N3)? mem[1219] : 
                          (N0)? mem[2819] : 1'b0;
  assign r_data_o[1218] = (N3)? mem[1218] : 
                          (N0)? mem[2818] : 1'b0;
  assign r_data_o[1217] = (N3)? mem[1217] : 
                          (N0)? mem[2817] : 1'b0;
  assign r_data_o[1216] = (N3)? mem[1216] : 
                          (N0)? mem[2816] : 1'b0;
  assign r_data_o[1215] = (N3)? mem[1215] : 
                          (N0)? mem[2815] : 1'b0;
  assign r_data_o[1214] = (N3)? mem[1214] : 
                          (N0)? mem[2814] : 1'b0;
  assign r_data_o[1213] = (N3)? mem[1213] : 
                          (N0)? mem[2813] : 1'b0;
  assign r_data_o[1212] = (N3)? mem[1212] : 
                          (N0)? mem[2812] : 1'b0;
  assign r_data_o[1211] = (N3)? mem[1211] : 
                          (N0)? mem[2811] : 1'b0;
  assign r_data_o[1210] = (N3)? mem[1210] : 
                          (N0)? mem[2810] : 1'b0;
  assign r_data_o[1209] = (N3)? mem[1209] : 
                          (N0)? mem[2809] : 1'b0;
  assign r_data_o[1208] = (N3)? mem[1208] : 
                          (N0)? mem[2808] : 1'b0;
  assign r_data_o[1207] = (N3)? mem[1207] : 
                          (N0)? mem[2807] : 1'b0;
  assign r_data_o[1206] = (N3)? mem[1206] : 
                          (N0)? mem[2806] : 1'b0;
  assign r_data_o[1205] = (N3)? mem[1205] : 
                          (N0)? mem[2805] : 1'b0;
  assign r_data_o[1204] = (N3)? mem[1204] : 
                          (N0)? mem[2804] : 1'b0;
  assign r_data_o[1203] = (N3)? mem[1203] : 
                          (N0)? mem[2803] : 1'b0;
  assign r_data_o[1202] = (N3)? mem[1202] : 
                          (N0)? mem[2802] : 1'b0;
  assign r_data_o[1201] = (N3)? mem[1201] : 
                          (N0)? mem[2801] : 1'b0;
  assign r_data_o[1200] = (N3)? mem[1200] : 
                          (N0)? mem[2800] : 1'b0;
  assign r_data_o[1199] = (N3)? mem[1199] : 
                          (N0)? mem[2799] : 1'b0;
  assign r_data_o[1198] = (N3)? mem[1198] : 
                          (N0)? mem[2798] : 1'b0;
  assign r_data_o[1197] = (N3)? mem[1197] : 
                          (N0)? mem[2797] : 1'b0;
  assign r_data_o[1196] = (N3)? mem[1196] : 
                          (N0)? mem[2796] : 1'b0;
  assign r_data_o[1195] = (N3)? mem[1195] : 
                          (N0)? mem[2795] : 1'b0;
  assign r_data_o[1194] = (N3)? mem[1194] : 
                          (N0)? mem[2794] : 1'b0;
  assign r_data_o[1193] = (N3)? mem[1193] : 
                          (N0)? mem[2793] : 1'b0;
  assign r_data_o[1192] = (N3)? mem[1192] : 
                          (N0)? mem[2792] : 1'b0;
  assign r_data_o[1191] = (N3)? mem[1191] : 
                          (N0)? mem[2791] : 1'b0;
  assign r_data_o[1190] = (N3)? mem[1190] : 
                          (N0)? mem[2790] : 1'b0;
  assign r_data_o[1189] = (N3)? mem[1189] : 
                          (N0)? mem[2789] : 1'b0;
  assign r_data_o[1188] = (N3)? mem[1188] : 
                          (N0)? mem[2788] : 1'b0;
  assign r_data_o[1187] = (N3)? mem[1187] : 
                          (N0)? mem[2787] : 1'b0;
  assign r_data_o[1186] = (N3)? mem[1186] : 
                          (N0)? mem[2786] : 1'b0;
  assign r_data_o[1185] = (N3)? mem[1185] : 
                          (N0)? mem[2785] : 1'b0;
  assign r_data_o[1184] = (N3)? mem[1184] : 
                          (N0)? mem[2784] : 1'b0;
  assign r_data_o[1183] = (N3)? mem[1183] : 
                          (N0)? mem[2783] : 1'b0;
  assign r_data_o[1182] = (N3)? mem[1182] : 
                          (N0)? mem[2782] : 1'b0;
  assign r_data_o[1181] = (N3)? mem[1181] : 
                          (N0)? mem[2781] : 1'b0;
  assign r_data_o[1180] = (N3)? mem[1180] : 
                          (N0)? mem[2780] : 1'b0;
  assign r_data_o[1179] = (N3)? mem[1179] : 
                          (N0)? mem[2779] : 1'b0;
  assign r_data_o[1178] = (N3)? mem[1178] : 
                          (N0)? mem[2778] : 1'b0;
  assign r_data_o[1177] = (N3)? mem[1177] : 
                          (N0)? mem[2777] : 1'b0;
  assign r_data_o[1176] = (N3)? mem[1176] : 
                          (N0)? mem[2776] : 1'b0;
  assign r_data_o[1175] = (N3)? mem[1175] : 
                          (N0)? mem[2775] : 1'b0;
  assign r_data_o[1174] = (N3)? mem[1174] : 
                          (N0)? mem[2774] : 1'b0;
  assign r_data_o[1173] = (N3)? mem[1173] : 
                          (N0)? mem[2773] : 1'b0;
  assign r_data_o[1172] = (N3)? mem[1172] : 
                          (N0)? mem[2772] : 1'b0;
  assign r_data_o[1171] = (N3)? mem[1171] : 
                          (N0)? mem[2771] : 1'b0;
  assign r_data_o[1170] = (N3)? mem[1170] : 
                          (N0)? mem[2770] : 1'b0;
  assign r_data_o[1169] = (N3)? mem[1169] : 
                          (N0)? mem[2769] : 1'b0;
  assign r_data_o[1168] = (N3)? mem[1168] : 
                          (N0)? mem[2768] : 1'b0;
  assign r_data_o[1167] = (N3)? mem[1167] : 
                          (N0)? mem[2767] : 1'b0;
  assign r_data_o[1166] = (N3)? mem[1166] : 
                          (N0)? mem[2766] : 1'b0;
  assign r_data_o[1165] = (N3)? mem[1165] : 
                          (N0)? mem[2765] : 1'b0;
  assign r_data_o[1164] = (N3)? mem[1164] : 
                          (N0)? mem[2764] : 1'b0;
  assign r_data_o[1163] = (N3)? mem[1163] : 
                          (N0)? mem[2763] : 1'b0;
  assign r_data_o[1162] = (N3)? mem[1162] : 
                          (N0)? mem[2762] : 1'b0;
  assign r_data_o[1161] = (N3)? mem[1161] : 
                          (N0)? mem[2761] : 1'b0;
  assign r_data_o[1160] = (N3)? mem[1160] : 
                          (N0)? mem[2760] : 1'b0;
  assign r_data_o[1159] = (N3)? mem[1159] : 
                          (N0)? mem[2759] : 1'b0;
  assign r_data_o[1158] = (N3)? mem[1158] : 
                          (N0)? mem[2758] : 1'b0;
  assign r_data_o[1157] = (N3)? mem[1157] : 
                          (N0)? mem[2757] : 1'b0;
  assign r_data_o[1156] = (N3)? mem[1156] : 
                          (N0)? mem[2756] : 1'b0;
  assign r_data_o[1155] = (N3)? mem[1155] : 
                          (N0)? mem[2755] : 1'b0;
  assign r_data_o[1154] = (N3)? mem[1154] : 
                          (N0)? mem[2754] : 1'b0;
  assign r_data_o[1153] = (N3)? mem[1153] : 
                          (N0)? mem[2753] : 1'b0;
  assign r_data_o[1152] = (N3)? mem[1152] : 
                          (N0)? mem[2752] : 1'b0;
  assign r_data_o[1151] = (N3)? mem[1151] : 
                          (N0)? mem[2751] : 1'b0;
  assign r_data_o[1150] = (N3)? mem[1150] : 
                          (N0)? mem[2750] : 1'b0;
  assign r_data_o[1149] = (N3)? mem[1149] : 
                          (N0)? mem[2749] : 1'b0;
  assign r_data_o[1148] = (N3)? mem[1148] : 
                          (N0)? mem[2748] : 1'b0;
  assign r_data_o[1147] = (N3)? mem[1147] : 
                          (N0)? mem[2747] : 1'b0;
  assign r_data_o[1146] = (N3)? mem[1146] : 
                          (N0)? mem[2746] : 1'b0;
  assign r_data_o[1145] = (N3)? mem[1145] : 
                          (N0)? mem[2745] : 1'b0;
  assign r_data_o[1144] = (N3)? mem[1144] : 
                          (N0)? mem[2744] : 1'b0;
  assign r_data_o[1143] = (N3)? mem[1143] : 
                          (N0)? mem[2743] : 1'b0;
  assign r_data_o[1142] = (N3)? mem[1142] : 
                          (N0)? mem[2742] : 1'b0;
  assign r_data_o[1141] = (N3)? mem[1141] : 
                          (N0)? mem[2741] : 1'b0;
  assign r_data_o[1140] = (N3)? mem[1140] : 
                          (N0)? mem[2740] : 1'b0;
  assign r_data_o[1139] = (N3)? mem[1139] : 
                          (N0)? mem[2739] : 1'b0;
  assign r_data_o[1138] = (N3)? mem[1138] : 
                          (N0)? mem[2738] : 1'b0;
  assign r_data_o[1137] = (N3)? mem[1137] : 
                          (N0)? mem[2737] : 1'b0;
  assign r_data_o[1136] = (N3)? mem[1136] : 
                          (N0)? mem[2736] : 1'b0;
  assign r_data_o[1135] = (N3)? mem[1135] : 
                          (N0)? mem[2735] : 1'b0;
  assign r_data_o[1134] = (N3)? mem[1134] : 
                          (N0)? mem[2734] : 1'b0;
  assign r_data_o[1133] = (N3)? mem[1133] : 
                          (N0)? mem[2733] : 1'b0;
  assign r_data_o[1132] = (N3)? mem[1132] : 
                          (N0)? mem[2732] : 1'b0;
  assign r_data_o[1131] = (N3)? mem[1131] : 
                          (N0)? mem[2731] : 1'b0;
  assign r_data_o[1130] = (N3)? mem[1130] : 
                          (N0)? mem[2730] : 1'b0;
  assign r_data_o[1129] = (N3)? mem[1129] : 
                          (N0)? mem[2729] : 1'b0;
  assign r_data_o[1128] = (N3)? mem[1128] : 
                          (N0)? mem[2728] : 1'b0;
  assign r_data_o[1127] = (N3)? mem[1127] : 
                          (N0)? mem[2727] : 1'b0;
  assign r_data_o[1126] = (N3)? mem[1126] : 
                          (N0)? mem[2726] : 1'b0;
  assign r_data_o[1125] = (N3)? mem[1125] : 
                          (N0)? mem[2725] : 1'b0;
  assign r_data_o[1124] = (N3)? mem[1124] : 
                          (N0)? mem[2724] : 1'b0;
  assign r_data_o[1123] = (N3)? mem[1123] : 
                          (N0)? mem[2723] : 1'b0;
  assign r_data_o[1122] = (N3)? mem[1122] : 
                          (N0)? mem[2722] : 1'b0;
  assign r_data_o[1121] = (N3)? mem[1121] : 
                          (N0)? mem[2721] : 1'b0;
  assign r_data_o[1120] = (N3)? mem[1120] : 
                          (N0)? mem[2720] : 1'b0;
  assign r_data_o[1119] = (N3)? mem[1119] : 
                          (N0)? mem[2719] : 1'b0;
  assign r_data_o[1118] = (N3)? mem[1118] : 
                          (N0)? mem[2718] : 1'b0;
  assign r_data_o[1117] = (N3)? mem[1117] : 
                          (N0)? mem[2717] : 1'b0;
  assign r_data_o[1116] = (N3)? mem[1116] : 
                          (N0)? mem[2716] : 1'b0;
  assign r_data_o[1115] = (N3)? mem[1115] : 
                          (N0)? mem[2715] : 1'b0;
  assign r_data_o[1114] = (N3)? mem[1114] : 
                          (N0)? mem[2714] : 1'b0;
  assign r_data_o[1113] = (N3)? mem[1113] : 
                          (N0)? mem[2713] : 1'b0;
  assign r_data_o[1112] = (N3)? mem[1112] : 
                          (N0)? mem[2712] : 1'b0;
  assign r_data_o[1111] = (N3)? mem[1111] : 
                          (N0)? mem[2711] : 1'b0;
  assign r_data_o[1110] = (N3)? mem[1110] : 
                          (N0)? mem[2710] : 1'b0;
  assign r_data_o[1109] = (N3)? mem[1109] : 
                          (N0)? mem[2709] : 1'b0;
  assign r_data_o[1108] = (N3)? mem[1108] : 
                          (N0)? mem[2708] : 1'b0;
  assign r_data_o[1107] = (N3)? mem[1107] : 
                          (N0)? mem[2707] : 1'b0;
  assign r_data_o[1106] = (N3)? mem[1106] : 
                          (N0)? mem[2706] : 1'b0;
  assign r_data_o[1105] = (N3)? mem[1105] : 
                          (N0)? mem[2705] : 1'b0;
  assign r_data_o[1104] = (N3)? mem[1104] : 
                          (N0)? mem[2704] : 1'b0;
  assign r_data_o[1103] = (N3)? mem[1103] : 
                          (N0)? mem[2703] : 1'b0;
  assign r_data_o[1102] = (N3)? mem[1102] : 
                          (N0)? mem[2702] : 1'b0;
  assign r_data_o[1101] = (N3)? mem[1101] : 
                          (N0)? mem[2701] : 1'b0;
  assign r_data_o[1100] = (N3)? mem[1100] : 
                          (N0)? mem[2700] : 1'b0;
  assign r_data_o[1099] = (N3)? mem[1099] : 
                          (N0)? mem[2699] : 1'b0;
  assign r_data_o[1098] = (N3)? mem[1098] : 
                          (N0)? mem[2698] : 1'b0;
  assign r_data_o[1097] = (N3)? mem[1097] : 
                          (N0)? mem[2697] : 1'b0;
  assign r_data_o[1096] = (N3)? mem[1096] : 
                          (N0)? mem[2696] : 1'b0;
  assign r_data_o[1095] = (N3)? mem[1095] : 
                          (N0)? mem[2695] : 1'b0;
  assign r_data_o[1094] = (N3)? mem[1094] : 
                          (N0)? mem[2694] : 1'b0;
  assign r_data_o[1093] = (N3)? mem[1093] : 
                          (N0)? mem[2693] : 1'b0;
  assign r_data_o[1092] = (N3)? mem[1092] : 
                          (N0)? mem[2692] : 1'b0;
  assign r_data_o[1091] = (N3)? mem[1091] : 
                          (N0)? mem[2691] : 1'b0;
  assign r_data_o[1090] = (N3)? mem[1090] : 
                          (N0)? mem[2690] : 1'b0;
  assign r_data_o[1089] = (N3)? mem[1089] : 
                          (N0)? mem[2689] : 1'b0;
  assign r_data_o[1088] = (N3)? mem[1088] : 
                          (N0)? mem[2688] : 1'b0;
  assign r_data_o[1087] = (N3)? mem[1087] : 
                          (N0)? mem[2687] : 1'b0;
  assign r_data_o[1086] = (N3)? mem[1086] : 
                          (N0)? mem[2686] : 1'b0;
  assign r_data_o[1085] = (N3)? mem[1085] : 
                          (N0)? mem[2685] : 1'b0;
  assign r_data_o[1084] = (N3)? mem[1084] : 
                          (N0)? mem[2684] : 1'b0;
  assign r_data_o[1083] = (N3)? mem[1083] : 
                          (N0)? mem[2683] : 1'b0;
  assign r_data_o[1082] = (N3)? mem[1082] : 
                          (N0)? mem[2682] : 1'b0;
  assign r_data_o[1081] = (N3)? mem[1081] : 
                          (N0)? mem[2681] : 1'b0;
  assign r_data_o[1080] = (N3)? mem[1080] : 
                          (N0)? mem[2680] : 1'b0;
  assign r_data_o[1079] = (N3)? mem[1079] : 
                          (N0)? mem[2679] : 1'b0;
  assign r_data_o[1078] = (N3)? mem[1078] : 
                          (N0)? mem[2678] : 1'b0;
  assign r_data_o[1077] = (N3)? mem[1077] : 
                          (N0)? mem[2677] : 1'b0;
  assign r_data_o[1076] = (N3)? mem[1076] : 
                          (N0)? mem[2676] : 1'b0;
  assign r_data_o[1075] = (N3)? mem[1075] : 
                          (N0)? mem[2675] : 1'b0;
  assign r_data_o[1074] = (N3)? mem[1074] : 
                          (N0)? mem[2674] : 1'b0;
  assign r_data_o[1073] = (N3)? mem[1073] : 
                          (N0)? mem[2673] : 1'b0;
  assign r_data_o[1072] = (N3)? mem[1072] : 
                          (N0)? mem[2672] : 1'b0;
  assign r_data_o[1071] = (N3)? mem[1071] : 
                          (N0)? mem[2671] : 1'b0;
  assign r_data_o[1070] = (N3)? mem[1070] : 
                          (N0)? mem[2670] : 1'b0;
  assign r_data_o[1069] = (N3)? mem[1069] : 
                          (N0)? mem[2669] : 1'b0;
  assign r_data_o[1068] = (N3)? mem[1068] : 
                          (N0)? mem[2668] : 1'b0;
  assign r_data_o[1067] = (N3)? mem[1067] : 
                          (N0)? mem[2667] : 1'b0;
  assign r_data_o[1066] = (N3)? mem[1066] : 
                          (N0)? mem[2666] : 1'b0;
  assign r_data_o[1065] = (N3)? mem[1065] : 
                          (N0)? mem[2665] : 1'b0;
  assign r_data_o[1064] = (N3)? mem[1064] : 
                          (N0)? mem[2664] : 1'b0;
  assign r_data_o[1063] = (N3)? mem[1063] : 
                          (N0)? mem[2663] : 1'b0;
  assign r_data_o[1062] = (N3)? mem[1062] : 
                          (N0)? mem[2662] : 1'b0;
  assign r_data_o[1061] = (N3)? mem[1061] : 
                          (N0)? mem[2661] : 1'b0;
  assign r_data_o[1060] = (N3)? mem[1060] : 
                          (N0)? mem[2660] : 1'b0;
  assign r_data_o[1059] = (N3)? mem[1059] : 
                          (N0)? mem[2659] : 1'b0;
  assign r_data_o[1058] = (N3)? mem[1058] : 
                          (N0)? mem[2658] : 1'b0;
  assign r_data_o[1057] = (N3)? mem[1057] : 
                          (N0)? mem[2657] : 1'b0;
  assign r_data_o[1056] = (N3)? mem[1056] : 
                          (N0)? mem[2656] : 1'b0;
  assign r_data_o[1055] = (N3)? mem[1055] : 
                          (N0)? mem[2655] : 1'b0;
  assign r_data_o[1054] = (N3)? mem[1054] : 
                          (N0)? mem[2654] : 1'b0;
  assign r_data_o[1053] = (N3)? mem[1053] : 
                          (N0)? mem[2653] : 1'b0;
  assign r_data_o[1052] = (N3)? mem[1052] : 
                          (N0)? mem[2652] : 1'b0;
  assign r_data_o[1051] = (N3)? mem[1051] : 
                          (N0)? mem[2651] : 1'b0;
  assign r_data_o[1050] = (N3)? mem[1050] : 
                          (N0)? mem[2650] : 1'b0;
  assign r_data_o[1049] = (N3)? mem[1049] : 
                          (N0)? mem[2649] : 1'b0;
  assign r_data_o[1048] = (N3)? mem[1048] : 
                          (N0)? mem[2648] : 1'b0;
  assign r_data_o[1047] = (N3)? mem[1047] : 
                          (N0)? mem[2647] : 1'b0;
  assign r_data_o[1046] = (N3)? mem[1046] : 
                          (N0)? mem[2646] : 1'b0;
  assign r_data_o[1045] = (N3)? mem[1045] : 
                          (N0)? mem[2645] : 1'b0;
  assign r_data_o[1044] = (N3)? mem[1044] : 
                          (N0)? mem[2644] : 1'b0;
  assign r_data_o[1043] = (N3)? mem[1043] : 
                          (N0)? mem[2643] : 1'b0;
  assign r_data_o[1042] = (N3)? mem[1042] : 
                          (N0)? mem[2642] : 1'b0;
  assign r_data_o[1041] = (N3)? mem[1041] : 
                          (N0)? mem[2641] : 1'b0;
  assign r_data_o[1040] = (N3)? mem[1040] : 
                          (N0)? mem[2640] : 1'b0;
  assign r_data_o[1039] = (N3)? mem[1039] : 
                          (N0)? mem[2639] : 1'b0;
  assign r_data_o[1038] = (N3)? mem[1038] : 
                          (N0)? mem[2638] : 1'b0;
  assign r_data_o[1037] = (N3)? mem[1037] : 
                          (N0)? mem[2637] : 1'b0;
  assign r_data_o[1036] = (N3)? mem[1036] : 
                          (N0)? mem[2636] : 1'b0;
  assign r_data_o[1035] = (N3)? mem[1035] : 
                          (N0)? mem[2635] : 1'b0;
  assign r_data_o[1034] = (N3)? mem[1034] : 
                          (N0)? mem[2634] : 1'b0;
  assign r_data_o[1033] = (N3)? mem[1033] : 
                          (N0)? mem[2633] : 1'b0;
  assign r_data_o[1032] = (N3)? mem[1032] : 
                          (N0)? mem[2632] : 1'b0;
  assign r_data_o[1031] = (N3)? mem[1031] : 
                          (N0)? mem[2631] : 1'b0;
  assign r_data_o[1030] = (N3)? mem[1030] : 
                          (N0)? mem[2630] : 1'b0;
  assign r_data_o[1029] = (N3)? mem[1029] : 
                          (N0)? mem[2629] : 1'b0;
  assign r_data_o[1028] = (N3)? mem[1028] : 
                          (N0)? mem[2628] : 1'b0;
  assign r_data_o[1027] = (N3)? mem[1027] : 
                          (N0)? mem[2627] : 1'b0;
  assign r_data_o[1026] = (N3)? mem[1026] : 
                          (N0)? mem[2626] : 1'b0;
  assign r_data_o[1025] = (N3)? mem[1025] : 
                          (N0)? mem[2625] : 1'b0;
  assign r_data_o[1024] = (N3)? mem[1024] : 
                          (N0)? mem[2624] : 1'b0;
  assign r_data_o[1023] = (N3)? mem[1023] : 
                          (N0)? mem[2623] : 1'b0;
  assign r_data_o[1022] = (N3)? mem[1022] : 
                          (N0)? mem[2622] : 1'b0;
  assign r_data_o[1021] = (N3)? mem[1021] : 
                          (N0)? mem[2621] : 1'b0;
  assign r_data_o[1020] = (N3)? mem[1020] : 
                          (N0)? mem[2620] : 1'b0;
  assign r_data_o[1019] = (N3)? mem[1019] : 
                          (N0)? mem[2619] : 1'b0;
  assign r_data_o[1018] = (N3)? mem[1018] : 
                          (N0)? mem[2618] : 1'b0;
  assign r_data_o[1017] = (N3)? mem[1017] : 
                          (N0)? mem[2617] : 1'b0;
  assign r_data_o[1016] = (N3)? mem[1016] : 
                          (N0)? mem[2616] : 1'b0;
  assign r_data_o[1015] = (N3)? mem[1015] : 
                          (N0)? mem[2615] : 1'b0;
  assign r_data_o[1014] = (N3)? mem[1014] : 
                          (N0)? mem[2614] : 1'b0;
  assign r_data_o[1013] = (N3)? mem[1013] : 
                          (N0)? mem[2613] : 1'b0;
  assign r_data_o[1012] = (N3)? mem[1012] : 
                          (N0)? mem[2612] : 1'b0;
  assign r_data_o[1011] = (N3)? mem[1011] : 
                          (N0)? mem[2611] : 1'b0;
  assign r_data_o[1010] = (N3)? mem[1010] : 
                          (N0)? mem[2610] : 1'b0;
  assign r_data_o[1009] = (N3)? mem[1009] : 
                          (N0)? mem[2609] : 1'b0;
  assign r_data_o[1008] = (N3)? mem[1008] : 
                          (N0)? mem[2608] : 1'b0;
  assign r_data_o[1007] = (N3)? mem[1007] : 
                          (N0)? mem[2607] : 1'b0;
  assign r_data_o[1006] = (N3)? mem[1006] : 
                          (N0)? mem[2606] : 1'b0;
  assign r_data_o[1005] = (N3)? mem[1005] : 
                          (N0)? mem[2605] : 1'b0;
  assign r_data_o[1004] = (N3)? mem[1004] : 
                          (N0)? mem[2604] : 1'b0;
  assign r_data_o[1003] = (N3)? mem[1003] : 
                          (N0)? mem[2603] : 1'b0;
  assign r_data_o[1002] = (N3)? mem[1002] : 
                          (N0)? mem[2602] : 1'b0;
  assign r_data_o[1001] = (N3)? mem[1001] : 
                          (N0)? mem[2601] : 1'b0;
  assign r_data_o[1000] = (N3)? mem[1000] : 
                          (N0)? mem[2600] : 1'b0;
  assign r_data_o[999] = (N3)? mem[999] : 
                         (N0)? mem[2599] : 1'b0;
  assign r_data_o[998] = (N3)? mem[998] : 
                         (N0)? mem[2598] : 1'b0;
  assign r_data_o[997] = (N3)? mem[997] : 
                         (N0)? mem[2597] : 1'b0;
  assign r_data_o[996] = (N3)? mem[996] : 
                         (N0)? mem[2596] : 1'b0;
  assign r_data_o[995] = (N3)? mem[995] : 
                         (N0)? mem[2595] : 1'b0;
  assign r_data_o[994] = (N3)? mem[994] : 
                         (N0)? mem[2594] : 1'b0;
  assign r_data_o[993] = (N3)? mem[993] : 
                         (N0)? mem[2593] : 1'b0;
  assign r_data_o[992] = (N3)? mem[992] : 
                         (N0)? mem[2592] : 1'b0;
  assign r_data_o[991] = (N3)? mem[991] : 
                         (N0)? mem[2591] : 1'b0;
  assign r_data_o[990] = (N3)? mem[990] : 
                         (N0)? mem[2590] : 1'b0;
  assign r_data_o[989] = (N3)? mem[989] : 
                         (N0)? mem[2589] : 1'b0;
  assign r_data_o[988] = (N3)? mem[988] : 
                         (N0)? mem[2588] : 1'b0;
  assign r_data_o[987] = (N3)? mem[987] : 
                         (N0)? mem[2587] : 1'b0;
  assign r_data_o[986] = (N3)? mem[986] : 
                         (N0)? mem[2586] : 1'b0;
  assign r_data_o[985] = (N3)? mem[985] : 
                         (N0)? mem[2585] : 1'b0;
  assign r_data_o[984] = (N3)? mem[984] : 
                         (N0)? mem[2584] : 1'b0;
  assign r_data_o[983] = (N3)? mem[983] : 
                         (N0)? mem[2583] : 1'b0;
  assign r_data_o[982] = (N3)? mem[982] : 
                         (N0)? mem[2582] : 1'b0;
  assign r_data_o[981] = (N3)? mem[981] : 
                         (N0)? mem[2581] : 1'b0;
  assign r_data_o[980] = (N3)? mem[980] : 
                         (N0)? mem[2580] : 1'b0;
  assign r_data_o[979] = (N3)? mem[979] : 
                         (N0)? mem[2579] : 1'b0;
  assign r_data_o[978] = (N3)? mem[978] : 
                         (N0)? mem[2578] : 1'b0;
  assign r_data_o[977] = (N3)? mem[977] : 
                         (N0)? mem[2577] : 1'b0;
  assign r_data_o[976] = (N3)? mem[976] : 
                         (N0)? mem[2576] : 1'b0;
  assign r_data_o[975] = (N3)? mem[975] : 
                         (N0)? mem[2575] : 1'b0;
  assign r_data_o[974] = (N3)? mem[974] : 
                         (N0)? mem[2574] : 1'b0;
  assign r_data_o[973] = (N3)? mem[973] : 
                         (N0)? mem[2573] : 1'b0;
  assign r_data_o[972] = (N3)? mem[972] : 
                         (N0)? mem[2572] : 1'b0;
  assign r_data_o[971] = (N3)? mem[971] : 
                         (N0)? mem[2571] : 1'b0;
  assign r_data_o[970] = (N3)? mem[970] : 
                         (N0)? mem[2570] : 1'b0;
  assign r_data_o[969] = (N3)? mem[969] : 
                         (N0)? mem[2569] : 1'b0;
  assign r_data_o[968] = (N3)? mem[968] : 
                         (N0)? mem[2568] : 1'b0;
  assign r_data_o[967] = (N3)? mem[967] : 
                         (N0)? mem[2567] : 1'b0;
  assign r_data_o[966] = (N3)? mem[966] : 
                         (N0)? mem[2566] : 1'b0;
  assign r_data_o[965] = (N3)? mem[965] : 
                         (N0)? mem[2565] : 1'b0;
  assign r_data_o[964] = (N3)? mem[964] : 
                         (N0)? mem[2564] : 1'b0;
  assign r_data_o[963] = (N3)? mem[963] : 
                         (N0)? mem[2563] : 1'b0;
  assign r_data_o[962] = (N3)? mem[962] : 
                         (N0)? mem[2562] : 1'b0;
  assign r_data_o[961] = (N3)? mem[961] : 
                         (N0)? mem[2561] : 1'b0;
  assign r_data_o[960] = (N3)? mem[960] : 
                         (N0)? mem[2560] : 1'b0;
  assign r_data_o[959] = (N3)? mem[959] : 
                         (N0)? mem[2559] : 1'b0;
  assign r_data_o[958] = (N3)? mem[958] : 
                         (N0)? mem[2558] : 1'b0;
  assign r_data_o[957] = (N3)? mem[957] : 
                         (N0)? mem[2557] : 1'b0;
  assign r_data_o[956] = (N3)? mem[956] : 
                         (N0)? mem[2556] : 1'b0;
  assign r_data_o[955] = (N3)? mem[955] : 
                         (N0)? mem[2555] : 1'b0;
  assign r_data_o[954] = (N3)? mem[954] : 
                         (N0)? mem[2554] : 1'b0;
  assign r_data_o[953] = (N3)? mem[953] : 
                         (N0)? mem[2553] : 1'b0;
  assign r_data_o[952] = (N3)? mem[952] : 
                         (N0)? mem[2552] : 1'b0;
  assign r_data_o[951] = (N3)? mem[951] : 
                         (N0)? mem[2551] : 1'b0;
  assign r_data_o[950] = (N3)? mem[950] : 
                         (N0)? mem[2550] : 1'b0;
  assign r_data_o[949] = (N3)? mem[949] : 
                         (N0)? mem[2549] : 1'b0;
  assign r_data_o[948] = (N3)? mem[948] : 
                         (N0)? mem[2548] : 1'b0;
  assign r_data_o[947] = (N3)? mem[947] : 
                         (N0)? mem[2547] : 1'b0;
  assign r_data_o[946] = (N3)? mem[946] : 
                         (N0)? mem[2546] : 1'b0;
  assign r_data_o[945] = (N3)? mem[945] : 
                         (N0)? mem[2545] : 1'b0;
  assign r_data_o[944] = (N3)? mem[944] : 
                         (N0)? mem[2544] : 1'b0;
  assign r_data_o[943] = (N3)? mem[943] : 
                         (N0)? mem[2543] : 1'b0;
  assign r_data_o[942] = (N3)? mem[942] : 
                         (N0)? mem[2542] : 1'b0;
  assign r_data_o[941] = (N3)? mem[941] : 
                         (N0)? mem[2541] : 1'b0;
  assign r_data_o[940] = (N3)? mem[940] : 
                         (N0)? mem[2540] : 1'b0;
  assign r_data_o[939] = (N3)? mem[939] : 
                         (N0)? mem[2539] : 1'b0;
  assign r_data_o[938] = (N3)? mem[938] : 
                         (N0)? mem[2538] : 1'b0;
  assign r_data_o[937] = (N3)? mem[937] : 
                         (N0)? mem[2537] : 1'b0;
  assign r_data_o[936] = (N3)? mem[936] : 
                         (N0)? mem[2536] : 1'b0;
  assign r_data_o[935] = (N3)? mem[935] : 
                         (N0)? mem[2535] : 1'b0;
  assign r_data_o[934] = (N3)? mem[934] : 
                         (N0)? mem[2534] : 1'b0;
  assign r_data_o[933] = (N3)? mem[933] : 
                         (N0)? mem[2533] : 1'b0;
  assign r_data_o[932] = (N3)? mem[932] : 
                         (N0)? mem[2532] : 1'b0;
  assign r_data_o[931] = (N3)? mem[931] : 
                         (N0)? mem[2531] : 1'b0;
  assign r_data_o[930] = (N3)? mem[930] : 
                         (N0)? mem[2530] : 1'b0;
  assign r_data_o[929] = (N3)? mem[929] : 
                         (N0)? mem[2529] : 1'b0;
  assign r_data_o[928] = (N3)? mem[928] : 
                         (N0)? mem[2528] : 1'b0;
  assign r_data_o[927] = (N3)? mem[927] : 
                         (N0)? mem[2527] : 1'b0;
  assign r_data_o[926] = (N3)? mem[926] : 
                         (N0)? mem[2526] : 1'b0;
  assign r_data_o[925] = (N3)? mem[925] : 
                         (N0)? mem[2525] : 1'b0;
  assign r_data_o[924] = (N3)? mem[924] : 
                         (N0)? mem[2524] : 1'b0;
  assign r_data_o[923] = (N3)? mem[923] : 
                         (N0)? mem[2523] : 1'b0;
  assign r_data_o[922] = (N3)? mem[922] : 
                         (N0)? mem[2522] : 1'b0;
  assign r_data_o[921] = (N3)? mem[921] : 
                         (N0)? mem[2521] : 1'b0;
  assign r_data_o[920] = (N3)? mem[920] : 
                         (N0)? mem[2520] : 1'b0;
  assign r_data_o[919] = (N3)? mem[919] : 
                         (N0)? mem[2519] : 1'b0;
  assign r_data_o[918] = (N3)? mem[918] : 
                         (N0)? mem[2518] : 1'b0;
  assign r_data_o[917] = (N3)? mem[917] : 
                         (N0)? mem[2517] : 1'b0;
  assign r_data_o[916] = (N3)? mem[916] : 
                         (N0)? mem[2516] : 1'b0;
  assign r_data_o[915] = (N3)? mem[915] : 
                         (N0)? mem[2515] : 1'b0;
  assign r_data_o[914] = (N3)? mem[914] : 
                         (N0)? mem[2514] : 1'b0;
  assign r_data_o[913] = (N3)? mem[913] : 
                         (N0)? mem[2513] : 1'b0;
  assign r_data_o[912] = (N3)? mem[912] : 
                         (N0)? mem[2512] : 1'b0;
  assign r_data_o[911] = (N3)? mem[911] : 
                         (N0)? mem[2511] : 1'b0;
  assign r_data_o[910] = (N3)? mem[910] : 
                         (N0)? mem[2510] : 1'b0;
  assign r_data_o[909] = (N3)? mem[909] : 
                         (N0)? mem[2509] : 1'b0;
  assign r_data_o[908] = (N3)? mem[908] : 
                         (N0)? mem[2508] : 1'b0;
  assign r_data_o[907] = (N3)? mem[907] : 
                         (N0)? mem[2507] : 1'b0;
  assign r_data_o[906] = (N3)? mem[906] : 
                         (N0)? mem[2506] : 1'b0;
  assign r_data_o[905] = (N3)? mem[905] : 
                         (N0)? mem[2505] : 1'b0;
  assign r_data_o[904] = (N3)? mem[904] : 
                         (N0)? mem[2504] : 1'b0;
  assign r_data_o[903] = (N3)? mem[903] : 
                         (N0)? mem[2503] : 1'b0;
  assign r_data_o[902] = (N3)? mem[902] : 
                         (N0)? mem[2502] : 1'b0;
  assign r_data_o[901] = (N3)? mem[901] : 
                         (N0)? mem[2501] : 1'b0;
  assign r_data_o[900] = (N3)? mem[900] : 
                         (N0)? mem[2500] : 1'b0;
  assign r_data_o[899] = (N3)? mem[899] : 
                         (N0)? mem[2499] : 1'b0;
  assign r_data_o[898] = (N3)? mem[898] : 
                         (N0)? mem[2498] : 1'b0;
  assign r_data_o[897] = (N3)? mem[897] : 
                         (N0)? mem[2497] : 1'b0;
  assign r_data_o[896] = (N3)? mem[896] : 
                         (N0)? mem[2496] : 1'b0;
  assign r_data_o[895] = (N3)? mem[895] : 
                         (N0)? mem[2495] : 1'b0;
  assign r_data_o[894] = (N3)? mem[894] : 
                         (N0)? mem[2494] : 1'b0;
  assign r_data_o[893] = (N3)? mem[893] : 
                         (N0)? mem[2493] : 1'b0;
  assign r_data_o[892] = (N3)? mem[892] : 
                         (N0)? mem[2492] : 1'b0;
  assign r_data_o[891] = (N3)? mem[891] : 
                         (N0)? mem[2491] : 1'b0;
  assign r_data_o[890] = (N3)? mem[890] : 
                         (N0)? mem[2490] : 1'b0;
  assign r_data_o[889] = (N3)? mem[889] : 
                         (N0)? mem[2489] : 1'b0;
  assign r_data_o[888] = (N3)? mem[888] : 
                         (N0)? mem[2488] : 1'b0;
  assign r_data_o[887] = (N3)? mem[887] : 
                         (N0)? mem[2487] : 1'b0;
  assign r_data_o[886] = (N3)? mem[886] : 
                         (N0)? mem[2486] : 1'b0;
  assign r_data_o[885] = (N3)? mem[885] : 
                         (N0)? mem[2485] : 1'b0;
  assign r_data_o[884] = (N3)? mem[884] : 
                         (N0)? mem[2484] : 1'b0;
  assign r_data_o[883] = (N3)? mem[883] : 
                         (N0)? mem[2483] : 1'b0;
  assign r_data_o[882] = (N3)? mem[882] : 
                         (N0)? mem[2482] : 1'b0;
  assign r_data_o[881] = (N3)? mem[881] : 
                         (N0)? mem[2481] : 1'b0;
  assign r_data_o[880] = (N3)? mem[880] : 
                         (N0)? mem[2480] : 1'b0;
  assign r_data_o[879] = (N3)? mem[879] : 
                         (N0)? mem[2479] : 1'b0;
  assign r_data_o[878] = (N3)? mem[878] : 
                         (N0)? mem[2478] : 1'b0;
  assign r_data_o[877] = (N3)? mem[877] : 
                         (N0)? mem[2477] : 1'b0;
  assign r_data_o[876] = (N3)? mem[876] : 
                         (N0)? mem[2476] : 1'b0;
  assign r_data_o[875] = (N3)? mem[875] : 
                         (N0)? mem[2475] : 1'b0;
  assign r_data_o[874] = (N3)? mem[874] : 
                         (N0)? mem[2474] : 1'b0;
  assign r_data_o[873] = (N3)? mem[873] : 
                         (N0)? mem[2473] : 1'b0;
  assign r_data_o[872] = (N3)? mem[872] : 
                         (N0)? mem[2472] : 1'b0;
  assign r_data_o[871] = (N3)? mem[871] : 
                         (N0)? mem[2471] : 1'b0;
  assign r_data_o[870] = (N3)? mem[870] : 
                         (N0)? mem[2470] : 1'b0;
  assign r_data_o[869] = (N3)? mem[869] : 
                         (N0)? mem[2469] : 1'b0;
  assign r_data_o[868] = (N3)? mem[868] : 
                         (N0)? mem[2468] : 1'b0;
  assign r_data_o[867] = (N3)? mem[867] : 
                         (N0)? mem[2467] : 1'b0;
  assign r_data_o[866] = (N3)? mem[866] : 
                         (N0)? mem[2466] : 1'b0;
  assign r_data_o[865] = (N3)? mem[865] : 
                         (N0)? mem[2465] : 1'b0;
  assign r_data_o[864] = (N3)? mem[864] : 
                         (N0)? mem[2464] : 1'b0;
  assign r_data_o[863] = (N3)? mem[863] : 
                         (N0)? mem[2463] : 1'b0;
  assign r_data_o[862] = (N3)? mem[862] : 
                         (N0)? mem[2462] : 1'b0;
  assign r_data_o[861] = (N3)? mem[861] : 
                         (N0)? mem[2461] : 1'b0;
  assign r_data_o[860] = (N3)? mem[860] : 
                         (N0)? mem[2460] : 1'b0;
  assign r_data_o[859] = (N3)? mem[859] : 
                         (N0)? mem[2459] : 1'b0;
  assign r_data_o[858] = (N3)? mem[858] : 
                         (N0)? mem[2458] : 1'b0;
  assign r_data_o[857] = (N3)? mem[857] : 
                         (N0)? mem[2457] : 1'b0;
  assign r_data_o[856] = (N3)? mem[856] : 
                         (N0)? mem[2456] : 1'b0;
  assign r_data_o[855] = (N3)? mem[855] : 
                         (N0)? mem[2455] : 1'b0;
  assign r_data_o[854] = (N3)? mem[854] : 
                         (N0)? mem[2454] : 1'b0;
  assign r_data_o[853] = (N3)? mem[853] : 
                         (N0)? mem[2453] : 1'b0;
  assign r_data_o[852] = (N3)? mem[852] : 
                         (N0)? mem[2452] : 1'b0;
  assign r_data_o[851] = (N3)? mem[851] : 
                         (N0)? mem[2451] : 1'b0;
  assign r_data_o[850] = (N3)? mem[850] : 
                         (N0)? mem[2450] : 1'b0;
  assign r_data_o[849] = (N3)? mem[849] : 
                         (N0)? mem[2449] : 1'b0;
  assign r_data_o[848] = (N3)? mem[848] : 
                         (N0)? mem[2448] : 1'b0;
  assign r_data_o[847] = (N3)? mem[847] : 
                         (N0)? mem[2447] : 1'b0;
  assign r_data_o[846] = (N3)? mem[846] : 
                         (N0)? mem[2446] : 1'b0;
  assign r_data_o[845] = (N3)? mem[845] : 
                         (N0)? mem[2445] : 1'b0;
  assign r_data_o[844] = (N3)? mem[844] : 
                         (N0)? mem[2444] : 1'b0;
  assign r_data_o[843] = (N3)? mem[843] : 
                         (N0)? mem[2443] : 1'b0;
  assign r_data_o[842] = (N3)? mem[842] : 
                         (N0)? mem[2442] : 1'b0;
  assign r_data_o[841] = (N3)? mem[841] : 
                         (N0)? mem[2441] : 1'b0;
  assign r_data_o[840] = (N3)? mem[840] : 
                         (N0)? mem[2440] : 1'b0;
  assign r_data_o[839] = (N3)? mem[839] : 
                         (N0)? mem[2439] : 1'b0;
  assign r_data_o[838] = (N3)? mem[838] : 
                         (N0)? mem[2438] : 1'b0;
  assign r_data_o[837] = (N3)? mem[837] : 
                         (N0)? mem[2437] : 1'b0;
  assign r_data_o[836] = (N3)? mem[836] : 
                         (N0)? mem[2436] : 1'b0;
  assign r_data_o[835] = (N3)? mem[835] : 
                         (N0)? mem[2435] : 1'b0;
  assign r_data_o[834] = (N3)? mem[834] : 
                         (N0)? mem[2434] : 1'b0;
  assign r_data_o[833] = (N3)? mem[833] : 
                         (N0)? mem[2433] : 1'b0;
  assign r_data_o[832] = (N3)? mem[832] : 
                         (N0)? mem[2432] : 1'b0;
  assign r_data_o[831] = (N3)? mem[831] : 
                         (N0)? mem[2431] : 1'b0;
  assign r_data_o[830] = (N3)? mem[830] : 
                         (N0)? mem[2430] : 1'b0;
  assign r_data_o[829] = (N3)? mem[829] : 
                         (N0)? mem[2429] : 1'b0;
  assign r_data_o[828] = (N3)? mem[828] : 
                         (N0)? mem[2428] : 1'b0;
  assign r_data_o[827] = (N3)? mem[827] : 
                         (N0)? mem[2427] : 1'b0;
  assign r_data_o[826] = (N3)? mem[826] : 
                         (N0)? mem[2426] : 1'b0;
  assign r_data_o[825] = (N3)? mem[825] : 
                         (N0)? mem[2425] : 1'b0;
  assign r_data_o[824] = (N3)? mem[824] : 
                         (N0)? mem[2424] : 1'b0;
  assign r_data_o[823] = (N3)? mem[823] : 
                         (N0)? mem[2423] : 1'b0;
  assign r_data_o[822] = (N3)? mem[822] : 
                         (N0)? mem[2422] : 1'b0;
  assign r_data_o[821] = (N3)? mem[821] : 
                         (N0)? mem[2421] : 1'b0;
  assign r_data_o[820] = (N3)? mem[820] : 
                         (N0)? mem[2420] : 1'b0;
  assign r_data_o[819] = (N3)? mem[819] : 
                         (N0)? mem[2419] : 1'b0;
  assign r_data_o[818] = (N3)? mem[818] : 
                         (N0)? mem[2418] : 1'b0;
  assign r_data_o[817] = (N3)? mem[817] : 
                         (N0)? mem[2417] : 1'b0;
  assign r_data_o[816] = (N3)? mem[816] : 
                         (N0)? mem[2416] : 1'b0;
  assign r_data_o[815] = (N3)? mem[815] : 
                         (N0)? mem[2415] : 1'b0;
  assign r_data_o[814] = (N3)? mem[814] : 
                         (N0)? mem[2414] : 1'b0;
  assign r_data_o[813] = (N3)? mem[813] : 
                         (N0)? mem[2413] : 1'b0;
  assign r_data_o[812] = (N3)? mem[812] : 
                         (N0)? mem[2412] : 1'b0;
  assign r_data_o[811] = (N3)? mem[811] : 
                         (N0)? mem[2411] : 1'b0;
  assign r_data_o[810] = (N3)? mem[810] : 
                         (N0)? mem[2410] : 1'b0;
  assign r_data_o[809] = (N3)? mem[809] : 
                         (N0)? mem[2409] : 1'b0;
  assign r_data_o[808] = (N3)? mem[808] : 
                         (N0)? mem[2408] : 1'b0;
  assign r_data_o[807] = (N3)? mem[807] : 
                         (N0)? mem[2407] : 1'b0;
  assign r_data_o[806] = (N3)? mem[806] : 
                         (N0)? mem[2406] : 1'b0;
  assign r_data_o[805] = (N3)? mem[805] : 
                         (N0)? mem[2405] : 1'b0;
  assign r_data_o[804] = (N3)? mem[804] : 
                         (N0)? mem[2404] : 1'b0;
  assign r_data_o[803] = (N3)? mem[803] : 
                         (N0)? mem[2403] : 1'b0;
  assign r_data_o[802] = (N3)? mem[802] : 
                         (N0)? mem[2402] : 1'b0;
  assign r_data_o[801] = (N3)? mem[801] : 
                         (N0)? mem[2401] : 1'b0;
  assign r_data_o[800] = (N3)? mem[800] : 
                         (N0)? mem[2400] : 1'b0;
  assign r_data_o[799] = (N3)? mem[799] : 
                         (N0)? mem[2399] : 1'b0;
  assign r_data_o[798] = (N3)? mem[798] : 
                         (N0)? mem[2398] : 1'b0;
  assign r_data_o[797] = (N3)? mem[797] : 
                         (N0)? mem[2397] : 1'b0;
  assign r_data_o[796] = (N3)? mem[796] : 
                         (N0)? mem[2396] : 1'b0;
  assign r_data_o[795] = (N3)? mem[795] : 
                         (N0)? mem[2395] : 1'b0;
  assign r_data_o[794] = (N3)? mem[794] : 
                         (N0)? mem[2394] : 1'b0;
  assign r_data_o[793] = (N3)? mem[793] : 
                         (N0)? mem[2393] : 1'b0;
  assign r_data_o[792] = (N3)? mem[792] : 
                         (N0)? mem[2392] : 1'b0;
  assign r_data_o[791] = (N3)? mem[791] : 
                         (N0)? mem[2391] : 1'b0;
  assign r_data_o[790] = (N3)? mem[790] : 
                         (N0)? mem[2390] : 1'b0;
  assign r_data_o[789] = (N3)? mem[789] : 
                         (N0)? mem[2389] : 1'b0;
  assign r_data_o[788] = (N3)? mem[788] : 
                         (N0)? mem[2388] : 1'b0;
  assign r_data_o[787] = (N3)? mem[787] : 
                         (N0)? mem[2387] : 1'b0;
  assign r_data_o[786] = (N3)? mem[786] : 
                         (N0)? mem[2386] : 1'b0;
  assign r_data_o[785] = (N3)? mem[785] : 
                         (N0)? mem[2385] : 1'b0;
  assign r_data_o[784] = (N3)? mem[784] : 
                         (N0)? mem[2384] : 1'b0;
  assign r_data_o[783] = (N3)? mem[783] : 
                         (N0)? mem[2383] : 1'b0;
  assign r_data_o[782] = (N3)? mem[782] : 
                         (N0)? mem[2382] : 1'b0;
  assign r_data_o[781] = (N3)? mem[781] : 
                         (N0)? mem[2381] : 1'b0;
  assign r_data_o[780] = (N3)? mem[780] : 
                         (N0)? mem[2380] : 1'b0;
  assign r_data_o[779] = (N3)? mem[779] : 
                         (N0)? mem[2379] : 1'b0;
  assign r_data_o[778] = (N3)? mem[778] : 
                         (N0)? mem[2378] : 1'b0;
  assign r_data_o[777] = (N3)? mem[777] : 
                         (N0)? mem[2377] : 1'b0;
  assign r_data_o[776] = (N3)? mem[776] : 
                         (N0)? mem[2376] : 1'b0;
  assign r_data_o[775] = (N3)? mem[775] : 
                         (N0)? mem[2375] : 1'b0;
  assign r_data_o[774] = (N3)? mem[774] : 
                         (N0)? mem[2374] : 1'b0;
  assign r_data_o[773] = (N3)? mem[773] : 
                         (N0)? mem[2373] : 1'b0;
  assign r_data_o[772] = (N3)? mem[772] : 
                         (N0)? mem[2372] : 1'b0;
  assign r_data_o[771] = (N3)? mem[771] : 
                         (N0)? mem[2371] : 1'b0;
  assign r_data_o[770] = (N3)? mem[770] : 
                         (N0)? mem[2370] : 1'b0;
  assign r_data_o[769] = (N3)? mem[769] : 
                         (N0)? mem[2369] : 1'b0;
  assign r_data_o[768] = (N3)? mem[768] : 
                         (N0)? mem[2368] : 1'b0;
  assign r_data_o[767] = (N3)? mem[767] : 
                         (N0)? mem[2367] : 1'b0;
  assign r_data_o[766] = (N3)? mem[766] : 
                         (N0)? mem[2366] : 1'b0;
  assign r_data_o[765] = (N3)? mem[765] : 
                         (N0)? mem[2365] : 1'b0;
  assign r_data_o[764] = (N3)? mem[764] : 
                         (N0)? mem[2364] : 1'b0;
  assign r_data_o[763] = (N3)? mem[763] : 
                         (N0)? mem[2363] : 1'b0;
  assign r_data_o[762] = (N3)? mem[762] : 
                         (N0)? mem[2362] : 1'b0;
  assign r_data_o[761] = (N3)? mem[761] : 
                         (N0)? mem[2361] : 1'b0;
  assign r_data_o[760] = (N3)? mem[760] : 
                         (N0)? mem[2360] : 1'b0;
  assign r_data_o[759] = (N3)? mem[759] : 
                         (N0)? mem[2359] : 1'b0;
  assign r_data_o[758] = (N3)? mem[758] : 
                         (N0)? mem[2358] : 1'b0;
  assign r_data_o[757] = (N3)? mem[757] : 
                         (N0)? mem[2357] : 1'b0;
  assign r_data_o[756] = (N3)? mem[756] : 
                         (N0)? mem[2356] : 1'b0;
  assign r_data_o[755] = (N3)? mem[755] : 
                         (N0)? mem[2355] : 1'b0;
  assign r_data_o[754] = (N3)? mem[754] : 
                         (N0)? mem[2354] : 1'b0;
  assign r_data_o[753] = (N3)? mem[753] : 
                         (N0)? mem[2353] : 1'b0;
  assign r_data_o[752] = (N3)? mem[752] : 
                         (N0)? mem[2352] : 1'b0;
  assign r_data_o[751] = (N3)? mem[751] : 
                         (N0)? mem[2351] : 1'b0;
  assign r_data_o[750] = (N3)? mem[750] : 
                         (N0)? mem[2350] : 1'b0;
  assign r_data_o[749] = (N3)? mem[749] : 
                         (N0)? mem[2349] : 1'b0;
  assign r_data_o[748] = (N3)? mem[748] : 
                         (N0)? mem[2348] : 1'b0;
  assign r_data_o[747] = (N3)? mem[747] : 
                         (N0)? mem[2347] : 1'b0;
  assign r_data_o[746] = (N3)? mem[746] : 
                         (N0)? mem[2346] : 1'b0;
  assign r_data_o[745] = (N3)? mem[745] : 
                         (N0)? mem[2345] : 1'b0;
  assign r_data_o[744] = (N3)? mem[744] : 
                         (N0)? mem[2344] : 1'b0;
  assign r_data_o[743] = (N3)? mem[743] : 
                         (N0)? mem[2343] : 1'b0;
  assign r_data_o[742] = (N3)? mem[742] : 
                         (N0)? mem[2342] : 1'b0;
  assign r_data_o[741] = (N3)? mem[741] : 
                         (N0)? mem[2341] : 1'b0;
  assign r_data_o[740] = (N3)? mem[740] : 
                         (N0)? mem[2340] : 1'b0;
  assign r_data_o[739] = (N3)? mem[739] : 
                         (N0)? mem[2339] : 1'b0;
  assign r_data_o[738] = (N3)? mem[738] : 
                         (N0)? mem[2338] : 1'b0;
  assign r_data_o[737] = (N3)? mem[737] : 
                         (N0)? mem[2337] : 1'b0;
  assign r_data_o[736] = (N3)? mem[736] : 
                         (N0)? mem[2336] : 1'b0;
  assign r_data_o[735] = (N3)? mem[735] : 
                         (N0)? mem[2335] : 1'b0;
  assign r_data_o[734] = (N3)? mem[734] : 
                         (N0)? mem[2334] : 1'b0;
  assign r_data_o[733] = (N3)? mem[733] : 
                         (N0)? mem[2333] : 1'b0;
  assign r_data_o[732] = (N3)? mem[732] : 
                         (N0)? mem[2332] : 1'b0;
  assign r_data_o[731] = (N3)? mem[731] : 
                         (N0)? mem[2331] : 1'b0;
  assign r_data_o[730] = (N3)? mem[730] : 
                         (N0)? mem[2330] : 1'b0;
  assign r_data_o[729] = (N3)? mem[729] : 
                         (N0)? mem[2329] : 1'b0;
  assign r_data_o[728] = (N3)? mem[728] : 
                         (N0)? mem[2328] : 1'b0;
  assign r_data_o[727] = (N3)? mem[727] : 
                         (N0)? mem[2327] : 1'b0;
  assign r_data_o[726] = (N3)? mem[726] : 
                         (N0)? mem[2326] : 1'b0;
  assign r_data_o[725] = (N3)? mem[725] : 
                         (N0)? mem[2325] : 1'b0;
  assign r_data_o[724] = (N3)? mem[724] : 
                         (N0)? mem[2324] : 1'b0;
  assign r_data_o[723] = (N3)? mem[723] : 
                         (N0)? mem[2323] : 1'b0;
  assign r_data_o[722] = (N3)? mem[722] : 
                         (N0)? mem[2322] : 1'b0;
  assign r_data_o[721] = (N3)? mem[721] : 
                         (N0)? mem[2321] : 1'b0;
  assign r_data_o[720] = (N3)? mem[720] : 
                         (N0)? mem[2320] : 1'b0;
  assign r_data_o[719] = (N3)? mem[719] : 
                         (N0)? mem[2319] : 1'b0;
  assign r_data_o[718] = (N3)? mem[718] : 
                         (N0)? mem[2318] : 1'b0;
  assign r_data_o[717] = (N3)? mem[717] : 
                         (N0)? mem[2317] : 1'b0;
  assign r_data_o[716] = (N3)? mem[716] : 
                         (N0)? mem[2316] : 1'b0;
  assign r_data_o[715] = (N3)? mem[715] : 
                         (N0)? mem[2315] : 1'b0;
  assign r_data_o[714] = (N3)? mem[714] : 
                         (N0)? mem[2314] : 1'b0;
  assign r_data_o[713] = (N3)? mem[713] : 
                         (N0)? mem[2313] : 1'b0;
  assign r_data_o[712] = (N3)? mem[712] : 
                         (N0)? mem[2312] : 1'b0;
  assign r_data_o[711] = (N3)? mem[711] : 
                         (N0)? mem[2311] : 1'b0;
  assign r_data_o[710] = (N3)? mem[710] : 
                         (N0)? mem[2310] : 1'b0;
  assign r_data_o[709] = (N3)? mem[709] : 
                         (N0)? mem[2309] : 1'b0;
  assign r_data_o[708] = (N3)? mem[708] : 
                         (N0)? mem[2308] : 1'b0;
  assign r_data_o[707] = (N3)? mem[707] : 
                         (N0)? mem[2307] : 1'b0;
  assign r_data_o[706] = (N3)? mem[706] : 
                         (N0)? mem[2306] : 1'b0;
  assign r_data_o[705] = (N3)? mem[705] : 
                         (N0)? mem[2305] : 1'b0;
  assign r_data_o[704] = (N3)? mem[704] : 
                         (N0)? mem[2304] : 1'b0;
  assign r_data_o[703] = (N3)? mem[703] : 
                         (N0)? mem[2303] : 1'b0;
  assign r_data_o[702] = (N3)? mem[702] : 
                         (N0)? mem[2302] : 1'b0;
  assign r_data_o[701] = (N3)? mem[701] : 
                         (N0)? mem[2301] : 1'b0;
  assign r_data_o[700] = (N3)? mem[700] : 
                         (N0)? mem[2300] : 1'b0;
  assign r_data_o[699] = (N3)? mem[699] : 
                         (N0)? mem[2299] : 1'b0;
  assign r_data_o[698] = (N3)? mem[698] : 
                         (N0)? mem[2298] : 1'b0;
  assign r_data_o[697] = (N3)? mem[697] : 
                         (N0)? mem[2297] : 1'b0;
  assign r_data_o[696] = (N3)? mem[696] : 
                         (N0)? mem[2296] : 1'b0;
  assign r_data_o[695] = (N3)? mem[695] : 
                         (N0)? mem[2295] : 1'b0;
  assign r_data_o[694] = (N3)? mem[694] : 
                         (N0)? mem[2294] : 1'b0;
  assign r_data_o[693] = (N3)? mem[693] : 
                         (N0)? mem[2293] : 1'b0;
  assign r_data_o[692] = (N3)? mem[692] : 
                         (N0)? mem[2292] : 1'b0;
  assign r_data_o[691] = (N3)? mem[691] : 
                         (N0)? mem[2291] : 1'b0;
  assign r_data_o[690] = (N3)? mem[690] : 
                         (N0)? mem[2290] : 1'b0;
  assign r_data_o[689] = (N3)? mem[689] : 
                         (N0)? mem[2289] : 1'b0;
  assign r_data_o[688] = (N3)? mem[688] : 
                         (N0)? mem[2288] : 1'b0;
  assign r_data_o[687] = (N3)? mem[687] : 
                         (N0)? mem[2287] : 1'b0;
  assign r_data_o[686] = (N3)? mem[686] : 
                         (N0)? mem[2286] : 1'b0;
  assign r_data_o[685] = (N3)? mem[685] : 
                         (N0)? mem[2285] : 1'b0;
  assign r_data_o[684] = (N3)? mem[684] : 
                         (N0)? mem[2284] : 1'b0;
  assign r_data_o[683] = (N3)? mem[683] : 
                         (N0)? mem[2283] : 1'b0;
  assign r_data_o[682] = (N3)? mem[682] : 
                         (N0)? mem[2282] : 1'b0;
  assign r_data_o[681] = (N3)? mem[681] : 
                         (N0)? mem[2281] : 1'b0;
  assign r_data_o[680] = (N3)? mem[680] : 
                         (N0)? mem[2280] : 1'b0;
  assign r_data_o[679] = (N3)? mem[679] : 
                         (N0)? mem[2279] : 1'b0;
  assign r_data_o[678] = (N3)? mem[678] : 
                         (N0)? mem[2278] : 1'b0;
  assign r_data_o[677] = (N3)? mem[677] : 
                         (N0)? mem[2277] : 1'b0;
  assign r_data_o[676] = (N3)? mem[676] : 
                         (N0)? mem[2276] : 1'b0;
  assign r_data_o[675] = (N3)? mem[675] : 
                         (N0)? mem[2275] : 1'b0;
  assign r_data_o[674] = (N3)? mem[674] : 
                         (N0)? mem[2274] : 1'b0;
  assign r_data_o[673] = (N3)? mem[673] : 
                         (N0)? mem[2273] : 1'b0;
  assign r_data_o[672] = (N3)? mem[672] : 
                         (N0)? mem[2272] : 1'b0;
  assign r_data_o[671] = (N3)? mem[671] : 
                         (N0)? mem[2271] : 1'b0;
  assign r_data_o[670] = (N3)? mem[670] : 
                         (N0)? mem[2270] : 1'b0;
  assign r_data_o[669] = (N3)? mem[669] : 
                         (N0)? mem[2269] : 1'b0;
  assign r_data_o[668] = (N3)? mem[668] : 
                         (N0)? mem[2268] : 1'b0;
  assign r_data_o[667] = (N3)? mem[667] : 
                         (N0)? mem[2267] : 1'b0;
  assign r_data_o[666] = (N3)? mem[666] : 
                         (N0)? mem[2266] : 1'b0;
  assign r_data_o[665] = (N3)? mem[665] : 
                         (N0)? mem[2265] : 1'b0;
  assign r_data_o[664] = (N3)? mem[664] : 
                         (N0)? mem[2264] : 1'b0;
  assign r_data_o[663] = (N3)? mem[663] : 
                         (N0)? mem[2263] : 1'b0;
  assign r_data_o[662] = (N3)? mem[662] : 
                         (N0)? mem[2262] : 1'b0;
  assign r_data_o[661] = (N3)? mem[661] : 
                         (N0)? mem[2261] : 1'b0;
  assign r_data_o[660] = (N3)? mem[660] : 
                         (N0)? mem[2260] : 1'b0;
  assign r_data_o[659] = (N3)? mem[659] : 
                         (N0)? mem[2259] : 1'b0;
  assign r_data_o[658] = (N3)? mem[658] : 
                         (N0)? mem[2258] : 1'b0;
  assign r_data_o[657] = (N3)? mem[657] : 
                         (N0)? mem[2257] : 1'b0;
  assign r_data_o[656] = (N3)? mem[656] : 
                         (N0)? mem[2256] : 1'b0;
  assign r_data_o[655] = (N3)? mem[655] : 
                         (N0)? mem[2255] : 1'b0;
  assign r_data_o[654] = (N3)? mem[654] : 
                         (N0)? mem[2254] : 1'b0;
  assign r_data_o[653] = (N3)? mem[653] : 
                         (N0)? mem[2253] : 1'b0;
  assign r_data_o[652] = (N3)? mem[652] : 
                         (N0)? mem[2252] : 1'b0;
  assign r_data_o[651] = (N3)? mem[651] : 
                         (N0)? mem[2251] : 1'b0;
  assign r_data_o[650] = (N3)? mem[650] : 
                         (N0)? mem[2250] : 1'b0;
  assign r_data_o[649] = (N3)? mem[649] : 
                         (N0)? mem[2249] : 1'b0;
  assign r_data_o[648] = (N3)? mem[648] : 
                         (N0)? mem[2248] : 1'b0;
  assign r_data_o[647] = (N3)? mem[647] : 
                         (N0)? mem[2247] : 1'b0;
  assign r_data_o[646] = (N3)? mem[646] : 
                         (N0)? mem[2246] : 1'b0;
  assign r_data_o[645] = (N3)? mem[645] : 
                         (N0)? mem[2245] : 1'b0;
  assign r_data_o[644] = (N3)? mem[644] : 
                         (N0)? mem[2244] : 1'b0;
  assign r_data_o[643] = (N3)? mem[643] : 
                         (N0)? mem[2243] : 1'b0;
  assign r_data_o[642] = (N3)? mem[642] : 
                         (N0)? mem[2242] : 1'b0;
  assign r_data_o[641] = (N3)? mem[641] : 
                         (N0)? mem[2241] : 1'b0;
  assign r_data_o[640] = (N3)? mem[640] : 
                         (N0)? mem[2240] : 1'b0;
  assign r_data_o[639] = (N3)? mem[639] : 
                         (N0)? mem[2239] : 1'b0;
  assign r_data_o[638] = (N3)? mem[638] : 
                         (N0)? mem[2238] : 1'b0;
  assign r_data_o[637] = (N3)? mem[637] : 
                         (N0)? mem[2237] : 1'b0;
  assign r_data_o[636] = (N3)? mem[636] : 
                         (N0)? mem[2236] : 1'b0;
  assign r_data_o[635] = (N3)? mem[635] : 
                         (N0)? mem[2235] : 1'b0;
  assign r_data_o[634] = (N3)? mem[634] : 
                         (N0)? mem[2234] : 1'b0;
  assign r_data_o[633] = (N3)? mem[633] : 
                         (N0)? mem[2233] : 1'b0;
  assign r_data_o[632] = (N3)? mem[632] : 
                         (N0)? mem[2232] : 1'b0;
  assign r_data_o[631] = (N3)? mem[631] : 
                         (N0)? mem[2231] : 1'b0;
  assign r_data_o[630] = (N3)? mem[630] : 
                         (N0)? mem[2230] : 1'b0;
  assign r_data_o[629] = (N3)? mem[629] : 
                         (N0)? mem[2229] : 1'b0;
  assign r_data_o[628] = (N3)? mem[628] : 
                         (N0)? mem[2228] : 1'b0;
  assign r_data_o[627] = (N3)? mem[627] : 
                         (N0)? mem[2227] : 1'b0;
  assign r_data_o[626] = (N3)? mem[626] : 
                         (N0)? mem[2226] : 1'b0;
  assign r_data_o[625] = (N3)? mem[625] : 
                         (N0)? mem[2225] : 1'b0;
  assign r_data_o[624] = (N3)? mem[624] : 
                         (N0)? mem[2224] : 1'b0;
  assign r_data_o[623] = (N3)? mem[623] : 
                         (N0)? mem[2223] : 1'b0;
  assign r_data_o[622] = (N3)? mem[622] : 
                         (N0)? mem[2222] : 1'b0;
  assign r_data_o[621] = (N3)? mem[621] : 
                         (N0)? mem[2221] : 1'b0;
  assign r_data_o[620] = (N3)? mem[620] : 
                         (N0)? mem[2220] : 1'b0;
  assign r_data_o[619] = (N3)? mem[619] : 
                         (N0)? mem[2219] : 1'b0;
  assign r_data_o[618] = (N3)? mem[618] : 
                         (N0)? mem[2218] : 1'b0;
  assign r_data_o[617] = (N3)? mem[617] : 
                         (N0)? mem[2217] : 1'b0;
  assign r_data_o[616] = (N3)? mem[616] : 
                         (N0)? mem[2216] : 1'b0;
  assign r_data_o[615] = (N3)? mem[615] : 
                         (N0)? mem[2215] : 1'b0;
  assign r_data_o[614] = (N3)? mem[614] : 
                         (N0)? mem[2214] : 1'b0;
  assign r_data_o[613] = (N3)? mem[613] : 
                         (N0)? mem[2213] : 1'b0;
  assign r_data_o[612] = (N3)? mem[612] : 
                         (N0)? mem[2212] : 1'b0;
  assign r_data_o[611] = (N3)? mem[611] : 
                         (N0)? mem[2211] : 1'b0;
  assign r_data_o[610] = (N3)? mem[610] : 
                         (N0)? mem[2210] : 1'b0;
  assign r_data_o[609] = (N3)? mem[609] : 
                         (N0)? mem[2209] : 1'b0;
  assign r_data_o[608] = (N3)? mem[608] : 
                         (N0)? mem[2208] : 1'b0;
  assign r_data_o[607] = (N3)? mem[607] : 
                         (N0)? mem[2207] : 1'b0;
  assign r_data_o[606] = (N3)? mem[606] : 
                         (N0)? mem[2206] : 1'b0;
  assign r_data_o[605] = (N3)? mem[605] : 
                         (N0)? mem[2205] : 1'b0;
  assign r_data_o[604] = (N3)? mem[604] : 
                         (N0)? mem[2204] : 1'b0;
  assign r_data_o[603] = (N3)? mem[603] : 
                         (N0)? mem[2203] : 1'b0;
  assign r_data_o[602] = (N3)? mem[602] : 
                         (N0)? mem[2202] : 1'b0;
  assign r_data_o[601] = (N3)? mem[601] : 
                         (N0)? mem[2201] : 1'b0;
  assign r_data_o[600] = (N3)? mem[600] : 
                         (N0)? mem[2200] : 1'b0;
  assign r_data_o[599] = (N3)? mem[599] : 
                         (N0)? mem[2199] : 1'b0;
  assign r_data_o[598] = (N3)? mem[598] : 
                         (N0)? mem[2198] : 1'b0;
  assign r_data_o[597] = (N3)? mem[597] : 
                         (N0)? mem[2197] : 1'b0;
  assign r_data_o[596] = (N3)? mem[596] : 
                         (N0)? mem[2196] : 1'b0;
  assign r_data_o[595] = (N3)? mem[595] : 
                         (N0)? mem[2195] : 1'b0;
  assign r_data_o[594] = (N3)? mem[594] : 
                         (N0)? mem[2194] : 1'b0;
  assign r_data_o[593] = (N3)? mem[593] : 
                         (N0)? mem[2193] : 1'b0;
  assign r_data_o[592] = (N3)? mem[592] : 
                         (N0)? mem[2192] : 1'b0;
  assign r_data_o[591] = (N3)? mem[591] : 
                         (N0)? mem[2191] : 1'b0;
  assign r_data_o[590] = (N3)? mem[590] : 
                         (N0)? mem[2190] : 1'b0;
  assign r_data_o[589] = (N3)? mem[589] : 
                         (N0)? mem[2189] : 1'b0;
  assign r_data_o[588] = (N3)? mem[588] : 
                         (N0)? mem[2188] : 1'b0;
  assign r_data_o[587] = (N3)? mem[587] : 
                         (N0)? mem[2187] : 1'b0;
  assign r_data_o[586] = (N3)? mem[586] : 
                         (N0)? mem[2186] : 1'b0;
  assign r_data_o[585] = (N3)? mem[585] : 
                         (N0)? mem[2185] : 1'b0;
  assign r_data_o[584] = (N3)? mem[584] : 
                         (N0)? mem[2184] : 1'b0;
  assign r_data_o[583] = (N3)? mem[583] : 
                         (N0)? mem[2183] : 1'b0;
  assign r_data_o[582] = (N3)? mem[582] : 
                         (N0)? mem[2182] : 1'b0;
  assign r_data_o[581] = (N3)? mem[581] : 
                         (N0)? mem[2181] : 1'b0;
  assign r_data_o[580] = (N3)? mem[580] : 
                         (N0)? mem[2180] : 1'b0;
  assign r_data_o[579] = (N3)? mem[579] : 
                         (N0)? mem[2179] : 1'b0;
  assign r_data_o[578] = (N3)? mem[578] : 
                         (N0)? mem[2178] : 1'b0;
  assign r_data_o[577] = (N3)? mem[577] : 
                         (N0)? mem[2177] : 1'b0;
  assign r_data_o[576] = (N3)? mem[576] : 
                         (N0)? mem[2176] : 1'b0;
  assign r_data_o[575] = (N3)? mem[575] : 
                         (N0)? mem[2175] : 1'b0;
  assign r_data_o[574] = (N3)? mem[574] : 
                         (N0)? mem[2174] : 1'b0;
  assign r_data_o[573] = (N3)? mem[573] : 
                         (N0)? mem[2173] : 1'b0;
  assign r_data_o[572] = (N3)? mem[572] : 
                         (N0)? mem[2172] : 1'b0;
  assign r_data_o[571] = (N3)? mem[571] : 
                         (N0)? mem[2171] : 1'b0;
  assign r_data_o[570] = (N3)? mem[570] : 
                         (N0)? mem[2170] : 1'b0;
  assign r_data_o[569] = (N3)? mem[569] : 
                         (N0)? mem[2169] : 1'b0;
  assign r_data_o[568] = (N3)? mem[568] : 
                         (N0)? mem[2168] : 1'b0;
  assign r_data_o[567] = (N3)? mem[567] : 
                         (N0)? mem[2167] : 1'b0;
  assign r_data_o[566] = (N3)? mem[566] : 
                         (N0)? mem[2166] : 1'b0;
  assign r_data_o[565] = (N3)? mem[565] : 
                         (N0)? mem[2165] : 1'b0;
  assign r_data_o[564] = (N3)? mem[564] : 
                         (N0)? mem[2164] : 1'b0;
  assign r_data_o[563] = (N3)? mem[563] : 
                         (N0)? mem[2163] : 1'b0;
  assign r_data_o[562] = (N3)? mem[562] : 
                         (N0)? mem[2162] : 1'b0;
  assign r_data_o[561] = (N3)? mem[561] : 
                         (N0)? mem[2161] : 1'b0;
  assign r_data_o[560] = (N3)? mem[560] : 
                         (N0)? mem[2160] : 1'b0;
  assign r_data_o[559] = (N3)? mem[559] : 
                         (N0)? mem[2159] : 1'b0;
  assign r_data_o[558] = (N3)? mem[558] : 
                         (N0)? mem[2158] : 1'b0;
  assign r_data_o[557] = (N3)? mem[557] : 
                         (N0)? mem[2157] : 1'b0;
  assign r_data_o[556] = (N3)? mem[556] : 
                         (N0)? mem[2156] : 1'b0;
  assign r_data_o[555] = (N3)? mem[555] : 
                         (N0)? mem[2155] : 1'b0;
  assign r_data_o[554] = (N3)? mem[554] : 
                         (N0)? mem[2154] : 1'b0;
  assign r_data_o[553] = (N3)? mem[553] : 
                         (N0)? mem[2153] : 1'b0;
  assign r_data_o[552] = (N3)? mem[552] : 
                         (N0)? mem[2152] : 1'b0;
  assign r_data_o[551] = (N3)? mem[551] : 
                         (N0)? mem[2151] : 1'b0;
  assign r_data_o[550] = (N3)? mem[550] : 
                         (N0)? mem[2150] : 1'b0;
  assign r_data_o[549] = (N3)? mem[549] : 
                         (N0)? mem[2149] : 1'b0;
  assign r_data_o[548] = (N3)? mem[548] : 
                         (N0)? mem[2148] : 1'b0;
  assign r_data_o[547] = (N3)? mem[547] : 
                         (N0)? mem[2147] : 1'b0;
  assign r_data_o[546] = (N3)? mem[546] : 
                         (N0)? mem[2146] : 1'b0;
  assign r_data_o[545] = (N3)? mem[545] : 
                         (N0)? mem[2145] : 1'b0;
  assign r_data_o[544] = (N3)? mem[544] : 
                         (N0)? mem[2144] : 1'b0;
  assign r_data_o[543] = (N3)? mem[543] : 
                         (N0)? mem[2143] : 1'b0;
  assign r_data_o[542] = (N3)? mem[542] : 
                         (N0)? mem[2142] : 1'b0;
  assign r_data_o[541] = (N3)? mem[541] : 
                         (N0)? mem[2141] : 1'b0;
  assign r_data_o[540] = (N3)? mem[540] : 
                         (N0)? mem[2140] : 1'b0;
  assign r_data_o[539] = (N3)? mem[539] : 
                         (N0)? mem[2139] : 1'b0;
  assign r_data_o[538] = (N3)? mem[538] : 
                         (N0)? mem[2138] : 1'b0;
  assign r_data_o[537] = (N3)? mem[537] : 
                         (N0)? mem[2137] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] : 
                         (N0)? mem[2136] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] : 
                         (N0)? mem[2135] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] : 
                         (N0)? mem[2134] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] : 
                         (N0)? mem[2133] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] : 
                         (N0)? mem[2132] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] : 
                         (N0)? mem[2131] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] : 
                         (N0)? mem[2130] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] : 
                         (N0)? mem[2129] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] : 
                         (N0)? mem[2128] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] : 
                         (N0)? mem[2127] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] : 
                         (N0)? mem[2126] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] : 
                         (N0)? mem[2125] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] : 
                         (N0)? mem[2124] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] : 
                         (N0)? mem[2123] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] : 
                         (N0)? mem[2122] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] : 
                         (N0)? mem[2121] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] : 
                         (N0)? mem[2120] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] : 
                         (N0)? mem[2119] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] : 
                         (N0)? mem[2118] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] : 
                         (N0)? mem[2117] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] : 
                         (N0)? mem[2116] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] : 
                         (N0)? mem[2115] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] : 
                         (N0)? mem[2114] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] : 
                         (N0)? mem[2113] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] : 
                         (N0)? mem[2112] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] : 
                         (N0)? mem[2111] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] : 
                         (N0)? mem[2110] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] : 
                         (N0)? mem[2109] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] : 
                         (N0)? mem[2108] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] : 
                         (N0)? mem[2107] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] : 
                         (N0)? mem[2106] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] : 
                         (N0)? mem[2105] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] : 
                         (N0)? mem[2104] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] : 
                         (N0)? mem[2103] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] : 
                         (N0)? mem[2102] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] : 
                         (N0)? mem[2101] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] : 
                         (N0)? mem[2100] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] : 
                         (N0)? mem[2099] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] : 
                         (N0)? mem[2098] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] : 
                         (N0)? mem[2097] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] : 
                         (N0)? mem[2096] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] : 
                         (N0)? mem[2095] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] : 
                         (N0)? mem[2094] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] : 
                         (N0)? mem[2093] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] : 
                         (N0)? mem[2092] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] : 
                         (N0)? mem[2091] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] : 
                         (N0)? mem[2090] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] : 
                         (N0)? mem[2089] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] : 
                         (N0)? mem[2088] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] : 
                         (N0)? mem[2087] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] : 
                         (N0)? mem[2086] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] : 
                         (N0)? mem[2085] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] : 
                         (N0)? mem[2084] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] : 
                         (N0)? mem[2083] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] : 
                         (N0)? mem[2082] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] : 
                         (N0)? mem[2081] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] : 
                         (N0)? mem[2080] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] : 
                         (N0)? mem[2079] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] : 
                         (N0)? mem[2078] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] : 
                         (N0)? mem[2077] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] : 
                         (N0)? mem[2076] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] : 
                         (N0)? mem[2075] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] : 
                         (N0)? mem[2074] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] : 
                         (N0)? mem[2073] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] : 
                         (N0)? mem[2072] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] : 
                         (N0)? mem[2071] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] : 
                         (N0)? mem[2070] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] : 
                         (N0)? mem[2069] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] : 
                         (N0)? mem[2068] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] : 
                         (N0)? mem[2067] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] : 
                         (N0)? mem[2066] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] : 
                         (N0)? mem[2065] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] : 
                         (N0)? mem[2064] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] : 
                         (N0)? mem[2063] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] : 
                         (N0)? mem[2062] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] : 
                         (N0)? mem[2061] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] : 
                         (N0)? mem[2060] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] : 
                         (N0)? mem[2059] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] : 
                         (N0)? mem[2058] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] : 
                         (N0)? mem[2057] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] : 
                         (N0)? mem[2056] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] : 
                         (N0)? mem[2055] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] : 
                         (N0)? mem[2054] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] : 
                         (N0)? mem[2053] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] : 
                         (N0)? mem[2052] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] : 
                         (N0)? mem[2051] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] : 
                         (N0)? mem[2050] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] : 
                         (N0)? mem[2049] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] : 
                         (N0)? mem[2048] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] : 
                         (N0)? mem[2047] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] : 
                         (N0)? mem[2046] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] : 
                         (N0)? mem[2045] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] : 
                         (N0)? mem[2044] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] : 
                         (N0)? mem[2043] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] : 
                         (N0)? mem[2042] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] : 
                         (N0)? mem[2041] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] : 
                         (N0)? mem[2040] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] : 
                         (N0)? mem[2039] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] : 
                         (N0)? mem[2038] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] : 
                         (N0)? mem[2037] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] : 
                         (N0)? mem[2036] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] : 
                         (N0)? mem[2035] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] : 
                         (N0)? mem[2034] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] : 
                         (N0)? mem[2033] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] : 
                         (N0)? mem[2032] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] : 
                         (N0)? mem[2031] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] : 
                         (N0)? mem[2030] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] : 
                         (N0)? mem[2029] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] : 
                         (N0)? mem[2028] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] : 
                         (N0)? mem[2027] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] : 
                         (N0)? mem[2026] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] : 
                         (N0)? mem[2025] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] : 
                         (N0)? mem[2024] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] : 
                         (N0)? mem[2023] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] : 
                         (N0)? mem[2022] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] : 
                         (N0)? mem[2021] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] : 
                         (N0)? mem[2020] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] : 
                         (N0)? mem[2019] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] : 
                         (N0)? mem[2018] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] : 
                         (N0)? mem[2017] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] : 
                         (N0)? mem[2016] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] : 
                         (N0)? mem[2015] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] : 
                         (N0)? mem[2014] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] : 
                         (N0)? mem[2013] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] : 
                         (N0)? mem[2012] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] : 
                         (N0)? mem[2011] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] : 
                         (N0)? mem[2010] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] : 
                         (N0)? mem[2009] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] : 
                         (N0)? mem[2008] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] : 
                         (N0)? mem[2007] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] : 
                         (N0)? mem[2006] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] : 
                         (N0)? mem[2005] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] : 
                         (N0)? mem[2004] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] : 
                         (N0)? mem[2003] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] : 
                         (N0)? mem[2002] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] : 
                         (N0)? mem[2001] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] : 
                         (N0)? mem[2000] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] : 
                         (N0)? mem[1999] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] : 
                         (N0)? mem[1998] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] : 
                         (N0)? mem[1997] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] : 
                         (N0)? mem[1996] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] : 
                         (N0)? mem[1995] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] : 
                         (N0)? mem[1994] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] : 
                         (N0)? mem[1993] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] : 
                         (N0)? mem[1992] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] : 
                         (N0)? mem[1991] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] : 
                         (N0)? mem[1990] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] : 
                         (N0)? mem[1989] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] : 
                         (N0)? mem[1988] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] : 
                         (N0)? mem[1987] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] : 
                         (N0)? mem[1986] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] : 
                         (N0)? mem[1985] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] : 
                         (N0)? mem[1984] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] : 
                         (N0)? mem[1983] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] : 
                         (N0)? mem[1982] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] : 
                         (N0)? mem[1981] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] : 
                         (N0)? mem[1980] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] : 
                         (N0)? mem[1979] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] : 
                         (N0)? mem[1978] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] : 
                         (N0)? mem[1977] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] : 
                         (N0)? mem[1976] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] : 
                         (N0)? mem[1975] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] : 
                         (N0)? mem[1974] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] : 
                         (N0)? mem[1973] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] : 
                         (N0)? mem[1972] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] : 
                         (N0)? mem[1971] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] : 
                         (N0)? mem[1970] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] : 
                         (N0)? mem[1969] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] : 
                         (N0)? mem[1968] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] : 
                         (N0)? mem[1967] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] : 
                         (N0)? mem[1966] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] : 
                         (N0)? mem[1965] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] : 
                         (N0)? mem[1964] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] : 
                         (N0)? mem[1963] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] : 
                         (N0)? mem[1962] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] : 
                         (N0)? mem[1961] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] : 
                         (N0)? mem[1960] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] : 
                         (N0)? mem[1959] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] : 
                         (N0)? mem[1958] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] : 
                         (N0)? mem[1957] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] : 
                         (N0)? mem[1956] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] : 
                         (N0)? mem[1955] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] : 
                         (N0)? mem[1954] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] : 
                         (N0)? mem[1953] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] : 
                         (N0)? mem[1952] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] : 
                         (N0)? mem[1951] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] : 
                         (N0)? mem[1950] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] : 
                         (N0)? mem[1949] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] : 
                         (N0)? mem[1948] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] : 
                         (N0)? mem[1947] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] : 
                         (N0)? mem[1946] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] : 
                         (N0)? mem[1945] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] : 
                         (N0)? mem[1944] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] : 
                         (N0)? mem[1943] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] : 
                         (N0)? mem[1942] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] : 
                         (N0)? mem[1941] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] : 
                         (N0)? mem[1940] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] : 
                         (N0)? mem[1939] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] : 
                         (N0)? mem[1938] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] : 
                         (N0)? mem[1937] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] : 
                         (N0)? mem[1936] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] : 
                         (N0)? mem[1935] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] : 
                         (N0)? mem[1934] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] : 
                         (N0)? mem[1933] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] : 
                         (N0)? mem[1932] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] : 
                         (N0)? mem[1931] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] : 
                         (N0)? mem[1930] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] : 
                         (N0)? mem[1929] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] : 
                         (N0)? mem[1928] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] : 
                         (N0)? mem[1927] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] : 
                         (N0)? mem[1926] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] : 
                         (N0)? mem[1925] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] : 
                         (N0)? mem[1924] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] : 
                         (N0)? mem[1923] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] : 
                         (N0)? mem[1922] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] : 
                         (N0)? mem[1921] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] : 
                         (N0)? mem[1920] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] : 
                         (N0)? mem[1919] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] : 
                         (N0)? mem[1918] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] : 
                         (N0)? mem[1917] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] : 
                         (N0)? mem[1916] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] : 
                         (N0)? mem[1915] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] : 
                         (N0)? mem[1914] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] : 
                         (N0)? mem[1913] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] : 
                         (N0)? mem[1912] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] : 
                         (N0)? mem[1911] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] : 
                         (N0)? mem[1910] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] : 
                         (N0)? mem[1909] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] : 
                         (N0)? mem[1908] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] : 
                         (N0)? mem[1907] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] : 
                         (N0)? mem[1906] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] : 
                         (N0)? mem[1905] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] : 
                         (N0)? mem[1904] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] : 
                         (N0)? mem[1903] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] : 
                         (N0)? mem[1902] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] : 
                         (N0)? mem[1901] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] : 
                         (N0)? mem[1900] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] : 
                         (N0)? mem[1899] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] : 
                         (N0)? mem[1898] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] : 
                         (N0)? mem[1897] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] : 
                         (N0)? mem[1896] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] : 
                         (N0)? mem[1895] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] : 
                         (N0)? mem[1894] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] : 
                         (N0)? mem[1893] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] : 
                         (N0)? mem[1892] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] : 
                         (N0)? mem[1891] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] : 
                         (N0)? mem[1890] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] : 
                         (N0)? mem[1889] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] : 
                         (N0)? mem[1888] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] : 
                         (N0)? mem[1887] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] : 
                         (N0)? mem[1886] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] : 
                         (N0)? mem[1885] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] : 
                         (N0)? mem[1884] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] : 
                         (N0)? mem[1883] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] : 
                         (N0)? mem[1882] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] : 
                         (N0)? mem[1881] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] : 
                         (N0)? mem[1880] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] : 
                         (N0)? mem[1879] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] : 
                         (N0)? mem[1878] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] : 
                         (N0)? mem[1877] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] : 
                         (N0)? mem[1876] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] : 
                         (N0)? mem[1875] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] : 
                         (N0)? mem[1874] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] : 
                         (N0)? mem[1873] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] : 
                         (N0)? mem[1872] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] : 
                         (N0)? mem[1871] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] : 
                         (N0)? mem[1870] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] : 
                         (N0)? mem[1869] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] : 
                         (N0)? mem[1868] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] : 
                         (N0)? mem[1867] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] : 
                         (N0)? mem[1866] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] : 
                         (N0)? mem[1865] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] : 
                         (N0)? mem[1864] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] : 
                         (N0)? mem[1863] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] : 
                         (N0)? mem[1862] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] : 
                         (N0)? mem[1861] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] : 
                         (N0)? mem[1860] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] : 
                         (N0)? mem[1859] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] : 
                         (N0)? mem[1858] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] : 
                         (N0)? mem[1857] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] : 
                         (N0)? mem[1856] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[1855] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[1854] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[1853] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[1852] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[1851] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[1850] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[1849] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[1848] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[1847] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[1846] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[1845] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[1844] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[1843] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[1842] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[1841] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[1840] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[1839] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[1838] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[1837] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[1836] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[1835] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[1834] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[1833] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[1832] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[1831] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[1830] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[1829] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[1828] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[1827] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[1826] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[1825] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[1824] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[1823] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[1822] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[1821] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[1820] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[1819] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[1818] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[1817] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[1816] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[1815] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[1814] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[1813] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[1812] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[1811] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[1810] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[1809] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[1808] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[1807] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[1806] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[1805] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[1804] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[1803] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[1802] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[1801] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[1800] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[1799] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[1798] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[1797] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[1796] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[1795] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[1794] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[1793] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[1792] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[1791] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[1790] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[1789] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[1788] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[1787] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[1786] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[1785] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[1784] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[1783] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[1782] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[1781] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[1780] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[1779] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[1778] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[1777] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[1776] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[1775] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[1774] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[1773] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[1772] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[1771] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[1770] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[1769] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[1768] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[1767] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[1766] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[1765] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[1764] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[1763] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[1762] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[1761] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[1760] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[1759] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[1758] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[1757] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[1756] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[1755] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[1754] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[1753] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[1752] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[1751] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[1750] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[1749] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[1748] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[1747] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[1746] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[1745] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[1744] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[1743] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[1742] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[1741] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[1740] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[1739] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[1738] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[1737] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[1736] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[1735] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[1734] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[1733] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[1732] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[1731] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[1730] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[1729] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[1728] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[1727] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[1726] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[1725] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[1724] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[1723] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[1722] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[1721] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[1720] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[1719] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[1718] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[1717] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[1716] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[1715] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[1714] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[1713] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[1712] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[1711] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[1710] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[1709] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[1708] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[1707] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[1706] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[1705] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[1704] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[1703] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[1702] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[1701] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[1700] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[1699] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[1698] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[1697] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[1696] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[1695] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[1694] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[1693] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[1692] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[1691] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[1690] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[1689] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[1688] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[1687] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[1686] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[1685] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[1684] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[1683] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[1682] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[1681] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[1680] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[1679] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[1678] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[1677] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[1676] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[1675] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[1674] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[1673] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[1672] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[1671] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[1670] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[1669] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[1668] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[1667] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[1666] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[1665] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[1664] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[1663] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[1662] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[1661] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[1660] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[1659] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[1658] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[1657] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[1656] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[1655] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[1654] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[1653] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[1652] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[1651] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[1650] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[1649] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[1648] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[1647] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[1646] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[1645] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[1644] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[1643] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[1642] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[1641] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[1640] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[1639] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[1638] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[1637] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[1636] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[1635] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[1634] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[1633] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[1632] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[1631] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[1630] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[1629] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[1628] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[1627] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[1626] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[1625] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[1624] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[1623] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[1622] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[1621] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[1620] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[1619] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[1618] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[1617] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[1616] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[1615] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[1614] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[1613] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[1612] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[1611] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[1610] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[1609] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[1608] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[1607] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[1606] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[1605] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[1604] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[1603] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[1602] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[1601] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[1600] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5 } : 
                                                                                                                                                                           (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N23) begin
      mem_3199_sv2v_reg <= w_data_i[1599];
      mem_3198_sv2v_reg <= w_data_i[1598];
      mem_3197_sv2v_reg <= w_data_i[1597];
      mem_3196_sv2v_reg <= w_data_i[1596];
      mem_3195_sv2v_reg <= w_data_i[1595];
      mem_3194_sv2v_reg <= w_data_i[1594];
      mem_3193_sv2v_reg <= w_data_i[1593];
      mem_3192_sv2v_reg <= w_data_i[1592];
      mem_3191_sv2v_reg <= w_data_i[1591];
      mem_3190_sv2v_reg <= w_data_i[1590];
      mem_3189_sv2v_reg <= w_data_i[1589];
      mem_3188_sv2v_reg <= w_data_i[1588];
      mem_3187_sv2v_reg <= w_data_i[1587];
      mem_3186_sv2v_reg <= w_data_i[1586];
      mem_3185_sv2v_reg <= w_data_i[1585];
      mem_3184_sv2v_reg <= w_data_i[1584];
      mem_3183_sv2v_reg <= w_data_i[1583];
      mem_3182_sv2v_reg <= w_data_i[1582];
      mem_3181_sv2v_reg <= w_data_i[1581];
      mem_3180_sv2v_reg <= w_data_i[1580];
      mem_3179_sv2v_reg <= w_data_i[1579];
      mem_3178_sv2v_reg <= w_data_i[1578];
      mem_3177_sv2v_reg <= w_data_i[1577];
      mem_3176_sv2v_reg <= w_data_i[1576];
      mem_3175_sv2v_reg <= w_data_i[1575];
      mem_3174_sv2v_reg <= w_data_i[1574];
      mem_3173_sv2v_reg <= w_data_i[1573];
      mem_3172_sv2v_reg <= w_data_i[1572];
      mem_3171_sv2v_reg <= w_data_i[1571];
      mem_3170_sv2v_reg <= w_data_i[1570];
      mem_3169_sv2v_reg <= w_data_i[1569];
      mem_3168_sv2v_reg <= w_data_i[1568];
      mem_3167_sv2v_reg <= w_data_i[1567];
      mem_3166_sv2v_reg <= w_data_i[1566];
      mem_3165_sv2v_reg <= w_data_i[1565];
      mem_3164_sv2v_reg <= w_data_i[1564];
      mem_3163_sv2v_reg <= w_data_i[1563];
      mem_3162_sv2v_reg <= w_data_i[1562];
      mem_3161_sv2v_reg <= w_data_i[1561];
      mem_3160_sv2v_reg <= w_data_i[1560];
      mem_3159_sv2v_reg <= w_data_i[1559];
      mem_3158_sv2v_reg <= w_data_i[1558];
      mem_3157_sv2v_reg <= w_data_i[1557];
      mem_3156_sv2v_reg <= w_data_i[1556];
      mem_3155_sv2v_reg <= w_data_i[1555];
      mem_3154_sv2v_reg <= w_data_i[1554];
      mem_3153_sv2v_reg <= w_data_i[1553];
      mem_3152_sv2v_reg <= w_data_i[1552];
      mem_3151_sv2v_reg <= w_data_i[1551];
      mem_3150_sv2v_reg <= w_data_i[1550];
      mem_3149_sv2v_reg <= w_data_i[1549];
      mem_3148_sv2v_reg <= w_data_i[1548];
      mem_3147_sv2v_reg <= w_data_i[1547];
      mem_3146_sv2v_reg <= w_data_i[1546];
      mem_3145_sv2v_reg <= w_data_i[1545];
      mem_3144_sv2v_reg <= w_data_i[1544];
      mem_3143_sv2v_reg <= w_data_i[1543];
      mem_3142_sv2v_reg <= w_data_i[1542];
      mem_3141_sv2v_reg <= w_data_i[1541];
      mem_3140_sv2v_reg <= w_data_i[1540];
      mem_3139_sv2v_reg <= w_data_i[1539];
      mem_3138_sv2v_reg <= w_data_i[1538];
      mem_3137_sv2v_reg <= w_data_i[1537];
      mem_3136_sv2v_reg <= w_data_i[1536];
      mem_3135_sv2v_reg <= w_data_i[1535];
      mem_3134_sv2v_reg <= w_data_i[1534];
      mem_3133_sv2v_reg <= w_data_i[1533];
      mem_3132_sv2v_reg <= w_data_i[1532];
      mem_3131_sv2v_reg <= w_data_i[1531];
      mem_3130_sv2v_reg <= w_data_i[1530];
      mem_3129_sv2v_reg <= w_data_i[1529];
      mem_3128_sv2v_reg <= w_data_i[1528];
      mem_3127_sv2v_reg <= w_data_i[1527];
      mem_3126_sv2v_reg <= w_data_i[1526];
      mem_3125_sv2v_reg <= w_data_i[1525];
      mem_3124_sv2v_reg <= w_data_i[1524];
      mem_3123_sv2v_reg <= w_data_i[1523];
      mem_3122_sv2v_reg <= w_data_i[1522];
      mem_3121_sv2v_reg <= w_data_i[1521];
      mem_3120_sv2v_reg <= w_data_i[1520];
      mem_3119_sv2v_reg <= w_data_i[1519];
      mem_3118_sv2v_reg <= w_data_i[1518];
      mem_3117_sv2v_reg <= w_data_i[1517];
      mem_3116_sv2v_reg <= w_data_i[1516];
      mem_3115_sv2v_reg <= w_data_i[1515];
      mem_3114_sv2v_reg <= w_data_i[1514];
      mem_3113_sv2v_reg <= w_data_i[1513];
      mem_3112_sv2v_reg <= w_data_i[1512];
      mem_3111_sv2v_reg <= w_data_i[1511];
      mem_3110_sv2v_reg <= w_data_i[1510];
      mem_3109_sv2v_reg <= w_data_i[1509];
      mem_3108_sv2v_reg <= w_data_i[1508];
      mem_3107_sv2v_reg <= w_data_i[1507];
      mem_3106_sv2v_reg <= w_data_i[1506];
      mem_3105_sv2v_reg <= w_data_i[1505];
      mem_3104_sv2v_reg <= w_data_i[1504];
      mem_3103_sv2v_reg <= w_data_i[1503];
      mem_3102_sv2v_reg <= w_data_i[1502];
      mem_3101_sv2v_reg <= w_data_i[1501];
      mem_1600_sv2v_reg <= w_data_i[0];
    end 
    if(N24) begin
      mem_3100_sv2v_reg <= w_data_i[1500];
      mem_3099_sv2v_reg <= w_data_i[1499];
      mem_3098_sv2v_reg <= w_data_i[1498];
      mem_3097_sv2v_reg <= w_data_i[1497];
      mem_3096_sv2v_reg <= w_data_i[1496];
      mem_3095_sv2v_reg <= w_data_i[1495];
      mem_3094_sv2v_reg <= w_data_i[1494];
      mem_3093_sv2v_reg <= w_data_i[1493];
      mem_3092_sv2v_reg <= w_data_i[1492];
      mem_3091_sv2v_reg <= w_data_i[1491];
      mem_3090_sv2v_reg <= w_data_i[1490];
      mem_3089_sv2v_reg <= w_data_i[1489];
      mem_3088_sv2v_reg <= w_data_i[1488];
      mem_3087_sv2v_reg <= w_data_i[1487];
      mem_3086_sv2v_reg <= w_data_i[1486];
      mem_3085_sv2v_reg <= w_data_i[1485];
      mem_3084_sv2v_reg <= w_data_i[1484];
      mem_3083_sv2v_reg <= w_data_i[1483];
      mem_3082_sv2v_reg <= w_data_i[1482];
      mem_3081_sv2v_reg <= w_data_i[1481];
      mem_3080_sv2v_reg <= w_data_i[1480];
      mem_3079_sv2v_reg <= w_data_i[1479];
      mem_3078_sv2v_reg <= w_data_i[1478];
      mem_3077_sv2v_reg <= w_data_i[1477];
      mem_3076_sv2v_reg <= w_data_i[1476];
      mem_3075_sv2v_reg <= w_data_i[1475];
      mem_3074_sv2v_reg <= w_data_i[1474];
      mem_3073_sv2v_reg <= w_data_i[1473];
      mem_3072_sv2v_reg <= w_data_i[1472];
      mem_3071_sv2v_reg <= w_data_i[1471];
      mem_3070_sv2v_reg <= w_data_i[1470];
      mem_3069_sv2v_reg <= w_data_i[1469];
      mem_3068_sv2v_reg <= w_data_i[1468];
      mem_3067_sv2v_reg <= w_data_i[1467];
      mem_3066_sv2v_reg <= w_data_i[1466];
      mem_3065_sv2v_reg <= w_data_i[1465];
      mem_3064_sv2v_reg <= w_data_i[1464];
      mem_3063_sv2v_reg <= w_data_i[1463];
      mem_3062_sv2v_reg <= w_data_i[1462];
      mem_3061_sv2v_reg <= w_data_i[1461];
      mem_3060_sv2v_reg <= w_data_i[1460];
      mem_3059_sv2v_reg <= w_data_i[1459];
      mem_3058_sv2v_reg <= w_data_i[1458];
      mem_3057_sv2v_reg <= w_data_i[1457];
      mem_3056_sv2v_reg <= w_data_i[1456];
      mem_3055_sv2v_reg <= w_data_i[1455];
      mem_3054_sv2v_reg <= w_data_i[1454];
      mem_3053_sv2v_reg <= w_data_i[1453];
      mem_3052_sv2v_reg <= w_data_i[1452];
      mem_3051_sv2v_reg <= w_data_i[1451];
      mem_3050_sv2v_reg <= w_data_i[1450];
      mem_3049_sv2v_reg <= w_data_i[1449];
      mem_3048_sv2v_reg <= w_data_i[1448];
      mem_3047_sv2v_reg <= w_data_i[1447];
      mem_3046_sv2v_reg <= w_data_i[1446];
      mem_3045_sv2v_reg <= w_data_i[1445];
      mem_3044_sv2v_reg <= w_data_i[1444];
      mem_3043_sv2v_reg <= w_data_i[1443];
      mem_3042_sv2v_reg <= w_data_i[1442];
      mem_3041_sv2v_reg <= w_data_i[1441];
      mem_3040_sv2v_reg <= w_data_i[1440];
      mem_3039_sv2v_reg <= w_data_i[1439];
      mem_3038_sv2v_reg <= w_data_i[1438];
      mem_3037_sv2v_reg <= w_data_i[1437];
      mem_3036_sv2v_reg <= w_data_i[1436];
      mem_3035_sv2v_reg <= w_data_i[1435];
      mem_3034_sv2v_reg <= w_data_i[1434];
      mem_3033_sv2v_reg <= w_data_i[1433];
      mem_3032_sv2v_reg <= w_data_i[1432];
      mem_3031_sv2v_reg <= w_data_i[1431];
      mem_3030_sv2v_reg <= w_data_i[1430];
      mem_3029_sv2v_reg <= w_data_i[1429];
      mem_3028_sv2v_reg <= w_data_i[1428];
      mem_3027_sv2v_reg <= w_data_i[1427];
      mem_3026_sv2v_reg <= w_data_i[1426];
      mem_3025_sv2v_reg <= w_data_i[1425];
      mem_3024_sv2v_reg <= w_data_i[1424];
      mem_3023_sv2v_reg <= w_data_i[1423];
      mem_3022_sv2v_reg <= w_data_i[1422];
      mem_3021_sv2v_reg <= w_data_i[1421];
      mem_3020_sv2v_reg <= w_data_i[1420];
      mem_3019_sv2v_reg <= w_data_i[1419];
      mem_3018_sv2v_reg <= w_data_i[1418];
      mem_3017_sv2v_reg <= w_data_i[1417];
      mem_3016_sv2v_reg <= w_data_i[1416];
      mem_3015_sv2v_reg <= w_data_i[1415];
      mem_3014_sv2v_reg <= w_data_i[1414];
      mem_3013_sv2v_reg <= w_data_i[1413];
      mem_3012_sv2v_reg <= w_data_i[1412];
      mem_3011_sv2v_reg <= w_data_i[1411];
      mem_3010_sv2v_reg <= w_data_i[1410];
      mem_3009_sv2v_reg <= w_data_i[1409];
      mem_3008_sv2v_reg <= w_data_i[1408];
      mem_3007_sv2v_reg <= w_data_i[1407];
      mem_3006_sv2v_reg <= w_data_i[1406];
      mem_3005_sv2v_reg <= w_data_i[1405];
      mem_3004_sv2v_reg <= w_data_i[1404];
      mem_3003_sv2v_reg <= w_data_i[1403];
      mem_3002_sv2v_reg <= w_data_i[1402];
      mem_1601_sv2v_reg <= w_data_i[1];
    end 
    if(N25) begin
      mem_3001_sv2v_reg <= w_data_i[1401];
      mem_3000_sv2v_reg <= w_data_i[1400];
      mem_2999_sv2v_reg <= w_data_i[1399];
      mem_2998_sv2v_reg <= w_data_i[1398];
      mem_2997_sv2v_reg <= w_data_i[1397];
      mem_2996_sv2v_reg <= w_data_i[1396];
      mem_2995_sv2v_reg <= w_data_i[1395];
      mem_2994_sv2v_reg <= w_data_i[1394];
      mem_2993_sv2v_reg <= w_data_i[1393];
      mem_2992_sv2v_reg <= w_data_i[1392];
      mem_2991_sv2v_reg <= w_data_i[1391];
      mem_2990_sv2v_reg <= w_data_i[1390];
      mem_2989_sv2v_reg <= w_data_i[1389];
      mem_2988_sv2v_reg <= w_data_i[1388];
      mem_2987_sv2v_reg <= w_data_i[1387];
      mem_2986_sv2v_reg <= w_data_i[1386];
      mem_2985_sv2v_reg <= w_data_i[1385];
      mem_2984_sv2v_reg <= w_data_i[1384];
      mem_2983_sv2v_reg <= w_data_i[1383];
      mem_2982_sv2v_reg <= w_data_i[1382];
      mem_2981_sv2v_reg <= w_data_i[1381];
      mem_2980_sv2v_reg <= w_data_i[1380];
      mem_2979_sv2v_reg <= w_data_i[1379];
      mem_2978_sv2v_reg <= w_data_i[1378];
      mem_2977_sv2v_reg <= w_data_i[1377];
      mem_2976_sv2v_reg <= w_data_i[1376];
      mem_2975_sv2v_reg <= w_data_i[1375];
      mem_2974_sv2v_reg <= w_data_i[1374];
      mem_2973_sv2v_reg <= w_data_i[1373];
      mem_2972_sv2v_reg <= w_data_i[1372];
      mem_2971_sv2v_reg <= w_data_i[1371];
      mem_2970_sv2v_reg <= w_data_i[1370];
      mem_2969_sv2v_reg <= w_data_i[1369];
      mem_2968_sv2v_reg <= w_data_i[1368];
      mem_2967_sv2v_reg <= w_data_i[1367];
      mem_2966_sv2v_reg <= w_data_i[1366];
      mem_2965_sv2v_reg <= w_data_i[1365];
      mem_2964_sv2v_reg <= w_data_i[1364];
      mem_2963_sv2v_reg <= w_data_i[1363];
      mem_2962_sv2v_reg <= w_data_i[1362];
      mem_2961_sv2v_reg <= w_data_i[1361];
      mem_2960_sv2v_reg <= w_data_i[1360];
      mem_2959_sv2v_reg <= w_data_i[1359];
      mem_2958_sv2v_reg <= w_data_i[1358];
      mem_2957_sv2v_reg <= w_data_i[1357];
      mem_2956_sv2v_reg <= w_data_i[1356];
      mem_2955_sv2v_reg <= w_data_i[1355];
      mem_2954_sv2v_reg <= w_data_i[1354];
      mem_2953_sv2v_reg <= w_data_i[1353];
      mem_2952_sv2v_reg <= w_data_i[1352];
      mem_2951_sv2v_reg <= w_data_i[1351];
      mem_2950_sv2v_reg <= w_data_i[1350];
      mem_2949_sv2v_reg <= w_data_i[1349];
      mem_2948_sv2v_reg <= w_data_i[1348];
      mem_2947_sv2v_reg <= w_data_i[1347];
      mem_2946_sv2v_reg <= w_data_i[1346];
      mem_2945_sv2v_reg <= w_data_i[1345];
      mem_2944_sv2v_reg <= w_data_i[1344];
      mem_2943_sv2v_reg <= w_data_i[1343];
      mem_2942_sv2v_reg <= w_data_i[1342];
      mem_2941_sv2v_reg <= w_data_i[1341];
      mem_2940_sv2v_reg <= w_data_i[1340];
      mem_2939_sv2v_reg <= w_data_i[1339];
      mem_2938_sv2v_reg <= w_data_i[1338];
      mem_2937_sv2v_reg <= w_data_i[1337];
      mem_2936_sv2v_reg <= w_data_i[1336];
      mem_2935_sv2v_reg <= w_data_i[1335];
      mem_2934_sv2v_reg <= w_data_i[1334];
      mem_2933_sv2v_reg <= w_data_i[1333];
      mem_2932_sv2v_reg <= w_data_i[1332];
      mem_2931_sv2v_reg <= w_data_i[1331];
      mem_2930_sv2v_reg <= w_data_i[1330];
      mem_2929_sv2v_reg <= w_data_i[1329];
      mem_2928_sv2v_reg <= w_data_i[1328];
      mem_2927_sv2v_reg <= w_data_i[1327];
      mem_2926_sv2v_reg <= w_data_i[1326];
      mem_2925_sv2v_reg <= w_data_i[1325];
      mem_2924_sv2v_reg <= w_data_i[1324];
      mem_2923_sv2v_reg <= w_data_i[1323];
      mem_2922_sv2v_reg <= w_data_i[1322];
      mem_2921_sv2v_reg <= w_data_i[1321];
      mem_2920_sv2v_reg <= w_data_i[1320];
      mem_2919_sv2v_reg <= w_data_i[1319];
      mem_2918_sv2v_reg <= w_data_i[1318];
      mem_2917_sv2v_reg <= w_data_i[1317];
      mem_2916_sv2v_reg <= w_data_i[1316];
      mem_2915_sv2v_reg <= w_data_i[1315];
      mem_2914_sv2v_reg <= w_data_i[1314];
      mem_2913_sv2v_reg <= w_data_i[1313];
      mem_2912_sv2v_reg <= w_data_i[1312];
      mem_2911_sv2v_reg <= w_data_i[1311];
      mem_2910_sv2v_reg <= w_data_i[1310];
      mem_2909_sv2v_reg <= w_data_i[1309];
      mem_2908_sv2v_reg <= w_data_i[1308];
      mem_2907_sv2v_reg <= w_data_i[1307];
      mem_2906_sv2v_reg <= w_data_i[1306];
      mem_2905_sv2v_reg <= w_data_i[1305];
      mem_2904_sv2v_reg <= w_data_i[1304];
      mem_2903_sv2v_reg <= w_data_i[1303];
      mem_1602_sv2v_reg <= w_data_i[2];
    end 
    if(N26) begin
      mem_2902_sv2v_reg <= w_data_i[1302];
      mem_2901_sv2v_reg <= w_data_i[1301];
      mem_2900_sv2v_reg <= w_data_i[1300];
      mem_2899_sv2v_reg <= w_data_i[1299];
      mem_2898_sv2v_reg <= w_data_i[1298];
      mem_2897_sv2v_reg <= w_data_i[1297];
      mem_2896_sv2v_reg <= w_data_i[1296];
      mem_2895_sv2v_reg <= w_data_i[1295];
      mem_2894_sv2v_reg <= w_data_i[1294];
      mem_2893_sv2v_reg <= w_data_i[1293];
      mem_2892_sv2v_reg <= w_data_i[1292];
      mem_2891_sv2v_reg <= w_data_i[1291];
      mem_2890_sv2v_reg <= w_data_i[1290];
      mem_2889_sv2v_reg <= w_data_i[1289];
      mem_2888_sv2v_reg <= w_data_i[1288];
      mem_2887_sv2v_reg <= w_data_i[1287];
      mem_2886_sv2v_reg <= w_data_i[1286];
      mem_2885_sv2v_reg <= w_data_i[1285];
      mem_2884_sv2v_reg <= w_data_i[1284];
      mem_2883_sv2v_reg <= w_data_i[1283];
      mem_2882_sv2v_reg <= w_data_i[1282];
      mem_2881_sv2v_reg <= w_data_i[1281];
      mem_2880_sv2v_reg <= w_data_i[1280];
      mem_2879_sv2v_reg <= w_data_i[1279];
      mem_2878_sv2v_reg <= w_data_i[1278];
      mem_2877_sv2v_reg <= w_data_i[1277];
      mem_2876_sv2v_reg <= w_data_i[1276];
      mem_2875_sv2v_reg <= w_data_i[1275];
      mem_2874_sv2v_reg <= w_data_i[1274];
      mem_2873_sv2v_reg <= w_data_i[1273];
      mem_2872_sv2v_reg <= w_data_i[1272];
      mem_2871_sv2v_reg <= w_data_i[1271];
      mem_2870_sv2v_reg <= w_data_i[1270];
      mem_2869_sv2v_reg <= w_data_i[1269];
      mem_2868_sv2v_reg <= w_data_i[1268];
      mem_2867_sv2v_reg <= w_data_i[1267];
      mem_2866_sv2v_reg <= w_data_i[1266];
      mem_2865_sv2v_reg <= w_data_i[1265];
      mem_2864_sv2v_reg <= w_data_i[1264];
      mem_2863_sv2v_reg <= w_data_i[1263];
      mem_2862_sv2v_reg <= w_data_i[1262];
      mem_2861_sv2v_reg <= w_data_i[1261];
      mem_2860_sv2v_reg <= w_data_i[1260];
      mem_2859_sv2v_reg <= w_data_i[1259];
      mem_2858_sv2v_reg <= w_data_i[1258];
      mem_2857_sv2v_reg <= w_data_i[1257];
      mem_2856_sv2v_reg <= w_data_i[1256];
      mem_2855_sv2v_reg <= w_data_i[1255];
      mem_2854_sv2v_reg <= w_data_i[1254];
      mem_2853_sv2v_reg <= w_data_i[1253];
      mem_2852_sv2v_reg <= w_data_i[1252];
      mem_2851_sv2v_reg <= w_data_i[1251];
      mem_2850_sv2v_reg <= w_data_i[1250];
      mem_2849_sv2v_reg <= w_data_i[1249];
      mem_2848_sv2v_reg <= w_data_i[1248];
      mem_2847_sv2v_reg <= w_data_i[1247];
      mem_2846_sv2v_reg <= w_data_i[1246];
      mem_2845_sv2v_reg <= w_data_i[1245];
      mem_2844_sv2v_reg <= w_data_i[1244];
      mem_2843_sv2v_reg <= w_data_i[1243];
      mem_2842_sv2v_reg <= w_data_i[1242];
      mem_2841_sv2v_reg <= w_data_i[1241];
      mem_2840_sv2v_reg <= w_data_i[1240];
      mem_2839_sv2v_reg <= w_data_i[1239];
      mem_2838_sv2v_reg <= w_data_i[1238];
      mem_2837_sv2v_reg <= w_data_i[1237];
      mem_2836_sv2v_reg <= w_data_i[1236];
      mem_2835_sv2v_reg <= w_data_i[1235];
      mem_2834_sv2v_reg <= w_data_i[1234];
      mem_2833_sv2v_reg <= w_data_i[1233];
      mem_2832_sv2v_reg <= w_data_i[1232];
      mem_2831_sv2v_reg <= w_data_i[1231];
      mem_2830_sv2v_reg <= w_data_i[1230];
      mem_2829_sv2v_reg <= w_data_i[1229];
      mem_2828_sv2v_reg <= w_data_i[1228];
      mem_2827_sv2v_reg <= w_data_i[1227];
      mem_2826_sv2v_reg <= w_data_i[1226];
      mem_2825_sv2v_reg <= w_data_i[1225];
      mem_2824_sv2v_reg <= w_data_i[1224];
      mem_2823_sv2v_reg <= w_data_i[1223];
      mem_2822_sv2v_reg <= w_data_i[1222];
      mem_2821_sv2v_reg <= w_data_i[1221];
      mem_2820_sv2v_reg <= w_data_i[1220];
      mem_2819_sv2v_reg <= w_data_i[1219];
      mem_2818_sv2v_reg <= w_data_i[1218];
      mem_2817_sv2v_reg <= w_data_i[1217];
      mem_2816_sv2v_reg <= w_data_i[1216];
      mem_2815_sv2v_reg <= w_data_i[1215];
      mem_2814_sv2v_reg <= w_data_i[1214];
      mem_2813_sv2v_reg <= w_data_i[1213];
      mem_2812_sv2v_reg <= w_data_i[1212];
      mem_2811_sv2v_reg <= w_data_i[1211];
      mem_2810_sv2v_reg <= w_data_i[1210];
      mem_2809_sv2v_reg <= w_data_i[1209];
      mem_2808_sv2v_reg <= w_data_i[1208];
      mem_2807_sv2v_reg <= w_data_i[1207];
      mem_2806_sv2v_reg <= w_data_i[1206];
      mem_2805_sv2v_reg <= w_data_i[1205];
      mem_2804_sv2v_reg <= w_data_i[1204];
      mem_1603_sv2v_reg <= w_data_i[3];
    end 
    if(N27) begin
      mem_2803_sv2v_reg <= w_data_i[1203];
      mem_2802_sv2v_reg <= w_data_i[1202];
      mem_2801_sv2v_reg <= w_data_i[1201];
      mem_2800_sv2v_reg <= w_data_i[1200];
      mem_2799_sv2v_reg <= w_data_i[1199];
      mem_2798_sv2v_reg <= w_data_i[1198];
      mem_2797_sv2v_reg <= w_data_i[1197];
      mem_2796_sv2v_reg <= w_data_i[1196];
      mem_2795_sv2v_reg <= w_data_i[1195];
      mem_2794_sv2v_reg <= w_data_i[1194];
      mem_2793_sv2v_reg <= w_data_i[1193];
      mem_2792_sv2v_reg <= w_data_i[1192];
      mem_2791_sv2v_reg <= w_data_i[1191];
      mem_2790_sv2v_reg <= w_data_i[1190];
      mem_2789_sv2v_reg <= w_data_i[1189];
      mem_2788_sv2v_reg <= w_data_i[1188];
      mem_2787_sv2v_reg <= w_data_i[1187];
      mem_2786_sv2v_reg <= w_data_i[1186];
      mem_2785_sv2v_reg <= w_data_i[1185];
      mem_2784_sv2v_reg <= w_data_i[1184];
      mem_2783_sv2v_reg <= w_data_i[1183];
      mem_2782_sv2v_reg <= w_data_i[1182];
      mem_2781_sv2v_reg <= w_data_i[1181];
      mem_2780_sv2v_reg <= w_data_i[1180];
      mem_2779_sv2v_reg <= w_data_i[1179];
      mem_2778_sv2v_reg <= w_data_i[1178];
      mem_2777_sv2v_reg <= w_data_i[1177];
      mem_2776_sv2v_reg <= w_data_i[1176];
      mem_2775_sv2v_reg <= w_data_i[1175];
      mem_2774_sv2v_reg <= w_data_i[1174];
      mem_2773_sv2v_reg <= w_data_i[1173];
      mem_2772_sv2v_reg <= w_data_i[1172];
      mem_2771_sv2v_reg <= w_data_i[1171];
      mem_2770_sv2v_reg <= w_data_i[1170];
      mem_2769_sv2v_reg <= w_data_i[1169];
      mem_2768_sv2v_reg <= w_data_i[1168];
      mem_2767_sv2v_reg <= w_data_i[1167];
      mem_2766_sv2v_reg <= w_data_i[1166];
      mem_2765_sv2v_reg <= w_data_i[1165];
      mem_2764_sv2v_reg <= w_data_i[1164];
      mem_2763_sv2v_reg <= w_data_i[1163];
      mem_2762_sv2v_reg <= w_data_i[1162];
      mem_2761_sv2v_reg <= w_data_i[1161];
      mem_2760_sv2v_reg <= w_data_i[1160];
      mem_2759_sv2v_reg <= w_data_i[1159];
      mem_2758_sv2v_reg <= w_data_i[1158];
      mem_2757_sv2v_reg <= w_data_i[1157];
      mem_2756_sv2v_reg <= w_data_i[1156];
      mem_2755_sv2v_reg <= w_data_i[1155];
      mem_2754_sv2v_reg <= w_data_i[1154];
      mem_2753_sv2v_reg <= w_data_i[1153];
      mem_2752_sv2v_reg <= w_data_i[1152];
      mem_2751_sv2v_reg <= w_data_i[1151];
      mem_2750_sv2v_reg <= w_data_i[1150];
      mem_2749_sv2v_reg <= w_data_i[1149];
      mem_2748_sv2v_reg <= w_data_i[1148];
      mem_2747_sv2v_reg <= w_data_i[1147];
      mem_2746_sv2v_reg <= w_data_i[1146];
      mem_2745_sv2v_reg <= w_data_i[1145];
      mem_2744_sv2v_reg <= w_data_i[1144];
      mem_2743_sv2v_reg <= w_data_i[1143];
      mem_2742_sv2v_reg <= w_data_i[1142];
      mem_2741_sv2v_reg <= w_data_i[1141];
      mem_2740_sv2v_reg <= w_data_i[1140];
      mem_2739_sv2v_reg <= w_data_i[1139];
      mem_2738_sv2v_reg <= w_data_i[1138];
      mem_2737_sv2v_reg <= w_data_i[1137];
      mem_2736_sv2v_reg <= w_data_i[1136];
      mem_2735_sv2v_reg <= w_data_i[1135];
      mem_2734_sv2v_reg <= w_data_i[1134];
      mem_2733_sv2v_reg <= w_data_i[1133];
      mem_2732_sv2v_reg <= w_data_i[1132];
      mem_2731_sv2v_reg <= w_data_i[1131];
      mem_2730_sv2v_reg <= w_data_i[1130];
      mem_2729_sv2v_reg <= w_data_i[1129];
      mem_2728_sv2v_reg <= w_data_i[1128];
      mem_2727_sv2v_reg <= w_data_i[1127];
      mem_2726_sv2v_reg <= w_data_i[1126];
      mem_2725_sv2v_reg <= w_data_i[1125];
      mem_2724_sv2v_reg <= w_data_i[1124];
      mem_2723_sv2v_reg <= w_data_i[1123];
      mem_2722_sv2v_reg <= w_data_i[1122];
      mem_2721_sv2v_reg <= w_data_i[1121];
      mem_2720_sv2v_reg <= w_data_i[1120];
      mem_2719_sv2v_reg <= w_data_i[1119];
      mem_2718_sv2v_reg <= w_data_i[1118];
      mem_2717_sv2v_reg <= w_data_i[1117];
      mem_2716_sv2v_reg <= w_data_i[1116];
      mem_2715_sv2v_reg <= w_data_i[1115];
      mem_2714_sv2v_reg <= w_data_i[1114];
      mem_2713_sv2v_reg <= w_data_i[1113];
      mem_2712_sv2v_reg <= w_data_i[1112];
      mem_2711_sv2v_reg <= w_data_i[1111];
      mem_2710_sv2v_reg <= w_data_i[1110];
      mem_2709_sv2v_reg <= w_data_i[1109];
      mem_2708_sv2v_reg <= w_data_i[1108];
      mem_2707_sv2v_reg <= w_data_i[1107];
      mem_2706_sv2v_reg <= w_data_i[1106];
      mem_2705_sv2v_reg <= w_data_i[1105];
      mem_1604_sv2v_reg <= w_data_i[4];
    end 
    if(N28) begin
      mem_2704_sv2v_reg <= w_data_i[1104];
      mem_2703_sv2v_reg <= w_data_i[1103];
      mem_2702_sv2v_reg <= w_data_i[1102];
      mem_2701_sv2v_reg <= w_data_i[1101];
      mem_2700_sv2v_reg <= w_data_i[1100];
      mem_2699_sv2v_reg <= w_data_i[1099];
      mem_2698_sv2v_reg <= w_data_i[1098];
      mem_2697_sv2v_reg <= w_data_i[1097];
      mem_2696_sv2v_reg <= w_data_i[1096];
      mem_2695_sv2v_reg <= w_data_i[1095];
      mem_2694_sv2v_reg <= w_data_i[1094];
      mem_2693_sv2v_reg <= w_data_i[1093];
      mem_2692_sv2v_reg <= w_data_i[1092];
      mem_2691_sv2v_reg <= w_data_i[1091];
      mem_2690_sv2v_reg <= w_data_i[1090];
      mem_2689_sv2v_reg <= w_data_i[1089];
      mem_2688_sv2v_reg <= w_data_i[1088];
      mem_2687_sv2v_reg <= w_data_i[1087];
      mem_2686_sv2v_reg <= w_data_i[1086];
      mem_2685_sv2v_reg <= w_data_i[1085];
      mem_2684_sv2v_reg <= w_data_i[1084];
      mem_2683_sv2v_reg <= w_data_i[1083];
      mem_2682_sv2v_reg <= w_data_i[1082];
      mem_2681_sv2v_reg <= w_data_i[1081];
      mem_2680_sv2v_reg <= w_data_i[1080];
      mem_2679_sv2v_reg <= w_data_i[1079];
      mem_2678_sv2v_reg <= w_data_i[1078];
      mem_2677_sv2v_reg <= w_data_i[1077];
      mem_2676_sv2v_reg <= w_data_i[1076];
      mem_2675_sv2v_reg <= w_data_i[1075];
      mem_2674_sv2v_reg <= w_data_i[1074];
      mem_2673_sv2v_reg <= w_data_i[1073];
      mem_2672_sv2v_reg <= w_data_i[1072];
      mem_2671_sv2v_reg <= w_data_i[1071];
      mem_2670_sv2v_reg <= w_data_i[1070];
      mem_2669_sv2v_reg <= w_data_i[1069];
      mem_2668_sv2v_reg <= w_data_i[1068];
      mem_2667_sv2v_reg <= w_data_i[1067];
      mem_2666_sv2v_reg <= w_data_i[1066];
      mem_2665_sv2v_reg <= w_data_i[1065];
      mem_2664_sv2v_reg <= w_data_i[1064];
      mem_2663_sv2v_reg <= w_data_i[1063];
      mem_2662_sv2v_reg <= w_data_i[1062];
      mem_2661_sv2v_reg <= w_data_i[1061];
      mem_2660_sv2v_reg <= w_data_i[1060];
      mem_2659_sv2v_reg <= w_data_i[1059];
      mem_2658_sv2v_reg <= w_data_i[1058];
      mem_2657_sv2v_reg <= w_data_i[1057];
      mem_2656_sv2v_reg <= w_data_i[1056];
      mem_2655_sv2v_reg <= w_data_i[1055];
      mem_2654_sv2v_reg <= w_data_i[1054];
      mem_2653_sv2v_reg <= w_data_i[1053];
      mem_2652_sv2v_reg <= w_data_i[1052];
      mem_2651_sv2v_reg <= w_data_i[1051];
      mem_2650_sv2v_reg <= w_data_i[1050];
      mem_2649_sv2v_reg <= w_data_i[1049];
      mem_2648_sv2v_reg <= w_data_i[1048];
      mem_2647_sv2v_reg <= w_data_i[1047];
      mem_2646_sv2v_reg <= w_data_i[1046];
      mem_2645_sv2v_reg <= w_data_i[1045];
      mem_2644_sv2v_reg <= w_data_i[1044];
      mem_2643_sv2v_reg <= w_data_i[1043];
      mem_2642_sv2v_reg <= w_data_i[1042];
      mem_2641_sv2v_reg <= w_data_i[1041];
      mem_2640_sv2v_reg <= w_data_i[1040];
      mem_2639_sv2v_reg <= w_data_i[1039];
      mem_2638_sv2v_reg <= w_data_i[1038];
      mem_2637_sv2v_reg <= w_data_i[1037];
      mem_2636_sv2v_reg <= w_data_i[1036];
      mem_2635_sv2v_reg <= w_data_i[1035];
      mem_2634_sv2v_reg <= w_data_i[1034];
      mem_2633_sv2v_reg <= w_data_i[1033];
      mem_2632_sv2v_reg <= w_data_i[1032];
      mem_2631_sv2v_reg <= w_data_i[1031];
      mem_2630_sv2v_reg <= w_data_i[1030];
      mem_2629_sv2v_reg <= w_data_i[1029];
      mem_2628_sv2v_reg <= w_data_i[1028];
      mem_2627_sv2v_reg <= w_data_i[1027];
      mem_2626_sv2v_reg <= w_data_i[1026];
      mem_2625_sv2v_reg <= w_data_i[1025];
      mem_2624_sv2v_reg <= w_data_i[1024];
      mem_2623_sv2v_reg <= w_data_i[1023];
      mem_2622_sv2v_reg <= w_data_i[1022];
      mem_2621_sv2v_reg <= w_data_i[1021];
      mem_2620_sv2v_reg <= w_data_i[1020];
      mem_2619_sv2v_reg <= w_data_i[1019];
      mem_2618_sv2v_reg <= w_data_i[1018];
      mem_2617_sv2v_reg <= w_data_i[1017];
      mem_2616_sv2v_reg <= w_data_i[1016];
      mem_2615_sv2v_reg <= w_data_i[1015];
      mem_2614_sv2v_reg <= w_data_i[1014];
      mem_2613_sv2v_reg <= w_data_i[1013];
      mem_2612_sv2v_reg <= w_data_i[1012];
      mem_2611_sv2v_reg <= w_data_i[1011];
      mem_2610_sv2v_reg <= w_data_i[1010];
      mem_2609_sv2v_reg <= w_data_i[1009];
      mem_2608_sv2v_reg <= w_data_i[1008];
      mem_2607_sv2v_reg <= w_data_i[1007];
      mem_2606_sv2v_reg <= w_data_i[1006];
      mem_1605_sv2v_reg <= w_data_i[5];
    end 
    if(N29) begin
      mem_2605_sv2v_reg <= w_data_i[1005];
      mem_2604_sv2v_reg <= w_data_i[1004];
      mem_2603_sv2v_reg <= w_data_i[1003];
      mem_2602_sv2v_reg <= w_data_i[1002];
      mem_2601_sv2v_reg <= w_data_i[1001];
      mem_2600_sv2v_reg <= w_data_i[1000];
      mem_2599_sv2v_reg <= w_data_i[999];
      mem_2598_sv2v_reg <= w_data_i[998];
      mem_2597_sv2v_reg <= w_data_i[997];
      mem_2596_sv2v_reg <= w_data_i[996];
      mem_2595_sv2v_reg <= w_data_i[995];
      mem_2594_sv2v_reg <= w_data_i[994];
      mem_2593_sv2v_reg <= w_data_i[993];
      mem_2592_sv2v_reg <= w_data_i[992];
      mem_2591_sv2v_reg <= w_data_i[991];
      mem_2590_sv2v_reg <= w_data_i[990];
      mem_2589_sv2v_reg <= w_data_i[989];
      mem_2588_sv2v_reg <= w_data_i[988];
      mem_2587_sv2v_reg <= w_data_i[987];
      mem_2586_sv2v_reg <= w_data_i[986];
      mem_2585_sv2v_reg <= w_data_i[985];
      mem_2584_sv2v_reg <= w_data_i[984];
      mem_2583_sv2v_reg <= w_data_i[983];
      mem_2582_sv2v_reg <= w_data_i[982];
      mem_2581_sv2v_reg <= w_data_i[981];
      mem_2580_sv2v_reg <= w_data_i[980];
      mem_2579_sv2v_reg <= w_data_i[979];
      mem_2578_sv2v_reg <= w_data_i[978];
      mem_2577_sv2v_reg <= w_data_i[977];
      mem_2576_sv2v_reg <= w_data_i[976];
      mem_2575_sv2v_reg <= w_data_i[975];
      mem_2574_sv2v_reg <= w_data_i[974];
      mem_2573_sv2v_reg <= w_data_i[973];
      mem_2572_sv2v_reg <= w_data_i[972];
      mem_2571_sv2v_reg <= w_data_i[971];
      mem_2570_sv2v_reg <= w_data_i[970];
      mem_2569_sv2v_reg <= w_data_i[969];
      mem_2568_sv2v_reg <= w_data_i[968];
      mem_2567_sv2v_reg <= w_data_i[967];
      mem_2566_sv2v_reg <= w_data_i[966];
      mem_2565_sv2v_reg <= w_data_i[965];
      mem_2564_sv2v_reg <= w_data_i[964];
      mem_2563_sv2v_reg <= w_data_i[963];
      mem_2562_sv2v_reg <= w_data_i[962];
      mem_2561_sv2v_reg <= w_data_i[961];
      mem_2560_sv2v_reg <= w_data_i[960];
      mem_2559_sv2v_reg <= w_data_i[959];
      mem_2558_sv2v_reg <= w_data_i[958];
      mem_2557_sv2v_reg <= w_data_i[957];
      mem_2556_sv2v_reg <= w_data_i[956];
      mem_2555_sv2v_reg <= w_data_i[955];
      mem_2554_sv2v_reg <= w_data_i[954];
      mem_2553_sv2v_reg <= w_data_i[953];
      mem_2552_sv2v_reg <= w_data_i[952];
      mem_2551_sv2v_reg <= w_data_i[951];
      mem_2550_sv2v_reg <= w_data_i[950];
      mem_2549_sv2v_reg <= w_data_i[949];
      mem_2548_sv2v_reg <= w_data_i[948];
      mem_2547_sv2v_reg <= w_data_i[947];
      mem_2546_sv2v_reg <= w_data_i[946];
      mem_2545_sv2v_reg <= w_data_i[945];
      mem_2544_sv2v_reg <= w_data_i[944];
      mem_2543_sv2v_reg <= w_data_i[943];
      mem_2542_sv2v_reg <= w_data_i[942];
      mem_2541_sv2v_reg <= w_data_i[941];
      mem_2540_sv2v_reg <= w_data_i[940];
      mem_2539_sv2v_reg <= w_data_i[939];
      mem_2538_sv2v_reg <= w_data_i[938];
      mem_2537_sv2v_reg <= w_data_i[937];
      mem_2536_sv2v_reg <= w_data_i[936];
      mem_2535_sv2v_reg <= w_data_i[935];
      mem_2534_sv2v_reg <= w_data_i[934];
      mem_2533_sv2v_reg <= w_data_i[933];
      mem_2532_sv2v_reg <= w_data_i[932];
      mem_2531_sv2v_reg <= w_data_i[931];
      mem_2530_sv2v_reg <= w_data_i[930];
      mem_2529_sv2v_reg <= w_data_i[929];
      mem_2528_sv2v_reg <= w_data_i[928];
      mem_2527_sv2v_reg <= w_data_i[927];
      mem_2526_sv2v_reg <= w_data_i[926];
      mem_2525_sv2v_reg <= w_data_i[925];
      mem_2524_sv2v_reg <= w_data_i[924];
      mem_2523_sv2v_reg <= w_data_i[923];
      mem_2522_sv2v_reg <= w_data_i[922];
      mem_2521_sv2v_reg <= w_data_i[921];
      mem_2520_sv2v_reg <= w_data_i[920];
      mem_2519_sv2v_reg <= w_data_i[919];
      mem_2518_sv2v_reg <= w_data_i[918];
      mem_2517_sv2v_reg <= w_data_i[917];
      mem_2516_sv2v_reg <= w_data_i[916];
      mem_2515_sv2v_reg <= w_data_i[915];
      mem_2514_sv2v_reg <= w_data_i[914];
      mem_2513_sv2v_reg <= w_data_i[913];
      mem_2512_sv2v_reg <= w_data_i[912];
      mem_2511_sv2v_reg <= w_data_i[911];
      mem_2510_sv2v_reg <= w_data_i[910];
      mem_2509_sv2v_reg <= w_data_i[909];
      mem_2508_sv2v_reg <= w_data_i[908];
      mem_2507_sv2v_reg <= w_data_i[907];
      mem_1606_sv2v_reg <= w_data_i[6];
    end 
    if(N30) begin
      mem_2506_sv2v_reg <= w_data_i[906];
      mem_2505_sv2v_reg <= w_data_i[905];
      mem_2504_sv2v_reg <= w_data_i[904];
      mem_2503_sv2v_reg <= w_data_i[903];
      mem_2502_sv2v_reg <= w_data_i[902];
      mem_2501_sv2v_reg <= w_data_i[901];
      mem_2500_sv2v_reg <= w_data_i[900];
      mem_2499_sv2v_reg <= w_data_i[899];
      mem_2498_sv2v_reg <= w_data_i[898];
      mem_2497_sv2v_reg <= w_data_i[897];
      mem_2496_sv2v_reg <= w_data_i[896];
      mem_2495_sv2v_reg <= w_data_i[895];
      mem_2494_sv2v_reg <= w_data_i[894];
      mem_2493_sv2v_reg <= w_data_i[893];
      mem_2492_sv2v_reg <= w_data_i[892];
      mem_2491_sv2v_reg <= w_data_i[891];
      mem_2490_sv2v_reg <= w_data_i[890];
      mem_2489_sv2v_reg <= w_data_i[889];
      mem_2488_sv2v_reg <= w_data_i[888];
      mem_2487_sv2v_reg <= w_data_i[887];
      mem_2486_sv2v_reg <= w_data_i[886];
      mem_2485_sv2v_reg <= w_data_i[885];
      mem_2484_sv2v_reg <= w_data_i[884];
      mem_2483_sv2v_reg <= w_data_i[883];
      mem_2482_sv2v_reg <= w_data_i[882];
      mem_2481_sv2v_reg <= w_data_i[881];
      mem_2480_sv2v_reg <= w_data_i[880];
      mem_2479_sv2v_reg <= w_data_i[879];
      mem_2478_sv2v_reg <= w_data_i[878];
      mem_2477_sv2v_reg <= w_data_i[877];
      mem_2476_sv2v_reg <= w_data_i[876];
      mem_2475_sv2v_reg <= w_data_i[875];
      mem_2474_sv2v_reg <= w_data_i[874];
      mem_2473_sv2v_reg <= w_data_i[873];
      mem_2472_sv2v_reg <= w_data_i[872];
      mem_2471_sv2v_reg <= w_data_i[871];
      mem_2470_sv2v_reg <= w_data_i[870];
      mem_2469_sv2v_reg <= w_data_i[869];
      mem_2468_sv2v_reg <= w_data_i[868];
      mem_2467_sv2v_reg <= w_data_i[867];
      mem_2466_sv2v_reg <= w_data_i[866];
      mem_2465_sv2v_reg <= w_data_i[865];
      mem_2464_sv2v_reg <= w_data_i[864];
      mem_2463_sv2v_reg <= w_data_i[863];
      mem_2462_sv2v_reg <= w_data_i[862];
      mem_2461_sv2v_reg <= w_data_i[861];
      mem_2460_sv2v_reg <= w_data_i[860];
      mem_2459_sv2v_reg <= w_data_i[859];
      mem_2458_sv2v_reg <= w_data_i[858];
      mem_2457_sv2v_reg <= w_data_i[857];
      mem_2456_sv2v_reg <= w_data_i[856];
      mem_2455_sv2v_reg <= w_data_i[855];
      mem_2454_sv2v_reg <= w_data_i[854];
      mem_2453_sv2v_reg <= w_data_i[853];
      mem_2452_sv2v_reg <= w_data_i[852];
      mem_2451_sv2v_reg <= w_data_i[851];
      mem_2450_sv2v_reg <= w_data_i[850];
      mem_2449_sv2v_reg <= w_data_i[849];
      mem_2448_sv2v_reg <= w_data_i[848];
      mem_2447_sv2v_reg <= w_data_i[847];
      mem_2446_sv2v_reg <= w_data_i[846];
      mem_2445_sv2v_reg <= w_data_i[845];
      mem_2444_sv2v_reg <= w_data_i[844];
      mem_2443_sv2v_reg <= w_data_i[843];
      mem_2442_sv2v_reg <= w_data_i[842];
      mem_2441_sv2v_reg <= w_data_i[841];
      mem_2440_sv2v_reg <= w_data_i[840];
      mem_2439_sv2v_reg <= w_data_i[839];
      mem_2438_sv2v_reg <= w_data_i[838];
      mem_2437_sv2v_reg <= w_data_i[837];
      mem_2436_sv2v_reg <= w_data_i[836];
      mem_2435_sv2v_reg <= w_data_i[835];
      mem_2434_sv2v_reg <= w_data_i[834];
      mem_2433_sv2v_reg <= w_data_i[833];
      mem_2432_sv2v_reg <= w_data_i[832];
      mem_2431_sv2v_reg <= w_data_i[831];
      mem_2430_sv2v_reg <= w_data_i[830];
      mem_2429_sv2v_reg <= w_data_i[829];
      mem_2428_sv2v_reg <= w_data_i[828];
      mem_2427_sv2v_reg <= w_data_i[827];
      mem_2426_sv2v_reg <= w_data_i[826];
      mem_2425_sv2v_reg <= w_data_i[825];
      mem_2424_sv2v_reg <= w_data_i[824];
      mem_2423_sv2v_reg <= w_data_i[823];
      mem_2422_sv2v_reg <= w_data_i[822];
      mem_2421_sv2v_reg <= w_data_i[821];
      mem_2420_sv2v_reg <= w_data_i[820];
      mem_2419_sv2v_reg <= w_data_i[819];
      mem_2418_sv2v_reg <= w_data_i[818];
      mem_2417_sv2v_reg <= w_data_i[817];
      mem_2416_sv2v_reg <= w_data_i[816];
      mem_2415_sv2v_reg <= w_data_i[815];
      mem_2414_sv2v_reg <= w_data_i[814];
      mem_2413_sv2v_reg <= w_data_i[813];
      mem_2412_sv2v_reg <= w_data_i[812];
      mem_2411_sv2v_reg <= w_data_i[811];
      mem_2410_sv2v_reg <= w_data_i[810];
      mem_2409_sv2v_reg <= w_data_i[809];
      mem_2408_sv2v_reg <= w_data_i[808];
      mem_1607_sv2v_reg <= w_data_i[7];
    end 
    if(N31) begin
      mem_2407_sv2v_reg <= w_data_i[807];
      mem_2406_sv2v_reg <= w_data_i[806];
      mem_2405_sv2v_reg <= w_data_i[805];
      mem_2404_sv2v_reg <= w_data_i[804];
      mem_2403_sv2v_reg <= w_data_i[803];
      mem_2402_sv2v_reg <= w_data_i[802];
      mem_2401_sv2v_reg <= w_data_i[801];
      mem_2400_sv2v_reg <= w_data_i[800];
      mem_2399_sv2v_reg <= w_data_i[799];
      mem_2398_sv2v_reg <= w_data_i[798];
      mem_2397_sv2v_reg <= w_data_i[797];
      mem_2396_sv2v_reg <= w_data_i[796];
      mem_2395_sv2v_reg <= w_data_i[795];
      mem_2394_sv2v_reg <= w_data_i[794];
      mem_2393_sv2v_reg <= w_data_i[793];
      mem_2392_sv2v_reg <= w_data_i[792];
      mem_2391_sv2v_reg <= w_data_i[791];
      mem_2390_sv2v_reg <= w_data_i[790];
      mem_2389_sv2v_reg <= w_data_i[789];
      mem_2388_sv2v_reg <= w_data_i[788];
      mem_2387_sv2v_reg <= w_data_i[787];
      mem_2386_sv2v_reg <= w_data_i[786];
      mem_2385_sv2v_reg <= w_data_i[785];
      mem_2384_sv2v_reg <= w_data_i[784];
      mem_2383_sv2v_reg <= w_data_i[783];
      mem_2382_sv2v_reg <= w_data_i[782];
      mem_2381_sv2v_reg <= w_data_i[781];
      mem_2380_sv2v_reg <= w_data_i[780];
      mem_2379_sv2v_reg <= w_data_i[779];
      mem_2378_sv2v_reg <= w_data_i[778];
      mem_2377_sv2v_reg <= w_data_i[777];
      mem_2376_sv2v_reg <= w_data_i[776];
      mem_2375_sv2v_reg <= w_data_i[775];
      mem_2374_sv2v_reg <= w_data_i[774];
      mem_2373_sv2v_reg <= w_data_i[773];
      mem_2372_sv2v_reg <= w_data_i[772];
      mem_2371_sv2v_reg <= w_data_i[771];
      mem_2370_sv2v_reg <= w_data_i[770];
      mem_2369_sv2v_reg <= w_data_i[769];
      mem_2368_sv2v_reg <= w_data_i[768];
      mem_2367_sv2v_reg <= w_data_i[767];
      mem_2366_sv2v_reg <= w_data_i[766];
      mem_2365_sv2v_reg <= w_data_i[765];
      mem_2364_sv2v_reg <= w_data_i[764];
      mem_2363_sv2v_reg <= w_data_i[763];
      mem_2362_sv2v_reg <= w_data_i[762];
      mem_2361_sv2v_reg <= w_data_i[761];
      mem_2360_sv2v_reg <= w_data_i[760];
      mem_2359_sv2v_reg <= w_data_i[759];
      mem_2358_sv2v_reg <= w_data_i[758];
      mem_2357_sv2v_reg <= w_data_i[757];
      mem_2356_sv2v_reg <= w_data_i[756];
      mem_2355_sv2v_reg <= w_data_i[755];
      mem_2354_sv2v_reg <= w_data_i[754];
      mem_2353_sv2v_reg <= w_data_i[753];
      mem_2352_sv2v_reg <= w_data_i[752];
      mem_2351_sv2v_reg <= w_data_i[751];
      mem_2350_sv2v_reg <= w_data_i[750];
      mem_2349_sv2v_reg <= w_data_i[749];
      mem_2348_sv2v_reg <= w_data_i[748];
      mem_2347_sv2v_reg <= w_data_i[747];
      mem_2346_sv2v_reg <= w_data_i[746];
      mem_2345_sv2v_reg <= w_data_i[745];
      mem_2344_sv2v_reg <= w_data_i[744];
      mem_2343_sv2v_reg <= w_data_i[743];
      mem_2342_sv2v_reg <= w_data_i[742];
      mem_2341_sv2v_reg <= w_data_i[741];
      mem_2340_sv2v_reg <= w_data_i[740];
      mem_2339_sv2v_reg <= w_data_i[739];
      mem_2338_sv2v_reg <= w_data_i[738];
      mem_2337_sv2v_reg <= w_data_i[737];
      mem_2336_sv2v_reg <= w_data_i[736];
      mem_2335_sv2v_reg <= w_data_i[735];
      mem_2334_sv2v_reg <= w_data_i[734];
      mem_2333_sv2v_reg <= w_data_i[733];
      mem_2332_sv2v_reg <= w_data_i[732];
      mem_2331_sv2v_reg <= w_data_i[731];
      mem_2330_sv2v_reg <= w_data_i[730];
      mem_2329_sv2v_reg <= w_data_i[729];
      mem_2328_sv2v_reg <= w_data_i[728];
      mem_2327_sv2v_reg <= w_data_i[727];
      mem_2326_sv2v_reg <= w_data_i[726];
      mem_2325_sv2v_reg <= w_data_i[725];
      mem_2324_sv2v_reg <= w_data_i[724];
      mem_2323_sv2v_reg <= w_data_i[723];
      mem_2322_sv2v_reg <= w_data_i[722];
      mem_2321_sv2v_reg <= w_data_i[721];
      mem_2320_sv2v_reg <= w_data_i[720];
      mem_2319_sv2v_reg <= w_data_i[719];
      mem_2318_sv2v_reg <= w_data_i[718];
      mem_2317_sv2v_reg <= w_data_i[717];
      mem_2316_sv2v_reg <= w_data_i[716];
      mem_2315_sv2v_reg <= w_data_i[715];
      mem_2314_sv2v_reg <= w_data_i[714];
      mem_2313_sv2v_reg <= w_data_i[713];
      mem_2312_sv2v_reg <= w_data_i[712];
      mem_2311_sv2v_reg <= w_data_i[711];
      mem_2310_sv2v_reg <= w_data_i[710];
      mem_2309_sv2v_reg <= w_data_i[709];
      mem_1608_sv2v_reg <= w_data_i[8];
    end 
    if(N32) begin
      mem_2308_sv2v_reg <= w_data_i[708];
      mem_2307_sv2v_reg <= w_data_i[707];
      mem_2306_sv2v_reg <= w_data_i[706];
      mem_2305_sv2v_reg <= w_data_i[705];
      mem_2304_sv2v_reg <= w_data_i[704];
      mem_2303_sv2v_reg <= w_data_i[703];
      mem_2302_sv2v_reg <= w_data_i[702];
      mem_2301_sv2v_reg <= w_data_i[701];
      mem_2300_sv2v_reg <= w_data_i[700];
      mem_2299_sv2v_reg <= w_data_i[699];
      mem_2298_sv2v_reg <= w_data_i[698];
      mem_2297_sv2v_reg <= w_data_i[697];
      mem_2296_sv2v_reg <= w_data_i[696];
      mem_2295_sv2v_reg <= w_data_i[695];
      mem_2294_sv2v_reg <= w_data_i[694];
      mem_2293_sv2v_reg <= w_data_i[693];
      mem_2292_sv2v_reg <= w_data_i[692];
      mem_2291_sv2v_reg <= w_data_i[691];
      mem_2290_sv2v_reg <= w_data_i[690];
      mem_2289_sv2v_reg <= w_data_i[689];
      mem_2288_sv2v_reg <= w_data_i[688];
      mem_2287_sv2v_reg <= w_data_i[687];
      mem_2286_sv2v_reg <= w_data_i[686];
      mem_2285_sv2v_reg <= w_data_i[685];
      mem_2284_sv2v_reg <= w_data_i[684];
      mem_2283_sv2v_reg <= w_data_i[683];
      mem_2282_sv2v_reg <= w_data_i[682];
      mem_2281_sv2v_reg <= w_data_i[681];
      mem_2280_sv2v_reg <= w_data_i[680];
      mem_2279_sv2v_reg <= w_data_i[679];
      mem_2278_sv2v_reg <= w_data_i[678];
      mem_2277_sv2v_reg <= w_data_i[677];
      mem_2276_sv2v_reg <= w_data_i[676];
      mem_2275_sv2v_reg <= w_data_i[675];
      mem_2274_sv2v_reg <= w_data_i[674];
      mem_2273_sv2v_reg <= w_data_i[673];
      mem_2272_sv2v_reg <= w_data_i[672];
      mem_2271_sv2v_reg <= w_data_i[671];
      mem_2270_sv2v_reg <= w_data_i[670];
      mem_2269_sv2v_reg <= w_data_i[669];
      mem_2268_sv2v_reg <= w_data_i[668];
      mem_2267_sv2v_reg <= w_data_i[667];
      mem_2266_sv2v_reg <= w_data_i[666];
      mem_2265_sv2v_reg <= w_data_i[665];
      mem_2264_sv2v_reg <= w_data_i[664];
      mem_2263_sv2v_reg <= w_data_i[663];
      mem_2262_sv2v_reg <= w_data_i[662];
      mem_2261_sv2v_reg <= w_data_i[661];
      mem_2260_sv2v_reg <= w_data_i[660];
      mem_2259_sv2v_reg <= w_data_i[659];
      mem_2258_sv2v_reg <= w_data_i[658];
      mem_2257_sv2v_reg <= w_data_i[657];
      mem_2256_sv2v_reg <= w_data_i[656];
      mem_2255_sv2v_reg <= w_data_i[655];
      mem_2254_sv2v_reg <= w_data_i[654];
      mem_2253_sv2v_reg <= w_data_i[653];
      mem_2252_sv2v_reg <= w_data_i[652];
      mem_2251_sv2v_reg <= w_data_i[651];
      mem_2250_sv2v_reg <= w_data_i[650];
      mem_2249_sv2v_reg <= w_data_i[649];
      mem_2248_sv2v_reg <= w_data_i[648];
      mem_2247_sv2v_reg <= w_data_i[647];
      mem_2246_sv2v_reg <= w_data_i[646];
      mem_2245_sv2v_reg <= w_data_i[645];
      mem_2244_sv2v_reg <= w_data_i[644];
      mem_2243_sv2v_reg <= w_data_i[643];
      mem_2242_sv2v_reg <= w_data_i[642];
      mem_2241_sv2v_reg <= w_data_i[641];
      mem_2240_sv2v_reg <= w_data_i[640];
      mem_2239_sv2v_reg <= w_data_i[639];
      mem_2238_sv2v_reg <= w_data_i[638];
      mem_2237_sv2v_reg <= w_data_i[637];
      mem_2236_sv2v_reg <= w_data_i[636];
      mem_2235_sv2v_reg <= w_data_i[635];
      mem_2234_sv2v_reg <= w_data_i[634];
      mem_2233_sv2v_reg <= w_data_i[633];
      mem_2232_sv2v_reg <= w_data_i[632];
      mem_2231_sv2v_reg <= w_data_i[631];
      mem_2230_sv2v_reg <= w_data_i[630];
      mem_2229_sv2v_reg <= w_data_i[629];
      mem_2228_sv2v_reg <= w_data_i[628];
      mem_2227_sv2v_reg <= w_data_i[627];
      mem_2226_sv2v_reg <= w_data_i[626];
      mem_2225_sv2v_reg <= w_data_i[625];
      mem_2224_sv2v_reg <= w_data_i[624];
      mem_2223_sv2v_reg <= w_data_i[623];
      mem_2222_sv2v_reg <= w_data_i[622];
      mem_2221_sv2v_reg <= w_data_i[621];
      mem_2220_sv2v_reg <= w_data_i[620];
      mem_2219_sv2v_reg <= w_data_i[619];
      mem_2218_sv2v_reg <= w_data_i[618];
      mem_2217_sv2v_reg <= w_data_i[617];
      mem_2216_sv2v_reg <= w_data_i[616];
      mem_2215_sv2v_reg <= w_data_i[615];
      mem_2214_sv2v_reg <= w_data_i[614];
      mem_2213_sv2v_reg <= w_data_i[613];
      mem_2212_sv2v_reg <= w_data_i[612];
      mem_2211_sv2v_reg <= w_data_i[611];
      mem_2210_sv2v_reg <= w_data_i[610];
      mem_1609_sv2v_reg <= w_data_i[9];
    end 
    if(N33) begin
      mem_2209_sv2v_reg <= w_data_i[609];
      mem_2208_sv2v_reg <= w_data_i[608];
      mem_2207_sv2v_reg <= w_data_i[607];
      mem_2206_sv2v_reg <= w_data_i[606];
      mem_2205_sv2v_reg <= w_data_i[605];
      mem_2204_sv2v_reg <= w_data_i[604];
      mem_2203_sv2v_reg <= w_data_i[603];
      mem_2202_sv2v_reg <= w_data_i[602];
      mem_2201_sv2v_reg <= w_data_i[601];
      mem_2200_sv2v_reg <= w_data_i[600];
      mem_2199_sv2v_reg <= w_data_i[599];
      mem_2198_sv2v_reg <= w_data_i[598];
      mem_2197_sv2v_reg <= w_data_i[597];
      mem_2196_sv2v_reg <= w_data_i[596];
      mem_2195_sv2v_reg <= w_data_i[595];
      mem_2194_sv2v_reg <= w_data_i[594];
      mem_2193_sv2v_reg <= w_data_i[593];
      mem_2192_sv2v_reg <= w_data_i[592];
      mem_2191_sv2v_reg <= w_data_i[591];
      mem_2190_sv2v_reg <= w_data_i[590];
      mem_2189_sv2v_reg <= w_data_i[589];
      mem_2188_sv2v_reg <= w_data_i[588];
      mem_2187_sv2v_reg <= w_data_i[587];
      mem_2186_sv2v_reg <= w_data_i[586];
      mem_2185_sv2v_reg <= w_data_i[585];
      mem_2184_sv2v_reg <= w_data_i[584];
      mem_2183_sv2v_reg <= w_data_i[583];
      mem_2182_sv2v_reg <= w_data_i[582];
      mem_2181_sv2v_reg <= w_data_i[581];
      mem_2180_sv2v_reg <= w_data_i[580];
      mem_2179_sv2v_reg <= w_data_i[579];
      mem_2178_sv2v_reg <= w_data_i[578];
      mem_2177_sv2v_reg <= w_data_i[577];
      mem_2176_sv2v_reg <= w_data_i[576];
      mem_2175_sv2v_reg <= w_data_i[575];
      mem_2174_sv2v_reg <= w_data_i[574];
      mem_2173_sv2v_reg <= w_data_i[573];
      mem_2172_sv2v_reg <= w_data_i[572];
      mem_2171_sv2v_reg <= w_data_i[571];
      mem_2170_sv2v_reg <= w_data_i[570];
      mem_2169_sv2v_reg <= w_data_i[569];
      mem_2168_sv2v_reg <= w_data_i[568];
      mem_2167_sv2v_reg <= w_data_i[567];
      mem_2166_sv2v_reg <= w_data_i[566];
      mem_2165_sv2v_reg <= w_data_i[565];
      mem_2164_sv2v_reg <= w_data_i[564];
      mem_2163_sv2v_reg <= w_data_i[563];
      mem_2162_sv2v_reg <= w_data_i[562];
      mem_2161_sv2v_reg <= w_data_i[561];
      mem_2160_sv2v_reg <= w_data_i[560];
      mem_2159_sv2v_reg <= w_data_i[559];
      mem_2158_sv2v_reg <= w_data_i[558];
      mem_2157_sv2v_reg <= w_data_i[557];
      mem_2156_sv2v_reg <= w_data_i[556];
      mem_2155_sv2v_reg <= w_data_i[555];
      mem_2154_sv2v_reg <= w_data_i[554];
      mem_2153_sv2v_reg <= w_data_i[553];
      mem_2152_sv2v_reg <= w_data_i[552];
      mem_2151_sv2v_reg <= w_data_i[551];
      mem_2150_sv2v_reg <= w_data_i[550];
      mem_2149_sv2v_reg <= w_data_i[549];
      mem_2148_sv2v_reg <= w_data_i[548];
      mem_2147_sv2v_reg <= w_data_i[547];
      mem_2146_sv2v_reg <= w_data_i[546];
      mem_2145_sv2v_reg <= w_data_i[545];
      mem_2144_sv2v_reg <= w_data_i[544];
      mem_2143_sv2v_reg <= w_data_i[543];
      mem_2142_sv2v_reg <= w_data_i[542];
      mem_2141_sv2v_reg <= w_data_i[541];
      mem_2140_sv2v_reg <= w_data_i[540];
      mem_2139_sv2v_reg <= w_data_i[539];
      mem_2138_sv2v_reg <= w_data_i[538];
      mem_2137_sv2v_reg <= w_data_i[537];
      mem_2136_sv2v_reg <= w_data_i[536];
      mem_2135_sv2v_reg <= w_data_i[535];
      mem_2134_sv2v_reg <= w_data_i[534];
      mem_2133_sv2v_reg <= w_data_i[533];
      mem_2132_sv2v_reg <= w_data_i[532];
      mem_2131_sv2v_reg <= w_data_i[531];
      mem_2130_sv2v_reg <= w_data_i[530];
      mem_2129_sv2v_reg <= w_data_i[529];
      mem_2128_sv2v_reg <= w_data_i[528];
      mem_2127_sv2v_reg <= w_data_i[527];
      mem_2126_sv2v_reg <= w_data_i[526];
      mem_2125_sv2v_reg <= w_data_i[525];
      mem_2124_sv2v_reg <= w_data_i[524];
      mem_2123_sv2v_reg <= w_data_i[523];
      mem_2122_sv2v_reg <= w_data_i[522];
      mem_2121_sv2v_reg <= w_data_i[521];
      mem_2120_sv2v_reg <= w_data_i[520];
      mem_2119_sv2v_reg <= w_data_i[519];
      mem_2118_sv2v_reg <= w_data_i[518];
      mem_2117_sv2v_reg <= w_data_i[517];
      mem_2116_sv2v_reg <= w_data_i[516];
      mem_2115_sv2v_reg <= w_data_i[515];
      mem_2114_sv2v_reg <= w_data_i[514];
      mem_2113_sv2v_reg <= w_data_i[513];
      mem_2112_sv2v_reg <= w_data_i[512];
      mem_2111_sv2v_reg <= w_data_i[511];
      mem_1610_sv2v_reg <= w_data_i[10];
    end 
    if(N34) begin
      mem_2110_sv2v_reg <= w_data_i[510];
      mem_2109_sv2v_reg <= w_data_i[509];
      mem_2108_sv2v_reg <= w_data_i[508];
      mem_2107_sv2v_reg <= w_data_i[507];
      mem_2106_sv2v_reg <= w_data_i[506];
      mem_2105_sv2v_reg <= w_data_i[505];
      mem_2104_sv2v_reg <= w_data_i[504];
      mem_2103_sv2v_reg <= w_data_i[503];
      mem_2102_sv2v_reg <= w_data_i[502];
      mem_2101_sv2v_reg <= w_data_i[501];
      mem_2100_sv2v_reg <= w_data_i[500];
      mem_2099_sv2v_reg <= w_data_i[499];
      mem_2098_sv2v_reg <= w_data_i[498];
      mem_2097_sv2v_reg <= w_data_i[497];
      mem_2096_sv2v_reg <= w_data_i[496];
      mem_2095_sv2v_reg <= w_data_i[495];
      mem_2094_sv2v_reg <= w_data_i[494];
      mem_2093_sv2v_reg <= w_data_i[493];
      mem_2092_sv2v_reg <= w_data_i[492];
      mem_2091_sv2v_reg <= w_data_i[491];
      mem_2090_sv2v_reg <= w_data_i[490];
      mem_2089_sv2v_reg <= w_data_i[489];
      mem_2088_sv2v_reg <= w_data_i[488];
      mem_2087_sv2v_reg <= w_data_i[487];
      mem_2086_sv2v_reg <= w_data_i[486];
      mem_2085_sv2v_reg <= w_data_i[485];
      mem_2084_sv2v_reg <= w_data_i[484];
      mem_2083_sv2v_reg <= w_data_i[483];
      mem_2082_sv2v_reg <= w_data_i[482];
      mem_2081_sv2v_reg <= w_data_i[481];
      mem_2080_sv2v_reg <= w_data_i[480];
      mem_2079_sv2v_reg <= w_data_i[479];
      mem_2078_sv2v_reg <= w_data_i[478];
      mem_2077_sv2v_reg <= w_data_i[477];
      mem_2076_sv2v_reg <= w_data_i[476];
      mem_2075_sv2v_reg <= w_data_i[475];
      mem_2074_sv2v_reg <= w_data_i[474];
      mem_2073_sv2v_reg <= w_data_i[473];
      mem_2072_sv2v_reg <= w_data_i[472];
      mem_2071_sv2v_reg <= w_data_i[471];
      mem_2070_sv2v_reg <= w_data_i[470];
      mem_2069_sv2v_reg <= w_data_i[469];
      mem_2068_sv2v_reg <= w_data_i[468];
      mem_2067_sv2v_reg <= w_data_i[467];
      mem_2066_sv2v_reg <= w_data_i[466];
      mem_2065_sv2v_reg <= w_data_i[465];
      mem_2064_sv2v_reg <= w_data_i[464];
      mem_2063_sv2v_reg <= w_data_i[463];
      mem_2062_sv2v_reg <= w_data_i[462];
      mem_2061_sv2v_reg <= w_data_i[461];
      mem_2060_sv2v_reg <= w_data_i[460];
      mem_2059_sv2v_reg <= w_data_i[459];
      mem_2058_sv2v_reg <= w_data_i[458];
      mem_2057_sv2v_reg <= w_data_i[457];
      mem_2056_sv2v_reg <= w_data_i[456];
      mem_2055_sv2v_reg <= w_data_i[455];
      mem_2054_sv2v_reg <= w_data_i[454];
      mem_2053_sv2v_reg <= w_data_i[453];
      mem_2052_sv2v_reg <= w_data_i[452];
      mem_2051_sv2v_reg <= w_data_i[451];
      mem_2050_sv2v_reg <= w_data_i[450];
      mem_2049_sv2v_reg <= w_data_i[449];
      mem_2048_sv2v_reg <= w_data_i[448];
      mem_2047_sv2v_reg <= w_data_i[447];
      mem_2046_sv2v_reg <= w_data_i[446];
      mem_2045_sv2v_reg <= w_data_i[445];
      mem_2044_sv2v_reg <= w_data_i[444];
      mem_2043_sv2v_reg <= w_data_i[443];
      mem_2042_sv2v_reg <= w_data_i[442];
      mem_2041_sv2v_reg <= w_data_i[441];
      mem_2040_sv2v_reg <= w_data_i[440];
      mem_2039_sv2v_reg <= w_data_i[439];
      mem_2038_sv2v_reg <= w_data_i[438];
      mem_2037_sv2v_reg <= w_data_i[437];
      mem_2036_sv2v_reg <= w_data_i[436];
      mem_2035_sv2v_reg <= w_data_i[435];
      mem_2034_sv2v_reg <= w_data_i[434];
      mem_2033_sv2v_reg <= w_data_i[433];
      mem_2032_sv2v_reg <= w_data_i[432];
      mem_2031_sv2v_reg <= w_data_i[431];
      mem_2030_sv2v_reg <= w_data_i[430];
      mem_2029_sv2v_reg <= w_data_i[429];
      mem_2028_sv2v_reg <= w_data_i[428];
      mem_2027_sv2v_reg <= w_data_i[427];
      mem_2026_sv2v_reg <= w_data_i[426];
      mem_2025_sv2v_reg <= w_data_i[425];
      mem_2024_sv2v_reg <= w_data_i[424];
      mem_2023_sv2v_reg <= w_data_i[423];
      mem_2022_sv2v_reg <= w_data_i[422];
      mem_2021_sv2v_reg <= w_data_i[421];
      mem_2020_sv2v_reg <= w_data_i[420];
      mem_2019_sv2v_reg <= w_data_i[419];
      mem_2018_sv2v_reg <= w_data_i[418];
      mem_2017_sv2v_reg <= w_data_i[417];
      mem_2016_sv2v_reg <= w_data_i[416];
      mem_2015_sv2v_reg <= w_data_i[415];
      mem_2014_sv2v_reg <= w_data_i[414];
      mem_2013_sv2v_reg <= w_data_i[413];
      mem_2012_sv2v_reg <= w_data_i[412];
      mem_1611_sv2v_reg <= w_data_i[11];
    end 
    if(N35) begin
      mem_2011_sv2v_reg <= w_data_i[411];
      mem_2010_sv2v_reg <= w_data_i[410];
      mem_2009_sv2v_reg <= w_data_i[409];
      mem_2008_sv2v_reg <= w_data_i[408];
      mem_2007_sv2v_reg <= w_data_i[407];
      mem_2006_sv2v_reg <= w_data_i[406];
      mem_2005_sv2v_reg <= w_data_i[405];
      mem_2004_sv2v_reg <= w_data_i[404];
      mem_2003_sv2v_reg <= w_data_i[403];
      mem_2002_sv2v_reg <= w_data_i[402];
      mem_2001_sv2v_reg <= w_data_i[401];
      mem_2000_sv2v_reg <= w_data_i[400];
      mem_1999_sv2v_reg <= w_data_i[399];
      mem_1998_sv2v_reg <= w_data_i[398];
      mem_1997_sv2v_reg <= w_data_i[397];
      mem_1996_sv2v_reg <= w_data_i[396];
      mem_1995_sv2v_reg <= w_data_i[395];
      mem_1994_sv2v_reg <= w_data_i[394];
      mem_1993_sv2v_reg <= w_data_i[393];
      mem_1992_sv2v_reg <= w_data_i[392];
      mem_1991_sv2v_reg <= w_data_i[391];
      mem_1990_sv2v_reg <= w_data_i[390];
      mem_1989_sv2v_reg <= w_data_i[389];
      mem_1988_sv2v_reg <= w_data_i[388];
      mem_1987_sv2v_reg <= w_data_i[387];
      mem_1986_sv2v_reg <= w_data_i[386];
      mem_1985_sv2v_reg <= w_data_i[385];
      mem_1984_sv2v_reg <= w_data_i[384];
      mem_1983_sv2v_reg <= w_data_i[383];
      mem_1982_sv2v_reg <= w_data_i[382];
      mem_1981_sv2v_reg <= w_data_i[381];
      mem_1980_sv2v_reg <= w_data_i[380];
      mem_1979_sv2v_reg <= w_data_i[379];
      mem_1978_sv2v_reg <= w_data_i[378];
      mem_1977_sv2v_reg <= w_data_i[377];
      mem_1976_sv2v_reg <= w_data_i[376];
      mem_1975_sv2v_reg <= w_data_i[375];
      mem_1974_sv2v_reg <= w_data_i[374];
      mem_1973_sv2v_reg <= w_data_i[373];
      mem_1972_sv2v_reg <= w_data_i[372];
      mem_1971_sv2v_reg <= w_data_i[371];
      mem_1970_sv2v_reg <= w_data_i[370];
      mem_1969_sv2v_reg <= w_data_i[369];
      mem_1968_sv2v_reg <= w_data_i[368];
      mem_1967_sv2v_reg <= w_data_i[367];
      mem_1966_sv2v_reg <= w_data_i[366];
      mem_1965_sv2v_reg <= w_data_i[365];
      mem_1964_sv2v_reg <= w_data_i[364];
      mem_1963_sv2v_reg <= w_data_i[363];
      mem_1962_sv2v_reg <= w_data_i[362];
      mem_1961_sv2v_reg <= w_data_i[361];
      mem_1960_sv2v_reg <= w_data_i[360];
      mem_1959_sv2v_reg <= w_data_i[359];
      mem_1958_sv2v_reg <= w_data_i[358];
      mem_1957_sv2v_reg <= w_data_i[357];
      mem_1956_sv2v_reg <= w_data_i[356];
      mem_1955_sv2v_reg <= w_data_i[355];
      mem_1954_sv2v_reg <= w_data_i[354];
      mem_1953_sv2v_reg <= w_data_i[353];
      mem_1952_sv2v_reg <= w_data_i[352];
      mem_1951_sv2v_reg <= w_data_i[351];
      mem_1950_sv2v_reg <= w_data_i[350];
      mem_1949_sv2v_reg <= w_data_i[349];
      mem_1948_sv2v_reg <= w_data_i[348];
      mem_1947_sv2v_reg <= w_data_i[347];
      mem_1946_sv2v_reg <= w_data_i[346];
      mem_1945_sv2v_reg <= w_data_i[345];
      mem_1944_sv2v_reg <= w_data_i[344];
      mem_1943_sv2v_reg <= w_data_i[343];
      mem_1942_sv2v_reg <= w_data_i[342];
      mem_1941_sv2v_reg <= w_data_i[341];
      mem_1940_sv2v_reg <= w_data_i[340];
      mem_1939_sv2v_reg <= w_data_i[339];
      mem_1938_sv2v_reg <= w_data_i[338];
      mem_1937_sv2v_reg <= w_data_i[337];
      mem_1936_sv2v_reg <= w_data_i[336];
      mem_1935_sv2v_reg <= w_data_i[335];
      mem_1934_sv2v_reg <= w_data_i[334];
      mem_1933_sv2v_reg <= w_data_i[333];
      mem_1932_sv2v_reg <= w_data_i[332];
      mem_1931_sv2v_reg <= w_data_i[331];
      mem_1930_sv2v_reg <= w_data_i[330];
      mem_1929_sv2v_reg <= w_data_i[329];
      mem_1928_sv2v_reg <= w_data_i[328];
      mem_1927_sv2v_reg <= w_data_i[327];
      mem_1926_sv2v_reg <= w_data_i[326];
      mem_1925_sv2v_reg <= w_data_i[325];
      mem_1924_sv2v_reg <= w_data_i[324];
      mem_1923_sv2v_reg <= w_data_i[323];
      mem_1922_sv2v_reg <= w_data_i[322];
      mem_1921_sv2v_reg <= w_data_i[321];
      mem_1920_sv2v_reg <= w_data_i[320];
      mem_1919_sv2v_reg <= w_data_i[319];
      mem_1918_sv2v_reg <= w_data_i[318];
      mem_1917_sv2v_reg <= w_data_i[317];
      mem_1916_sv2v_reg <= w_data_i[316];
      mem_1915_sv2v_reg <= w_data_i[315];
      mem_1914_sv2v_reg <= w_data_i[314];
      mem_1913_sv2v_reg <= w_data_i[313];
      mem_1612_sv2v_reg <= w_data_i[12];
    end 
    if(N36) begin
      mem_1912_sv2v_reg <= w_data_i[312];
      mem_1911_sv2v_reg <= w_data_i[311];
      mem_1910_sv2v_reg <= w_data_i[310];
      mem_1909_sv2v_reg <= w_data_i[309];
      mem_1908_sv2v_reg <= w_data_i[308];
      mem_1907_sv2v_reg <= w_data_i[307];
      mem_1906_sv2v_reg <= w_data_i[306];
      mem_1905_sv2v_reg <= w_data_i[305];
      mem_1904_sv2v_reg <= w_data_i[304];
      mem_1903_sv2v_reg <= w_data_i[303];
      mem_1902_sv2v_reg <= w_data_i[302];
      mem_1901_sv2v_reg <= w_data_i[301];
      mem_1900_sv2v_reg <= w_data_i[300];
      mem_1899_sv2v_reg <= w_data_i[299];
      mem_1898_sv2v_reg <= w_data_i[298];
      mem_1897_sv2v_reg <= w_data_i[297];
      mem_1896_sv2v_reg <= w_data_i[296];
      mem_1895_sv2v_reg <= w_data_i[295];
      mem_1894_sv2v_reg <= w_data_i[294];
      mem_1893_sv2v_reg <= w_data_i[293];
      mem_1892_sv2v_reg <= w_data_i[292];
      mem_1891_sv2v_reg <= w_data_i[291];
      mem_1890_sv2v_reg <= w_data_i[290];
      mem_1889_sv2v_reg <= w_data_i[289];
      mem_1888_sv2v_reg <= w_data_i[288];
      mem_1887_sv2v_reg <= w_data_i[287];
      mem_1886_sv2v_reg <= w_data_i[286];
      mem_1885_sv2v_reg <= w_data_i[285];
      mem_1884_sv2v_reg <= w_data_i[284];
      mem_1883_sv2v_reg <= w_data_i[283];
      mem_1882_sv2v_reg <= w_data_i[282];
      mem_1881_sv2v_reg <= w_data_i[281];
      mem_1880_sv2v_reg <= w_data_i[280];
      mem_1879_sv2v_reg <= w_data_i[279];
      mem_1878_sv2v_reg <= w_data_i[278];
      mem_1877_sv2v_reg <= w_data_i[277];
      mem_1876_sv2v_reg <= w_data_i[276];
      mem_1875_sv2v_reg <= w_data_i[275];
      mem_1874_sv2v_reg <= w_data_i[274];
      mem_1873_sv2v_reg <= w_data_i[273];
      mem_1872_sv2v_reg <= w_data_i[272];
      mem_1871_sv2v_reg <= w_data_i[271];
      mem_1870_sv2v_reg <= w_data_i[270];
      mem_1869_sv2v_reg <= w_data_i[269];
      mem_1868_sv2v_reg <= w_data_i[268];
      mem_1867_sv2v_reg <= w_data_i[267];
      mem_1866_sv2v_reg <= w_data_i[266];
      mem_1865_sv2v_reg <= w_data_i[265];
      mem_1864_sv2v_reg <= w_data_i[264];
      mem_1863_sv2v_reg <= w_data_i[263];
      mem_1862_sv2v_reg <= w_data_i[262];
      mem_1861_sv2v_reg <= w_data_i[261];
      mem_1860_sv2v_reg <= w_data_i[260];
      mem_1859_sv2v_reg <= w_data_i[259];
      mem_1858_sv2v_reg <= w_data_i[258];
      mem_1857_sv2v_reg <= w_data_i[257];
      mem_1856_sv2v_reg <= w_data_i[256];
      mem_1855_sv2v_reg <= w_data_i[255];
      mem_1854_sv2v_reg <= w_data_i[254];
      mem_1853_sv2v_reg <= w_data_i[253];
      mem_1852_sv2v_reg <= w_data_i[252];
      mem_1851_sv2v_reg <= w_data_i[251];
      mem_1850_sv2v_reg <= w_data_i[250];
      mem_1849_sv2v_reg <= w_data_i[249];
      mem_1848_sv2v_reg <= w_data_i[248];
      mem_1847_sv2v_reg <= w_data_i[247];
      mem_1846_sv2v_reg <= w_data_i[246];
      mem_1845_sv2v_reg <= w_data_i[245];
      mem_1844_sv2v_reg <= w_data_i[244];
      mem_1843_sv2v_reg <= w_data_i[243];
      mem_1842_sv2v_reg <= w_data_i[242];
      mem_1841_sv2v_reg <= w_data_i[241];
      mem_1840_sv2v_reg <= w_data_i[240];
      mem_1839_sv2v_reg <= w_data_i[239];
      mem_1838_sv2v_reg <= w_data_i[238];
      mem_1837_sv2v_reg <= w_data_i[237];
      mem_1836_sv2v_reg <= w_data_i[236];
      mem_1835_sv2v_reg <= w_data_i[235];
      mem_1834_sv2v_reg <= w_data_i[234];
      mem_1833_sv2v_reg <= w_data_i[233];
      mem_1832_sv2v_reg <= w_data_i[232];
      mem_1831_sv2v_reg <= w_data_i[231];
      mem_1830_sv2v_reg <= w_data_i[230];
      mem_1829_sv2v_reg <= w_data_i[229];
      mem_1828_sv2v_reg <= w_data_i[228];
      mem_1827_sv2v_reg <= w_data_i[227];
      mem_1826_sv2v_reg <= w_data_i[226];
      mem_1825_sv2v_reg <= w_data_i[225];
      mem_1824_sv2v_reg <= w_data_i[224];
      mem_1823_sv2v_reg <= w_data_i[223];
      mem_1822_sv2v_reg <= w_data_i[222];
      mem_1821_sv2v_reg <= w_data_i[221];
      mem_1820_sv2v_reg <= w_data_i[220];
      mem_1819_sv2v_reg <= w_data_i[219];
      mem_1818_sv2v_reg <= w_data_i[218];
      mem_1817_sv2v_reg <= w_data_i[217];
      mem_1816_sv2v_reg <= w_data_i[216];
      mem_1815_sv2v_reg <= w_data_i[215];
      mem_1814_sv2v_reg <= w_data_i[214];
      mem_1613_sv2v_reg <= w_data_i[13];
    end 
    if(N37) begin
      mem_1813_sv2v_reg <= w_data_i[213];
      mem_1812_sv2v_reg <= w_data_i[212];
      mem_1811_sv2v_reg <= w_data_i[211];
      mem_1810_sv2v_reg <= w_data_i[210];
      mem_1809_sv2v_reg <= w_data_i[209];
      mem_1808_sv2v_reg <= w_data_i[208];
      mem_1807_sv2v_reg <= w_data_i[207];
      mem_1806_sv2v_reg <= w_data_i[206];
      mem_1805_sv2v_reg <= w_data_i[205];
      mem_1804_sv2v_reg <= w_data_i[204];
      mem_1803_sv2v_reg <= w_data_i[203];
      mem_1802_sv2v_reg <= w_data_i[202];
      mem_1801_sv2v_reg <= w_data_i[201];
      mem_1800_sv2v_reg <= w_data_i[200];
      mem_1799_sv2v_reg <= w_data_i[199];
      mem_1798_sv2v_reg <= w_data_i[198];
      mem_1797_sv2v_reg <= w_data_i[197];
      mem_1796_sv2v_reg <= w_data_i[196];
      mem_1795_sv2v_reg <= w_data_i[195];
      mem_1794_sv2v_reg <= w_data_i[194];
      mem_1793_sv2v_reg <= w_data_i[193];
      mem_1792_sv2v_reg <= w_data_i[192];
      mem_1791_sv2v_reg <= w_data_i[191];
      mem_1790_sv2v_reg <= w_data_i[190];
      mem_1789_sv2v_reg <= w_data_i[189];
      mem_1788_sv2v_reg <= w_data_i[188];
      mem_1787_sv2v_reg <= w_data_i[187];
      mem_1786_sv2v_reg <= w_data_i[186];
      mem_1785_sv2v_reg <= w_data_i[185];
      mem_1784_sv2v_reg <= w_data_i[184];
      mem_1783_sv2v_reg <= w_data_i[183];
      mem_1782_sv2v_reg <= w_data_i[182];
      mem_1781_sv2v_reg <= w_data_i[181];
      mem_1780_sv2v_reg <= w_data_i[180];
      mem_1779_sv2v_reg <= w_data_i[179];
      mem_1778_sv2v_reg <= w_data_i[178];
      mem_1777_sv2v_reg <= w_data_i[177];
      mem_1776_sv2v_reg <= w_data_i[176];
      mem_1775_sv2v_reg <= w_data_i[175];
      mem_1774_sv2v_reg <= w_data_i[174];
      mem_1773_sv2v_reg <= w_data_i[173];
      mem_1772_sv2v_reg <= w_data_i[172];
      mem_1771_sv2v_reg <= w_data_i[171];
      mem_1770_sv2v_reg <= w_data_i[170];
      mem_1769_sv2v_reg <= w_data_i[169];
      mem_1768_sv2v_reg <= w_data_i[168];
      mem_1767_sv2v_reg <= w_data_i[167];
      mem_1766_sv2v_reg <= w_data_i[166];
      mem_1765_sv2v_reg <= w_data_i[165];
      mem_1764_sv2v_reg <= w_data_i[164];
      mem_1763_sv2v_reg <= w_data_i[163];
      mem_1762_sv2v_reg <= w_data_i[162];
      mem_1761_sv2v_reg <= w_data_i[161];
      mem_1760_sv2v_reg <= w_data_i[160];
      mem_1759_sv2v_reg <= w_data_i[159];
      mem_1758_sv2v_reg <= w_data_i[158];
      mem_1757_sv2v_reg <= w_data_i[157];
      mem_1756_sv2v_reg <= w_data_i[156];
      mem_1755_sv2v_reg <= w_data_i[155];
      mem_1754_sv2v_reg <= w_data_i[154];
      mem_1753_sv2v_reg <= w_data_i[153];
      mem_1752_sv2v_reg <= w_data_i[152];
      mem_1751_sv2v_reg <= w_data_i[151];
      mem_1750_sv2v_reg <= w_data_i[150];
      mem_1749_sv2v_reg <= w_data_i[149];
      mem_1748_sv2v_reg <= w_data_i[148];
      mem_1747_sv2v_reg <= w_data_i[147];
      mem_1746_sv2v_reg <= w_data_i[146];
      mem_1745_sv2v_reg <= w_data_i[145];
      mem_1744_sv2v_reg <= w_data_i[144];
      mem_1743_sv2v_reg <= w_data_i[143];
      mem_1742_sv2v_reg <= w_data_i[142];
      mem_1741_sv2v_reg <= w_data_i[141];
      mem_1740_sv2v_reg <= w_data_i[140];
      mem_1739_sv2v_reg <= w_data_i[139];
      mem_1738_sv2v_reg <= w_data_i[138];
      mem_1737_sv2v_reg <= w_data_i[137];
      mem_1736_sv2v_reg <= w_data_i[136];
      mem_1735_sv2v_reg <= w_data_i[135];
      mem_1734_sv2v_reg <= w_data_i[134];
      mem_1733_sv2v_reg <= w_data_i[133];
      mem_1732_sv2v_reg <= w_data_i[132];
      mem_1731_sv2v_reg <= w_data_i[131];
      mem_1730_sv2v_reg <= w_data_i[130];
      mem_1729_sv2v_reg <= w_data_i[129];
      mem_1728_sv2v_reg <= w_data_i[128];
      mem_1727_sv2v_reg <= w_data_i[127];
      mem_1726_sv2v_reg <= w_data_i[126];
      mem_1725_sv2v_reg <= w_data_i[125];
      mem_1724_sv2v_reg <= w_data_i[124];
      mem_1723_sv2v_reg <= w_data_i[123];
      mem_1722_sv2v_reg <= w_data_i[122];
      mem_1721_sv2v_reg <= w_data_i[121];
      mem_1720_sv2v_reg <= w_data_i[120];
      mem_1719_sv2v_reg <= w_data_i[119];
      mem_1718_sv2v_reg <= w_data_i[118];
      mem_1717_sv2v_reg <= w_data_i[117];
      mem_1716_sv2v_reg <= w_data_i[116];
      mem_1715_sv2v_reg <= w_data_i[115];
      mem_1614_sv2v_reg <= w_data_i[14];
    end 
    if(N38) begin
      mem_1714_sv2v_reg <= w_data_i[114];
      mem_1713_sv2v_reg <= w_data_i[113];
      mem_1712_sv2v_reg <= w_data_i[112];
      mem_1711_sv2v_reg <= w_data_i[111];
      mem_1710_sv2v_reg <= w_data_i[110];
      mem_1709_sv2v_reg <= w_data_i[109];
      mem_1708_sv2v_reg <= w_data_i[108];
      mem_1707_sv2v_reg <= w_data_i[107];
      mem_1706_sv2v_reg <= w_data_i[106];
      mem_1705_sv2v_reg <= w_data_i[105];
      mem_1704_sv2v_reg <= w_data_i[104];
      mem_1703_sv2v_reg <= w_data_i[103];
      mem_1702_sv2v_reg <= w_data_i[102];
      mem_1701_sv2v_reg <= w_data_i[101];
      mem_1700_sv2v_reg <= w_data_i[100];
      mem_1699_sv2v_reg <= w_data_i[99];
      mem_1698_sv2v_reg <= w_data_i[98];
      mem_1697_sv2v_reg <= w_data_i[97];
      mem_1696_sv2v_reg <= w_data_i[96];
      mem_1695_sv2v_reg <= w_data_i[95];
      mem_1694_sv2v_reg <= w_data_i[94];
      mem_1693_sv2v_reg <= w_data_i[93];
      mem_1692_sv2v_reg <= w_data_i[92];
      mem_1691_sv2v_reg <= w_data_i[91];
      mem_1690_sv2v_reg <= w_data_i[90];
      mem_1689_sv2v_reg <= w_data_i[89];
      mem_1688_sv2v_reg <= w_data_i[88];
      mem_1687_sv2v_reg <= w_data_i[87];
      mem_1686_sv2v_reg <= w_data_i[86];
      mem_1685_sv2v_reg <= w_data_i[85];
      mem_1684_sv2v_reg <= w_data_i[84];
      mem_1683_sv2v_reg <= w_data_i[83];
      mem_1682_sv2v_reg <= w_data_i[82];
      mem_1681_sv2v_reg <= w_data_i[81];
      mem_1680_sv2v_reg <= w_data_i[80];
      mem_1679_sv2v_reg <= w_data_i[79];
      mem_1678_sv2v_reg <= w_data_i[78];
      mem_1677_sv2v_reg <= w_data_i[77];
      mem_1676_sv2v_reg <= w_data_i[76];
      mem_1675_sv2v_reg <= w_data_i[75];
      mem_1674_sv2v_reg <= w_data_i[74];
      mem_1673_sv2v_reg <= w_data_i[73];
      mem_1672_sv2v_reg <= w_data_i[72];
      mem_1671_sv2v_reg <= w_data_i[71];
      mem_1670_sv2v_reg <= w_data_i[70];
      mem_1669_sv2v_reg <= w_data_i[69];
      mem_1668_sv2v_reg <= w_data_i[68];
      mem_1667_sv2v_reg <= w_data_i[67];
      mem_1666_sv2v_reg <= w_data_i[66];
      mem_1665_sv2v_reg <= w_data_i[65];
      mem_1664_sv2v_reg <= w_data_i[64];
      mem_1663_sv2v_reg <= w_data_i[63];
      mem_1662_sv2v_reg <= w_data_i[62];
      mem_1661_sv2v_reg <= w_data_i[61];
      mem_1660_sv2v_reg <= w_data_i[60];
      mem_1659_sv2v_reg <= w_data_i[59];
      mem_1658_sv2v_reg <= w_data_i[58];
      mem_1657_sv2v_reg <= w_data_i[57];
      mem_1656_sv2v_reg <= w_data_i[56];
      mem_1655_sv2v_reg <= w_data_i[55];
      mem_1654_sv2v_reg <= w_data_i[54];
      mem_1653_sv2v_reg <= w_data_i[53];
      mem_1652_sv2v_reg <= w_data_i[52];
      mem_1651_sv2v_reg <= w_data_i[51];
      mem_1650_sv2v_reg <= w_data_i[50];
      mem_1649_sv2v_reg <= w_data_i[49];
      mem_1648_sv2v_reg <= w_data_i[48];
      mem_1647_sv2v_reg <= w_data_i[47];
      mem_1646_sv2v_reg <= w_data_i[46];
      mem_1645_sv2v_reg <= w_data_i[45];
      mem_1644_sv2v_reg <= w_data_i[44];
      mem_1643_sv2v_reg <= w_data_i[43];
      mem_1642_sv2v_reg <= w_data_i[42];
      mem_1641_sv2v_reg <= w_data_i[41];
      mem_1640_sv2v_reg <= w_data_i[40];
      mem_1639_sv2v_reg <= w_data_i[39];
      mem_1638_sv2v_reg <= w_data_i[38];
      mem_1637_sv2v_reg <= w_data_i[37];
      mem_1636_sv2v_reg <= w_data_i[36];
      mem_1635_sv2v_reg <= w_data_i[35];
      mem_1634_sv2v_reg <= w_data_i[34];
      mem_1633_sv2v_reg <= w_data_i[33];
      mem_1632_sv2v_reg <= w_data_i[32];
      mem_1631_sv2v_reg <= w_data_i[31];
      mem_1630_sv2v_reg <= w_data_i[30];
      mem_1629_sv2v_reg <= w_data_i[29];
      mem_1628_sv2v_reg <= w_data_i[28];
      mem_1627_sv2v_reg <= w_data_i[27];
      mem_1626_sv2v_reg <= w_data_i[26];
      mem_1625_sv2v_reg <= w_data_i[25];
      mem_1624_sv2v_reg <= w_data_i[24];
      mem_1623_sv2v_reg <= w_data_i[23];
      mem_1622_sv2v_reg <= w_data_i[22];
      mem_1621_sv2v_reg <= w_data_i[21];
      mem_1620_sv2v_reg <= w_data_i[20];
      mem_1619_sv2v_reg <= w_data_i[19];
      mem_1618_sv2v_reg <= w_data_i[18];
      mem_1617_sv2v_reg <= w_data_i[17];
      mem_1616_sv2v_reg <= w_data_i[16];
      mem_1615_sv2v_reg <= w_data_i[15];
    end 
    if(N7) begin
      mem_1599_sv2v_reg <= w_data_i[1599];
      mem_1598_sv2v_reg <= w_data_i[1598];
      mem_1597_sv2v_reg <= w_data_i[1597];
      mem_1596_sv2v_reg <= w_data_i[1596];
      mem_1595_sv2v_reg <= w_data_i[1595];
      mem_1594_sv2v_reg <= w_data_i[1594];
      mem_1593_sv2v_reg <= w_data_i[1593];
      mem_1592_sv2v_reg <= w_data_i[1592];
      mem_1591_sv2v_reg <= w_data_i[1591];
      mem_1590_sv2v_reg <= w_data_i[1590];
      mem_1589_sv2v_reg <= w_data_i[1589];
      mem_1588_sv2v_reg <= w_data_i[1588];
      mem_1587_sv2v_reg <= w_data_i[1587];
      mem_1586_sv2v_reg <= w_data_i[1586];
      mem_1585_sv2v_reg <= w_data_i[1585];
      mem_1584_sv2v_reg <= w_data_i[1584];
      mem_1583_sv2v_reg <= w_data_i[1583];
      mem_1582_sv2v_reg <= w_data_i[1582];
      mem_1581_sv2v_reg <= w_data_i[1581];
      mem_1580_sv2v_reg <= w_data_i[1580];
      mem_1579_sv2v_reg <= w_data_i[1579];
      mem_1578_sv2v_reg <= w_data_i[1578];
      mem_1577_sv2v_reg <= w_data_i[1577];
      mem_1576_sv2v_reg <= w_data_i[1576];
      mem_1575_sv2v_reg <= w_data_i[1575];
      mem_1574_sv2v_reg <= w_data_i[1574];
      mem_1573_sv2v_reg <= w_data_i[1573];
      mem_1572_sv2v_reg <= w_data_i[1572];
      mem_1571_sv2v_reg <= w_data_i[1571];
      mem_1570_sv2v_reg <= w_data_i[1570];
      mem_1569_sv2v_reg <= w_data_i[1569];
      mem_1568_sv2v_reg <= w_data_i[1568];
      mem_1567_sv2v_reg <= w_data_i[1567];
      mem_1566_sv2v_reg <= w_data_i[1566];
      mem_1565_sv2v_reg <= w_data_i[1565];
      mem_1564_sv2v_reg <= w_data_i[1564];
      mem_1563_sv2v_reg <= w_data_i[1563];
      mem_1562_sv2v_reg <= w_data_i[1562];
      mem_1561_sv2v_reg <= w_data_i[1561];
      mem_1560_sv2v_reg <= w_data_i[1560];
      mem_1559_sv2v_reg <= w_data_i[1559];
      mem_1558_sv2v_reg <= w_data_i[1558];
      mem_1557_sv2v_reg <= w_data_i[1557];
      mem_1556_sv2v_reg <= w_data_i[1556];
      mem_1555_sv2v_reg <= w_data_i[1555];
      mem_1554_sv2v_reg <= w_data_i[1554];
      mem_1553_sv2v_reg <= w_data_i[1553];
      mem_1552_sv2v_reg <= w_data_i[1552];
      mem_1551_sv2v_reg <= w_data_i[1551];
      mem_1550_sv2v_reg <= w_data_i[1550];
      mem_1549_sv2v_reg <= w_data_i[1549];
      mem_1548_sv2v_reg <= w_data_i[1548];
      mem_1547_sv2v_reg <= w_data_i[1547];
      mem_1546_sv2v_reg <= w_data_i[1546];
      mem_1545_sv2v_reg <= w_data_i[1545];
      mem_1544_sv2v_reg <= w_data_i[1544];
      mem_1543_sv2v_reg <= w_data_i[1543];
      mem_1542_sv2v_reg <= w_data_i[1542];
      mem_1541_sv2v_reg <= w_data_i[1541];
      mem_1540_sv2v_reg <= w_data_i[1540];
      mem_1539_sv2v_reg <= w_data_i[1539];
      mem_1538_sv2v_reg <= w_data_i[1538];
      mem_1537_sv2v_reg <= w_data_i[1537];
      mem_1536_sv2v_reg <= w_data_i[1536];
      mem_1535_sv2v_reg <= w_data_i[1535];
      mem_1534_sv2v_reg <= w_data_i[1534];
      mem_1533_sv2v_reg <= w_data_i[1533];
      mem_1532_sv2v_reg <= w_data_i[1532];
      mem_1531_sv2v_reg <= w_data_i[1531];
      mem_1530_sv2v_reg <= w_data_i[1530];
      mem_1529_sv2v_reg <= w_data_i[1529];
      mem_1528_sv2v_reg <= w_data_i[1528];
      mem_1527_sv2v_reg <= w_data_i[1527];
      mem_1526_sv2v_reg <= w_data_i[1526];
      mem_1525_sv2v_reg <= w_data_i[1525];
      mem_1524_sv2v_reg <= w_data_i[1524];
      mem_1523_sv2v_reg <= w_data_i[1523];
      mem_1522_sv2v_reg <= w_data_i[1522];
      mem_1521_sv2v_reg <= w_data_i[1521];
      mem_1520_sv2v_reg <= w_data_i[1520];
      mem_1519_sv2v_reg <= w_data_i[1519];
      mem_1518_sv2v_reg <= w_data_i[1518];
      mem_1517_sv2v_reg <= w_data_i[1517];
      mem_1516_sv2v_reg <= w_data_i[1516];
      mem_1515_sv2v_reg <= w_data_i[1515];
      mem_1514_sv2v_reg <= w_data_i[1514];
      mem_1513_sv2v_reg <= w_data_i[1513];
      mem_1512_sv2v_reg <= w_data_i[1512];
      mem_1511_sv2v_reg <= w_data_i[1511];
      mem_1510_sv2v_reg <= w_data_i[1510];
      mem_1509_sv2v_reg <= w_data_i[1509];
      mem_1508_sv2v_reg <= w_data_i[1508];
      mem_1507_sv2v_reg <= w_data_i[1507];
      mem_1506_sv2v_reg <= w_data_i[1506];
      mem_1505_sv2v_reg <= w_data_i[1505];
      mem_1504_sv2v_reg <= w_data_i[1504];
      mem_1503_sv2v_reg <= w_data_i[1503];
      mem_1502_sv2v_reg <= w_data_i[1502];
      mem_1501_sv2v_reg <= w_data_i[1501];
      mem_0_sv2v_reg <= w_data_i[0];
    end 
    if(N8) begin
      mem_1500_sv2v_reg <= w_data_i[1500];
      mem_1499_sv2v_reg <= w_data_i[1499];
      mem_1498_sv2v_reg <= w_data_i[1498];
      mem_1497_sv2v_reg <= w_data_i[1497];
      mem_1496_sv2v_reg <= w_data_i[1496];
      mem_1495_sv2v_reg <= w_data_i[1495];
      mem_1494_sv2v_reg <= w_data_i[1494];
      mem_1493_sv2v_reg <= w_data_i[1493];
      mem_1492_sv2v_reg <= w_data_i[1492];
      mem_1491_sv2v_reg <= w_data_i[1491];
      mem_1490_sv2v_reg <= w_data_i[1490];
      mem_1489_sv2v_reg <= w_data_i[1489];
      mem_1488_sv2v_reg <= w_data_i[1488];
      mem_1487_sv2v_reg <= w_data_i[1487];
      mem_1486_sv2v_reg <= w_data_i[1486];
      mem_1485_sv2v_reg <= w_data_i[1485];
      mem_1484_sv2v_reg <= w_data_i[1484];
      mem_1483_sv2v_reg <= w_data_i[1483];
      mem_1482_sv2v_reg <= w_data_i[1482];
      mem_1481_sv2v_reg <= w_data_i[1481];
      mem_1480_sv2v_reg <= w_data_i[1480];
      mem_1479_sv2v_reg <= w_data_i[1479];
      mem_1478_sv2v_reg <= w_data_i[1478];
      mem_1477_sv2v_reg <= w_data_i[1477];
      mem_1476_sv2v_reg <= w_data_i[1476];
      mem_1475_sv2v_reg <= w_data_i[1475];
      mem_1474_sv2v_reg <= w_data_i[1474];
      mem_1473_sv2v_reg <= w_data_i[1473];
      mem_1472_sv2v_reg <= w_data_i[1472];
      mem_1471_sv2v_reg <= w_data_i[1471];
      mem_1470_sv2v_reg <= w_data_i[1470];
      mem_1469_sv2v_reg <= w_data_i[1469];
      mem_1468_sv2v_reg <= w_data_i[1468];
      mem_1467_sv2v_reg <= w_data_i[1467];
      mem_1466_sv2v_reg <= w_data_i[1466];
      mem_1465_sv2v_reg <= w_data_i[1465];
      mem_1464_sv2v_reg <= w_data_i[1464];
      mem_1463_sv2v_reg <= w_data_i[1463];
      mem_1462_sv2v_reg <= w_data_i[1462];
      mem_1461_sv2v_reg <= w_data_i[1461];
      mem_1460_sv2v_reg <= w_data_i[1460];
      mem_1459_sv2v_reg <= w_data_i[1459];
      mem_1458_sv2v_reg <= w_data_i[1458];
      mem_1457_sv2v_reg <= w_data_i[1457];
      mem_1456_sv2v_reg <= w_data_i[1456];
      mem_1455_sv2v_reg <= w_data_i[1455];
      mem_1454_sv2v_reg <= w_data_i[1454];
      mem_1453_sv2v_reg <= w_data_i[1453];
      mem_1452_sv2v_reg <= w_data_i[1452];
      mem_1451_sv2v_reg <= w_data_i[1451];
      mem_1450_sv2v_reg <= w_data_i[1450];
      mem_1449_sv2v_reg <= w_data_i[1449];
      mem_1448_sv2v_reg <= w_data_i[1448];
      mem_1447_sv2v_reg <= w_data_i[1447];
      mem_1446_sv2v_reg <= w_data_i[1446];
      mem_1445_sv2v_reg <= w_data_i[1445];
      mem_1444_sv2v_reg <= w_data_i[1444];
      mem_1443_sv2v_reg <= w_data_i[1443];
      mem_1442_sv2v_reg <= w_data_i[1442];
      mem_1441_sv2v_reg <= w_data_i[1441];
      mem_1440_sv2v_reg <= w_data_i[1440];
      mem_1439_sv2v_reg <= w_data_i[1439];
      mem_1438_sv2v_reg <= w_data_i[1438];
      mem_1437_sv2v_reg <= w_data_i[1437];
      mem_1436_sv2v_reg <= w_data_i[1436];
      mem_1435_sv2v_reg <= w_data_i[1435];
      mem_1434_sv2v_reg <= w_data_i[1434];
      mem_1433_sv2v_reg <= w_data_i[1433];
      mem_1432_sv2v_reg <= w_data_i[1432];
      mem_1431_sv2v_reg <= w_data_i[1431];
      mem_1430_sv2v_reg <= w_data_i[1430];
      mem_1429_sv2v_reg <= w_data_i[1429];
      mem_1428_sv2v_reg <= w_data_i[1428];
      mem_1427_sv2v_reg <= w_data_i[1427];
      mem_1426_sv2v_reg <= w_data_i[1426];
      mem_1425_sv2v_reg <= w_data_i[1425];
      mem_1424_sv2v_reg <= w_data_i[1424];
      mem_1423_sv2v_reg <= w_data_i[1423];
      mem_1422_sv2v_reg <= w_data_i[1422];
      mem_1421_sv2v_reg <= w_data_i[1421];
      mem_1420_sv2v_reg <= w_data_i[1420];
      mem_1419_sv2v_reg <= w_data_i[1419];
      mem_1418_sv2v_reg <= w_data_i[1418];
      mem_1417_sv2v_reg <= w_data_i[1417];
      mem_1416_sv2v_reg <= w_data_i[1416];
      mem_1415_sv2v_reg <= w_data_i[1415];
      mem_1414_sv2v_reg <= w_data_i[1414];
      mem_1413_sv2v_reg <= w_data_i[1413];
      mem_1412_sv2v_reg <= w_data_i[1412];
      mem_1411_sv2v_reg <= w_data_i[1411];
      mem_1410_sv2v_reg <= w_data_i[1410];
      mem_1409_sv2v_reg <= w_data_i[1409];
      mem_1408_sv2v_reg <= w_data_i[1408];
      mem_1407_sv2v_reg <= w_data_i[1407];
      mem_1406_sv2v_reg <= w_data_i[1406];
      mem_1405_sv2v_reg <= w_data_i[1405];
      mem_1404_sv2v_reg <= w_data_i[1404];
      mem_1403_sv2v_reg <= w_data_i[1403];
      mem_1402_sv2v_reg <= w_data_i[1402];
      mem_1_sv2v_reg <= w_data_i[1];
    end 
    if(N9) begin
      mem_1401_sv2v_reg <= w_data_i[1401];
      mem_1400_sv2v_reg <= w_data_i[1400];
      mem_1399_sv2v_reg <= w_data_i[1399];
      mem_1398_sv2v_reg <= w_data_i[1398];
      mem_1397_sv2v_reg <= w_data_i[1397];
      mem_1396_sv2v_reg <= w_data_i[1396];
      mem_1395_sv2v_reg <= w_data_i[1395];
      mem_1394_sv2v_reg <= w_data_i[1394];
      mem_1393_sv2v_reg <= w_data_i[1393];
      mem_1392_sv2v_reg <= w_data_i[1392];
      mem_1391_sv2v_reg <= w_data_i[1391];
      mem_1390_sv2v_reg <= w_data_i[1390];
      mem_1389_sv2v_reg <= w_data_i[1389];
      mem_1388_sv2v_reg <= w_data_i[1388];
      mem_1387_sv2v_reg <= w_data_i[1387];
      mem_1386_sv2v_reg <= w_data_i[1386];
      mem_1385_sv2v_reg <= w_data_i[1385];
      mem_1384_sv2v_reg <= w_data_i[1384];
      mem_1383_sv2v_reg <= w_data_i[1383];
      mem_1382_sv2v_reg <= w_data_i[1382];
      mem_1381_sv2v_reg <= w_data_i[1381];
      mem_1380_sv2v_reg <= w_data_i[1380];
      mem_1379_sv2v_reg <= w_data_i[1379];
      mem_1378_sv2v_reg <= w_data_i[1378];
      mem_1377_sv2v_reg <= w_data_i[1377];
      mem_1376_sv2v_reg <= w_data_i[1376];
      mem_1375_sv2v_reg <= w_data_i[1375];
      mem_1374_sv2v_reg <= w_data_i[1374];
      mem_1373_sv2v_reg <= w_data_i[1373];
      mem_1372_sv2v_reg <= w_data_i[1372];
      mem_1371_sv2v_reg <= w_data_i[1371];
      mem_1370_sv2v_reg <= w_data_i[1370];
      mem_1369_sv2v_reg <= w_data_i[1369];
      mem_1368_sv2v_reg <= w_data_i[1368];
      mem_1367_sv2v_reg <= w_data_i[1367];
      mem_1366_sv2v_reg <= w_data_i[1366];
      mem_1365_sv2v_reg <= w_data_i[1365];
      mem_1364_sv2v_reg <= w_data_i[1364];
      mem_1363_sv2v_reg <= w_data_i[1363];
      mem_1362_sv2v_reg <= w_data_i[1362];
      mem_1361_sv2v_reg <= w_data_i[1361];
      mem_1360_sv2v_reg <= w_data_i[1360];
      mem_1359_sv2v_reg <= w_data_i[1359];
      mem_1358_sv2v_reg <= w_data_i[1358];
      mem_1357_sv2v_reg <= w_data_i[1357];
      mem_1356_sv2v_reg <= w_data_i[1356];
      mem_1355_sv2v_reg <= w_data_i[1355];
      mem_1354_sv2v_reg <= w_data_i[1354];
      mem_1353_sv2v_reg <= w_data_i[1353];
      mem_1352_sv2v_reg <= w_data_i[1352];
      mem_1351_sv2v_reg <= w_data_i[1351];
      mem_1350_sv2v_reg <= w_data_i[1350];
      mem_1349_sv2v_reg <= w_data_i[1349];
      mem_1348_sv2v_reg <= w_data_i[1348];
      mem_1347_sv2v_reg <= w_data_i[1347];
      mem_1346_sv2v_reg <= w_data_i[1346];
      mem_1345_sv2v_reg <= w_data_i[1345];
      mem_1344_sv2v_reg <= w_data_i[1344];
      mem_1343_sv2v_reg <= w_data_i[1343];
      mem_1342_sv2v_reg <= w_data_i[1342];
      mem_1341_sv2v_reg <= w_data_i[1341];
      mem_1340_sv2v_reg <= w_data_i[1340];
      mem_1339_sv2v_reg <= w_data_i[1339];
      mem_1338_sv2v_reg <= w_data_i[1338];
      mem_1337_sv2v_reg <= w_data_i[1337];
      mem_1336_sv2v_reg <= w_data_i[1336];
      mem_1335_sv2v_reg <= w_data_i[1335];
      mem_1334_sv2v_reg <= w_data_i[1334];
      mem_1333_sv2v_reg <= w_data_i[1333];
      mem_1332_sv2v_reg <= w_data_i[1332];
      mem_1331_sv2v_reg <= w_data_i[1331];
      mem_1330_sv2v_reg <= w_data_i[1330];
      mem_1329_sv2v_reg <= w_data_i[1329];
      mem_1328_sv2v_reg <= w_data_i[1328];
      mem_1327_sv2v_reg <= w_data_i[1327];
      mem_1326_sv2v_reg <= w_data_i[1326];
      mem_1325_sv2v_reg <= w_data_i[1325];
      mem_1324_sv2v_reg <= w_data_i[1324];
      mem_1323_sv2v_reg <= w_data_i[1323];
      mem_1322_sv2v_reg <= w_data_i[1322];
      mem_1321_sv2v_reg <= w_data_i[1321];
      mem_1320_sv2v_reg <= w_data_i[1320];
      mem_1319_sv2v_reg <= w_data_i[1319];
      mem_1318_sv2v_reg <= w_data_i[1318];
      mem_1317_sv2v_reg <= w_data_i[1317];
      mem_1316_sv2v_reg <= w_data_i[1316];
      mem_1315_sv2v_reg <= w_data_i[1315];
      mem_1314_sv2v_reg <= w_data_i[1314];
      mem_1313_sv2v_reg <= w_data_i[1313];
      mem_1312_sv2v_reg <= w_data_i[1312];
      mem_1311_sv2v_reg <= w_data_i[1311];
      mem_1310_sv2v_reg <= w_data_i[1310];
      mem_1309_sv2v_reg <= w_data_i[1309];
      mem_1308_sv2v_reg <= w_data_i[1308];
      mem_1307_sv2v_reg <= w_data_i[1307];
      mem_1306_sv2v_reg <= w_data_i[1306];
      mem_1305_sv2v_reg <= w_data_i[1305];
      mem_1304_sv2v_reg <= w_data_i[1304];
      mem_1303_sv2v_reg <= w_data_i[1303];
      mem_2_sv2v_reg <= w_data_i[2];
    end 
    if(N10) begin
      mem_1302_sv2v_reg <= w_data_i[1302];
      mem_1301_sv2v_reg <= w_data_i[1301];
      mem_1300_sv2v_reg <= w_data_i[1300];
      mem_1299_sv2v_reg <= w_data_i[1299];
      mem_1298_sv2v_reg <= w_data_i[1298];
      mem_1297_sv2v_reg <= w_data_i[1297];
      mem_1296_sv2v_reg <= w_data_i[1296];
      mem_1295_sv2v_reg <= w_data_i[1295];
      mem_1294_sv2v_reg <= w_data_i[1294];
      mem_1293_sv2v_reg <= w_data_i[1293];
      mem_1292_sv2v_reg <= w_data_i[1292];
      mem_1291_sv2v_reg <= w_data_i[1291];
      mem_1290_sv2v_reg <= w_data_i[1290];
      mem_1289_sv2v_reg <= w_data_i[1289];
      mem_1288_sv2v_reg <= w_data_i[1288];
      mem_1287_sv2v_reg <= w_data_i[1287];
      mem_1286_sv2v_reg <= w_data_i[1286];
      mem_1285_sv2v_reg <= w_data_i[1285];
      mem_1284_sv2v_reg <= w_data_i[1284];
      mem_1283_sv2v_reg <= w_data_i[1283];
      mem_1282_sv2v_reg <= w_data_i[1282];
      mem_1281_sv2v_reg <= w_data_i[1281];
      mem_1280_sv2v_reg <= w_data_i[1280];
      mem_1279_sv2v_reg <= w_data_i[1279];
      mem_1278_sv2v_reg <= w_data_i[1278];
      mem_1277_sv2v_reg <= w_data_i[1277];
      mem_1276_sv2v_reg <= w_data_i[1276];
      mem_1275_sv2v_reg <= w_data_i[1275];
      mem_1274_sv2v_reg <= w_data_i[1274];
      mem_1273_sv2v_reg <= w_data_i[1273];
      mem_1272_sv2v_reg <= w_data_i[1272];
      mem_1271_sv2v_reg <= w_data_i[1271];
      mem_1270_sv2v_reg <= w_data_i[1270];
      mem_1269_sv2v_reg <= w_data_i[1269];
      mem_1268_sv2v_reg <= w_data_i[1268];
      mem_1267_sv2v_reg <= w_data_i[1267];
      mem_1266_sv2v_reg <= w_data_i[1266];
      mem_1265_sv2v_reg <= w_data_i[1265];
      mem_1264_sv2v_reg <= w_data_i[1264];
      mem_1263_sv2v_reg <= w_data_i[1263];
      mem_1262_sv2v_reg <= w_data_i[1262];
      mem_1261_sv2v_reg <= w_data_i[1261];
      mem_1260_sv2v_reg <= w_data_i[1260];
      mem_1259_sv2v_reg <= w_data_i[1259];
      mem_1258_sv2v_reg <= w_data_i[1258];
      mem_1257_sv2v_reg <= w_data_i[1257];
      mem_1256_sv2v_reg <= w_data_i[1256];
      mem_1255_sv2v_reg <= w_data_i[1255];
      mem_1254_sv2v_reg <= w_data_i[1254];
      mem_1253_sv2v_reg <= w_data_i[1253];
      mem_1252_sv2v_reg <= w_data_i[1252];
      mem_1251_sv2v_reg <= w_data_i[1251];
      mem_1250_sv2v_reg <= w_data_i[1250];
      mem_1249_sv2v_reg <= w_data_i[1249];
      mem_1248_sv2v_reg <= w_data_i[1248];
      mem_1247_sv2v_reg <= w_data_i[1247];
      mem_1246_sv2v_reg <= w_data_i[1246];
      mem_1245_sv2v_reg <= w_data_i[1245];
      mem_1244_sv2v_reg <= w_data_i[1244];
      mem_1243_sv2v_reg <= w_data_i[1243];
      mem_1242_sv2v_reg <= w_data_i[1242];
      mem_1241_sv2v_reg <= w_data_i[1241];
      mem_1240_sv2v_reg <= w_data_i[1240];
      mem_1239_sv2v_reg <= w_data_i[1239];
      mem_1238_sv2v_reg <= w_data_i[1238];
      mem_1237_sv2v_reg <= w_data_i[1237];
      mem_1236_sv2v_reg <= w_data_i[1236];
      mem_1235_sv2v_reg <= w_data_i[1235];
      mem_1234_sv2v_reg <= w_data_i[1234];
      mem_1233_sv2v_reg <= w_data_i[1233];
      mem_1232_sv2v_reg <= w_data_i[1232];
      mem_1231_sv2v_reg <= w_data_i[1231];
      mem_1230_sv2v_reg <= w_data_i[1230];
      mem_1229_sv2v_reg <= w_data_i[1229];
      mem_1228_sv2v_reg <= w_data_i[1228];
      mem_1227_sv2v_reg <= w_data_i[1227];
      mem_1226_sv2v_reg <= w_data_i[1226];
      mem_1225_sv2v_reg <= w_data_i[1225];
      mem_1224_sv2v_reg <= w_data_i[1224];
      mem_1223_sv2v_reg <= w_data_i[1223];
      mem_1222_sv2v_reg <= w_data_i[1222];
      mem_1221_sv2v_reg <= w_data_i[1221];
      mem_1220_sv2v_reg <= w_data_i[1220];
      mem_1219_sv2v_reg <= w_data_i[1219];
      mem_1218_sv2v_reg <= w_data_i[1218];
      mem_1217_sv2v_reg <= w_data_i[1217];
      mem_1216_sv2v_reg <= w_data_i[1216];
      mem_1215_sv2v_reg <= w_data_i[1215];
      mem_1214_sv2v_reg <= w_data_i[1214];
      mem_1213_sv2v_reg <= w_data_i[1213];
      mem_1212_sv2v_reg <= w_data_i[1212];
      mem_1211_sv2v_reg <= w_data_i[1211];
      mem_1210_sv2v_reg <= w_data_i[1210];
      mem_1209_sv2v_reg <= w_data_i[1209];
      mem_1208_sv2v_reg <= w_data_i[1208];
      mem_1207_sv2v_reg <= w_data_i[1207];
      mem_1206_sv2v_reg <= w_data_i[1206];
      mem_1205_sv2v_reg <= w_data_i[1205];
      mem_1204_sv2v_reg <= w_data_i[1204];
      mem_3_sv2v_reg <= w_data_i[3];
    end 
    if(N11) begin
      mem_1203_sv2v_reg <= w_data_i[1203];
      mem_1202_sv2v_reg <= w_data_i[1202];
      mem_1201_sv2v_reg <= w_data_i[1201];
      mem_1200_sv2v_reg <= w_data_i[1200];
      mem_1199_sv2v_reg <= w_data_i[1199];
      mem_1198_sv2v_reg <= w_data_i[1198];
      mem_1197_sv2v_reg <= w_data_i[1197];
      mem_1196_sv2v_reg <= w_data_i[1196];
      mem_1195_sv2v_reg <= w_data_i[1195];
      mem_1194_sv2v_reg <= w_data_i[1194];
      mem_1193_sv2v_reg <= w_data_i[1193];
      mem_1192_sv2v_reg <= w_data_i[1192];
      mem_1191_sv2v_reg <= w_data_i[1191];
      mem_1190_sv2v_reg <= w_data_i[1190];
      mem_1189_sv2v_reg <= w_data_i[1189];
      mem_1188_sv2v_reg <= w_data_i[1188];
      mem_1187_sv2v_reg <= w_data_i[1187];
      mem_1186_sv2v_reg <= w_data_i[1186];
      mem_1185_sv2v_reg <= w_data_i[1185];
      mem_1184_sv2v_reg <= w_data_i[1184];
      mem_1183_sv2v_reg <= w_data_i[1183];
      mem_1182_sv2v_reg <= w_data_i[1182];
      mem_1181_sv2v_reg <= w_data_i[1181];
      mem_1180_sv2v_reg <= w_data_i[1180];
      mem_1179_sv2v_reg <= w_data_i[1179];
      mem_1178_sv2v_reg <= w_data_i[1178];
      mem_1177_sv2v_reg <= w_data_i[1177];
      mem_1176_sv2v_reg <= w_data_i[1176];
      mem_1175_sv2v_reg <= w_data_i[1175];
      mem_1174_sv2v_reg <= w_data_i[1174];
      mem_1173_sv2v_reg <= w_data_i[1173];
      mem_1172_sv2v_reg <= w_data_i[1172];
      mem_1171_sv2v_reg <= w_data_i[1171];
      mem_1170_sv2v_reg <= w_data_i[1170];
      mem_1169_sv2v_reg <= w_data_i[1169];
      mem_1168_sv2v_reg <= w_data_i[1168];
      mem_1167_sv2v_reg <= w_data_i[1167];
      mem_1166_sv2v_reg <= w_data_i[1166];
      mem_1165_sv2v_reg <= w_data_i[1165];
      mem_1164_sv2v_reg <= w_data_i[1164];
      mem_1163_sv2v_reg <= w_data_i[1163];
      mem_1162_sv2v_reg <= w_data_i[1162];
      mem_1161_sv2v_reg <= w_data_i[1161];
      mem_1160_sv2v_reg <= w_data_i[1160];
      mem_1159_sv2v_reg <= w_data_i[1159];
      mem_1158_sv2v_reg <= w_data_i[1158];
      mem_1157_sv2v_reg <= w_data_i[1157];
      mem_1156_sv2v_reg <= w_data_i[1156];
      mem_1155_sv2v_reg <= w_data_i[1155];
      mem_1154_sv2v_reg <= w_data_i[1154];
      mem_1153_sv2v_reg <= w_data_i[1153];
      mem_1152_sv2v_reg <= w_data_i[1152];
      mem_1151_sv2v_reg <= w_data_i[1151];
      mem_1150_sv2v_reg <= w_data_i[1150];
      mem_1149_sv2v_reg <= w_data_i[1149];
      mem_1148_sv2v_reg <= w_data_i[1148];
      mem_1147_sv2v_reg <= w_data_i[1147];
      mem_1146_sv2v_reg <= w_data_i[1146];
      mem_1145_sv2v_reg <= w_data_i[1145];
      mem_1144_sv2v_reg <= w_data_i[1144];
      mem_1143_sv2v_reg <= w_data_i[1143];
      mem_1142_sv2v_reg <= w_data_i[1142];
      mem_1141_sv2v_reg <= w_data_i[1141];
      mem_1140_sv2v_reg <= w_data_i[1140];
      mem_1139_sv2v_reg <= w_data_i[1139];
      mem_1138_sv2v_reg <= w_data_i[1138];
      mem_1137_sv2v_reg <= w_data_i[1137];
      mem_1136_sv2v_reg <= w_data_i[1136];
      mem_1135_sv2v_reg <= w_data_i[1135];
      mem_1134_sv2v_reg <= w_data_i[1134];
      mem_1133_sv2v_reg <= w_data_i[1133];
      mem_1132_sv2v_reg <= w_data_i[1132];
      mem_1131_sv2v_reg <= w_data_i[1131];
      mem_1130_sv2v_reg <= w_data_i[1130];
      mem_1129_sv2v_reg <= w_data_i[1129];
      mem_1128_sv2v_reg <= w_data_i[1128];
      mem_1127_sv2v_reg <= w_data_i[1127];
      mem_1126_sv2v_reg <= w_data_i[1126];
      mem_1125_sv2v_reg <= w_data_i[1125];
      mem_1124_sv2v_reg <= w_data_i[1124];
      mem_1123_sv2v_reg <= w_data_i[1123];
      mem_1122_sv2v_reg <= w_data_i[1122];
      mem_1121_sv2v_reg <= w_data_i[1121];
      mem_1120_sv2v_reg <= w_data_i[1120];
      mem_1119_sv2v_reg <= w_data_i[1119];
      mem_1118_sv2v_reg <= w_data_i[1118];
      mem_1117_sv2v_reg <= w_data_i[1117];
      mem_1116_sv2v_reg <= w_data_i[1116];
      mem_1115_sv2v_reg <= w_data_i[1115];
      mem_1114_sv2v_reg <= w_data_i[1114];
      mem_1113_sv2v_reg <= w_data_i[1113];
      mem_1112_sv2v_reg <= w_data_i[1112];
      mem_1111_sv2v_reg <= w_data_i[1111];
      mem_1110_sv2v_reg <= w_data_i[1110];
      mem_1109_sv2v_reg <= w_data_i[1109];
      mem_1108_sv2v_reg <= w_data_i[1108];
      mem_1107_sv2v_reg <= w_data_i[1107];
      mem_1106_sv2v_reg <= w_data_i[1106];
      mem_1105_sv2v_reg <= w_data_i[1105];
      mem_4_sv2v_reg <= w_data_i[4];
    end 
    if(N12) begin
      mem_1104_sv2v_reg <= w_data_i[1104];
      mem_1103_sv2v_reg <= w_data_i[1103];
      mem_1102_sv2v_reg <= w_data_i[1102];
      mem_1101_sv2v_reg <= w_data_i[1101];
      mem_1100_sv2v_reg <= w_data_i[1100];
      mem_1099_sv2v_reg <= w_data_i[1099];
      mem_1098_sv2v_reg <= w_data_i[1098];
      mem_1097_sv2v_reg <= w_data_i[1097];
      mem_1096_sv2v_reg <= w_data_i[1096];
      mem_1095_sv2v_reg <= w_data_i[1095];
      mem_1094_sv2v_reg <= w_data_i[1094];
      mem_1093_sv2v_reg <= w_data_i[1093];
      mem_1092_sv2v_reg <= w_data_i[1092];
      mem_1091_sv2v_reg <= w_data_i[1091];
      mem_1090_sv2v_reg <= w_data_i[1090];
      mem_1089_sv2v_reg <= w_data_i[1089];
      mem_1088_sv2v_reg <= w_data_i[1088];
      mem_1087_sv2v_reg <= w_data_i[1087];
      mem_1086_sv2v_reg <= w_data_i[1086];
      mem_1085_sv2v_reg <= w_data_i[1085];
      mem_1084_sv2v_reg <= w_data_i[1084];
      mem_1083_sv2v_reg <= w_data_i[1083];
      mem_1082_sv2v_reg <= w_data_i[1082];
      mem_1081_sv2v_reg <= w_data_i[1081];
      mem_1080_sv2v_reg <= w_data_i[1080];
      mem_1079_sv2v_reg <= w_data_i[1079];
      mem_1078_sv2v_reg <= w_data_i[1078];
      mem_1077_sv2v_reg <= w_data_i[1077];
      mem_1076_sv2v_reg <= w_data_i[1076];
      mem_1075_sv2v_reg <= w_data_i[1075];
      mem_1074_sv2v_reg <= w_data_i[1074];
      mem_1073_sv2v_reg <= w_data_i[1073];
      mem_1072_sv2v_reg <= w_data_i[1072];
      mem_1071_sv2v_reg <= w_data_i[1071];
      mem_1070_sv2v_reg <= w_data_i[1070];
      mem_1069_sv2v_reg <= w_data_i[1069];
      mem_1068_sv2v_reg <= w_data_i[1068];
      mem_1067_sv2v_reg <= w_data_i[1067];
      mem_1066_sv2v_reg <= w_data_i[1066];
      mem_1065_sv2v_reg <= w_data_i[1065];
      mem_1064_sv2v_reg <= w_data_i[1064];
      mem_1063_sv2v_reg <= w_data_i[1063];
      mem_1062_sv2v_reg <= w_data_i[1062];
      mem_1061_sv2v_reg <= w_data_i[1061];
      mem_1060_sv2v_reg <= w_data_i[1060];
      mem_1059_sv2v_reg <= w_data_i[1059];
      mem_1058_sv2v_reg <= w_data_i[1058];
      mem_1057_sv2v_reg <= w_data_i[1057];
      mem_1056_sv2v_reg <= w_data_i[1056];
      mem_1055_sv2v_reg <= w_data_i[1055];
      mem_1054_sv2v_reg <= w_data_i[1054];
      mem_1053_sv2v_reg <= w_data_i[1053];
      mem_1052_sv2v_reg <= w_data_i[1052];
      mem_1051_sv2v_reg <= w_data_i[1051];
      mem_1050_sv2v_reg <= w_data_i[1050];
      mem_1049_sv2v_reg <= w_data_i[1049];
      mem_1048_sv2v_reg <= w_data_i[1048];
      mem_1047_sv2v_reg <= w_data_i[1047];
      mem_1046_sv2v_reg <= w_data_i[1046];
      mem_1045_sv2v_reg <= w_data_i[1045];
      mem_1044_sv2v_reg <= w_data_i[1044];
      mem_1043_sv2v_reg <= w_data_i[1043];
      mem_1042_sv2v_reg <= w_data_i[1042];
      mem_1041_sv2v_reg <= w_data_i[1041];
      mem_1040_sv2v_reg <= w_data_i[1040];
      mem_1039_sv2v_reg <= w_data_i[1039];
      mem_1038_sv2v_reg <= w_data_i[1038];
      mem_1037_sv2v_reg <= w_data_i[1037];
      mem_1036_sv2v_reg <= w_data_i[1036];
      mem_1035_sv2v_reg <= w_data_i[1035];
      mem_1034_sv2v_reg <= w_data_i[1034];
      mem_1033_sv2v_reg <= w_data_i[1033];
      mem_1032_sv2v_reg <= w_data_i[1032];
      mem_1031_sv2v_reg <= w_data_i[1031];
      mem_1030_sv2v_reg <= w_data_i[1030];
      mem_1029_sv2v_reg <= w_data_i[1029];
      mem_1028_sv2v_reg <= w_data_i[1028];
      mem_1027_sv2v_reg <= w_data_i[1027];
      mem_1026_sv2v_reg <= w_data_i[1026];
      mem_1025_sv2v_reg <= w_data_i[1025];
      mem_1024_sv2v_reg <= w_data_i[1024];
      mem_1023_sv2v_reg <= w_data_i[1023];
      mem_1022_sv2v_reg <= w_data_i[1022];
      mem_1021_sv2v_reg <= w_data_i[1021];
      mem_1020_sv2v_reg <= w_data_i[1020];
      mem_1019_sv2v_reg <= w_data_i[1019];
      mem_1018_sv2v_reg <= w_data_i[1018];
      mem_1017_sv2v_reg <= w_data_i[1017];
      mem_1016_sv2v_reg <= w_data_i[1016];
      mem_1015_sv2v_reg <= w_data_i[1015];
      mem_1014_sv2v_reg <= w_data_i[1014];
      mem_1013_sv2v_reg <= w_data_i[1013];
      mem_1012_sv2v_reg <= w_data_i[1012];
      mem_1011_sv2v_reg <= w_data_i[1011];
      mem_1010_sv2v_reg <= w_data_i[1010];
      mem_1009_sv2v_reg <= w_data_i[1009];
      mem_1008_sv2v_reg <= w_data_i[1008];
      mem_1007_sv2v_reg <= w_data_i[1007];
      mem_1006_sv2v_reg <= w_data_i[1006];
      mem_5_sv2v_reg <= w_data_i[5];
    end 
    if(N13) begin
      mem_1005_sv2v_reg <= w_data_i[1005];
      mem_1004_sv2v_reg <= w_data_i[1004];
      mem_1003_sv2v_reg <= w_data_i[1003];
      mem_1002_sv2v_reg <= w_data_i[1002];
      mem_1001_sv2v_reg <= w_data_i[1001];
      mem_1000_sv2v_reg <= w_data_i[1000];
      mem_999_sv2v_reg <= w_data_i[999];
      mem_998_sv2v_reg <= w_data_i[998];
      mem_997_sv2v_reg <= w_data_i[997];
      mem_996_sv2v_reg <= w_data_i[996];
      mem_995_sv2v_reg <= w_data_i[995];
      mem_994_sv2v_reg <= w_data_i[994];
      mem_993_sv2v_reg <= w_data_i[993];
      mem_992_sv2v_reg <= w_data_i[992];
      mem_991_sv2v_reg <= w_data_i[991];
      mem_990_sv2v_reg <= w_data_i[990];
      mem_989_sv2v_reg <= w_data_i[989];
      mem_988_sv2v_reg <= w_data_i[988];
      mem_987_sv2v_reg <= w_data_i[987];
      mem_986_sv2v_reg <= w_data_i[986];
      mem_985_sv2v_reg <= w_data_i[985];
      mem_984_sv2v_reg <= w_data_i[984];
      mem_983_sv2v_reg <= w_data_i[983];
      mem_982_sv2v_reg <= w_data_i[982];
      mem_981_sv2v_reg <= w_data_i[981];
      mem_980_sv2v_reg <= w_data_i[980];
      mem_979_sv2v_reg <= w_data_i[979];
      mem_978_sv2v_reg <= w_data_i[978];
      mem_977_sv2v_reg <= w_data_i[977];
      mem_976_sv2v_reg <= w_data_i[976];
      mem_975_sv2v_reg <= w_data_i[975];
      mem_974_sv2v_reg <= w_data_i[974];
      mem_973_sv2v_reg <= w_data_i[973];
      mem_972_sv2v_reg <= w_data_i[972];
      mem_971_sv2v_reg <= w_data_i[971];
      mem_970_sv2v_reg <= w_data_i[970];
      mem_969_sv2v_reg <= w_data_i[969];
      mem_968_sv2v_reg <= w_data_i[968];
      mem_967_sv2v_reg <= w_data_i[967];
      mem_966_sv2v_reg <= w_data_i[966];
      mem_965_sv2v_reg <= w_data_i[965];
      mem_964_sv2v_reg <= w_data_i[964];
      mem_963_sv2v_reg <= w_data_i[963];
      mem_962_sv2v_reg <= w_data_i[962];
      mem_961_sv2v_reg <= w_data_i[961];
      mem_960_sv2v_reg <= w_data_i[960];
      mem_959_sv2v_reg <= w_data_i[959];
      mem_958_sv2v_reg <= w_data_i[958];
      mem_957_sv2v_reg <= w_data_i[957];
      mem_956_sv2v_reg <= w_data_i[956];
      mem_955_sv2v_reg <= w_data_i[955];
      mem_954_sv2v_reg <= w_data_i[954];
      mem_953_sv2v_reg <= w_data_i[953];
      mem_952_sv2v_reg <= w_data_i[952];
      mem_951_sv2v_reg <= w_data_i[951];
      mem_950_sv2v_reg <= w_data_i[950];
      mem_949_sv2v_reg <= w_data_i[949];
      mem_948_sv2v_reg <= w_data_i[948];
      mem_947_sv2v_reg <= w_data_i[947];
      mem_946_sv2v_reg <= w_data_i[946];
      mem_945_sv2v_reg <= w_data_i[945];
      mem_944_sv2v_reg <= w_data_i[944];
      mem_943_sv2v_reg <= w_data_i[943];
      mem_942_sv2v_reg <= w_data_i[942];
      mem_941_sv2v_reg <= w_data_i[941];
      mem_940_sv2v_reg <= w_data_i[940];
      mem_939_sv2v_reg <= w_data_i[939];
      mem_938_sv2v_reg <= w_data_i[938];
      mem_937_sv2v_reg <= w_data_i[937];
      mem_936_sv2v_reg <= w_data_i[936];
      mem_935_sv2v_reg <= w_data_i[935];
      mem_934_sv2v_reg <= w_data_i[934];
      mem_933_sv2v_reg <= w_data_i[933];
      mem_932_sv2v_reg <= w_data_i[932];
      mem_931_sv2v_reg <= w_data_i[931];
      mem_930_sv2v_reg <= w_data_i[930];
      mem_929_sv2v_reg <= w_data_i[929];
      mem_928_sv2v_reg <= w_data_i[928];
      mem_927_sv2v_reg <= w_data_i[927];
      mem_926_sv2v_reg <= w_data_i[926];
      mem_925_sv2v_reg <= w_data_i[925];
      mem_924_sv2v_reg <= w_data_i[924];
      mem_923_sv2v_reg <= w_data_i[923];
      mem_922_sv2v_reg <= w_data_i[922];
      mem_921_sv2v_reg <= w_data_i[921];
      mem_920_sv2v_reg <= w_data_i[920];
      mem_919_sv2v_reg <= w_data_i[919];
      mem_918_sv2v_reg <= w_data_i[918];
      mem_917_sv2v_reg <= w_data_i[917];
      mem_916_sv2v_reg <= w_data_i[916];
      mem_915_sv2v_reg <= w_data_i[915];
      mem_914_sv2v_reg <= w_data_i[914];
      mem_913_sv2v_reg <= w_data_i[913];
      mem_912_sv2v_reg <= w_data_i[912];
      mem_911_sv2v_reg <= w_data_i[911];
      mem_910_sv2v_reg <= w_data_i[910];
      mem_909_sv2v_reg <= w_data_i[909];
      mem_908_sv2v_reg <= w_data_i[908];
      mem_907_sv2v_reg <= w_data_i[907];
      mem_6_sv2v_reg <= w_data_i[6];
    end 
    if(N14) begin
      mem_906_sv2v_reg <= w_data_i[906];
      mem_905_sv2v_reg <= w_data_i[905];
      mem_904_sv2v_reg <= w_data_i[904];
      mem_903_sv2v_reg <= w_data_i[903];
      mem_902_sv2v_reg <= w_data_i[902];
      mem_901_sv2v_reg <= w_data_i[901];
      mem_900_sv2v_reg <= w_data_i[900];
      mem_899_sv2v_reg <= w_data_i[899];
      mem_898_sv2v_reg <= w_data_i[898];
      mem_897_sv2v_reg <= w_data_i[897];
      mem_896_sv2v_reg <= w_data_i[896];
      mem_895_sv2v_reg <= w_data_i[895];
      mem_894_sv2v_reg <= w_data_i[894];
      mem_893_sv2v_reg <= w_data_i[893];
      mem_892_sv2v_reg <= w_data_i[892];
      mem_891_sv2v_reg <= w_data_i[891];
      mem_890_sv2v_reg <= w_data_i[890];
      mem_889_sv2v_reg <= w_data_i[889];
      mem_888_sv2v_reg <= w_data_i[888];
      mem_887_sv2v_reg <= w_data_i[887];
      mem_886_sv2v_reg <= w_data_i[886];
      mem_885_sv2v_reg <= w_data_i[885];
      mem_884_sv2v_reg <= w_data_i[884];
      mem_883_sv2v_reg <= w_data_i[883];
      mem_882_sv2v_reg <= w_data_i[882];
      mem_881_sv2v_reg <= w_data_i[881];
      mem_880_sv2v_reg <= w_data_i[880];
      mem_879_sv2v_reg <= w_data_i[879];
      mem_878_sv2v_reg <= w_data_i[878];
      mem_877_sv2v_reg <= w_data_i[877];
      mem_876_sv2v_reg <= w_data_i[876];
      mem_875_sv2v_reg <= w_data_i[875];
      mem_874_sv2v_reg <= w_data_i[874];
      mem_873_sv2v_reg <= w_data_i[873];
      mem_872_sv2v_reg <= w_data_i[872];
      mem_871_sv2v_reg <= w_data_i[871];
      mem_870_sv2v_reg <= w_data_i[870];
      mem_869_sv2v_reg <= w_data_i[869];
      mem_868_sv2v_reg <= w_data_i[868];
      mem_867_sv2v_reg <= w_data_i[867];
      mem_866_sv2v_reg <= w_data_i[866];
      mem_865_sv2v_reg <= w_data_i[865];
      mem_864_sv2v_reg <= w_data_i[864];
      mem_863_sv2v_reg <= w_data_i[863];
      mem_862_sv2v_reg <= w_data_i[862];
      mem_861_sv2v_reg <= w_data_i[861];
      mem_860_sv2v_reg <= w_data_i[860];
      mem_859_sv2v_reg <= w_data_i[859];
      mem_858_sv2v_reg <= w_data_i[858];
      mem_857_sv2v_reg <= w_data_i[857];
      mem_856_sv2v_reg <= w_data_i[856];
      mem_855_sv2v_reg <= w_data_i[855];
      mem_854_sv2v_reg <= w_data_i[854];
      mem_853_sv2v_reg <= w_data_i[853];
      mem_852_sv2v_reg <= w_data_i[852];
      mem_851_sv2v_reg <= w_data_i[851];
      mem_850_sv2v_reg <= w_data_i[850];
      mem_849_sv2v_reg <= w_data_i[849];
      mem_848_sv2v_reg <= w_data_i[848];
      mem_847_sv2v_reg <= w_data_i[847];
      mem_846_sv2v_reg <= w_data_i[846];
      mem_845_sv2v_reg <= w_data_i[845];
      mem_844_sv2v_reg <= w_data_i[844];
      mem_843_sv2v_reg <= w_data_i[843];
      mem_842_sv2v_reg <= w_data_i[842];
      mem_841_sv2v_reg <= w_data_i[841];
      mem_840_sv2v_reg <= w_data_i[840];
      mem_839_sv2v_reg <= w_data_i[839];
      mem_838_sv2v_reg <= w_data_i[838];
      mem_837_sv2v_reg <= w_data_i[837];
      mem_836_sv2v_reg <= w_data_i[836];
      mem_835_sv2v_reg <= w_data_i[835];
      mem_834_sv2v_reg <= w_data_i[834];
      mem_833_sv2v_reg <= w_data_i[833];
      mem_832_sv2v_reg <= w_data_i[832];
      mem_831_sv2v_reg <= w_data_i[831];
      mem_830_sv2v_reg <= w_data_i[830];
      mem_829_sv2v_reg <= w_data_i[829];
      mem_828_sv2v_reg <= w_data_i[828];
      mem_827_sv2v_reg <= w_data_i[827];
      mem_826_sv2v_reg <= w_data_i[826];
      mem_825_sv2v_reg <= w_data_i[825];
      mem_824_sv2v_reg <= w_data_i[824];
      mem_823_sv2v_reg <= w_data_i[823];
      mem_822_sv2v_reg <= w_data_i[822];
      mem_821_sv2v_reg <= w_data_i[821];
      mem_820_sv2v_reg <= w_data_i[820];
      mem_819_sv2v_reg <= w_data_i[819];
      mem_818_sv2v_reg <= w_data_i[818];
      mem_817_sv2v_reg <= w_data_i[817];
      mem_816_sv2v_reg <= w_data_i[816];
      mem_815_sv2v_reg <= w_data_i[815];
      mem_814_sv2v_reg <= w_data_i[814];
      mem_813_sv2v_reg <= w_data_i[813];
      mem_812_sv2v_reg <= w_data_i[812];
      mem_811_sv2v_reg <= w_data_i[811];
      mem_810_sv2v_reg <= w_data_i[810];
      mem_809_sv2v_reg <= w_data_i[809];
      mem_808_sv2v_reg <= w_data_i[808];
      mem_7_sv2v_reg <= w_data_i[7];
    end 
    if(N15) begin
      mem_807_sv2v_reg <= w_data_i[807];
      mem_806_sv2v_reg <= w_data_i[806];
      mem_805_sv2v_reg <= w_data_i[805];
      mem_804_sv2v_reg <= w_data_i[804];
      mem_803_sv2v_reg <= w_data_i[803];
      mem_802_sv2v_reg <= w_data_i[802];
      mem_801_sv2v_reg <= w_data_i[801];
      mem_800_sv2v_reg <= w_data_i[800];
      mem_799_sv2v_reg <= w_data_i[799];
      mem_798_sv2v_reg <= w_data_i[798];
      mem_797_sv2v_reg <= w_data_i[797];
      mem_796_sv2v_reg <= w_data_i[796];
      mem_795_sv2v_reg <= w_data_i[795];
      mem_794_sv2v_reg <= w_data_i[794];
      mem_793_sv2v_reg <= w_data_i[793];
      mem_792_sv2v_reg <= w_data_i[792];
      mem_791_sv2v_reg <= w_data_i[791];
      mem_790_sv2v_reg <= w_data_i[790];
      mem_789_sv2v_reg <= w_data_i[789];
      mem_788_sv2v_reg <= w_data_i[788];
      mem_787_sv2v_reg <= w_data_i[787];
      mem_786_sv2v_reg <= w_data_i[786];
      mem_785_sv2v_reg <= w_data_i[785];
      mem_784_sv2v_reg <= w_data_i[784];
      mem_783_sv2v_reg <= w_data_i[783];
      mem_782_sv2v_reg <= w_data_i[782];
      mem_781_sv2v_reg <= w_data_i[781];
      mem_780_sv2v_reg <= w_data_i[780];
      mem_779_sv2v_reg <= w_data_i[779];
      mem_778_sv2v_reg <= w_data_i[778];
      mem_777_sv2v_reg <= w_data_i[777];
      mem_776_sv2v_reg <= w_data_i[776];
      mem_775_sv2v_reg <= w_data_i[775];
      mem_774_sv2v_reg <= w_data_i[774];
      mem_773_sv2v_reg <= w_data_i[773];
      mem_772_sv2v_reg <= w_data_i[772];
      mem_771_sv2v_reg <= w_data_i[771];
      mem_770_sv2v_reg <= w_data_i[770];
      mem_769_sv2v_reg <= w_data_i[769];
      mem_768_sv2v_reg <= w_data_i[768];
      mem_767_sv2v_reg <= w_data_i[767];
      mem_766_sv2v_reg <= w_data_i[766];
      mem_765_sv2v_reg <= w_data_i[765];
      mem_764_sv2v_reg <= w_data_i[764];
      mem_763_sv2v_reg <= w_data_i[763];
      mem_762_sv2v_reg <= w_data_i[762];
      mem_761_sv2v_reg <= w_data_i[761];
      mem_760_sv2v_reg <= w_data_i[760];
      mem_759_sv2v_reg <= w_data_i[759];
      mem_758_sv2v_reg <= w_data_i[758];
      mem_757_sv2v_reg <= w_data_i[757];
      mem_756_sv2v_reg <= w_data_i[756];
      mem_755_sv2v_reg <= w_data_i[755];
      mem_754_sv2v_reg <= w_data_i[754];
      mem_753_sv2v_reg <= w_data_i[753];
      mem_752_sv2v_reg <= w_data_i[752];
      mem_751_sv2v_reg <= w_data_i[751];
      mem_750_sv2v_reg <= w_data_i[750];
      mem_749_sv2v_reg <= w_data_i[749];
      mem_748_sv2v_reg <= w_data_i[748];
      mem_747_sv2v_reg <= w_data_i[747];
      mem_746_sv2v_reg <= w_data_i[746];
      mem_745_sv2v_reg <= w_data_i[745];
      mem_744_sv2v_reg <= w_data_i[744];
      mem_743_sv2v_reg <= w_data_i[743];
      mem_742_sv2v_reg <= w_data_i[742];
      mem_741_sv2v_reg <= w_data_i[741];
      mem_740_sv2v_reg <= w_data_i[740];
      mem_739_sv2v_reg <= w_data_i[739];
      mem_738_sv2v_reg <= w_data_i[738];
      mem_737_sv2v_reg <= w_data_i[737];
      mem_736_sv2v_reg <= w_data_i[736];
      mem_735_sv2v_reg <= w_data_i[735];
      mem_734_sv2v_reg <= w_data_i[734];
      mem_733_sv2v_reg <= w_data_i[733];
      mem_732_sv2v_reg <= w_data_i[732];
      mem_731_sv2v_reg <= w_data_i[731];
      mem_730_sv2v_reg <= w_data_i[730];
      mem_729_sv2v_reg <= w_data_i[729];
      mem_728_sv2v_reg <= w_data_i[728];
      mem_727_sv2v_reg <= w_data_i[727];
      mem_726_sv2v_reg <= w_data_i[726];
      mem_725_sv2v_reg <= w_data_i[725];
      mem_724_sv2v_reg <= w_data_i[724];
      mem_723_sv2v_reg <= w_data_i[723];
      mem_722_sv2v_reg <= w_data_i[722];
      mem_721_sv2v_reg <= w_data_i[721];
      mem_720_sv2v_reg <= w_data_i[720];
      mem_719_sv2v_reg <= w_data_i[719];
      mem_718_sv2v_reg <= w_data_i[718];
      mem_717_sv2v_reg <= w_data_i[717];
      mem_716_sv2v_reg <= w_data_i[716];
      mem_715_sv2v_reg <= w_data_i[715];
      mem_714_sv2v_reg <= w_data_i[714];
      mem_713_sv2v_reg <= w_data_i[713];
      mem_712_sv2v_reg <= w_data_i[712];
      mem_711_sv2v_reg <= w_data_i[711];
      mem_710_sv2v_reg <= w_data_i[710];
      mem_709_sv2v_reg <= w_data_i[709];
      mem_8_sv2v_reg <= w_data_i[8];
    end 
    if(N16) begin
      mem_708_sv2v_reg <= w_data_i[708];
      mem_707_sv2v_reg <= w_data_i[707];
      mem_706_sv2v_reg <= w_data_i[706];
      mem_705_sv2v_reg <= w_data_i[705];
      mem_704_sv2v_reg <= w_data_i[704];
      mem_703_sv2v_reg <= w_data_i[703];
      mem_702_sv2v_reg <= w_data_i[702];
      mem_701_sv2v_reg <= w_data_i[701];
      mem_700_sv2v_reg <= w_data_i[700];
      mem_699_sv2v_reg <= w_data_i[699];
      mem_698_sv2v_reg <= w_data_i[698];
      mem_697_sv2v_reg <= w_data_i[697];
      mem_696_sv2v_reg <= w_data_i[696];
      mem_695_sv2v_reg <= w_data_i[695];
      mem_694_sv2v_reg <= w_data_i[694];
      mem_693_sv2v_reg <= w_data_i[693];
      mem_692_sv2v_reg <= w_data_i[692];
      mem_691_sv2v_reg <= w_data_i[691];
      mem_690_sv2v_reg <= w_data_i[690];
      mem_689_sv2v_reg <= w_data_i[689];
      mem_688_sv2v_reg <= w_data_i[688];
      mem_687_sv2v_reg <= w_data_i[687];
      mem_686_sv2v_reg <= w_data_i[686];
      mem_685_sv2v_reg <= w_data_i[685];
      mem_684_sv2v_reg <= w_data_i[684];
      mem_683_sv2v_reg <= w_data_i[683];
      mem_682_sv2v_reg <= w_data_i[682];
      mem_681_sv2v_reg <= w_data_i[681];
      mem_680_sv2v_reg <= w_data_i[680];
      mem_679_sv2v_reg <= w_data_i[679];
      mem_678_sv2v_reg <= w_data_i[678];
      mem_677_sv2v_reg <= w_data_i[677];
      mem_676_sv2v_reg <= w_data_i[676];
      mem_675_sv2v_reg <= w_data_i[675];
      mem_674_sv2v_reg <= w_data_i[674];
      mem_673_sv2v_reg <= w_data_i[673];
      mem_672_sv2v_reg <= w_data_i[672];
      mem_671_sv2v_reg <= w_data_i[671];
      mem_670_sv2v_reg <= w_data_i[670];
      mem_669_sv2v_reg <= w_data_i[669];
      mem_668_sv2v_reg <= w_data_i[668];
      mem_667_sv2v_reg <= w_data_i[667];
      mem_666_sv2v_reg <= w_data_i[666];
      mem_665_sv2v_reg <= w_data_i[665];
      mem_664_sv2v_reg <= w_data_i[664];
      mem_663_sv2v_reg <= w_data_i[663];
      mem_662_sv2v_reg <= w_data_i[662];
      mem_661_sv2v_reg <= w_data_i[661];
      mem_660_sv2v_reg <= w_data_i[660];
      mem_659_sv2v_reg <= w_data_i[659];
      mem_658_sv2v_reg <= w_data_i[658];
      mem_657_sv2v_reg <= w_data_i[657];
      mem_656_sv2v_reg <= w_data_i[656];
      mem_655_sv2v_reg <= w_data_i[655];
      mem_654_sv2v_reg <= w_data_i[654];
      mem_653_sv2v_reg <= w_data_i[653];
      mem_652_sv2v_reg <= w_data_i[652];
      mem_651_sv2v_reg <= w_data_i[651];
      mem_650_sv2v_reg <= w_data_i[650];
      mem_649_sv2v_reg <= w_data_i[649];
      mem_648_sv2v_reg <= w_data_i[648];
      mem_647_sv2v_reg <= w_data_i[647];
      mem_646_sv2v_reg <= w_data_i[646];
      mem_645_sv2v_reg <= w_data_i[645];
      mem_644_sv2v_reg <= w_data_i[644];
      mem_643_sv2v_reg <= w_data_i[643];
      mem_642_sv2v_reg <= w_data_i[642];
      mem_641_sv2v_reg <= w_data_i[641];
      mem_640_sv2v_reg <= w_data_i[640];
      mem_639_sv2v_reg <= w_data_i[639];
      mem_638_sv2v_reg <= w_data_i[638];
      mem_637_sv2v_reg <= w_data_i[637];
      mem_636_sv2v_reg <= w_data_i[636];
      mem_635_sv2v_reg <= w_data_i[635];
      mem_634_sv2v_reg <= w_data_i[634];
      mem_633_sv2v_reg <= w_data_i[633];
      mem_632_sv2v_reg <= w_data_i[632];
      mem_631_sv2v_reg <= w_data_i[631];
      mem_630_sv2v_reg <= w_data_i[630];
      mem_629_sv2v_reg <= w_data_i[629];
      mem_628_sv2v_reg <= w_data_i[628];
      mem_627_sv2v_reg <= w_data_i[627];
      mem_626_sv2v_reg <= w_data_i[626];
      mem_625_sv2v_reg <= w_data_i[625];
      mem_624_sv2v_reg <= w_data_i[624];
      mem_623_sv2v_reg <= w_data_i[623];
      mem_622_sv2v_reg <= w_data_i[622];
      mem_621_sv2v_reg <= w_data_i[621];
      mem_620_sv2v_reg <= w_data_i[620];
      mem_619_sv2v_reg <= w_data_i[619];
      mem_618_sv2v_reg <= w_data_i[618];
      mem_617_sv2v_reg <= w_data_i[617];
      mem_616_sv2v_reg <= w_data_i[616];
      mem_615_sv2v_reg <= w_data_i[615];
      mem_614_sv2v_reg <= w_data_i[614];
      mem_613_sv2v_reg <= w_data_i[613];
      mem_612_sv2v_reg <= w_data_i[612];
      mem_611_sv2v_reg <= w_data_i[611];
      mem_610_sv2v_reg <= w_data_i[610];
      mem_9_sv2v_reg <= w_data_i[9];
    end 
    if(N17) begin
      mem_609_sv2v_reg <= w_data_i[609];
      mem_608_sv2v_reg <= w_data_i[608];
      mem_607_sv2v_reg <= w_data_i[607];
      mem_606_sv2v_reg <= w_data_i[606];
      mem_605_sv2v_reg <= w_data_i[605];
      mem_604_sv2v_reg <= w_data_i[604];
      mem_603_sv2v_reg <= w_data_i[603];
      mem_602_sv2v_reg <= w_data_i[602];
      mem_601_sv2v_reg <= w_data_i[601];
      mem_600_sv2v_reg <= w_data_i[600];
      mem_599_sv2v_reg <= w_data_i[599];
      mem_598_sv2v_reg <= w_data_i[598];
      mem_597_sv2v_reg <= w_data_i[597];
      mem_596_sv2v_reg <= w_data_i[596];
      mem_595_sv2v_reg <= w_data_i[595];
      mem_594_sv2v_reg <= w_data_i[594];
      mem_593_sv2v_reg <= w_data_i[593];
      mem_592_sv2v_reg <= w_data_i[592];
      mem_591_sv2v_reg <= w_data_i[591];
      mem_590_sv2v_reg <= w_data_i[590];
      mem_589_sv2v_reg <= w_data_i[589];
      mem_588_sv2v_reg <= w_data_i[588];
      mem_587_sv2v_reg <= w_data_i[587];
      mem_586_sv2v_reg <= w_data_i[586];
      mem_585_sv2v_reg <= w_data_i[585];
      mem_584_sv2v_reg <= w_data_i[584];
      mem_583_sv2v_reg <= w_data_i[583];
      mem_582_sv2v_reg <= w_data_i[582];
      mem_581_sv2v_reg <= w_data_i[581];
      mem_580_sv2v_reg <= w_data_i[580];
      mem_579_sv2v_reg <= w_data_i[579];
      mem_578_sv2v_reg <= w_data_i[578];
      mem_577_sv2v_reg <= w_data_i[577];
      mem_576_sv2v_reg <= w_data_i[576];
      mem_575_sv2v_reg <= w_data_i[575];
      mem_574_sv2v_reg <= w_data_i[574];
      mem_573_sv2v_reg <= w_data_i[573];
      mem_572_sv2v_reg <= w_data_i[572];
      mem_571_sv2v_reg <= w_data_i[571];
      mem_570_sv2v_reg <= w_data_i[570];
      mem_569_sv2v_reg <= w_data_i[569];
      mem_568_sv2v_reg <= w_data_i[568];
      mem_567_sv2v_reg <= w_data_i[567];
      mem_566_sv2v_reg <= w_data_i[566];
      mem_565_sv2v_reg <= w_data_i[565];
      mem_564_sv2v_reg <= w_data_i[564];
      mem_563_sv2v_reg <= w_data_i[563];
      mem_562_sv2v_reg <= w_data_i[562];
      mem_561_sv2v_reg <= w_data_i[561];
      mem_560_sv2v_reg <= w_data_i[560];
      mem_559_sv2v_reg <= w_data_i[559];
      mem_558_sv2v_reg <= w_data_i[558];
      mem_557_sv2v_reg <= w_data_i[557];
      mem_556_sv2v_reg <= w_data_i[556];
      mem_555_sv2v_reg <= w_data_i[555];
      mem_554_sv2v_reg <= w_data_i[554];
      mem_553_sv2v_reg <= w_data_i[553];
      mem_552_sv2v_reg <= w_data_i[552];
      mem_551_sv2v_reg <= w_data_i[551];
      mem_550_sv2v_reg <= w_data_i[550];
      mem_549_sv2v_reg <= w_data_i[549];
      mem_548_sv2v_reg <= w_data_i[548];
      mem_547_sv2v_reg <= w_data_i[547];
      mem_546_sv2v_reg <= w_data_i[546];
      mem_545_sv2v_reg <= w_data_i[545];
      mem_544_sv2v_reg <= w_data_i[544];
      mem_543_sv2v_reg <= w_data_i[543];
      mem_542_sv2v_reg <= w_data_i[542];
      mem_541_sv2v_reg <= w_data_i[541];
      mem_540_sv2v_reg <= w_data_i[540];
      mem_539_sv2v_reg <= w_data_i[539];
      mem_538_sv2v_reg <= w_data_i[538];
      mem_537_sv2v_reg <= w_data_i[537];
      mem_536_sv2v_reg <= w_data_i[536];
      mem_535_sv2v_reg <= w_data_i[535];
      mem_534_sv2v_reg <= w_data_i[534];
      mem_533_sv2v_reg <= w_data_i[533];
      mem_532_sv2v_reg <= w_data_i[532];
      mem_531_sv2v_reg <= w_data_i[531];
      mem_530_sv2v_reg <= w_data_i[530];
      mem_529_sv2v_reg <= w_data_i[529];
      mem_528_sv2v_reg <= w_data_i[528];
      mem_527_sv2v_reg <= w_data_i[527];
      mem_526_sv2v_reg <= w_data_i[526];
      mem_525_sv2v_reg <= w_data_i[525];
      mem_524_sv2v_reg <= w_data_i[524];
      mem_523_sv2v_reg <= w_data_i[523];
      mem_522_sv2v_reg <= w_data_i[522];
      mem_521_sv2v_reg <= w_data_i[521];
      mem_520_sv2v_reg <= w_data_i[520];
      mem_519_sv2v_reg <= w_data_i[519];
      mem_518_sv2v_reg <= w_data_i[518];
      mem_517_sv2v_reg <= w_data_i[517];
      mem_516_sv2v_reg <= w_data_i[516];
      mem_515_sv2v_reg <= w_data_i[515];
      mem_514_sv2v_reg <= w_data_i[514];
      mem_513_sv2v_reg <= w_data_i[513];
      mem_512_sv2v_reg <= w_data_i[512];
      mem_511_sv2v_reg <= w_data_i[511];
      mem_10_sv2v_reg <= w_data_i[10];
    end 
    if(N18) begin
      mem_510_sv2v_reg <= w_data_i[510];
      mem_509_sv2v_reg <= w_data_i[509];
      mem_508_sv2v_reg <= w_data_i[508];
      mem_507_sv2v_reg <= w_data_i[507];
      mem_506_sv2v_reg <= w_data_i[506];
      mem_505_sv2v_reg <= w_data_i[505];
      mem_504_sv2v_reg <= w_data_i[504];
      mem_503_sv2v_reg <= w_data_i[503];
      mem_502_sv2v_reg <= w_data_i[502];
      mem_501_sv2v_reg <= w_data_i[501];
      mem_500_sv2v_reg <= w_data_i[500];
      mem_499_sv2v_reg <= w_data_i[499];
      mem_498_sv2v_reg <= w_data_i[498];
      mem_497_sv2v_reg <= w_data_i[497];
      mem_496_sv2v_reg <= w_data_i[496];
      mem_495_sv2v_reg <= w_data_i[495];
      mem_494_sv2v_reg <= w_data_i[494];
      mem_493_sv2v_reg <= w_data_i[493];
      mem_492_sv2v_reg <= w_data_i[492];
      mem_491_sv2v_reg <= w_data_i[491];
      mem_490_sv2v_reg <= w_data_i[490];
      mem_489_sv2v_reg <= w_data_i[489];
      mem_488_sv2v_reg <= w_data_i[488];
      mem_487_sv2v_reg <= w_data_i[487];
      mem_486_sv2v_reg <= w_data_i[486];
      mem_485_sv2v_reg <= w_data_i[485];
      mem_484_sv2v_reg <= w_data_i[484];
      mem_483_sv2v_reg <= w_data_i[483];
      mem_482_sv2v_reg <= w_data_i[482];
      mem_481_sv2v_reg <= w_data_i[481];
      mem_480_sv2v_reg <= w_data_i[480];
      mem_479_sv2v_reg <= w_data_i[479];
      mem_478_sv2v_reg <= w_data_i[478];
      mem_477_sv2v_reg <= w_data_i[477];
      mem_476_sv2v_reg <= w_data_i[476];
      mem_475_sv2v_reg <= w_data_i[475];
      mem_474_sv2v_reg <= w_data_i[474];
      mem_473_sv2v_reg <= w_data_i[473];
      mem_472_sv2v_reg <= w_data_i[472];
      mem_471_sv2v_reg <= w_data_i[471];
      mem_470_sv2v_reg <= w_data_i[470];
      mem_469_sv2v_reg <= w_data_i[469];
      mem_468_sv2v_reg <= w_data_i[468];
      mem_467_sv2v_reg <= w_data_i[467];
      mem_466_sv2v_reg <= w_data_i[466];
      mem_465_sv2v_reg <= w_data_i[465];
      mem_464_sv2v_reg <= w_data_i[464];
      mem_463_sv2v_reg <= w_data_i[463];
      mem_462_sv2v_reg <= w_data_i[462];
      mem_461_sv2v_reg <= w_data_i[461];
      mem_460_sv2v_reg <= w_data_i[460];
      mem_459_sv2v_reg <= w_data_i[459];
      mem_458_sv2v_reg <= w_data_i[458];
      mem_457_sv2v_reg <= w_data_i[457];
      mem_456_sv2v_reg <= w_data_i[456];
      mem_455_sv2v_reg <= w_data_i[455];
      mem_454_sv2v_reg <= w_data_i[454];
      mem_453_sv2v_reg <= w_data_i[453];
      mem_452_sv2v_reg <= w_data_i[452];
      mem_451_sv2v_reg <= w_data_i[451];
      mem_450_sv2v_reg <= w_data_i[450];
      mem_449_sv2v_reg <= w_data_i[449];
      mem_448_sv2v_reg <= w_data_i[448];
      mem_447_sv2v_reg <= w_data_i[447];
      mem_446_sv2v_reg <= w_data_i[446];
      mem_445_sv2v_reg <= w_data_i[445];
      mem_444_sv2v_reg <= w_data_i[444];
      mem_443_sv2v_reg <= w_data_i[443];
      mem_442_sv2v_reg <= w_data_i[442];
      mem_441_sv2v_reg <= w_data_i[441];
      mem_440_sv2v_reg <= w_data_i[440];
      mem_439_sv2v_reg <= w_data_i[439];
      mem_438_sv2v_reg <= w_data_i[438];
      mem_437_sv2v_reg <= w_data_i[437];
      mem_436_sv2v_reg <= w_data_i[436];
      mem_435_sv2v_reg <= w_data_i[435];
      mem_434_sv2v_reg <= w_data_i[434];
      mem_433_sv2v_reg <= w_data_i[433];
      mem_432_sv2v_reg <= w_data_i[432];
      mem_431_sv2v_reg <= w_data_i[431];
      mem_430_sv2v_reg <= w_data_i[430];
      mem_429_sv2v_reg <= w_data_i[429];
      mem_428_sv2v_reg <= w_data_i[428];
      mem_427_sv2v_reg <= w_data_i[427];
      mem_426_sv2v_reg <= w_data_i[426];
      mem_425_sv2v_reg <= w_data_i[425];
      mem_424_sv2v_reg <= w_data_i[424];
      mem_423_sv2v_reg <= w_data_i[423];
      mem_422_sv2v_reg <= w_data_i[422];
      mem_421_sv2v_reg <= w_data_i[421];
      mem_420_sv2v_reg <= w_data_i[420];
      mem_419_sv2v_reg <= w_data_i[419];
      mem_418_sv2v_reg <= w_data_i[418];
      mem_417_sv2v_reg <= w_data_i[417];
      mem_416_sv2v_reg <= w_data_i[416];
      mem_415_sv2v_reg <= w_data_i[415];
      mem_414_sv2v_reg <= w_data_i[414];
      mem_413_sv2v_reg <= w_data_i[413];
      mem_412_sv2v_reg <= w_data_i[412];
      mem_11_sv2v_reg <= w_data_i[11];
    end 
    if(N19) begin
      mem_411_sv2v_reg <= w_data_i[411];
      mem_410_sv2v_reg <= w_data_i[410];
      mem_409_sv2v_reg <= w_data_i[409];
      mem_408_sv2v_reg <= w_data_i[408];
      mem_407_sv2v_reg <= w_data_i[407];
      mem_406_sv2v_reg <= w_data_i[406];
      mem_405_sv2v_reg <= w_data_i[405];
      mem_404_sv2v_reg <= w_data_i[404];
      mem_403_sv2v_reg <= w_data_i[403];
      mem_402_sv2v_reg <= w_data_i[402];
      mem_401_sv2v_reg <= w_data_i[401];
      mem_400_sv2v_reg <= w_data_i[400];
      mem_399_sv2v_reg <= w_data_i[399];
      mem_398_sv2v_reg <= w_data_i[398];
      mem_397_sv2v_reg <= w_data_i[397];
      mem_396_sv2v_reg <= w_data_i[396];
      mem_395_sv2v_reg <= w_data_i[395];
      mem_394_sv2v_reg <= w_data_i[394];
      mem_393_sv2v_reg <= w_data_i[393];
      mem_392_sv2v_reg <= w_data_i[392];
      mem_391_sv2v_reg <= w_data_i[391];
      mem_390_sv2v_reg <= w_data_i[390];
      mem_389_sv2v_reg <= w_data_i[389];
      mem_388_sv2v_reg <= w_data_i[388];
      mem_387_sv2v_reg <= w_data_i[387];
      mem_386_sv2v_reg <= w_data_i[386];
      mem_385_sv2v_reg <= w_data_i[385];
      mem_384_sv2v_reg <= w_data_i[384];
      mem_383_sv2v_reg <= w_data_i[383];
      mem_382_sv2v_reg <= w_data_i[382];
      mem_381_sv2v_reg <= w_data_i[381];
      mem_380_sv2v_reg <= w_data_i[380];
      mem_379_sv2v_reg <= w_data_i[379];
      mem_378_sv2v_reg <= w_data_i[378];
      mem_377_sv2v_reg <= w_data_i[377];
      mem_376_sv2v_reg <= w_data_i[376];
      mem_375_sv2v_reg <= w_data_i[375];
      mem_374_sv2v_reg <= w_data_i[374];
      mem_373_sv2v_reg <= w_data_i[373];
      mem_372_sv2v_reg <= w_data_i[372];
      mem_371_sv2v_reg <= w_data_i[371];
      mem_370_sv2v_reg <= w_data_i[370];
      mem_369_sv2v_reg <= w_data_i[369];
      mem_368_sv2v_reg <= w_data_i[368];
      mem_367_sv2v_reg <= w_data_i[367];
      mem_366_sv2v_reg <= w_data_i[366];
      mem_365_sv2v_reg <= w_data_i[365];
      mem_364_sv2v_reg <= w_data_i[364];
      mem_363_sv2v_reg <= w_data_i[363];
      mem_362_sv2v_reg <= w_data_i[362];
      mem_361_sv2v_reg <= w_data_i[361];
      mem_360_sv2v_reg <= w_data_i[360];
      mem_359_sv2v_reg <= w_data_i[359];
      mem_358_sv2v_reg <= w_data_i[358];
      mem_357_sv2v_reg <= w_data_i[357];
      mem_356_sv2v_reg <= w_data_i[356];
      mem_355_sv2v_reg <= w_data_i[355];
      mem_354_sv2v_reg <= w_data_i[354];
      mem_353_sv2v_reg <= w_data_i[353];
      mem_352_sv2v_reg <= w_data_i[352];
      mem_351_sv2v_reg <= w_data_i[351];
      mem_350_sv2v_reg <= w_data_i[350];
      mem_349_sv2v_reg <= w_data_i[349];
      mem_348_sv2v_reg <= w_data_i[348];
      mem_347_sv2v_reg <= w_data_i[347];
      mem_346_sv2v_reg <= w_data_i[346];
      mem_345_sv2v_reg <= w_data_i[345];
      mem_344_sv2v_reg <= w_data_i[344];
      mem_343_sv2v_reg <= w_data_i[343];
      mem_342_sv2v_reg <= w_data_i[342];
      mem_341_sv2v_reg <= w_data_i[341];
      mem_340_sv2v_reg <= w_data_i[340];
      mem_339_sv2v_reg <= w_data_i[339];
      mem_338_sv2v_reg <= w_data_i[338];
      mem_337_sv2v_reg <= w_data_i[337];
      mem_336_sv2v_reg <= w_data_i[336];
      mem_335_sv2v_reg <= w_data_i[335];
      mem_334_sv2v_reg <= w_data_i[334];
      mem_333_sv2v_reg <= w_data_i[333];
      mem_332_sv2v_reg <= w_data_i[332];
      mem_331_sv2v_reg <= w_data_i[331];
      mem_330_sv2v_reg <= w_data_i[330];
      mem_329_sv2v_reg <= w_data_i[329];
      mem_328_sv2v_reg <= w_data_i[328];
      mem_327_sv2v_reg <= w_data_i[327];
      mem_326_sv2v_reg <= w_data_i[326];
      mem_325_sv2v_reg <= w_data_i[325];
      mem_324_sv2v_reg <= w_data_i[324];
      mem_323_sv2v_reg <= w_data_i[323];
      mem_322_sv2v_reg <= w_data_i[322];
      mem_321_sv2v_reg <= w_data_i[321];
      mem_320_sv2v_reg <= w_data_i[320];
      mem_319_sv2v_reg <= w_data_i[319];
      mem_318_sv2v_reg <= w_data_i[318];
      mem_317_sv2v_reg <= w_data_i[317];
      mem_316_sv2v_reg <= w_data_i[316];
      mem_315_sv2v_reg <= w_data_i[315];
      mem_314_sv2v_reg <= w_data_i[314];
      mem_313_sv2v_reg <= w_data_i[313];
      mem_12_sv2v_reg <= w_data_i[12];
    end 
    if(N20) begin
      mem_312_sv2v_reg <= w_data_i[312];
      mem_311_sv2v_reg <= w_data_i[311];
      mem_310_sv2v_reg <= w_data_i[310];
      mem_309_sv2v_reg <= w_data_i[309];
      mem_308_sv2v_reg <= w_data_i[308];
      mem_307_sv2v_reg <= w_data_i[307];
      mem_306_sv2v_reg <= w_data_i[306];
      mem_305_sv2v_reg <= w_data_i[305];
      mem_304_sv2v_reg <= w_data_i[304];
      mem_303_sv2v_reg <= w_data_i[303];
      mem_302_sv2v_reg <= w_data_i[302];
      mem_301_sv2v_reg <= w_data_i[301];
      mem_300_sv2v_reg <= w_data_i[300];
      mem_299_sv2v_reg <= w_data_i[299];
      mem_298_sv2v_reg <= w_data_i[298];
      mem_297_sv2v_reg <= w_data_i[297];
      mem_296_sv2v_reg <= w_data_i[296];
      mem_295_sv2v_reg <= w_data_i[295];
      mem_294_sv2v_reg <= w_data_i[294];
      mem_293_sv2v_reg <= w_data_i[293];
      mem_292_sv2v_reg <= w_data_i[292];
      mem_291_sv2v_reg <= w_data_i[291];
      mem_290_sv2v_reg <= w_data_i[290];
      mem_289_sv2v_reg <= w_data_i[289];
      mem_288_sv2v_reg <= w_data_i[288];
      mem_287_sv2v_reg <= w_data_i[287];
      mem_286_sv2v_reg <= w_data_i[286];
      mem_285_sv2v_reg <= w_data_i[285];
      mem_284_sv2v_reg <= w_data_i[284];
      mem_283_sv2v_reg <= w_data_i[283];
      mem_282_sv2v_reg <= w_data_i[282];
      mem_281_sv2v_reg <= w_data_i[281];
      mem_280_sv2v_reg <= w_data_i[280];
      mem_279_sv2v_reg <= w_data_i[279];
      mem_278_sv2v_reg <= w_data_i[278];
      mem_277_sv2v_reg <= w_data_i[277];
      mem_276_sv2v_reg <= w_data_i[276];
      mem_275_sv2v_reg <= w_data_i[275];
      mem_274_sv2v_reg <= w_data_i[274];
      mem_273_sv2v_reg <= w_data_i[273];
      mem_272_sv2v_reg <= w_data_i[272];
      mem_271_sv2v_reg <= w_data_i[271];
      mem_270_sv2v_reg <= w_data_i[270];
      mem_269_sv2v_reg <= w_data_i[269];
      mem_268_sv2v_reg <= w_data_i[268];
      mem_267_sv2v_reg <= w_data_i[267];
      mem_266_sv2v_reg <= w_data_i[266];
      mem_265_sv2v_reg <= w_data_i[265];
      mem_264_sv2v_reg <= w_data_i[264];
      mem_263_sv2v_reg <= w_data_i[263];
      mem_262_sv2v_reg <= w_data_i[262];
      mem_261_sv2v_reg <= w_data_i[261];
      mem_260_sv2v_reg <= w_data_i[260];
      mem_259_sv2v_reg <= w_data_i[259];
      mem_258_sv2v_reg <= w_data_i[258];
      mem_257_sv2v_reg <= w_data_i[257];
      mem_256_sv2v_reg <= w_data_i[256];
      mem_255_sv2v_reg <= w_data_i[255];
      mem_254_sv2v_reg <= w_data_i[254];
      mem_253_sv2v_reg <= w_data_i[253];
      mem_252_sv2v_reg <= w_data_i[252];
      mem_251_sv2v_reg <= w_data_i[251];
      mem_250_sv2v_reg <= w_data_i[250];
      mem_249_sv2v_reg <= w_data_i[249];
      mem_248_sv2v_reg <= w_data_i[248];
      mem_247_sv2v_reg <= w_data_i[247];
      mem_246_sv2v_reg <= w_data_i[246];
      mem_245_sv2v_reg <= w_data_i[245];
      mem_244_sv2v_reg <= w_data_i[244];
      mem_243_sv2v_reg <= w_data_i[243];
      mem_242_sv2v_reg <= w_data_i[242];
      mem_241_sv2v_reg <= w_data_i[241];
      mem_240_sv2v_reg <= w_data_i[240];
      mem_239_sv2v_reg <= w_data_i[239];
      mem_238_sv2v_reg <= w_data_i[238];
      mem_237_sv2v_reg <= w_data_i[237];
      mem_236_sv2v_reg <= w_data_i[236];
      mem_235_sv2v_reg <= w_data_i[235];
      mem_234_sv2v_reg <= w_data_i[234];
      mem_233_sv2v_reg <= w_data_i[233];
      mem_232_sv2v_reg <= w_data_i[232];
      mem_231_sv2v_reg <= w_data_i[231];
      mem_230_sv2v_reg <= w_data_i[230];
      mem_229_sv2v_reg <= w_data_i[229];
      mem_228_sv2v_reg <= w_data_i[228];
      mem_227_sv2v_reg <= w_data_i[227];
      mem_226_sv2v_reg <= w_data_i[226];
      mem_225_sv2v_reg <= w_data_i[225];
      mem_224_sv2v_reg <= w_data_i[224];
      mem_223_sv2v_reg <= w_data_i[223];
      mem_222_sv2v_reg <= w_data_i[222];
      mem_221_sv2v_reg <= w_data_i[221];
      mem_220_sv2v_reg <= w_data_i[220];
      mem_219_sv2v_reg <= w_data_i[219];
      mem_218_sv2v_reg <= w_data_i[218];
      mem_217_sv2v_reg <= w_data_i[217];
      mem_216_sv2v_reg <= w_data_i[216];
      mem_215_sv2v_reg <= w_data_i[215];
      mem_214_sv2v_reg <= w_data_i[214];
      mem_13_sv2v_reg <= w_data_i[13];
    end 
    if(N21) begin
      mem_213_sv2v_reg <= w_data_i[213];
      mem_212_sv2v_reg <= w_data_i[212];
      mem_211_sv2v_reg <= w_data_i[211];
      mem_210_sv2v_reg <= w_data_i[210];
      mem_209_sv2v_reg <= w_data_i[209];
      mem_208_sv2v_reg <= w_data_i[208];
      mem_207_sv2v_reg <= w_data_i[207];
      mem_206_sv2v_reg <= w_data_i[206];
      mem_205_sv2v_reg <= w_data_i[205];
      mem_204_sv2v_reg <= w_data_i[204];
      mem_203_sv2v_reg <= w_data_i[203];
      mem_202_sv2v_reg <= w_data_i[202];
      mem_201_sv2v_reg <= w_data_i[201];
      mem_200_sv2v_reg <= w_data_i[200];
      mem_199_sv2v_reg <= w_data_i[199];
      mem_198_sv2v_reg <= w_data_i[198];
      mem_197_sv2v_reg <= w_data_i[197];
      mem_196_sv2v_reg <= w_data_i[196];
      mem_195_sv2v_reg <= w_data_i[195];
      mem_194_sv2v_reg <= w_data_i[194];
      mem_193_sv2v_reg <= w_data_i[193];
      mem_192_sv2v_reg <= w_data_i[192];
      mem_191_sv2v_reg <= w_data_i[191];
      mem_190_sv2v_reg <= w_data_i[190];
      mem_189_sv2v_reg <= w_data_i[189];
      mem_188_sv2v_reg <= w_data_i[188];
      mem_187_sv2v_reg <= w_data_i[187];
      mem_186_sv2v_reg <= w_data_i[186];
      mem_185_sv2v_reg <= w_data_i[185];
      mem_184_sv2v_reg <= w_data_i[184];
      mem_183_sv2v_reg <= w_data_i[183];
      mem_182_sv2v_reg <= w_data_i[182];
      mem_181_sv2v_reg <= w_data_i[181];
      mem_180_sv2v_reg <= w_data_i[180];
      mem_179_sv2v_reg <= w_data_i[179];
      mem_178_sv2v_reg <= w_data_i[178];
      mem_177_sv2v_reg <= w_data_i[177];
      mem_176_sv2v_reg <= w_data_i[176];
      mem_175_sv2v_reg <= w_data_i[175];
      mem_174_sv2v_reg <= w_data_i[174];
      mem_173_sv2v_reg <= w_data_i[173];
      mem_172_sv2v_reg <= w_data_i[172];
      mem_171_sv2v_reg <= w_data_i[171];
      mem_170_sv2v_reg <= w_data_i[170];
      mem_169_sv2v_reg <= w_data_i[169];
      mem_168_sv2v_reg <= w_data_i[168];
      mem_167_sv2v_reg <= w_data_i[167];
      mem_166_sv2v_reg <= w_data_i[166];
      mem_165_sv2v_reg <= w_data_i[165];
      mem_164_sv2v_reg <= w_data_i[164];
      mem_163_sv2v_reg <= w_data_i[163];
      mem_162_sv2v_reg <= w_data_i[162];
      mem_161_sv2v_reg <= w_data_i[161];
      mem_160_sv2v_reg <= w_data_i[160];
      mem_159_sv2v_reg <= w_data_i[159];
      mem_158_sv2v_reg <= w_data_i[158];
      mem_157_sv2v_reg <= w_data_i[157];
      mem_156_sv2v_reg <= w_data_i[156];
      mem_155_sv2v_reg <= w_data_i[155];
      mem_154_sv2v_reg <= w_data_i[154];
      mem_153_sv2v_reg <= w_data_i[153];
      mem_152_sv2v_reg <= w_data_i[152];
      mem_151_sv2v_reg <= w_data_i[151];
      mem_150_sv2v_reg <= w_data_i[150];
      mem_149_sv2v_reg <= w_data_i[149];
      mem_148_sv2v_reg <= w_data_i[148];
      mem_147_sv2v_reg <= w_data_i[147];
      mem_146_sv2v_reg <= w_data_i[146];
      mem_145_sv2v_reg <= w_data_i[145];
      mem_144_sv2v_reg <= w_data_i[144];
      mem_143_sv2v_reg <= w_data_i[143];
      mem_142_sv2v_reg <= w_data_i[142];
      mem_141_sv2v_reg <= w_data_i[141];
      mem_140_sv2v_reg <= w_data_i[140];
      mem_139_sv2v_reg <= w_data_i[139];
      mem_138_sv2v_reg <= w_data_i[138];
      mem_137_sv2v_reg <= w_data_i[137];
      mem_136_sv2v_reg <= w_data_i[136];
      mem_135_sv2v_reg <= w_data_i[135];
      mem_134_sv2v_reg <= w_data_i[134];
      mem_133_sv2v_reg <= w_data_i[133];
      mem_132_sv2v_reg <= w_data_i[132];
      mem_131_sv2v_reg <= w_data_i[131];
      mem_130_sv2v_reg <= w_data_i[130];
      mem_129_sv2v_reg <= w_data_i[129];
      mem_128_sv2v_reg <= w_data_i[128];
      mem_127_sv2v_reg <= w_data_i[127];
      mem_126_sv2v_reg <= w_data_i[126];
      mem_125_sv2v_reg <= w_data_i[125];
      mem_124_sv2v_reg <= w_data_i[124];
      mem_123_sv2v_reg <= w_data_i[123];
      mem_122_sv2v_reg <= w_data_i[122];
      mem_121_sv2v_reg <= w_data_i[121];
      mem_120_sv2v_reg <= w_data_i[120];
      mem_119_sv2v_reg <= w_data_i[119];
      mem_118_sv2v_reg <= w_data_i[118];
      mem_117_sv2v_reg <= w_data_i[117];
      mem_116_sv2v_reg <= w_data_i[116];
      mem_115_sv2v_reg <= w_data_i[115];
      mem_14_sv2v_reg <= w_data_i[14];
    end 
    if(N22) begin
      mem_114_sv2v_reg <= w_data_i[114];
      mem_113_sv2v_reg <= w_data_i[113];
      mem_112_sv2v_reg <= w_data_i[112];
      mem_111_sv2v_reg <= w_data_i[111];
      mem_110_sv2v_reg <= w_data_i[110];
      mem_109_sv2v_reg <= w_data_i[109];
      mem_108_sv2v_reg <= w_data_i[108];
      mem_107_sv2v_reg <= w_data_i[107];
      mem_106_sv2v_reg <= w_data_i[106];
      mem_105_sv2v_reg <= w_data_i[105];
      mem_104_sv2v_reg <= w_data_i[104];
      mem_103_sv2v_reg <= w_data_i[103];
      mem_102_sv2v_reg <= w_data_i[102];
      mem_101_sv2v_reg <= w_data_i[101];
      mem_100_sv2v_reg <= w_data_i[100];
      mem_99_sv2v_reg <= w_data_i[99];
      mem_98_sv2v_reg <= w_data_i[98];
      mem_97_sv2v_reg <= w_data_i[97];
      mem_96_sv2v_reg <= w_data_i[96];
      mem_95_sv2v_reg <= w_data_i[95];
      mem_94_sv2v_reg <= w_data_i[94];
      mem_93_sv2v_reg <= w_data_i[93];
      mem_92_sv2v_reg <= w_data_i[92];
      mem_91_sv2v_reg <= w_data_i[91];
      mem_90_sv2v_reg <= w_data_i[90];
      mem_89_sv2v_reg <= w_data_i[89];
      mem_88_sv2v_reg <= w_data_i[88];
      mem_87_sv2v_reg <= w_data_i[87];
      mem_86_sv2v_reg <= w_data_i[86];
      mem_85_sv2v_reg <= w_data_i[85];
      mem_84_sv2v_reg <= w_data_i[84];
      mem_83_sv2v_reg <= w_data_i[83];
      mem_82_sv2v_reg <= w_data_i[82];
      mem_81_sv2v_reg <= w_data_i[81];
      mem_80_sv2v_reg <= w_data_i[80];
      mem_79_sv2v_reg <= w_data_i[79];
      mem_78_sv2v_reg <= w_data_i[78];
      mem_77_sv2v_reg <= w_data_i[77];
      mem_76_sv2v_reg <= w_data_i[76];
      mem_75_sv2v_reg <= w_data_i[75];
      mem_74_sv2v_reg <= w_data_i[74];
      mem_73_sv2v_reg <= w_data_i[73];
      mem_72_sv2v_reg <= w_data_i[72];
      mem_71_sv2v_reg <= w_data_i[71];
      mem_70_sv2v_reg <= w_data_i[70];
      mem_69_sv2v_reg <= w_data_i[69];
      mem_68_sv2v_reg <= w_data_i[68];
      mem_67_sv2v_reg <= w_data_i[67];
      mem_66_sv2v_reg <= w_data_i[66];
      mem_65_sv2v_reg <= w_data_i[65];
      mem_64_sv2v_reg <= w_data_i[64];
      mem_63_sv2v_reg <= w_data_i[63];
      mem_62_sv2v_reg <= w_data_i[62];
      mem_61_sv2v_reg <= w_data_i[61];
      mem_60_sv2v_reg <= w_data_i[60];
      mem_59_sv2v_reg <= w_data_i[59];
      mem_58_sv2v_reg <= w_data_i[58];
      mem_57_sv2v_reg <= w_data_i[57];
      mem_56_sv2v_reg <= w_data_i[56];
      mem_55_sv2v_reg <= w_data_i[55];
      mem_54_sv2v_reg <= w_data_i[54];
      mem_53_sv2v_reg <= w_data_i[53];
      mem_52_sv2v_reg <= w_data_i[52];
      mem_51_sv2v_reg <= w_data_i[51];
      mem_50_sv2v_reg <= w_data_i[50];
      mem_49_sv2v_reg <= w_data_i[49];
      mem_48_sv2v_reg <= w_data_i[48];
      mem_47_sv2v_reg <= w_data_i[47];
      mem_46_sv2v_reg <= w_data_i[46];
      mem_45_sv2v_reg <= w_data_i[45];
      mem_44_sv2v_reg <= w_data_i[44];
      mem_43_sv2v_reg <= w_data_i[43];
      mem_42_sv2v_reg <= w_data_i[42];
      mem_41_sv2v_reg <= w_data_i[41];
      mem_40_sv2v_reg <= w_data_i[40];
      mem_39_sv2v_reg <= w_data_i[39];
      mem_38_sv2v_reg <= w_data_i[38];
      mem_37_sv2v_reg <= w_data_i[37];
      mem_36_sv2v_reg <= w_data_i[36];
      mem_35_sv2v_reg <= w_data_i[35];
      mem_34_sv2v_reg <= w_data_i[34];
      mem_33_sv2v_reg <= w_data_i[33];
      mem_32_sv2v_reg <= w_data_i[32];
      mem_31_sv2v_reg <= w_data_i[31];
      mem_30_sv2v_reg <= w_data_i[30];
      mem_29_sv2v_reg <= w_data_i[29];
      mem_28_sv2v_reg <= w_data_i[28];
      mem_27_sv2v_reg <= w_data_i[27];
      mem_26_sv2v_reg <= w_data_i[26];
      mem_25_sv2v_reg <= w_data_i[25];
      mem_24_sv2v_reg <= w_data_i[24];
      mem_23_sv2v_reg <= w_data_i[23];
      mem_22_sv2v_reg <= w_data_i[22];
      mem_21_sv2v_reg <= w_data_i[21];
      mem_20_sv2v_reg <= w_data_i[20];
      mem_19_sv2v_reg <= w_data_i[19];
      mem_18_sv2v_reg <= w_data_i[18];
      mem_17_sv2v_reg <= w_data_i[17];
      mem_16_sv2v_reg <= w_data_i[16];
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p1600_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [1599:0] w_data_i;
  input [0:0] r_addr_i;
  output [1599:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [1599:0] r_data_o;

  bsg_mem_1r1w_synth_width_p1600_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p1600
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [1599:0] data_i;
  output [1599:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [1599:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p1600_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p49_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [5:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [5:0] count_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12;
  reg count_o_5_sv2v_reg,count_o_4_sv2v_reg,count_o_3_sv2v_reg,count_o_2_sv2v_reg,
  count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[5] = count_o_5_sv2v_reg;
  assign count_o[4] = count_o_4_sv2v_reg;
  assign count_o[3] = count_o_3_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N12 = reset_i | clear_i;
  assign { N10, N9, N8, N7, N6, N5 } = count_o + up_i;
  assign N11 = (N0)? up_i : 
               (N1)? N5 : 1'b0;
  assign N0 = clear_i;
  assign N1 = N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;

  always @(posedge clk_i) begin
    if(N12) begin
      count_o_5_sv2v_reg <= 1'b0;
      count_o_4_sv2v_reg <= 1'b0;
      count_o_3_sv2v_reg <= 1'b0;
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_5_sv2v_reg <= N10;
      count_o_4_sv2v_reg <= N9;
      count_o_3_sv2v_reg <= N8;
      count_o_2_sv2v_reg <= N7;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      count_o_0_sv2v_reg <= N11;
    end 
  end


endmodule



module bsg_mux_width_p32_els_p50
(
  data_i,
  sel_i,
  data_o
);

  input [1599:0] data_i;
  input [5:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312;
  assign N0 = N4 & N5;
  assign N1 = N0 & N6;
  assign N2 = N1 & N7;
  assign N3 = N2 & N8;
  assign N263 = N3 & N9;
  assign N4 = ~sel_i[5];
  assign N5 = ~sel_i[4];
  assign N6 = ~sel_i[3];
  assign N7 = ~sel_i[2];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = sel_i[5] & N14;
  assign N11 = N10 & N15;
  assign N12 = N11 & N16;
  assign N13 = N12 & N17;
  assign N264 = N13 & N18;
  assign N14 = ~sel_i[4];
  assign N15 = ~sel_i[3];
  assign N16 = ~sel_i[2];
  assign N17 = ~sel_i[0];
  assign N18 = ~sel_i[1];
  assign N19 = N23 & N24;
  assign N20 = N19 & N25;
  assign N21 = N20 & N26;
  assign N22 = N21 & sel_i[0];
  assign N265 = N22 & N27;
  assign N23 = ~sel_i[5];
  assign N24 = ~sel_i[4];
  assign N25 = ~sel_i[3];
  assign N26 = ~sel_i[2];
  assign N27 = ~sel_i[1];
  assign N28 = N32 & N33;
  assign N29 = N28 & N34;
  assign N30 = N29 & N35;
  assign N31 = N30 & N36;
  assign N267 = N31 & sel_i[1];
  assign N32 = ~sel_i[5];
  assign N33 = ~sel_i[4];
  assign N34 = ~sel_i[3];
  assign N35 = ~sel_i[2];
  assign N36 = ~sel_i[0];
  assign N37 = N41 & N42;
  assign N38 = N37 & N43;
  assign N39 = N38 & N44;
  assign N40 = N39 & sel_i[0];
  assign N269 = N40 & sel_i[1];
  assign N41 = ~sel_i[5];
  assign N42 = ~sel_i[4];
  assign N43 = ~sel_i[3];
  assign N44 = ~sel_i[2];
  assign N45 = N49 & N50;
  assign N46 = N45 & N51;
  assign N47 = N46 & sel_i[2];
  assign N48 = N47 & N52;
  assign N271 = N48 & N53;
  assign N49 = ~sel_i[5];
  assign N50 = ~sel_i[4];
  assign N51 = ~sel_i[3];
  assign N52 = ~sel_i[0];
  assign N53 = ~sel_i[1];
  assign N54 = N58 & N59;
  assign N55 = N54 & N60;
  assign N56 = N55 & sel_i[2];
  assign N57 = N56 & sel_i[0];
  assign N273 = N57 & N61;
  assign N58 = ~sel_i[5];
  assign N59 = ~sel_i[4];
  assign N60 = ~sel_i[3];
  assign N61 = ~sel_i[1];
  assign N62 = N66 & N67;
  assign N63 = N62 & N68;
  assign N64 = N63 & sel_i[2];
  assign N65 = N64 & N69;
  assign N275 = N65 & sel_i[1];
  assign N66 = ~sel_i[5];
  assign N67 = ~sel_i[4];
  assign N68 = ~sel_i[3];
  assign N69 = ~sel_i[0];
  assign N70 = N74 & N75;
  assign N71 = N70 & N76;
  assign N72 = N71 & sel_i[2];
  assign N73 = N72 & sel_i[0];
  assign N277 = N73 & sel_i[1];
  assign N74 = ~sel_i[5];
  assign N75 = ~sel_i[4];
  assign N76 = ~sel_i[3];
  assign N77 = N81 & N82;
  assign N78 = N77 & sel_i[3];
  assign N79 = N78 & N83;
  assign N80 = N79 & N84;
  assign N279 = N80 & N85;
  assign N81 = ~sel_i[5];
  assign N82 = ~sel_i[4];
  assign N83 = ~sel_i[2];
  assign N84 = ~sel_i[0];
  assign N85 = ~sel_i[1];
  assign N86 = N90 & N91;
  assign N87 = N86 & sel_i[3];
  assign N88 = N87 & N92;
  assign N89 = N88 & sel_i[0];
  assign N281 = N89 & N93;
  assign N90 = ~sel_i[5];
  assign N91 = ~sel_i[4];
  assign N92 = ~sel_i[2];
  assign N93 = ~sel_i[1];
  assign N94 = N98 & N99;
  assign N95 = N94 & sel_i[3];
  assign N96 = N95 & N100;
  assign N97 = N96 & N101;
  assign N283 = N97 & sel_i[1];
  assign N98 = ~sel_i[5];
  assign N99 = ~sel_i[4];
  assign N100 = ~sel_i[2];
  assign N101 = ~sel_i[0];
  assign N102 = N106 & N107;
  assign N103 = N102 & sel_i[3];
  assign N104 = N103 & N108;
  assign N105 = N104 & sel_i[0];
  assign N285 = N105 & sel_i[1];
  assign N106 = ~sel_i[5];
  assign N107 = ~sel_i[4];
  assign N108 = ~sel_i[2];
  assign N109 = N113 & N114;
  assign N110 = N109 & sel_i[3];
  assign N111 = N110 & sel_i[2];
  assign N112 = N111 & N115;
  assign N287 = N112 & N116;
  assign N113 = ~sel_i[5];
  assign N114 = ~sel_i[4];
  assign N115 = ~sel_i[0];
  assign N116 = ~sel_i[1];
  assign N117 = N121 & N122;
  assign N118 = N117 & sel_i[3];
  assign N119 = N118 & sel_i[2];
  assign N120 = N119 & sel_i[0];
  assign N289 = N120 & N123;
  assign N121 = ~sel_i[5];
  assign N122 = ~sel_i[4];
  assign N123 = ~sel_i[1];
  assign N124 = N128 & N129;
  assign N125 = N124 & sel_i[3];
  assign N126 = N125 & sel_i[2];
  assign N127 = N126 & N130;
  assign N291 = N127 & sel_i[1];
  assign N128 = ~sel_i[5];
  assign N129 = ~sel_i[4];
  assign N130 = ~sel_i[0];
  assign N131 = N135 & N136;
  assign N132 = N131 & sel_i[3];
  assign N133 = N132 & sel_i[2];
  assign N134 = N133 & sel_i[0];
  assign N293 = N134 & sel_i[1];
  assign N135 = ~sel_i[5];
  assign N136 = ~sel_i[4];
  assign N137 = N141 & sel_i[4];
  assign N138 = N137 & N142;
  assign N139 = N138 & N143;
  assign N140 = N139 & N144;
  assign N295 = N140 & N145;
  assign N141 = ~sel_i[5];
  assign N142 = ~sel_i[3];
  assign N143 = ~sel_i[2];
  assign N144 = ~sel_i[0];
  assign N145 = ~sel_i[1];
  assign N146 = N150 & sel_i[4];
  assign N147 = N146 & N151;
  assign N148 = N147 & N152;
  assign N149 = N148 & sel_i[0];
  assign N297 = N149 & N153;
  assign N150 = ~sel_i[5];
  assign N151 = ~sel_i[3];
  assign N152 = ~sel_i[2];
  assign N153 = ~sel_i[1];
  assign N299 = sel_i[4] & N154 & (N155 & N156) & sel_i[1];
  assign N154 = ~sel_i[3];
  assign N155 = ~sel_i[2];
  assign N156 = ~sel_i[0];
  assign N300 = sel_i[4] & N157 & (N158 & sel_i[0]) & sel_i[1];
  assign N157 = ~sel_i[3];
  assign N158 = ~sel_i[2];
  assign N301 = sel_i[4] & N159 & (sel_i[2] & N160) & N161;
  assign N159 = ~sel_i[3];
  assign N160 = ~sel_i[0];
  assign N161 = ~sel_i[1];
  assign N302 = sel_i[4] & N162 & (sel_i[2] & sel_i[0]) & N163;
  assign N162 = ~sel_i[3];
  assign N163 = ~sel_i[1];
  assign N303 = sel_i[4] & N164 & (sel_i[2] & N165) & sel_i[1];
  assign N164 = ~sel_i[3];
  assign N165 = ~sel_i[0];
  assign N304 = sel_i[4] & N166 & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N166 = ~sel_i[3];
  assign N305 = sel_i[4] & sel_i[3] & (N167 & N168) & N169;
  assign N167 = ~sel_i[2];
  assign N168 = ~sel_i[0];
  assign N169 = ~sel_i[1];
  assign N306 = sel_i[4] & sel_i[3] & (N170 & sel_i[0]) & N171;
  assign N170 = ~sel_i[2];
  assign N171 = ~sel_i[1];
  assign N307 = sel_i[4] & sel_i[3] & (N172 & N173) & sel_i[1];
  assign N172 = ~sel_i[2];
  assign N173 = ~sel_i[0];
  assign N308 = sel_i[4] & sel_i[3] & (N174 & sel_i[0]) & sel_i[1];
  assign N174 = ~sel_i[2];
  assign N309 = sel_i[4] & sel_i[3] & (sel_i[2] & N175) & N176;
  assign N175 = ~sel_i[0];
  assign N176 = ~sel_i[1];
  assign N310 = sel_i[4] & sel_i[3] & (sel_i[2] & sel_i[0]) & N177;
  assign N177 = ~sel_i[1];
  assign N311 = sel_i[4] & sel_i[3] & (sel_i[2] & N178) & sel_i[1];
  assign N178 = ~sel_i[0];
  assign N312 = sel_i[4] & sel_i[3] & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N179 = sel_i[5] & N183;
  assign N180 = N179 & N184;
  assign N181 = N180 & N185;
  assign N182 = N181 & sel_i[0];
  assign N266 = N182 & N186;
  assign N183 = ~sel_i[4];
  assign N184 = ~sel_i[3];
  assign N185 = ~sel_i[2];
  assign N186 = ~sel_i[1];
  assign N268 = sel_i[5] & N187 & (N188 & N189) & sel_i[1];
  assign N187 = ~sel_i[3];
  assign N188 = ~sel_i[2];
  assign N189 = ~sel_i[0];
  assign N270 = sel_i[5] & N190 & (N191 & sel_i[0]) & sel_i[1];
  assign N190 = ~sel_i[3];
  assign N191 = ~sel_i[2];
  assign N272 = sel_i[5] & N192 & (sel_i[2] & N193) & N194;
  assign N192 = ~sel_i[3];
  assign N193 = ~sel_i[0];
  assign N194 = ~sel_i[1];
  assign N274 = sel_i[5] & N195 & (sel_i[2] & sel_i[0]) & N196;
  assign N195 = ~sel_i[3];
  assign N196 = ~sel_i[1];
  assign N276 = sel_i[5] & N197 & (sel_i[2] & N198) & sel_i[1];
  assign N197 = ~sel_i[3];
  assign N198 = ~sel_i[0];
  assign N278 = sel_i[5] & N199 & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N199 = ~sel_i[3];
  assign N280 = sel_i[5] & sel_i[3] & (N200 & N201) & N202;
  assign N200 = ~sel_i[2];
  assign N201 = ~sel_i[0];
  assign N202 = ~sel_i[1];
  assign N282 = sel_i[5] & sel_i[3] & (N203 & sel_i[0]) & N204;
  assign N203 = ~sel_i[2];
  assign N204 = ~sel_i[1];
  assign N284 = sel_i[5] & sel_i[3] & (N205 & N206) & sel_i[1];
  assign N205 = ~sel_i[2];
  assign N206 = ~sel_i[0];
  assign N286 = sel_i[5] & sel_i[3] & (N207 & sel_i[0]) & sel_i[1];
  assign N207 = ~sel_i[2];
  assign N288 = sel_i[5] & sel_i[3] & (sel_i[2] & N208) & N209;
  assign N208 = ~sel_i[0];
  assign N209 = ~sel_i[1];
  assign N290 = sel_i[5] & sel_i[3] & (sel_i[2] & sel_i[0]) & N210;
  assign N210 = ~sel_i[1];
  assign N292 = sel_i[5] & sel_i[3] & (sel_i[2] & N211) & sel_i[1];
  assign N211 = ~sel_i[0];
  assign N294 = sel_i[5] & sel_i[3] & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N296 = sel_i[5] & sel_i[4] & N212;
  assign N212 = ~sel_i[0];
  assign N298 = sel_i[5] & sel_i[4] & sel_i[0];
  assign data_o[31] = (N213)? data_i[31] : 
                      (N214)? data_i[63] : 
                      (N215)? data_i[95] : 
                      (N216)? data_i[127] : 
                      (N217)? data_i[159] : 
                      (N218)? data_i[191] : 
                      (N219)? data_i[223] : 
                      (N220)? data_i[255] : 
                      (N221)? data_i[287] : 
                      (N222)? data_i[319] : 
                      (N223)? data_i[351] : 
                      (N224)? data_i[383] : 
                      (N225)? data_i[415] : 
                      (N226)? data_i[447] : 
                      (N227)? data_i[479] : 
                      (N228)? data_i[511] : 
                      (N229)? data_i[543] : 
                      (N230)? data_i[575] : 
                      (N231)? data_i[607] : 
                      (N232)? data_i[639] : 
                      (N233)? data_i[671] : 
                      (N234)? data_i[703] : 
                      (N235)? data_i[735] : 
                      (N236)? data_i[767] : 
                      (N237)? data_i[799] : 
                      (N238)? data_i[831] : 
                      (N239)? data_i[863] : 
                      (N240)? data_i[895] : 
                      (N241)? data_i[927] : 
                      (N242)? data_i[959] : 
                      (N243)? data_i[991] : 
                      (N244)? data_i[1023] : 
                      (N245)? data_i[1055] : 
                      (N246)? data_i[1087] : 
                      (N247)? data_i[1119] : 
                      (N248)? data_i[1151] : 
                      (N249)? data_i[1183] : 
                      (N250)? data_i[1215] : 
                      (N251)? data_i[1247] : 
                      (N252)? data_i[1279] : 
                      (N253)? data_i[1311] : 
                      (N254)? data_i[1343] : 
                      (N255)? data_i[1375] : 
                      (N256)? data_i[1407] : 
                      (N257)? data_i[1439] : 
                      (N258)? data_i[1471] : 
                      (N259)? data_i[1503] : 
                      (N260)? data_i[1535] : 
                      (N261)? data_i[1567] : 
                      (N262)? data_i[1599] : 1'b0;
  assign N213 = N263;
  assign N214 = N265;
  assign N215 = N267;
  assign N216 = N269;
  assign N217 = N271;
  assign N218 = N273;
  assign N219 = N275;
  assign N220 = N277;
  assign N221 = N279;
  assign N222 = N281;
  assign N223 = N283;
  assign N224 = N285;
  assign N225 = N287;
  assign N226 = N289;
  assign N227 = N291;
  assign N228 = N293;
  assign N229 = N295;
  assign N230 = N297;
  assign N231 = N299;
  assign N232 = N300;
  assign N233 = N301;
  assign N234 = N302;
  assign N235 = N303;
  assign N236 = N304;
  assign N237 = N305;
  assign N238 = N306;
  assign N239 = N307;
  assign N240 = N308;
  assign N241 = N309;
  assign N242 = N310;
  assign N243 = N311;
  assign N244 = N312;
  assign N245 = N264;
  assign N246 = N266;
  assign N247 = N268;
  assign N248 = N270;
  assign N249 = N272;
  assign N250 = N274;
  assign N251 = N276;
  assign N252 = N278;
  assign N253 = N280;
  assign N254 = N282;
  assign N255 = N284;
  assign N256 = N286;
  assign N257 = N288;
  assign N258 = N290;
  assign N259 = N292;
  assign N260 = N294;
  assign N261 = N296;
  assign N262 = N298;
  assign data_o[30] = (N213)? data_i[30] : 
                      (N214)? data_i[62] : 
                      (N215)? data_i[94] : 
                      (N216)? data_i[126] : 
                      (N217)? data_i[158] : 
                      (N218)? data_i[190] : 
                      (N219)? data_i[222] : 
                      (N220)? data_i[254] : 
                      (N221)? data_i[286] : 
                      (N222)? data_i[318] : 
                      (N223)? data_i[350] : 
                      (N224)? data_i[382] : 
                      (N225)? data_i[414] : 
                      (N226)? data_i[446] : 
                      (N227)? data_i[478] : 
                      (N228)? data_i[510] : 
                      (N229)? data_i[542] : 
                      (N230)? data_i[574] : 
                      (N231)? data_i[606] : 
                      (N232)? data_i[638] : 
                      (N233)? data_i[670] : 
                      (N234)? data_i[702] : 
                      (N235)? data_i[734] : 
                      (N236)? data_i[766] : 
                      (N237)? data_i[798] : 
                      (N238)? data_i[830] : 
                      (N239)? data_i[862] : 
                      (N240)? data_i[894] : 
                      (N241)? data_i[926] : 
                      (N242)? data_i[958] : 
                      (N243)? data_i[990] : 
                      (N244)? data_i[1022] : 
                      (N245)? data_i[1054] : 
                      (N246)? data_i[1086] : 
                      (N247)? data_i[1118] : 
                      (N248)? data_i[1150] : 
                      (N249)? data_i[1182] : 
                      (N250)? data_i[1214] : 
                      (N251)? data_i[1246] : 
                      (N252)? data_i[1278] : 
                      (N253)? data_i[1310] : 
                      (N254)? data_i[1342] : 
                      (N255)? data_i[1374] : 
                      (N256)? data_i[1406] : 
                      (N257)? data_i[1438] : 
                      (N258)? data_i[1470] : 
                      (N259)? data_i[1502] : 
                      (N260)? data_i[1534] : 
                      (N261)? data_i[1566] : 
                      (N262)? data_i[1598] : 1'b0;
  assign data_o[29] = (N213)? data_i[29] : 
                      (N214)? data_i[61] : 
                      (N215)? data_i[93] : 
                      (N216)? data_i[125] : 
                      (N217)? data_i[157] : 
                      (N218)? data_i[189] : 
                      (N219)? data_i[221] : 
                      (N220)? data_i[253] : 
                      (N221)? data_i[285] : 
                      (N222)? data_i[317] : 
                      (N223)? data_i[349] : 
                      (N224)? data_i[381] : 
                      (N225)? data_i[413] : 
                      (N226)? data_i[445] : 
                      (N227)? data_i[477] : 
                      (N228)? data_i[509] : 
                      (N229)? data_i[541] : 
                      (N230)? data_i[573] : 
                      (N231)? data_i[605] : 
                      (N232)? data_i[637] : 
                      (N233)? data_i[669] : 
                      (N234)? data_i[701] : 
                      (N235)? data_i[733] : 
                      (N236)? data_i[765] : 
                      (N237)? data_i[797] : 
                      (N238)? data_i[829] : 
                      (N239)? data_i[861] : 
                      (N240)? data_i[893] : 
                      (N241)? data_i[925] : 
                      (N242)? data_i[957] : 
                      (N243)? data_i[989] : 
                      (N244)? data_i[1021] : 
                      (N245)? data_i[1053] : 
                      (N246)? data_i[1085] : 
                      (N247)? data_i[1117] : 
                      (N248)? data_i[1149] : 
                      (N249)? data_i[1181] : 
                      (N250)? data_i[1213] : 
                      (N251)? data_i[1245] : 
                      (N252)? data_i[1277] : 
                      (N253)? data_i[1309] : 
                      (N254)? data_i[1341] : 
                      (N255)? data_i[1373] : 
                      (N256)? data_i[1405] : 
                      (N257)? data_i[1437] : 
                      (N258)? data_i[1469] : 
                      (N259)? data_i[1501] : 
                      (N260)? data_i[1533] : 
                      (N261)? data_i[1565] : 
                      (N262)? data_i[1597] : 1'b0;
  assign data_o[28] = (N213)? data_i[28] : 
                      (N214)? data_i[60] : 
                      (N215)? data_i[92] : 
                      (N216)? data_i[124] : 
                      (N217)? data_i[156] : 
                      (N218)? data_i[188] : 
                      (N219)? data_i[220] : 
                      (N220)? data_i[252] : 
                      (N221)? data_i[284] : 
                      (N222)? data_i[316] : 
                      (N223)? data_i[348] : 
                      (N224)? data_i[380] : 
                      (N225)? data_i[412] : 
                      (N226)? data_i[444] : 
                      (N227)? data_i[476] : 
                      (N228)? data_i[508] : 
                      (N229)? data_i[540] : 
                      (N230)? data_i[572] : 
                      (N231)? data_i[604] : 
                      (N232)? data_i[636] : 
                      (N233)? data_i[668] : 
                      (N234)? data_i[700] : 
                      (N235)? data_i[732] : 
                      (N236)? data_i[764] : 
                      (N237)? data_i[796] : 
                      (N238)? data_i[828] : 
                      (N239)? data_i[860] : 
                      (N240)? data_i[892] : 
                      (N241)? data_i[924] : 
                      (N242)? data_i[956] : 
                      (N243)? data_i[988] : 
                      (N244)? data_i[1020] : 
                      (N245)? data_i[1052] : 
                      (N246)? data_i[1084] : 
                      (N247)? data_i[1116] : 
                      (N248)? data_i[1148] : 
                      (N249)? data_i[1180] : 
                      (N250)? data_i[1212] : 
                      (N251)? data_i[1244] : 
                      (N252)? data_i[1276] : 
                      (N253)? data_i[1308] : 
                      (N254)? data_i[1340] : 
                      (N255)? data_i[1372] : 
                      (N256)? data_i[1404] : 
                      (N257)? data_i[1436] : 
                      (N258)? data_i[1468] : 
                      (N259)? data_i[1500] : 
                      (N260)? data_i[1532] : 
                      (N261)? data_i[1564] : 
                      (N262)? data_i[1596] : 1'b0;
  assign data_o[27] = (N213)? data_i[27] : 
                      (N214)? data_i[59] : 
                      (N215)? data_i[91] : 
                      (N216)? data_i[123] : 
                      (N217)? data_i[155] : 
                      (N218)? data_i[187] : 
                      (N219)? data_i[219] : 
                      (N220)? data_i[251] : 
                      (N221)? data_i[283] : 
                      (N222)? data_i[315] : 
                      (N223)? data_i[347] : 
                      (N224)? data_i[379] : 
                      (N225)? data_i[411] : 
                      (N226)? data_i[443] : 
                      (N227)? data_i[475] : 
                      (N228)? data_i[507] : 
                      (N229)? data_i[539] : 
                      (N230)? data_i[571] : 
                      (N231)? data_i[603] : 
                      (N232)? data_i[635] : 
                      (N233)? data_i[667] : 
                      (N234)? data_i[699] : 
                      (N235)? data_i[731] : 
                      (N236)? data_i[763] : 
                      (N237)? data_i[795] : 
                      (N238)? data_i[827] : 
                      (N239)? data_i[859] : 
                      (N240)? data_i[891] : 
                      (N241)? data_i[923] : 
                      (N242)? data_i[955] : 
                      (N243)? data_i[987] : 
                      (N244)? data_i[1019] : 
                      (N245)? data_i[1051] : 
                      (N246)? data_i[1083] : 
                      (N247)? data_i[1115] : 
                      (N248)? data_i[1147] : 
                      (N249)? data_i[1179] : 
                      (N250)? data_i[1211] : 
                      (N251)? data_i[1243] : 
                      (N252)? data_i[1275] : 
                      (N253)? data_i[1307] : 
                      (N254)? data_i[1339] : 
                      (N255)? data_i[1371] : 
                      (N256)? data_i[1403] : 
                      (N257)? data_i[1435] : 
                      (N258)? data_i[1467] : 
                      (N259)? data_i[1499] : 
                      (N260)? data_i[1531] : 
                      (N261)? data_i[1563] : 
                      (N262)? data_i[1595] : 1'b0;
  assign data_o[26] = (N213)? data_i[26] : 
                      (N214)? data_i[58] : 
                      (N215)? data_i[90] : 
                      (N216)? data_i[122] : 
                      (N217)? data_i[154] : 
                      (N218)? data_i[186] : 
                      (N219)? data_i[218] : 
                      (N220)? data_i[250] : 
                      (N221)? data_i[282] : 
                      (N222)? data_i[314] : 
                      (N223)? data_i[346] : 
                      (N224)? data_i[378] : 
                      (N225)? data_i[410] : 
                      (N226)? data_i[442] : 
                      (N227)? data_i[474] : 
                      (N228)? data_i[506] : 
                      (N229)? data_i[538] : 
                      (N230)? data_i[570] : 
                      (N231)? data_i[602] : 
                      (N232)? data_i[634] : 
                      (N233)? data_i[666] : 
                      (N234)? data_i[698] : 
                      (N235)? data_i[730] : 
                      (N236)? data_i[762] : 
                      (N237)? data_i[794] : 
                      (N238)? data_i[826] : 
                      (N239)? data_i[858] : 
                      (N240)? data_i[890] : 
                      (N241)? data_i[922] : 
                      (N242)? data_i[954] : 
                      (N243)? data_i[986] : 
                      (N244)? data_i[1018] : 
                      (N245)? data_i[1050] : 
                      (N246)? data_i[1082] : 
                      (N247)? data_i[1114] : 
                      (N248)? data_i[1146] : 
                      (N249)? data_i[1178] : 
                      (N250)? data_i[1210] : 
                      (N251)? data_i[1242] : 
                      (N252)? data_i[1274] : 
                      (N253)? data_i[1306] : 
                      (N254)? data_i[1338] : 
                      (N255)? data_i[1370] : 
                      (N256)? data_i[1402] : 
                      (N257)? data_i[1434] : 
                      (N258)? data_i[1466] : 
                      (N259)? data_i[1498] : 
                      (N260)? data_i[1530] : 
                      (N261)? data_i[1562] : 
                      (N262)? data_i[1594] : 1'b0;
  assign data_o[25] = (N213)? data_i[25] : 
                      (N214)? data_i[57] : 
                      (N215)? data_i[89] : 
                      (N216)? data_i[121] : 
                      (N217)? data_i[153] : 
                      (N218)? data_i[185] : 
                      (N219)? data_i[217] : 
                      (N220)? data_i[249] : 
                      (N221)? data_i[281] : 
                      (N222)? data_i[313] : 
                      (N223)? data_i[345] : 
                      (N224)? data_i[377] : 
                      (N225)? data_i[409] : 
                      (N226)? data_i[441] : 
                      (N227)? data_i[473] : 
                      (N228)? data_i[505] : 
                      (N229)? data_i[537] : 
                      (N230)? data_i[569] : 
                      (N231)? data_i[601] : 
                      (N232)? data_i[633] : 
                      (N233)? data_i[665] : 
                      (N234)? data_i[697] : 
                      (N235)? data_i[729] : 
                      (N236)? data_i[761] : 
                      (N237)? data_i[793] : 
                      (N238)? data_i[825] : 
                      (N239)? data_i[857] : 
                      (N240)? data_i[889] : 
                      (N241)? data_i[921] : 
                      (N242)? data_i[953] : 
                      (N243)? data_i[985] : 
                      (N244)? data_i[1017] : 
                      (N245)? data_i[1049] : 
                      (N246)? data_i[1081] : 
                      (N247)? data_i[1113] : 
                      (N248)? data_i[1145] : 
                      (N249)? data_i[1177] : 
                      (N250)? data_i[1209] : 
                      (N251)? data_i[1241] : 
                      (N252)? data_i[1273] : 
                      (N253)? data_i[1305] : 
                      (N254)? data_i[1337] : 
                      (N255)? data_i[1369] : 
                      (N256)? data_i[1401] : 
                      (N257)? data_i[1433] : 
                      (N258)? data_i[1465] : 
                      (N259)? data_i[1497] : 
                      (N260)? data_i[1529] : 
                      (N261)? data_i[1561] : 
                      (N262)? data_i[1593] : 1'b0;
  assign data_o[24] = (N213)? data_i[24] : 
                      (N214)? data_i[56] : 
                      (N215)? data_i[88] : 
                      (N216)? data_i[120] : 
                      (N217)? data_i[152] : 
                      (N218)? data_i[184] : 
                      (N219)? data_i[216] : 
                      (N220)? data_i[248] : 
                      (N221)? data_i[280] : 
                      (N222)? data_i[312] : 
                      (N223)? data_i[344] : 
                      (N224)? data_i[376] : 
                      (N225)? data_i[408] : 
                      (N226)? data_i[440] : 
                      (N227)? data_i[472] : 
                      (N228)? data_i[504] : 
                      (N229)? data_i[536] : 
                      (N230)? data_i[568] : 
                      (N231)? data_i[600] : 
                      (N232)? data_i[632] : 
                      (N233)? data_i[664] : 
                      (N234)? data_i[696] : 
                      (N235)? data_i[728] : 
                      (N236)? data_i[760] : 
                      (N237)? data_i[792] : 
                      (N238)? data_i[824] : 
                      (N239)? data_i[856] : 
                      (N240)? data_i[888] : 
                      (N241)? data_i[920] : 
                      (N242)? data_i[952] : 
                      (N243)? data_i[984] : 
                      (N244)? data_i[1016] : 
                      (N245)? data_i[1048] : 
                      (N246)? data_i[1080] : 
                      (N247)? data_i[1112] : 
                      (N248)? data_i[1144] : 
                      (N249)? data_i[1176] : 
                      (N250)? data_i[1208] : 
                      (N251)? data_i[1240] : 
                      (N252)? data_i[1272] : 
                      (N253)? data_i[1304] : 
                      (N254)? data_i[1336] : 
                      (N255)? data_i[1368] : 
                      (N256)? data_i[1400] : 
                      (N257)? data_i[1432] : 
                      (N258)? data_i[1464] : 
                      (N259)? data_i[1496] : 
                      (N260)? data_i[1528] : 
                      (N261)? data_i[1560] : 
                      (N262)? data_i[1592] : 1'b0;
  assign data_o[23] = (N213)? data_i[23] : 
                      (N214)? data_i[55] : 
                      (N215)? data_i[87] : 
                      (N216)? data_i[119] : 
                      (N217)? data_i[151] : 
                      (N218)? data_i[183] : 
                      (N219)? data_i[215] : 
                      (N220)? data_i[247] : 
                      (N221)? data_i[279] : 
                      (N222)? data_i[311] : 
                      (N223)? data_i[343] : 
                      (N224)? data_i[375] : 
                      (N225)? data_i[407] : 
                      (N226)? data_i[439] : 
                      (N227)? data_i[471] : 
                      (N228)? data_i[503] : 
                      (N229)? data_i[535] : 
                      (N230)? data_i[567] : 
                      (N231)? data_i[599] : 
                      (N232)? data_i[631] : 
                      (N233)? data_i[663] : 
                      (N234)? data_i[695] : 
                      (N235)? data_i[727] : 
                      (N236)? data_i[759] : 
                      (N237)? data_i[791] : 
                      (N238)? data_i[823] : 
                      (N239)? data_i[855] : 
                      (N240)? data_i[887] : 
                      (N241)? data_i[919] : 
                      (N242)? data_i[951] : 
                      (N243)? data_i[983] : 
                      (N244)? data_i[1015] : 
                      (N245)? data_i[1047] : 
                      (N246)? data_i[1079] : 
                      (N247)? data_i[1111] : 
                      (N248)? data_i[1143] : 
                      (N249)? data_i[1175] : 
                      (N250)? data_i[1207] : 
                      (N251)? data_i[1239] : 
                      (N252)? data_i[1271] : 
                      (N253)? data_i[1303] : 
                      (N254)? data_i[1335] : 
                      (N255)? data_i[1367] : 
                      (N256)? data_i[1399] : 
                      (N257)? data_i[1431] : 
                      (N258)? data_i[1463] : 
                      (N259)? data_i[1495] : 
                      (N260)? data_i[1527] : 
                      (N261)? data_i[1559] : 
                      (N262)? data_i[1591] : 1'b0;
  assign data_o[22] = (N213)? data_i[22] : 
                      (N214)? data_i[54] : 
                      (N215)? data_i[86] : 
                      (N216)? data_i[118] : 
                      (N217)? data_i[150] : 
                      (N218)? data_i[182] : 
                      (N219)? data_i[214] : 
                      (N220)? data_i[246] : 
                      (N221)? data_i[278] : 
                      (N222)? data_i[310] : 
                      (N223)? data_i[342] : 
                      (N224)? data_i[374] : 
                      (N225)? data_i[406] : 
                      (N226)? data_i[438] : 
                      (N227)? data_i[470] : 
                      (N228)? data_i[502] : 
                      (N229)? data_i[534] : 
                      (N230)? data_i[566] : 
                      (N231)? data_i[598] : 
                      (N232)? data_i[630] : 
                      (N233)? data_i[662] : 
                      (N234)? data_i[694] : 
                      (N235)? data_i[726] : 
                      (N236)? data_i[758] : 
                      (N237)? data_i[790] : 
                      (N238)? data_i[822] : 
                      (N239)? data_i[854] : 
                      (N240)? data_i[886] : 
                      (N241)? data_i[918] : 
                      (N242)? data_i[950] : 
                      (N243)? data_i[982] : 
                      (N244)? data_i[1014] : 
                      (N245)? data_i[1046] : 
                      (N246)? data_i[1078] : 
                      (N247)? data_i[1110] : 
                      (N248)? data_i[1142] : 
                      (N249)? data_i[1174] : 
                      (N250)? data_i[1206] : 
                      (N251)? data_i[1238] : 
                      (N252)? data_i[1270] : 
                      (N253)? data_i[1302] : 
                      (N254)? data_i[1334] : 
                      (N255)? data_i[1366] : 
                      (N256)? data_i[1398] : 
                      (N257)? data_i[1430] : 
                      (N258)? data_i[1462] : 
                      (N259)? data_i[1494] : 
                      (N260)? data_i[1526] : 
                      (N261)? data_i[1558] : 
                      (N262)? data_i[1590] : 1'b0;
  assign data_o[21] = (N213)? data_i[21] : 
                      (N214)? data_i[53] : 
                      (N215)? data_i[85] : 
                      (N216)? data_i[117] : 
                      (N217)? data_i[149] : 
                      (N218)? data_i[181] : 
                      (N219)? data_i[213] : 
                      (N220)? data_i[245] : 
                      (N221)? data_i[277] : 
                      (N222)? data_i[309] : 
                      (N223)? data_i[341] : 
                      (N224)? data_i[373] : 
                      (N225)? data_i[405] : 
                      (N226)? data_i[437] : 
                      (N227)? data_i[469] : 
                      (N228)? data_i[501] : 
                      (N229)? data_i[533] : 
                      (N230)? data_i[565] : 
                      (N231)? data_i[597] : 
                      (N232)? data_i[629] : 
                      (N233)? data_i[661] : 
                      (N234)? data_i[693] : 
                      (N235)? data_i[725] : 
                      (N236)? data_i[757] : 
                      (N237)? data_i[789] : 
                      (N238)? data_i[821] : 
                      (N239)? data_i[853] : 
                      (N240)? data_i[885] : 
                      (N241)? data_i[917] : 
                      (N242)? data_i[949] : 
                      (N243)? data_i[981] : 
                      (N244)? data_i[1013] : 
                      (N245)? data_i[1045] : 
                      (N246)? data_i[1077] : 
                      (N247)? data_i[1109] : 
                      (N248)? data_i[1141] : 
                      (N249)? data_i[1173] : 
                      (N250)? data_i[1205] : 
                      (N251)? data_i[1237] : 
                      (N252)? data_i[1269] : 
                      (N253)? data_i[1301] : 
                      (N254)? data_i[1333] : 
                      (N255)? data_i[1365] : 
                      (N256)? data_i[1397] : 
                      (N257)? data_i[1429] : 
                      (N258)? data_i[1461] : 
                      (N259)? data_i[1493] : 
                      (N260)? data_i[1525] : 
                      (N261)? data_i[1557] : 
                      (N262)? data_i[1589] : 1'b0;
  assign data_o[20] = (N213)? data_i[20] : 
                      (N214)? data_i[52] : 
                      (N215)? data_i[84] : 
                      (N216)? data_i[116] : 
                      (N217)? data_i[148] : 
                      (N218)? data_i[180] : 
                      (N219)? data_i[212] : 
                      (N220)? data_i[244] : 
                      (N221)? data_i[276] : 
                      (N222)? data_i[308] : 
                      (N223)? data_i[340] : 
                      (N224)? data_i[372] : 
                      (N225)? data_i[404] : 
                      (N226)? data_i[436] : 
                      (N227)? data_i[468] : 
                      (N228)? data_i[500] : 
                      (N229)? data_i[532] : 
                      (N230)? data_i[564] : 
                      (N231)? data_i[596] : 
                      (N232)? data_i[628] : 
                      (N233)? data_i[660] : 
                      (N234)? data_i[692] : 
                      (N235)? data_i[724] : 
                      (N236)? data_i[756] : 
                      (N237)? data_i[788] : 
                      (N238)? data_i[820] : 
                      (N239)? data_i[852] : 
                      (N240)? data_i[884] : 
                      (N241)? data_i[916] : 
                      (N242)? data_i[948] : 
                      (N243)? data_i[980] : 
                      (N244)? data_i[1012] : 
                      (N245)? data_i[1044] : 
                      (N246)? data_i[1076] : 
                      (N247)? data_i[1108] : 
                      (N248)? data_i[1140] : 
                      (N249)? data_i[1172] : 
                      (N250)? data_i[1204] : 
                      (N251)? data_i[1236] : 
                      (N252)? data_i[1268] : 
                      (N253)? data_i[1300] : 
                      (N254)? data_i[1332] : 
                      (N255)? data_i[1364] : 
                      (N256)? data_i[1396] : 
                      (N257)? data_i[1428] : 
                      (N258)? data_i[1460] : 
                      (N259)? data_i[1492] : 
                      (N260)? data_i[1524] : 
                      (N261)? data_i[1556] : 
                      (N262)? data_i[1588] : 1'b0;
  assign data_o[19] = (N213)? data_i[19] : 
                      (N214)? data_i[51] : 
                      (N215)? data_i[83] : 
                      (N216)? data_i[115] : 
                      (N217)? data_i[147] : 
                      (N218)? data_i[179] : 
                      (N219)? data_i[211] : 
                      (N220)? data_i[243] : 
                      (N221)? data_i[275] : 
                      (N222)? data_i[307] : 
                      (N223)? data_i[339] : 
                      (N224)? data_i[371] : 
                      (N225)? data_i[403] : 
                      (N226)? data_i[435] : 
                      (N227)? data_i[467] : 
                      (N228)? data_i[499] : 
                      (N229)? data_i[531] : 
                      (N230)? data_i[563] : 
                      (N231)? data_i[595] : 
                      (N232)? data_i[627] : 
                      (N233)? data_i[659] : 
                      (N234)? data_i[691] : 
                      (N235)? data_i[723] : 
                      (N236)? data_i[755] : 
                      (N237)? data_i[787] : 
                      (N238)? data_i[819] : 
                      (N239)? data_i[851] : 
                      (N240)? data_i[883] : 
                      (N241)? data_i[915] : 
                      (N242)? data_i[947] : 
                      (N243)? data_i[979] : 
                      (N244)? data_i[1011] : 
                      (N245)? data_i[1043] : 
                      (N246)? data_i[1075] : 
                      (N247)? data_i[1107] : 
                      (N248)? data_i[1139] : 
                      (N249)? data_i[1171] : 
                      (N250)? data_i[1203] : 
                      (N251)? data_i[1235] : 
                      (N252)? data_i[1267] : 
                      (N253)? data_i[1299] : 
                      (N254)? data_i[1331] : 
                      (N255)? data_i[1363] : 
                      (N256)? data_i[1395] : 
                      (N257)? data_i[1427] : 
                      (N258)? data_i[1459] : 
                      (N259)? data_i[1491] : 
                      (N260)? data_i[1523] : 
                      (N261)? data_i[1555] : 
                      (N262)? data_i[1587] : 1'b0;
  assign data_o[18] = (N213)? data_i[18] : 
                      (N214)? data_i[50] : 
                      (N215)? data_i[82] : 
                      (N216)? data_i[114] : 
                      (N217)? data_i[146] : 
                      (N218)? data_i[178] : 
                      (N219)? data_i[210] : 
                      (N220)? data_i[242] : 
                      (N221)? data_i[274] : 
                      (N222)? data_i[306] : 
                      (N223)? data_i[338] : 
                      (N224)? data_i[370] : 
                      (N225)? data_i[402] : 
                      (N226)? data_i[434] : 
                      (N227)? data_i[466] : 
                      (N228)? data_i[498] : 
                      (N229)? data_i[530] : 
                      (N230)? data_i[562] : 
                      (N231)? data_i[594] : 
                      (N232)? data_i[626] : 
                      (N233)? data_i[658] : 
                      (N234)? data_i[690] : 
                      (N235)? data_i[722] : 
                      (N236)? data_i[754] : 
                      (N237)? data_i[786] : 
                      (N238)? data_i[818] : 
                      (N239)? data_i[850] : 
                      (N240)? data_i[882] : 
                      (N241)? data_i[914] : 
                      (N242)? data_i[946] : 
                      (N243)? data_i[978] : 
                      (N244)? data_i[1010] : 
                      (N245)? data_i[1042] : 
                      (N246)? data_i[1074] : 
                      (N247)? data_i[1106] : 
                      (N248)? data_i[1138] : 
                      (N249)? data_i[1170] : 
                      (N250)? data_i[1202] : 
                      (N251)? data_i[1234] : 
                      (N252)? data_i[1266] : 
                      (N253)? data_i[1298] : 
                      (N254)? data_i[1330] : 
                      (N255)? data_i[1362] : 
                      (N256)? data_i[1394] : 
                      (N257)? data_i[1426] : 
                      (N258)? data_i[1458] : 
                      (N259)? data_i[1490] : 
                      (N260)? data_i[1522] : 
                      (N261)? data_i[1554] : 
                      (N262)? data_i[1586] : 1'b0;
  assign data_o[17] = (N213)? data_i[17] : 
                      (N214)? data_i[49] : 
                      (N215)? data_i[81] : 
                      (N216)? data_i[113] : 
                      (N217)? data_i[145] : 
                      (N218)? data_i[177] : 
                      (N219)? data_i[209] : 
                      (N220)? data_i[241] : 
                      (N221)? data_i[273] : 
                      (N222)? data_i[305] : 
                      (N223)? data_i[337] : 
                      (N224)? data_i[369] : 
                      (N225)? data_i[401] : 
                      (N226)? data_i[433] : 
                      (N227)? data_i[465] : 
                      (N228)? data_i[497] : 
                      (N229)? data_i[529] : 
                      (N230)? data_i[561] : 
                      (N231)? data_i[593] : 
                      (N232)? data_i[625] : 
                      (N233)? data_i[657] : 
                      (N234)? data_i[689] : 
                      (N235)? data_i[721] : 
                      (N236)? data_i[753] : 
                      (N237)? data_i[785] : 
                      (N238)? data_i[817] : 
                      (N239)? data_i[849] : 
                      (N240)? data_i[881] : 
                      (N241)? data_i[913] : 
                      (N242)? data_i[945] : 
                      (N243)? data_i[977] : 
                      (N244)? data_i[1009] : 
                      (N245)? data_i[1041] : 
                      (N246)? data_i[1073] : 
                      (N247)? data_i[1105] : 
                      (N248)? data_i[1137] : 
                      (N249)? data_i[1169] : 
                      (N250)? data_i[1201] : 
                      (N251)? data_i[1233] : 
                      (N252)? data_i[1265] : 
                      (N253)? data_i[1297] : 
                      (N254)? data_i[1329] : 
                      (N255)? data_i[1361] : 
                      (N256)? data_i[1393] : 
                      (N257)? data_i[1425] : 
                      (N258)? data_i[1457] : 
                      (N259)? data_i[1489] : 
                      (N260)? data_i[1521] : 
                      (N261)? data_i[1553] : 
                      (N262)? data_i[1585] : 1'b0;
  assign data_o[16] = (N213)? data_i[16] : 
                      (N214)? data_i[48] : 
                      (N215)? data_i[80] : 
                      (N216)? data_i[112] : 
                      (N217)? data_i[144] : 
                      (N218)? data_i[176] : 
                      (N219)? data_i[208] : 
                      (N220)? data_i[240] : 
                      (N221)? data_i[272] : 
                      (N222)? data_i[304] : 
                      (N223)? data_i[336] : 
                      (N224)? data_i[368] : 
                      (N225)? data_i[400] : 
                      (N226)? data_i[432] : 
                      (N227)? data_i[464] : 
                      (N228)? data_i[496] : 
                      (N229)? data_i[528] : 
                      (N230)? data_i[560] : 
                      (N231)? data_i[592] : 
                      (N232)? data_i[624] : 
                      (N233)? data_i[656] : 
                      (N234)? data_i[688] : 
                      (N235)? data_i[720] : 
                      (N236)? data_i[752] : 
                      (N237)? data_i[784] : 
                      (N238)? data_i[816] : 
                      (N239)? data_i[848] : 
                      (N240)? data_i[880] : 
                      (N241)? data_i[912] : 
                      (N242)? data_i[944] : 
                      (N243)? data_i[976] : 
                      (N244)? data_i[1008] : 
                      (N245)? data_i[1040] : 
                      (N246)? data_i[1072] : 
                      (N247)? data_i[1104] : 
                      (N248)? data_i[1136] : 
                      (N249)? data_i[1168] : 
                      (N250)? data_i[1200] : 
                      (N251)? data_i[1232] : 
                      (N252)? data_i[1264] : 
                      (N253)? data_i[1296] : 
                      (N254)? data_i[1328] : 
                      (N255)? data_i[1360] : 
                      (N256)? data_i[1392] : 
                      (N257)? data_i[1424] : 
                      (N258)? data_i[1456] : 
                      (N259)? data_i[1488] : 
                      (N260)? data_i[1520] : 
                      (N261)? data_i[1552] : 
                      (N262)? data_i[1584] : 1'b0;
  assign data_o[15] = (N213)? data_i[15] : 
                      (N214)? data_i[47] : 
                      (N215)? data_i[79] : 
                      (N216)? data_i[111] : 
                      (N217)? data_i[143] : 
                      (N218)? data_i[175] : 
                      (N219)? data_i[207] : 
                      (N220)? data_i[239] : 
                      (N221)? data_i[271] : 
                      (N222)? data_i[303] : 
                      (N223)? data_i[335] : 
                      (N224)? data_i[367] : 
                      (N225)? data_i[399] : 
                      (N226)? data_i[431] : 
                      (N227)? data_i[463] : 
                      (N228)? data_i[495] : 
                      (N229)? data_i[527] : 
                      (N230)? data_i[559] : 
                      (N231)? data_i[591] : 
                      (N232)? data_i[623] : 
                      (N233)? data_i[655] : 
                      (N234)? data_i[687] : 
                      (N235)? data_i[719] : 
                      (N236)? data_i[751] : 
                      (N237)? data_i[783] : 
                      (N238)? data_i[815] : 
                      (N239)? data_i[847] : 
                      (N240)? data_i[879] : 
                      (N241)? data_i[911] : 
                      (N242)? data_i[943] : 
                      (N243)? data_i[975] : 
                      (N244)? data_i[1007] : 
                      (N245)? data_i[1039] : 
                      (N246)? data_i[1071] : 
                      (N247)? data_i[1103] : 
                      (N248)? data_i[1135] : 
                      (N249)? data_i[1167] : 
                      (N250)? data_i[1199] : 
                      (N251)? data_i[1231] : 
                      (N252)? data_i[1263] : 
                      (N253)? data_i[1295] : 
                      (N254)? data_i[1327] : 
                      (N255)? data_i[1359] : 
                      (N256)? data_i[1391] : 
                      (N257)? data_i[1423] : 
                      (N258)? data_i[1455] : 
                      (N259)? data_i[1487] : 
                      (N260)? data_i[1519] : 
                      (N261)? data_i[1551] : 
                      (N262)? data_i[1583] : 1'b0;
  assign data_o[14] = (N213)? data_i[14] : 
                      (N214)? data_i[46] : 
                      (N215)? data_i[78] : 
                      (N216)? data_i[110] : 
                      (N217)? data_i[142] : 
                      (N218)? data_i[174] : 
                      (N219)? data_i[206] : 
                      (N220)? data_i[238] : 
                      (N221)? data_i[270] : 
                      (N222)? data_i[302] : 
                      (N223)? data_i[334] : 
                      (N224)? data_i[366] : 
                      (N225)? data_i[398] : 
                      (N226)? data_i[430] : 
                      (N227)? data_i[462] : 
                      (N228)? data_i[494] : 
                      (N229)? data_i[526] : 
                      (N230)? data_i[558] : 
                      (N231)? data_i[590] : 
                      (N232)? data_i[622] : 
                      (N233)? data_i[654] : 
                      (N234)? data_i[686] : 
                      (N235)? data_i[718] : 
                      (N236)? data_i[750] : 
                      (N237)? data_i[782] : 
                      (N238)? data_i[814] : 
                      (N239)? data_i[846] : 
                      (N240)? data_i[878] : 
                      (N241)? data_i[910] : 
                      (N242)? data_i[942] : 
                      (N243)? data_i[974] : 
                      (N244)? data_i[1006] : 
                      (N245)? data_i[1038] : 
                      (N246)? data_i[1070] : 
                      (N247)? data_i[1102] : 
                      (N248)? data_i[1134] : 
                      (N249)? data_i[1166] : 
                      (N250)? data_i[1198] : 
                      (N251)? data_i[1230] : 
                      (N252)? data_i[1262] : 
                      (N253)? data_i[1294] : 
                      (N254)? data_i[1326] : 
                      (N255)? data_i[1358] : 
                      (N256)? data_i[1390] : 
                      (N257)? data_i[1422] : 
                      (N258)? data_i[1454] : 
                      (N259)? data_i[1486] : 
                      (N260)? data_i[1518] : 
                      (N261)? data_i[1550] : 
                      (N262)? data_i[1582] : 1'b0;
  assign data_o[13] = (N213)? data_i[13] : 
                      (N214)? data_i[45] : 
                      (N215)? data_i[77] : 
                      (N216)? data_i[109] : 
                      (N217)? data_i[141] : 
                      (N218)? data_i[173] : 
                      (N219)? data_i[205] : 
                      (N220)? data_i[237] : 
                      (N221)? data_i[269] : 
                      (N222)? data_i[301] : 
                      (N223)? data_i[333] : 
                      (N224)? data_i[365] : 
                      (N225)? data_i[397] : 
                      (N226)? data_i[429] : 
                      (N227)? data_i[461] : 
                      (N228)? data_i[493] : 
                      (N229)? data_i[525] : 
                      (N230)? data_i[557] : 
                      (N231)? data_i[589] : 
                      (N232)? data_i[621] : 
                      (N233)? data_i[653] : 
                      (N234)? data_i[685] : 
                      (N235)? data_i[717] : 
                      (N236)? data_i[749] : 
                      (N237)? data_i[781] : 
                      (N238)? data_i[813] : 
                      (N239)? data_i[845] : 
                      (N240)? data_i[877] : 
                      (N241)? data_i[909] : 
                      (N242)? data_i[941] : 
                      (N243)? data_i[973] : 
                      (N244)? data_i[1005] : 
                      (N245)? data_i[1037] : 
                      (N246)? data_i[1069] : 
                      (N247)? data_i[1101] : 
                      (N248)? data_i[1133] : 
                      (N249)? data_i[1165] : 
                      (N250)? data_i[1197] : 
                      (N251)? data_i[1229] : 
                      (N252)? data_i[1261] : 
                      (N253)? data_i[1293] : 
                      (N254)? data_i[1325] : 
                      (N255)? data_i[1357] : 
                      (N256)? data_i[1389] : 
                      (N257)? data_i[1421] : 
                      (N258)? data_i[1453] : 
                      (N259)? data_i[1485] : 
                      (N260)? data_i[1517] : 
                      (N261)? data_i[1549] : 
                      (N262)? data_i[1581] : 1'b0;
  assign data_o[12] = (N213)? data_i[12] : 
                      (N214)? data_i[44] : 
                      (N215)? data_i[76] : 
                      (N216)? data_i[108] : 
                      (N217)? data_i[140] : 
                      (N218)? data_i[172] : 
                      (N219)? data_i[204] : 
                      (N220)? data_i[236] : 
                      (N221)? data_i[268] : 
                      (N222)? data_i[300] : 
                      (N223)? data_i[332] : 
                      (N224)? data_i[364] : 
                      (N225)? data_i[396] : 
                      (N226)? data_i[428] : 
                      (N227)? data_i[460] : 
                      (N228)? data_i[492] : 
                      (N229)? data_i[524] : 
                      (N230)? data_i[556] : 
                      (N231)? data_i[588] : 
                      (N232)? data_i[620] : 
                      (N233)? data_i[652] : 
                      (N234)? data_i[684] : 
                      (N235)? data_i[716] : 
                      (N236)? data_i[748] : 
                      (N237)? data_i[780] : 
                      (N238)? data_i[812] : 
                      (N239)? data_i[844] : 
                      (N240)? data_i[876] : 
                      (N241)? data_i[908] : 
                      (N242)? data_i[940] : 
                      (N243)? data_i[972] : 
                      (N244)? data_i[1004] : 
                      (N245)? data_i[1036] : 
                      (N246)? data_i[1068] : 
                      (N247)? data_i[1100] : 
                      (N248)? data_i[1132] : 
                      (N249)? data_i[1164] : 
                      (N250)? data_i[1196] : 
                      (N251)? data_i[1228] : 
                      (N252)? data_i[1260] : 
                      (N253)? data_i[1292] : 
                      (N254)? data_i[1324] : 
                      (N255)? data_i[1356] : 
                      (N256)? data_i[1388] : 
                      (N257)? data_i[1420] : 
                      (N258)? data_i[1452] : 
                      (N259)? data_i[1484] : 
                      (N260)? data_i[1516] : 
                      (N261)? data_i[1548] : 
                      (N262)? data_i[1580] : 1'b0;
  assign data_o[11] = (N213)? data_i[11] : 
                      (N214)? data_i[43] : 
                      (N215)? data_i[75] : 
                      (N216)? data_i[107] : 
                      (N217)? data_i[139] : 
                      (N218)? data_i[171] : 
                      (N219)? data_i[203] : 
                      (N220)? data_i[235] : 
                      (N221)? data_i[267] : 
                      (N222)? data_i[299] : 
                      (N223)? data_i[331] : 
                      (N224)? data_i[363] : 
                      (N225)? data_i[395] : 
                      (N226)? data_i[427] : 
                      (N227)? data_i[459] : 
                      (N228)? data_i[491] : 
                      (N229)? data_i[523] : 
                      (N230)? data_i[555] : 
                      (N231)? data_i[587] : 
                      (N232)? data_i[619] : 
                      (N233)? data_i[651] : 
                      (N234)? data_i[683] : 
                      (N235)? data_i[715] : 
                      (N236)? data_i[747] : 
                      (N237)? data_i[779] : 
                      (N238)? data_i[811] : 
                      (N239)? data_i[843] : 
                      (N240)? data_i[875] : 
                      (N241)? data_i[907] : 
                      (N242)? data_i[939] : 
                      (N243)? data_i[971] : 
                      (N244)? data_i[1003] : 
                      (N245)? data_i[1035] : 
                      (N246)? data_i[1067] : 
                      (N247)? data_i[1099] : 
                      (N248)? data_i[1131] : 
                      (N249)? data_i[1163] : 
                      (N250)? data_i[1195] : 
                      (N251)? data_i[1227] : 
                      (N252)? data_i[1259] : 
                      (N253)? data_i[1291] : 
                      (N254)? data_i[1323] : 
                      (N255)? data_i[1355] : 
                      (N256)? data_i[1387] : 
                      (N257)? data_i[1419] : 
                      (N258)? data_i[1451] : 
                      (N259)? data_i[1483] : 
                      (N260)? data_i[1515] : 
                      (N261)? data_i[1547] : 
                      (N262)? data_i[1579] : 1'b0;
  assign data_o[10] = (N213)? data_i[10] : 
                      (N214)? data_i[42] : 
                      (N215)? data_i[74] : 
                      (N216)? data_i[106] : 
                      (N217)? data_i[138] : 
                      (N218)? data_i[170] : 
                      (N219)? data_i[202] : 
                      (N220)? data_i[234] : 
                      (N221)? data_i[266] : 
                      (N222)? data_i[298] : 
                      (N223)? data_i[330] : 
                      (N224)? data_i[362] : 
                      (N225)? data_i[394] : 
                      (N226)? data_i[426] : 
                      (N227)? data_i[458] : 
                      (N228)? data_i[490] : 
                      (N229)? data_i[522] : 
                      (N230)? data_i[554] : 
                      (N231)? data_i[586] : 
                      (N232)? data_i[618] : 
                      (N233)? data_i[650] : 
                      (N234)? data_i[682] : 
                      (N235)? data_i[714] : 
                      (N236)? data_i[746] : 
                      (N237)? data_i[778] : 
                      (N238)? data_i[810] : 
                      (N239)? data_i[842] : 
                      (N240)? data_i[874] : 
                      (N241)? data_i[906] : 
                      (N242)? data_i[938] : 
                      (N243)? data_i[970] : 
                      (N244)? data_i[1002] : 
                      (N245)? data_i[1034] : 
                      (N246)? data_i[1066] : 
                      (N247)? data_i[1098] : 
                      (N248)? data_i[1130] : 
                      (N249)? data_i[1162] : 
                      (N250)? data_i[1194] : 
                      (N251)? data_i[1226] : 
                      (N252)? data_i[1258] : 
                      (N253)? data_i[1290] : 
                      (N254)? data_i[1322] : 
                      (N255)? data_i[1354] : 
                      (N256)? data_i[1386] : 
                      (N257)? data_i[1418] : 
                      (N258)? data_i[1450] : 
                      (N259)? data_i[1482] : 
                      (N260)? data_i[1514] : 
                      (N261)? data_i[1546] : 
                      (N262)? data_i[1578] : 1'b0;
  assign data_o[9] = (N213)? data_i[9] : 
                     (N214)? data_i[41] : 
                     (N215)? data_i[73] : 
                     (N216)? data_i[105] : 
                     (N217)? data_i[137] : 
                     (N218)? data_i[169] : 
                     (N219)? data_i[201] : 
                     (N220)? data_i[233] : 
                     (N221)? data_i[265] : 
                     (N222)? data_i[297] : 
                     (N223)? data_i[329] : 
                     (N224)? data_i[361] : 
                     (N225)? data_i[393] : 
                     (N226)? data_i[425] : 
                     (N227)? data_i[457] : 
                     (N228)? data_i[489] : 
                     (N229)? data_i[521] : 
                     (N230)? data_i[553] : 
                     (N231)? data_i[585] : 
                     (N232)? data_i[617] : 
                     (N233)? data_i[649] : 
                     (N234)? data_i[681] : 
                     (N235)? data_i[713] : 
                     (N236)? data_i[745] : 
                     (N237)? data_i[777] : 
                     (N238)? data_i[809] : 
                     (N239)? data_i[841] : 
                     (N240)? data_i[873] : 
                     (N241)? data_i[905] : 
                     (N242)? data_i[937] : 
                     (N243)? data_i[969] : 
                     (N244)? data_i[1001] : 
                     (N245)? data_i[1033] : 
                     (N246)? data_i[1065] : 
                     (N247)? data_i[1097] : 
                     (N248)? data_i[1129] : 
                     (N249)? data_i[1161] : 
                     (N250)? data_i[1193] : 
                     (N251)? data_i[1225] : 
                     (N252)? data_i[1257] : 
                     (N253)? data_i[1289] : 
                     (N254)? data_i[1321] : 
                     (N255)? data_i[1353] : 
                     (N256)? data_i[1385] : 
                     (N257)? data_i[1417] : 
                     (N258)? data_i[1449] : 
                     (N259)? data_i[1481] : 
                     (N260)? data_i[1513] : 
                     (N261)? data_i[1545] : 
                     (N262)? data_i[1577] : 1'b0;
  assign data_o[8] = (N213)? data_i[8] : 
                     (N214)? data_i[40] : 
                     (N215)? data_i[72] : 
                     (N216)? data_i[104] : 
                     (N217)? data_i[136] : 
                     (N218)? data_i[168] : 
                     (N219)? data_i[200] : 
                     (N220)? data_i[232] : 
                     (N221)? data_i[264] : 
                     (N222)? data_i[296] : 
                     (N223)? data_i[328] : 
                     (N224)? data_i[360] : 
                     (N225)? data_i[392] : 
                     (N226)? data_i[424] : 
                     (N227)? data_i[456] : 
                     (N228)? data_i[488] : 
                     (N229)? data_i[520] : 
                     (N230)? data_i[552] : 
                     (N231)? data_i[584] : 
                     (N232)? data_i[616] : 
                     (N233)? data_i[648] : 
                     (N234)? data_i[680] : 
                     (N235)? data_i[712] : 
                     (N236)? data_i[744] : 
                     (N237)? data_i[776] : 
                     (N238)? data_i[808] : 
                     (N239)? data_i[840] : 
                     (N240)? data_i[872] : 
                     (N241)? data_i[904] : 
                     (N242)? data_i[936] : 
                     (N243)? data_i[968] : 
                     (N244)? data_i[1000] : 
                     (N245)? data_i[1032] : 
                     (N246)? data_i[1064] : 
                     (N247)? data_i[1096] : 
                     (N248)? data_i[1128] : 
                     (N249)? data_i[1160] : 
                     (N250)? data_i[1192] : 
                     (N251)? data_i[1224] : 
                     (N252)? data_i[1256] : 
                     (N253)? data_i[1288] : 
                     (N254)? data_i[1320] : 
                     (N255)? data_i[1352] : 
                     (N256)? data_i[1384] : 
                     (N257)? data_i[1416] : 
                     (N258)? data_i[1448] : 
                     (N259)? data_i[1480] : 
                     (N260)? data_i[1512] : 
                     (N261)? data_i[1544] : 
                     (N262)? data_i[1576] : 1'b0;
  assign data_o[7] = (N213)? data_i[7] : 
                     (N214)? data_i[39] : 
                     (N215)? data_i[71] : 
                     (N216)? data_i[103] : 
                     (N217)? data_i[135] : 
                     (N218)? data_i[167] : 
                     (N219)? data_i[199] : 
                     (N220)? data_i[231] : 
                     (N221)? data_i[263] : 
                     (N222)? data_i[295] : 
                     (N223)? data_i[327] : 
                     (N224)? data_i[359] : 
                     (N225)? data_i[391] : 
                     (N226)? data_i[423] : 
                     (N227)? data_i[455] : 
                     (N228)? data_i[487] : 
                     (N229)? data_i[519] : 
                     (N230)? data_i[551] : 
                     (N231)? data_i[583] : 
                     (N232)? data_i[615] : 
                     (N233)? data_i[647] : 
                     (N234)? data_i[679] : 
                     (N235)? data_i[711] : 
                     (N236)? data_i[743] : 
                     (N237)? data_i[775] : 
                     (N238)? data_i[807] : 
                     (N239)? data_i[839] : 
                     (N240)? data_i[871] : 
                     (N241)? data_i[903] : 
                     (N242)? data_i[935] : 
                     (N243)? data_i[967] : 
                     (N244)? data_i[999] : 
                     (N245)? data_i[1031] : 
                     (N246)? data_i[1063] : 
                     (N247)? data_i[1095] : 
                     (N248)? data_i[1127] : 
                     (N249)? data_i[1159] : 
                     (N250)? data_i[1191] : 
                     (N251)? data_i[1223] : 
                     (N252)? data_i[1255] : 
                     (N253)? data_i[1287] : 
                     (N254)? data_i[1319] : 
                     (N255)? data_i[1351] : 
                     (N256)? data_i[1383] : 
                     (N257)? data_i[1415] : 
                     (N258)? data_i[1447] : 
                     (N259)? data_i[1479] : 
                     (N260)? data_i[1511] : 
                     (N261)? data_i[1543] : 
                     (N262)? data_i[1575] : 1'b0;
  assign data_o[6] = (N213)? data_i[6] : 
                     (N214)? data_i[38] : 
                     (N215)? data_i[70] : 
                     (N216)? data_i[102] : 
                     (N217)? data_i[134] : 
                     (N218)? data_i[166] : 
                     (N219)? data_i[198] : 
                     (N220)? data_i[230] : 
                     (N221)? data_i[262] : 
                     (N222)? data_i[294] : 
                     (N223)? data_i[326] : 
                     (N224)? data_i[358] : 
                     (N225)? data_i[390] : 
                     (N226)? data_i[422] : 
                     (N227)? data_i[454] : 
                     (N228)? data_i[486] : 
                     (N229)? data_i[518] : 
                     (N230)? data_i[550] : 
                     (N231)? data_i[582] : 
                     (N232)? data_i[614] : 
                     (N233)? data_i[646] : 
                     (N234)? data_i[678] : 
                     (N235)? data_i[710] : 
                     (N236)? data_i[742] : 
                     (N237)? data_i[774] : 
                     (N238)? data_i[806] : 
                     (N239)? data_i[838] : 
                     (N240)? data_i[870] : 
                     (N241)? data_i[902] : 
                     (N242)? data_i[934] : 
                     (N243)? data_i[966] : 
                     (N244)? data_i[998] : 
                     (N245)? data_i[1030] : 
                     (N246)? data_i[1062] : 
                     (N247)? data_i[1094] : 
                     (N248)? data_i[1126] : 
                     (N249)? data_i[1158] : 
                     (N250)? data_i[1190] : 
                     (N251)? data_i[1222] : 
                     (N252)? data_i[1254] : 
                     (N253)? data_i[1286] : 
                     (N254)? data_i[1318] : 
                     (N255)? data_i[1350] : 
                     (N256)? data_i[1382] : 
                     (N257)? data_i[1414] : 
                     (N258)? data_i[1446] : 
                     (N259)? data_i[1478] : 
                     (N260)? data_i[1510] : 
                     (N261)? data_i[1542] : 
                     (N262)? data_i[1574] : 1'b0;
  assign data_o[5] = (N213)? data_i[5] : 
                     (N214)? data_i[37] : 
                     (N215)? data_i[69] : 
                     (N216)? data_i[101] : 
                     (N217)? data_i[133] : 
                     (N218)? data_i[165] : 
                     (N219)? data_i[197] : 
                     (N220)? data_i[229] : 
                     (N221)? data_i[261] : 
                     (N222)? data_i[293] : 
                     (N223)? data_i[325] : 
                     (N224)? data_i[357] : 
                     (N225)? data_i[389] : 
                     (N226)? data_i[421] : 
                     (N227)? data_i[453] : 
                     (N228)? data_i[485] : 
                     (N229)? data_i[517] : 
                     (N230)? data_i[549] : 
                     (N231)? data_i[581] : 
                     (N232)? data_i[613] : 
                     (N233)? data_i[645] : 
                     (N234)? data_i[677] : 
                     (N235)? data_i[709] : 
                     (N236)? data_i[741] : 
                     (N237)? data_i[773] : 
                     (N238)? data_i[805] : 
                     (N239)? data_i[837] : 
                     (N240)? data_i[869] : 
                     (N241)? data_i[901] : 
                     (N242)? data_i[933] : 
                     (N243)? data_i[965] : 
                     (N244)? data_i[997] : 
                     (N245)? data_i[1029] : 
                     (N246)? data_i[1061] : 
                     (N247)? data_i[1093] : 
                     (N248)? data_i[1125] : 
                     (N249)? data_i[1157] : 
                     (N250)? data_i[1189] : 
                     (N251)? data_i[1221] : 
                     (N252)? data_i[1253] : 
                     (N253)? data_i[1285] : 
                     (N254)? data_i[1317] : 
                     (N255)? data_i[1349] : 
                     (N256)? data_i[1381] : 
                     (N257)? data_i[1413] : 
                     (N258)? data_i[1445] : 
                     (N259)? data_i[1477] : 
                     (N260)? data_i[1509] : 
                     (N261)? data_i[1541] : 
                     (N262)? data_i[1573] : 1'b0;
  assign data_o[4] = (N213)? data_i[4] : 
                     (N214)? data_i[36] : 
                     (N215)? data_i[68] : 
                     (N216)? data_i[100] : 
                     (N217)? data_i[132] : 
                     (N218)? data_i[164] : 
                     (N219)? data_i[196] : 
                     (N220)? data_i[228] : 
                     (N221)? data_i[260] : 
                     (N222)? data_i[292] : 
                     (N223)? data_i[324] : 
                     (N224)? data_i[356] : 
                     (N225)? data_i[388] : 
                     (N226)? data_i[420] : 
                     (N227)? data_i[452] : 
                     (N228)? data_i[484] : 
                     (N229)? data_i[516] : 
                     (N230)? data_i[548] : 
                     (N231)? data_i[580] : 
                     (N232)? data_i[612] : 
                     (N233)? data_i[644] : 
                     (N234)? data_i[676] : 
                     (N235)? data_i[708] : 
                     (N236)? data_i[740] : 
                     (N237)? data_i[772] : 
                     (N238)? data_i[804] : 
                     (N239)? data_i[836] : 
                     (N240)? data_i[868] : 
                     (N241)? data_i[900] : 
                     (N242)? data_i[932] : 
                     (N243)? data_i[964] : 
                     (N244)? data_i[996] : 
                     (N245)? data_i[1028] : 
                     (N246)? data_i[1060] : 
                     (N247)? data_i[1092] : 
                     (N248)? data_i[1124] : 
                     (N249)? data_i[1156] : 
                     (N250)? data_i[1188] : 
                     (N251)? data_i[1220] : 
                     (N252)? data_i[1252] : 
                     (N253)? data_i[1284] : 
                     (N254)? data_i[1316] : 
                     (N255)? data_i[1348] : 
                     (N256)? data_i[1380] : 
                     (N257)? data_i[1412] : 
                     (N258)? data_i[1444] : 
                     (N259)? data_i[1476] : 
                     (N260)? data_i[1508] : 
                     (N261)? data_i[1540] : 
                     (N262)? data_i[1572] : 1'b0;
  assign data_o[3] = (N213)? data_i[3] : 
                     (N214)? data_i[35] : 
                     (N215)? data_i[67] : 
                     (N216)? data_i[99] : 
                     (N217)? data_i[131] : 
                     (N218)? data_i[163] : 
                     (N219)? data_i[195] : 
                     (N220)? data_i[227] : 
                     (N221)? data_i[259] : 
                     (N222)? data_i[291] : 
                     (N223)? data_i[323] : 
                     (N224)? data_i[355] : 
                     (N225)? data_i[387] : 
                     (N226)? data_i[419] : 
                     (N227)? data_i[451] : 
                     (N228)? data_i[483] : 
                     (N229)? data_i[515] : 
                     (N230)? data_i[547] : 
                     (N231)? data_i[579] : 
                     (N232)? data_i[611] : 
                     (N233)? data_i[643] : 
                     (N234)? data_i[675] : 
                     (N235)? data_i[707] : 
                     (N236)? data_i[739] : 
                     (N237)? data_i[771] : 
                     (N238)? data_i[803] : 
                     (N239)? data_i[835] : 
                     (N240)? data_i[867] : 
                     (N241)? data_i[899] : 
                     (N242)? data_i[931] : 
                     (N243)? data_i[963] : 
                     (N244)? data_i[995] : 
                     (N245)? data_i[1027] : 
                     (N246)? data_i[1059] : 
                     (N247)? data_i[1091] : 
                     (N248)? data_i[1123] : 
                     (N249)? data_i[1155] : 
                     (N250)? data_i[1187] : 
                     (N251)? data_i[1219] : 
                     (N252)? data_i[1251] : 
                     (N253)? data_i[1283] : 
                     (N254)? data_i[1315] : 
                     (N255)? data_i[1347] : 
                     (N256)? data_i[1379] : 
                     (N257)? data_i[1411] : 
                     (N258)? data_i[1443] : 
                     (N259)? data_i[1475] : 
                     (N260)? data_i[1507] : 
                     (N261)? data_i[1539] : 
                     (N262)? data_i[1571] : 1'b0;
  assign data_o[2] = (N213)? data_i[2] : 
                     (N214)? data_i[34] : 
                     (N215)? data_i[66] : 
                     (N216)? data_i[98] : 
                     (N217)? data_i[130] : 
                     (N218)? data_i[162] : 
                     (N219)? data_i[194] : 
                     (N220)? data_i[226] : 
                     (N221)? data_i[258] : 
                     (N222)? data_i[290] : 
                     (N223)? data_i[322] : 
                     (N224)? data_i[354] : 
                     (N225)? data_i[386] : 
                     (N226)? data_i[418] : 
                     (N227)? data_i[450] : 
                     (N228)? data_i[482] : 
                     (N229)? data_i[514] : 
                     (N230)? data_i[546] : 
                     (N231)? data_i[578] : 
                     (N232)? data_i[610] : 
                     (N233)? data_i[642] : 
                     (N234)? data_i[674] : 
                     (N235)? data_i[706] : 
                     (N236)? data_i[738] : 
                     (N237)? data_i[770] : 
                     (N238)? data_i[802] : 
                     (N239)? data_i[834] : 
                     (N240)? data_i[866] : 
                     (N241)? data_i[898] : 
                     (N242)? data_i[930] : 
                     (N243)? data_i[962] : 
                     (N244)? data_i[994] : 
                     (N245)? data_i[1026] : 
                     (N246)? data_i[1058] : 
                     (N247)? data_i[1090] : 
                     (N248)? data_i[1122] : 
                     (N249)? data_i[1154] : 
                     (N250)? data_i[1186] : 
                     (N251)? data_i[1218] : 
                     (N252)? data_i[1250] : 
                     (N253)? data_i[1282] : 
                     (N254)? data_i[1314] : 
                     (N255)? data_i[1346] : 
                     (N256)? data_i[1378] : 
                     (N257)? data_i[1410] : 
                     (N258)? data_i[1442] : 
                     (N259)? data_i[1474] : 
                     (N260)? data_i[1506] : 
                     (N261)? data_i[1538] : 
                     (N262)? data_i[1570] : 1'b0;
  assign data_o[1] = (N213)? data_i[1] : 
                     (N214)? data_i[33] : 
                     (N215)? data_i[65] : 
                     (N216)? data_i[97] : 
                     (N217)? data_i[129] : 
                     (N218)? data_i[161] : 
                     (N219)? data_i[193] : 
                     (N220)? data_i[225] : 
                     (N221)? data_i[257] : 
                     (N222)? data_i[289] : 
                     (N223)? data_i[321] : 
                     (N224)? data_i[353] : 
                     (N225)? data_i[385] : 
                     (N226)? data_i[417] : 
                     (N227)? data_i[449] : 
                     (N228)? data_i[481] : 
                     (N229)? data_i[513] : 
                     (N230)? data_i[545] : 
                     (N231)? data_i[577] : 
                     (N232)? data_i[609] : 
                     (N233)? data_i[641] : 
                     (N234)? data_i[673] : 
                     (N235)? data_i[705] : 
                     (N236)? data_i[737] : 
                     (N237)? data_i[769] : 
                     (N238)? data_i[801] : 
                     (N239)? data_i[833] : 
                     (N240)? data_i[865] : 
                     (N241)? data_i[897] : 
                     (N242)? data_i[929] : 
                     (N243)? data_i[961] : 
                     (N244)? data_i[993] : 
                     (N245)? data_i[1025] : 
                     (N246)? data_i[1057] : 
                     (N247)? data_i[1089] : 
                     (N248)? data_i[1121] : 
                     (N249)? data_i[1153] : 
                     (N250)? data_i[1185] : 
                     (N251)? data_i[1217] : 
                     (N252)? data_i[1249] : 
                     (N253)? data_i[1281] : 
                     (N254)? data_i[1313] : 
                     (N255)? data_i[1345] : 
                     (N256)? data_i[1377] : 
                     (N257)? data_i[1409] : 
                     (N258)? data_i[1441] : 
                     (N259)? data_i[1473] : 
                     (N260)? data_i[1505] : 
                     (N261)? data_i[1537] : 
                     (N262)? data_i[1569] : 1'b0;
  assign data_o[0] = (N213)? data_i[0] : 
                     (N214)? data_i[32] : 
                     (N215)? data_i[64] : 
                     (N216)? data_i[96] : 
                     (N217)? data_i[128] : 
                     (N218)? data_i[160] : 
                     (N219)? data_i[192] : 
                     (N220)? data_i[224] : 
                     (N221)? data_i[256] : 
                     (N222)? data_i[288] : 
                     (N223)? data_i[320] : 
                     (N224)? data_i[352] : 
                     (N225)? data_i[384] : 
                     (N226)? data_i[416] : 
                     (N227)? data_i[448] : 
                     (N228)? data_i[480] : 
                     (N229)? data_i[512] : 
                     (N230)? data_i[544] : 
                     (N231)? data_i[576] : 
                     (N232)? data_i[608] : 
                     (N233)? data_i[640] : 
                     (N234)? data_i[672] : 
                     (N235)? data_i[704] : 
                     (N236)? data_i[736] : 
                     (N237)? data_i[768] : 
                     (N238)? data_i[800] : 
                     (N239)? data_i[832] : 
                     (N240)? data_i[864] : 
                     (N241)? data_i[896] : 
                     (N242)? data_i[928] : 
                     (N243)? data_i[960] : 
                     (N244)? data_i[992] : 
                     (N245)? data_i[1024] : 
                     (N246)? data_i[1056] : 
                     (N247)? data_i[1088] : 
                     (N248)? data_i[1120] : 
                     (N249)? data_i[1152] : 
                     (N250)? data_i[1184] : 
                     (N251)? data_i[1216] : 
                     (N252)? data_i[1248] : 
                     (N253)? data_i[1280] : 
                     (N254)? data_i[1312] : 
                     (N255)? data_i[1344] : 
                     (N256)? data_i[1376] : 
                     (N257)? data_i[1408] : 
                     (N258)? data_i[1440] : 
                     (N259)? data_i[1472] : 
                     (N260)? data_i[1504] : 
                     (N261)? data_i[1536] : 
                     (N262)? data_i[1568] : 1'b0;

endmodule



module bsg_parallel_in_serial_out_dynamic
(
  clk_i,
  reset_i,
  v_i,
  len_i,
  data_i,
  ready_o,
  v_o,
  len_v_o,
  data_o,
  yumi_i
);

  input [5:0] len_i;
  input [1599:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output len_v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,len_v_o,count_r_is_last,up_li,clear_li,N0,N1,N2,N3,N4,N6;
  wire [5:0] len_lo,count_lo;
  wire [1599:0] fifo_data_lo;

  bsg_two_fifo_width_p6
  go_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(len_i),
    .v_i(v_i),
    .v_o(v_o),
    .data_o(len_lo),
    .yumi_i(clear_li)
  );


  bsg_two_fifo_width_p1600
  data_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(v_i),
    .data_o(fifo_data_lo),
    .yumi_i(clear_li)
  );

  assign count_r_is_last = count_lo == len_lo;

  bsg_counter_clear_up_max_val_p49_init_val_p0
  ctr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(clear_li),
    .up_i(up_li),
    .count_o(count_lo)
  );


  bsg_mux_width_p32_els_p50
  data_mux
  (
    .data_i(fifo_data_lo),
    .sel_i(count_lo),
    .data_o(data_o)
  );

  assign N0 = count_lo[4] | count_lo[5];
  assign N1 = count_lo[3] | N0;
  assign N2 = count_lo[2] | N1;
  assign N3 = count_lo[1] | N2;
  assign N4 = count_lo[0] | N3;
  assign len_v_o = ~N4;
  assign up_li = yumi_i & N6;
  assign N6 = ~count_r_is_last;
  assign clear_li = yumi_i & count_r_is_last;

endmodule

