

module top
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  yumi_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [69:0] cache_pkt_i;
  output [31:0] data_o;
  output [32:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output yumi_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;

  bsg_cache
  wrapper
  (
    .cache_pkt_i(cache_pkt_i),
    .data_o(data_o),
    .dma_pkt_o(dma_pkt_o),
    .dma_data_i(dma_data_i),
    .dma_data_o(dma_data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_yumi_i(dma_data_yumi_i),
    .yumi_o(yumi_o),
    .v_o(v_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_v_o(dma_data_v_o),
    .v_we_o(v_we_o)
  );


endmodule



module bsg_cache_decode
(
  opcode_i,
  decode_o
);

  input [5:0] opcode_i;
  output [20:0] decode_o;
  wire [20:0] decode_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N146,N147,N148,N150,N152,
  N153,N154,N155,N156,N158,N160,N161,N163,N165,N166,N167,N168,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297;
  assign N17 = N80 | N138;
  assign N18 = opcode_i[3] | opcode_i[2];
  assign N19 = opcode_i[1] | opcode_i[0];
  assign N20 = N17 | N18;
  assign N21 = N20 | N19;
  assign N22 = opcode_i[1] | N139;
  assign N23 = N20 | N22;
  assign N24 = N146 | N139;
  assign N25 = N20 | N24;
  assign N26 = opcode_i[3] | N165;
  assign N27 = N17 | N26;
  assign N28 = N27 | N19;
  assign N29 = N146 | opcode_i[0];
  assign N30 = N20 | N29;
  assign N31 = N27 | N22;
  assign N32 = N27 | N29;
  assign N33 = N27 | N24;
  assign N34 = N152 | opcode_i[2];
  assign N35 = N17 | N34;
  assign N36 = N35 | N19;
  assign N37 = opcode_i[5] | opcode_i[4];
  assign N38 = N37 | N18;
  assign N39 = N38 | N24;
  assign N40 = N37 | N34;
  assign N41 = N40 | N24;
  assign N42 = N37 | N26;
  assign N43 = N42 | N24;
  assign N45 = N80 | opcode_i[4];
  assign N46 = N45 | N18;
  assign N47 = N46 | N19;
  assign N48 = N46 | N22;
  assign N49 = N46 | N24;
  assign N50 = N45 | N26;
  assign N51 = N50 | N19;
  assign N52 = N46 | N29;
  assign N53 = N50 | N22;
  assign N54 = N50 | N29;
  assign N55 = N50 | N24;
  assign N56 = N45 | N34;
  assign N57 = N56 | N19;
  assign N58 = N38 | N29;
  assign N59 = N40 | N29;
  assign N60 = N42 | N29;
  assign N62 = N38 | N22;
  assign N63 = N40 | N22;
  assign N64 = N42 | N22;
  assign N66 = N80 & N138;
  assign N67 = N152 & N165;
  assign N68 = N146 & N139;
  assign N69 = N66 & N67;
  assign N70 = N69 & N68;
  assign N71 = N40 | N19;
  assign N72 = N42 | N19;
  assign N74 = opcode_i[5] & opcode_i[3];
  assign N75 = N74 & opcode_i[0];
  assign N76 = N74 & opcode_i[1];
  assign N77 = opcode_i[3] & opcode_i[2];
  assign N78 = N80 & opcode_i[4];
  assign N81 = N138 & N152;
  assign N82 = N165 & N146;
  assign N83 = N81 & N82;
  assign N84 = N83 & N139;
  assign N85 = N138 | opcode_i[3];
  assign N86 = opcode_i[2] | opcode_i[1];
  assign N87 = N85 | N86;
  assign N88 = N87 | opcode_i[0];
  assign N90 = opcode_i[4] | opcode_i[3];
  assign N91 = N90 | N86;
  assign N92 = N91 | N139;
  assign N93 = N87 | N139;
  assign N95 = opcode_i[2] | N146;
  assign N96 = N90 | N95;
  assign N97 = N96 | opcode_i[0];
  assign N98 = N85 | N95;
  assign N99 = N98 | opcode_i[0];
  assign N101 = N96 | N139;
  assign N102 = N98 | N139;
  assign N104 = N165 | opcode_i[1];
  assign N105 = N90 | N104;
  assign N106 = N105 | opcode_i[0];
  assign N107 = N85 | N104;
  assign N108 = N107 | opcode_i[0];
  assign N110 = N105 | N139;
  assign N111 = N107 | N139;
  assign N113 = N165 | N146;
  assign N114 = N90 | N113;
  assign N115 = N114 | opcode_i[0];
  assign N116 = N85 | N113;
  assign N117 = N116 | opcode_i[0];
  assign N119 = N114 | N139;
  assign N120 = N116 | N139;
  assign N122 = opcode_i[4] | N152;
  assign N123 = N122 | N86;
  assign N124 = N123 | opcode_i[0];
  assign N125 = N138 | N152;
  assign N126 = N125 | N86;
  assign N127 = N126 | opcode_i[0];
  assign N129 = opcode_i[3] & opcode_i[0];
  assign N130 = opcode_i[3] & opcode_i[1];
  assign N138 = ~opcode_i[4];
  assign N139 = ~opcode_i[0];
  assign N140 = N138 | opcode_i[5];
  assign N141 = opcode_i[3] | N140;
  assign N142 = opcode_i[2] | N141;
  assign N143 = opcode_i[1] | N142;
  assign N144 = N139 | N143;
  assign decode_o[13] = ~N144;
  assign N146 = ~opcode_i[1];
  assign N147 = N146 | N142;
  assign N148 = opcode_i[0] | N147;
  assign decode_o[12] = ~N148;
  assign N150 = N139 | N147;
  assign decode_o[11] = ~N150;
  assign N152 = ~opcode_i[3];
  assign N153 = N152 | N140;
  assign N154 = opcode_i[2] | N153;
  assign N155 = opcode_i[1] | N154;
  assign N156 = opcode_i[0] | N155;
  assign decode_o[10] = ~N156;
  assign N158 = N139 | N155;
  assign decode_o[9] = ~N158;
  assign N160 = N146 | N154;
  assign N161 = opcode_i[0] | N160;
  assign decode_o[8] = ~N161;
  assign N163 = N139 | N160;
  assign decode_o[7] = ~N163;
  assign N165 = ~opcode_i[2];
  assign N166 = N165 | N153;
  assign N167 = opcode_i[1] | N166;
  assign N168 = opcode_i[0] | N167;
  assign decode_o[6] = ~N168;
  assign N170 = opcode_i[4] | opcode_i[5];
  assign N171 = opcode_i[3] | N170;
  assign N172 = opcode_i[2] | N171;
  assign N173 = opcode_i[1] | N172;
  assign N174 = opcode_i[0] | N173;
  assign N175 = ~N174;
  assign N176 = N139 | N173;
  assign N177 = ~N176;
  assign N178 = N146 | N172;
  assign N179 = opcode_i[0] | N178;
  assign N180 = ~N179;
  assign N181 = N139 | N178;
  assign N182 = ~N181;
  assign N183 = N152 | N170;
  assign N184 = N165 | N183;
  assign N185 = opcode_i[1] | N184;
  assign N186 = opcode_i[0] | N185;
  assign N187 = ~N186;
  assign N188 = N139 | N185;
  assign N189 = ~N188;
  assign N190 = N165 | N171;
  assign N191 = opcode_i[1] | N190;
  assign N192 = opcode_i[0] | N191;
  assign N193 = ~N192;
  assign N194 = N139 | N191;
  assign N195 = ~N194;
  assign N196 = N146 | N190;
  assign N197 = opcode_i[0] | N196;
  assign N198 = ~N197;
  assign N199 = N139 | N196;
  assign N200 = ~N199;
  assign N201 = opcode_i[2] | N183;
  assign N202 = opcode_i[1] | N201;
  assign N203 = opcode_i[0] | N202;
  assign N204 = ~N203;
  assign N205 = N139 | N202;
  assign N206 = ~N205;
  assign N207 = N146 | N201;
  assign N208 = opcode_i[0] | N207;
  assign N209 = ~N208;
  assign N210 = N139 | N207;
  assign N211 = ~N210;
  assign N212 = opcode_i[0] | N143;
  assign decode_o[14] = ~N212;
  assign decode_o[20:19] = (N0)? { 1'b1, 1'b1 } : 
                           (N1)? { 1'b1, 1'b0 } : 
                           (N2)? { 1'b0, 1'b1 } : 
                           (N3)? { 1'b0, 1'b0 } : 
                           (N4)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = N44;
  assign N1 = N61;
  assign N2 = N65;
  assign N3 = N73;
  assign N4 = N79;
  assign { N135, N134, N133, N132 } = (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                      (N6)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                      (N7)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                      (N8)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                      (N9)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                      (N10)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                      (N11)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                      (N12)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                      (N13)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                      (N14)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N89;
  assign N6 = N94;
  assign N7 = N100;
  assign N8 = N103;
  assign N9 = N109;
  assign N10 = N112;
  assign N11 = N118;
  assign N12 = N121;
  assign N13 = N128;
  assign N14 = N131;
  assign decode_o[4:0] = (N15)? { N137, N135, N134, N133, N132 } : 
                         (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = opcode_i[5];
  assign N16 = N80;
  assign N44 = N234 | N235;
  assign N234 = N232 | N233;
  assign N232 = N230 | N231;
  assign N230 = N228 | N229;
  assign N228 = N226 | N227;
  assign N226 = N224 | N225;
  assign N224 = N222 | N223;
  assign N222 = N220 | N221;
  assign N220 = N218 | N219;
  assign N218 = N216 | N217;
  assign N216 = N214 | N215;
  assign N214 = ~N21;
  assign N215 = ~N23;
  assign N217 = ~N25;
  assign N219 = ~N28;
  assign N221 = ~N30;
  assign N223 = ~N31;
  assign N225 = ~N32;
  assign N227 = ~N33;
  assign N229 = ~N36;
  assign N231 = ~N39;
  assign N233 = ~N41;
  assign N235 = ~N43;
  assign N61 = N256 | N257;
  assign N256 = N254 | N255;
  assign N254 = N252 | N253;
  assign N252 = N250 | N251;
  assign N250 = N248 | N249;
  assign N248 = N246 | N247;
  assign N246 = N244 | N245;
  assign N244 = N242 | N243;
  assign N242 = N240 | N241;
  assign N240 = N238 | N239;
  assign N238 = N236 | N237;
  assign N236 = ~N47;
  assign N237 = ~N48;
  assign N239 = ~N49;
  assign N241 = ~N51;
  assign N243 = ~N52;
  assign N245 = ~N53;
  assign N247 = ~N54;
  assign N249 = ~N55;
  assign N251 = ~N57;
  assign N253 = ~N58;
  assign N255 = ~N59;
  assign N257 = ~N60;
  assign N65 = N260 | N261;
  assign N260 = N258 | N259;
  assign N258 = ~N62;
  assign N259 = ~N63;
  assign N261 = ~N64;
  assign N73 = N263 | N264;
  assign N263 = N70 | N262;
  assign N262 = ~N71;
  assign N264 = ~N72;
  assign N79 = N75 | N266;
  assign N266 = N76 | N265;
  assign N265 = N77 | N78;
  assign decode_o[17] = N187 | N189;
  assign decode_o[18] = N269 | decode_o[4];
  assign N269 = N268 | N182;
  assign N268 = N267 | N180;
  assign N267 = N175 | N177;
  assign decode_o[16] = N276 | N187;
  assign N276 = N275 | N200;
  assign N275 = N274 | N198;
  assign N274 = N273 | N195;
  assign N273 = N272 | N193;
  assign N272 = N271 | N182;
  assign N271 = N270 | N180;
  assign N270 = N175 | N177;
  assign decode_o[15] = N279 | N189;
  assign N279 = N278 | N211;
  assign N278 = N277 | N209;
  assign N277 = N204 | N206;
  assign decode_o[5] = ~decode_o[14];
  assign N80 = ~opcode_i[5];
  assign N89 = N84 | N280;
  assign N280 = ~N88;
  assign N94 = N281 | N282;
  assign N281 = ~N92;
  assign N282 = ~N93;
  assign N100 = N283 | N284;
  assign N283 = ~N97;
  assign N284 = ~N99;
  assign N103 = N285 | N286;
  assign N285 = ~N101;
  assign N286 = ~N102;
  assign N109 = N287 | N288;
  assign N287 = ~N106;
  assign N288 = ~N108;
  assign N112 = N289 | N290;
  assign N289 = ~N110;
  assign N290 = ~N111;
  assign N118 = N291 | N292;
  assign N291 = ~N115;
  assign N292 = ~N117;
  assign N121 = N293 | N294;
  assign N293 = ~N119;
  assign N294 = ~N120;
  assign N128 = N295 | N296;
  assign N295 = ~N124;
  assign N296 = ~N127;
  assign N131 = N129 | N297;
  assign N297 = N130 | N77;
  assign N136 = ~N131;
  assign N137 = N136;

endmodule



module bsg_dff_width_p1
(
  clk_i,
  data_i,
  data_o
);

  input [0:0] data_i;
  output [0:0] data_o;
  input clk_i;
  wire [0:0] data_o;
  reg data_o_0_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_width_p40_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input en_i;
  wire [39:0] data_o;
  reg data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_39_sv2v_reg <= data_i[39];
      data_o_38_sv2v_reg <= data_i[38];
      data_o_37_sv2v_reg <= data_i[37];
      data_o_36_sv2v_reg <= data_i[36];
      data_o_35_sv2v_reg <= data_i[35];
      data_o_34_sv2v_reg <= data_i[34];
      data_o_33_sv2v_reg <= data_i[33];
      data_o_32_sv2v_reg <= data_i[32];
      data_o_31_sv2v_reg <= data_i[31];
      data_o_30_sv2v_reg <= data_i[30];
      data_o_29_sv2v_reg <= data_i[29];
      data_o_28_sv2v_reg <= data_i[28];
      data_o_27_sv2v_reg <= data_i[27];
      data_o_26_sv2v_reg <= data_i[26];
      data_o_25_sv2v_reg <= data_i[25];
      data_o_24_sv2v_reg <= data_i[24];
      data_o_23_sv2v_reg <= data_i[23];
      data_o_22_sv2v_reg <= data_i[22];
      data_o_21_sv2v_reg <= data_i[21];
      data_o_20_sv2v_reg <= data_i[20];
      data_o_19_sv2v_reg <= data_i[19];
      data_o_18_sv2v_reg <= data_i[18];
      data_o_17_sv2v_reg <= data_i[17];
      data_o_16_sv2v_reg <= data_i[16];
      data_o_15_sv2v_reg <= data_i[15];
      data_o_14_sv2v_reg <= data_i[14];
      data_o_13_sv2v_reg <= data_i[13];
      data_o_12_sv2v_reg <= data_i[12];
      data_o_11_sv2v_reg <= data_i[11];
      data_o_10_sv2v_reg <= data_i[10];
      data_o_9_sv2v_reg <= data_i[9];
      data_o_8_sv2v_reg <= data_i[8];
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p40
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [39:0] data_i;
  output [39:0] data_o;
  input clk_i;
  input en_i;
  wire [39:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p40_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p40_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [39:0] data_i;
  input [5:0] addr_i;
  input [39:0] w_mask_i;
  output [39:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [39:0] data_o,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,\nz.read_en ,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  \nz.llr.read_en_r ,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,
  N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,
  N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,
  N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,
  N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,
  N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,
  N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,
  N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
  N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,
  N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,
  N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
  N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,
  N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,
  N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
  N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,
  N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,
  N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
  N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,
  N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,
  N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
  N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,
  N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,
  N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
  N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,
  N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,
  N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
  N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,
  N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,
  N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
  N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,
  N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,
  N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
  N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,
  N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,
  N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
  N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,
  N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,
  N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
  N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,
  N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,
  N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
  N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,
  N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,
  N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
  N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,
  N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,
  N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
  N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,
  N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,
  N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
  N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,
  N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,
  N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
  N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,
  N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,
  N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
  N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,
  N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,
  N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
  N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,
  N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,
  N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
  N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,
  N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,
  N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
  N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,
  N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,
  N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
  N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,
  N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,
  N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
  N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,
  N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,
  N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
  N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,
  N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,
  N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
  N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,
  N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,
  N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
  N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,
  N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,
  N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
  N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,
  N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,
  N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
  N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,
  N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,
  N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
  N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,
  N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,
  N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
  N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
  N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,
  N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
  N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,
  N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,
  N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
  N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,
  N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,
  N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
  N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,
  N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,
  N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
  N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,
  N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,
  N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
  N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,
  N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,
  N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
  N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,
  N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,
  N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
  N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,
  N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,
  N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
  N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,
  N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,
  N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
  N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,
  N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,
  N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
  N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,
  N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,
  N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
  N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,
  N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,
  N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
  N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,
  N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,
  N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
  N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,
  N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,
  N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
  N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,
  N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,
  N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
  N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,
  N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,
  N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
  N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,
  N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,
  N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
  N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,
  N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,
  N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
  N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,
  N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,
  N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
  N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,
  N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
  N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
  N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,
  N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,
  N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
  N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,
  N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,
  N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
  N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,
  N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,
  N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
  N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,
  N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,
  N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
  N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,
  N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,
  N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
  N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,
  N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,
  N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
  N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,
  N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,
  N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
  N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,
  N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,
  N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
  N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,
  N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,
  N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
  N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,
  N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,
  N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
  N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,
  N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,
  N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
  N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,
  N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,
  N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
  N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,
  N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,
  N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
  N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,
  N4193,N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,
  N4206,N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,
  N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,
  N4233,N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,
  N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,
  N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,
  N4273,N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,
  N4286,N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,
  N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,
  N4313,N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,
  N4326,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,
  N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,
  N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,
  N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,
  N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,
  N4393,N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,
  N4406,N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,
  N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,
  N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,
  N4446,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,
  N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,
  N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,
  N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,
  N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,
  N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,
  N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,
  N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,
  N4553,N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,
  N4566,N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,
  N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,
  N4593,N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,
  N4606,N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,
  N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,
  N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,
  N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,
  N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,
  N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,
  N4686,N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,
  N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,
  N4713,N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,
  N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,
  N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,
  N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,
  N4766,N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,
  N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,
  N4793,N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,
  N4806,N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,
  N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,
  N4833,N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,
  N4846,N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,
  N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,
  N4873,N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,
  N4886,N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,
  N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,
  N4913,N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,
  N4926,N4927,N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,
  N4939,N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,
  N4953,N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,
  N4966,N4967,N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,
  N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,
  N4993,N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,
  N5006,N5007,N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,
  N5019,N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,
  N5033,N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,
  N5046,N5047,N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,
  N5059,N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,
  N5073,N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,
  N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,
  N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,
  N5113,N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,
  N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,
  N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,
  N5153,N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,
  N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,
  N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,
  N5193,N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,
  N5206,N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,
  N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,
  N5233,N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,
  N5246,N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,
  N5259,N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,
  N5273,N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,
  N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,
  N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,
  N5313,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,
  N5326,N5327,N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,
  N5339,N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,
  N5353,N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,
  N5366,N5367,N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,
  N5379,N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,
  N5393,N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,
  N5406,N5407,N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,
  N5419,N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,
  N5433,N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,
  N5446,N5447,N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,
  N5459,N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,
  N5473,N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,
  N5486,N5487,N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,
  N5499,N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,
  N5513,N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,
  N5526,N5527,N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,
  N5539,N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,
  N5553,N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,
  N5566,N5567,N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,
  N5579,N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,
  N5593,N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,
  N5606,N5607,N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,
  N5619,N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,
  N5633,N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,
  N5646,N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,
  N5659,N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,
  N5673,N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,
  N5686,N5687,N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,
  N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,
  N5713,N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,
  N5726,N5727,N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,
  N5739,N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,
  N5753,N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,
  N5766,N5767,N5768,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,
  N5779,N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,
  N5793,N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,
  N5806,N5807,N5808,N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,
  N5819,N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,
  N5833,N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,
  N5846,N5847,N5848,N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,
  N5859,N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,
  N5873,N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,
  N5886,N5887,N5888,N5889,N5890,N5891,N5892,N5893;
  wire [5:0] \nz.addr_r ;
  wire [2559:0] \nz.mem ;
  reg \nz.addr_r_5_sv2v_reg ,\nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,
  \nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,
  \nz.mem_2559_sv2v_reg ,\nz.mem_2558_sv2v_reg ,\nz.mem_2557_sv2v_reg ,\nz.mem_2556_sv2v_reg ,
  \nz.mem_2555_sv2v_reg ,\nz.mem_2554_sv2v_reg ,\nz.mem_2553_sv2v_reg ,
  \nz.mem_2552_sv2v_reg ,\nz.mem_2551_sv2v_reg ,\nz.mem_2550_sv2v_reg ,\nz.mem_2549_sv2v_reg ,
  \nz.mem_2548_sv2v_reg ,\nz.mem_2547_sv2v_reg ,\nz.mem_2546_sv2v_reg ,
  \nz.mem_2545_sv2v_reg ,\nz.mem_2544_sv2v_reg ,\nz.mem_2543_sv2v_reg ,\nz.mem_2542_sv2v_reg ,
  \nz.mem_2541_sv2v_reg ,\nz.mem_2540_sv2v_reg ,\nz.mem_2539_sv2v_reg ,
  \nz.mem_2538_sv2v_reg ,\nz.mem_2537_sv2v_reg ,\nz.mem_2536_sv2v_reg ,\nz.mem_2535_sv2v_reg ,
  \nz.mem_2534_sv2v_reg ,\nz.mem_2533_sv2v_reg ,\nz.mem_2532_sv2v_reg ,
  \nz.mem_2531_sv2v_reg ,\nz.mem_2530_sv2v_reg ,\nz.mem_2529_sv2v_reg ,\nz.mem_2528_sv2v_reg ,
  \nz.mem_2527_sv2v_reg ,\nz.mem_2526_sv2v_reg ,\nz.mem_2525_sv2v_reg ,
  \nz.mem_2524_sv2v_reg ,\nz.mem_2523_sv2v_reg ,\nz.mem_2522_sv2v_reg ,\nz.mem_2521_sv2v_reg ,
  \nz.mem_2520_sv2v_reg ,\nz.mem_2519_sv2v_reg ,\nz.mem_2518_sv2v_reg ,
  \nz.mem_2517_sv2v_reg ,\nz.mem_2516_sv2v_reg ,\nz.mem_2515_sv2v_reg ,\nz.mem_2514_sv2v_reg ,
  \nz.mem_2513_sv2v_reg ,\nz.mem_2512_sv2v_reg ,\nz.mem_2511_sv2v_reg ,
  \nz.mem_2510_sv2v_reg ,\nz.mem_2509_sv2v_reg ,\nz.mem_2508_sv2v_reg ,\nz.mem_2507_sv2v_reg ,
  \nz.mem_2506_sv2v_reg ,\nz.mem_2505_sv2v_reg ,\nz.mem_2504_sv2v_reg ,
  \nz.mem_2503_sv2v_reg ,\nz.mem_2502_sv2v_reg ,\nz.mem_2501_sv2v_reg ,\nz.mem_2500_sv2v_reg ,
  \nz.mem_2499_sv2v_reg ,\nz.mem_2498_sv2v_reg ,\nz.mem_2497_sv2v_reg ,
  \nz.mem_2496_sv2v_reg ,\nz.mem_2495_sv2v_reg ,\nz.mem_2494_sv2v_reg ,\nz.mem_2493_sv2v_reg ,
  \nz.mem_2492_sv2v_reg ,\nz.mem_2491_sv2v_reg ,\nz.mem_2490_sv2v_reg ,
  \nz.mem_2489_sv2v_reg ,\nz.mem_2488_sv2v_reg ,\nz.mem_2487_sv2v_reg ,\nz.mem_2486_sv2v_reg ,
  \nz.mem_2485_sv2v_reg ,\nz.mem_2484_sv2v_reg ,\nz.mem_2483_sv2v_reg ,
  \nz.mem_2482_sv2v_reg ,\nz.mem_2481_sv2v_reg ,\nz.mem_2480_sv2v_reg ,
  \nz.mem_2479_sv2v_reg ,\nz.mem_2478_sv2v_reg ,\nz.mem_2477_sv2v_reg ,\nz.mem_2476_sv2v_reg ,
  \nz.mem_2475_sv2v_reg ,\nz.mem_2474_sv2v_reg ,\nz.mem_2473_sv2v_reg ,
  \nz.mem_2472_sv2v_reg ,\nz.mem_2471_sv2v_reg ,\nz.mem_2470_sv2v_reg ,\nz.mem_2469_sv2v_reg ,
  \nz.mem_2468_sv2v_reg ,\nz.mem_2467_sv2v_reg ,\nz.mem_2466_sv2v_reg ,
  \nz.mem_2465_sv2v_reg ,\nz.mem_2464_sv2v_reg ,\nz.mem_2463_sv2v_reg ,\nz.mem_2462_sv2v_reg ,
  \nz.mem_2461_sv2v_reg ,\nz.mem_2460_sv2v_reg ,\nz.mem_2459_sv2v_reg ,
  \nz.mem_2458_sv2v_reg ,\nz.mem_2457_sv2v_reg ,\nz.mem_2456_sv2v_reg ,\nz.mem_2455_sv2v_reg ,
  \nz.mem_2454_sv2v_reg ,\nz.mem_2453_sv2v_reg ,\nz.mem_2452_sv2v_reg ,
  \nz.mem_2451_sv2v_reg ,\nz.mem_2450_sv2v_reg ,\nz.mem_2449_sv2v_reg ,\nz.mem_2448_sv2v_reg ,
  \nz.mem_2447_sv2v_reg ,\nz.mem_2446_sv2v_reg ,\nz.mem_2445_sv2v_reg ,
  \nz.mem_2444_sv2v_reg ,\nz.mem_2443_sv2v_reg ,\nz.mem_2442_sv2v_reg ,\nz.mem_2441_sv2v_reg ,
  \nz.mem_2440_sv2v_reg ,\nz.mem_2439_sv2v_reg ,\nz.mem_2438_sv2v_reg ,
  \nz.mem_2437_sv2v_reg ,\nz.mem_2436_sv2v_reg ,\nz.mem_2435_sv2v_reg ,\nz.mem_2434_sv2v_reg ,
  \nz.mem_2433_sv2v_reg ,\nz.mem_2432_sv2v_reg ,\nz.mem_2431_sv2v_reg ,
  \nz.mem_2430_sv2v_reg ,\nz.mem_2429_sv2v_reg ,\nz.mem_2428_sv2v_reg ,\nz.mem_2427_sv2v_reg ,
  \nz.mem_2426_sv2v_reg ,\nz.mem_2425_sv2v_reg ,\nz.mem_2424_sv2v_reg ,
  \nz.mem_2423_sv2v_reg ,\nz.mem_2422_sv2v_reg ,\nz.mem_2421_sv2v_reg ,\nz.mem_2420_sv2v_reg ,
  \nz.mem_2419_sv2v_reg ,\nz.mem_2418_sv2v_reg ,\nz.mem_2417_sv2v_reg ,
  \nz.mem_2416_sv2v_reg ,\nz.mem_2415_sv2v_reg ,\nz.mem_2414_sv2v_reg ,\nz.mem_2413_sv2v_reg ,
  \nz.mem_2412_sv2v_reg ,\nz.mem_2411_sv2v_reg ,\nz.mem_2410_sv2v_reg ,
  \nz.mem_2409_sv2v_reg ,\nz.mem_2408_sv2v_reg ,\nz.mem_2407_sv2v_reg ,\nz.mem_2406_sv2v_reg ,
  \nz.mem_2405_sv2v_reg ,\nz.mem_2404_sv2v_reg ,\nz.mem_2403_sv2v_reg ,
  \nz.mem_2402_sv2v_reg ,\nz.mem_2401_sv2v_reg ,\nz.mem_2400_sv2v_reg ,
  \nz.mem_2399_sv2v_reg ,\nz.mem_2398_sv2v_reg ,\nz.mem_2397_sv2v_reg ,\nz.mem_2396_sv2v_reg ,
  \nz.mem_2395_sv2v_reg ,\nz.mem_2394_sv2v_reg ,\nz.mem_2393_sv2v_reg ,
  \nz.mem_2392_sv2v_reg ,\nz.mem_2391_sv2v_reg ,\nz.mem_2390_sv2v_reg ,\nz.mem_2389_sv2v_reg ,
  \nz.mem_2388_sv2v_reg ,\nz.mem_2387_sv2v_reg ,\nz.mem_2386_sv2v_reg ,
  \nz.mem_2385_sv2v_reg ,\nz.mem_2384_sv2v_reg ,\nz.mem_2383_sv2v_reg ,\nz.mem_2382_sv2v_reg ,
  \nz.mem_2381_sv2v_reg ,\nz.mem_2380_sv2v_reg ,\nz.mem_2379_sv2v_reg ,
  \nz.mem_2378_sv2v_reg ,\nz.mem_2377_sv2v_reg ,\nz.mem_2376_sv2v_reg ,\nz.mem_2375_sv2v_reg ,
  \nz.mem_2374_sv2v_reg ,\nz.mem_2373_sv2v_reg ,\nz.mem_2372_sv2v_reg ,
  \nz.mem_2371_sv2v_reg ,\nz.mem_2370_sv2v_reg ,\nz.mem_2369_sv2v_reg ,\nz.mem_2368_sv2v_reg ,
  \nz.mem_2367_sv2v_reg ,\nz.mem_2366_sv2v_reg ,\nz.mem_2365_sv2v_reg ,
  \nz.mem_2364_sv2v_reg ,\nz.mem_2363_sv2v_reg ,\nz.mem_2362_sv2v_reg ,\nz.mem_2361_sv2v_reg ,
  \nz.mem_2360_sv2v_reg ,\nz.mem_2359_sv2v_reg ,\nz.mem_2358_sv2v_reg ,
  \nz.mem_2357_sv2v_reg ,\nz.mem_2356_sv2v_reg ,\nz.mem_2355_sv2v_reg ,\nz.mem_2354_sv2v_reg ,
  \nz.mem_2353_sv2v_reg ,\nz.mem_2352_sv2v_reg ,\nz.mem_2351_sv2v_reg ,
  \nz.mem_2350_sv2v_reg ,\nz.mem_2349_sv2v_reg ,\nz.mem_2348_sv2v_reg ,\nz.mem_2347_sv2v_reg ,
  \nz.mem_2346_sv2v_reg ,\nz.mem_2345_sv2v_reg ,\nz.mem_2344_sv2v_reg ,
  \nz.mem_2343_sv2v_reg ,\nz.mem_2342_sv2v_reg ,\nz.mem_2341_sv2v_reg ,\nz.mem_2340_sv2v_reg ,
  \nz.mem_2339_sv2v_reg ,\nz.mem_2338_sv2v_reg ,\nz.mem_2337_sv2v_reg ,
  \nz.mem_2336_sv2v_reg ,\nz.mem_2335_sv2v_reg ,\nz.mem_2334_sv2v_reg ,\nz.mem_2333_sv2v_reg ,
  \nz.mem_2332_sv2v_reg ,\nz.mem_2331_sv2v_reg ,\nz.mem_2330_sv2v_reg ,
  \nz.mem_2329_sv2v_reg ,\nz.mem_2328_sv2v_reg ,\nz.mem_2327_sv2v_reg ,\nz.mem_2326_sv2v_reg ,
  \nz.mem_2325_sv2v_reg ,\nz.mem_2324_sv2v_reg ,\nz.mem_2323_sv2v_reg ,
  \nz.mem_2322_sv2v_reg ,\nz.mem_2321_sv2v_reg ,\nz.mem_2320_sv2v_reg ,
  \nz.mem_2319_sv2v_reg ,\nz.mem_2318_sv2v_reg ,\nz.mem_2317_sv2v_reg ,\nz.mem_2316_sv2v_reg ,
  \nz.mem_2315_sv2v_reg ,\nz.mem_2314_sv2v_reg ,\nz.mem_2313_sv2v_reg ,
  \nz.mem_2312_sv2v_reg ,\nz.mem_2311_sv2v_reg ,\nz.mem_2310_sv2v_reg ,\nz.mem_2309_sv2v_reg ,
  \nz.mem_2308_sv2v_reg ,\nz.mem_2307_sv2v_reg ,\nz.mem_2306_sv2v_reg ,
  \nz.mem_2305_sv2v_reg ,\nz.mem_2304_sv2v_reg ,\nz.mem_2303_sv2v_reg ,\nz.mem_2302_sv2v_reg ,
  \nz.mem_2301_sv2v_reg ,\nz.mem_2300_sv2v_reg ,\nz.mem_2299_sv2v_reg ,
  \nz.mem_2298_sv2v_reg ,\nz.mem_2297_sv2v_reg ,\nz.mem_2296_sv2v_reg ,\nz.mem_2295_sv2v_reg ,
  \nz.mem_2294_sv2v_reg ,\nz.mem_2293_sv2v_reg ,\nz.mem_2292_sv2v_reg ,
  \nz.mem_2291_sv2v_reg ,\nz.mem_2290_sv2v_reg ,\nz.mem_2289_sv2v_reg ,\nz.mem_2288_sv2v_reg ,
  \nz.mem_2287_sv2v_reg ,\nz.mem_2286_sv2v_reg ,\nz.mem_2285_sv2v_reg ,
  \nz.mem_2284_sv2v_reg ,\nz.mem_2283_sv2v_reg ,\nz.mem_2282_sv2v_reg ,\nz.mem_2281_sv2v_reg ,
  \nz.mem_2280_sv2v_reg ,\nz.mem_2279_sv2v_reg ,\nz.mem_2278_sv2v_reg ,
  \nz.mem_2277_sv2v_reg ,\nz.mem_2276_sv2v_reg ,\nz.mem_2275_sv2v_reg ,\nz.mem_2274_sv2v_reg ,
  \nz.mem_2273_sv2v_reg ,\nz.mem_2272_sv2v_reg ,\nz.mem_2271_sv2v_reg ,
  \nz.mem_2270_sv2v_reg ,\nz.mem_2269_sv2v_reg ,\nz.mem_2268_sv2v_reg ,\nz.mem_2267_sv2v_reg ,
  \nz.mem_2266_sv2v_reg ,\nz.mem_2265_sv2v_reg ,\nz.mem_2264_sv2v_reg ,
  \nz.mem_2263_sv2v_reg ,\nz.mem_2262_sv2v_reg ,\nz.mem_2261_sv2v_reg ,\nz.mem_2260_sv2v_reg ,
  \nz.mem_2259_sv2v_reg ,\nz.mem_2258_sv2v_reg ,\nz.mem_2257_sv2v_reg ,
  \nz.mem_2256_sv2v_reg ,\nz.mem_2255_sv2v_reg ,\nz.mem_2254_sv2v_reg ,\nz.mem_2253_sv2v_reg ,
  \nz.mem_2252_sv2v_reg ,\nz.mem_2251_sv2v_reg ,\nz.mem_2250_sv2v_reg ,
  \nz.mem_2249_sv2v_reg ,\nz.mem_2248_sv2v_reg ,\nz.mem_2247_sv2v_reg ,\nz.mem_2246_sv2v_reg ,
  \nz.mem_2245_sv2v_reg ,\nz.mem_2244_sv2v_reg ,\nz.mem_2243_sv2v_reg ,
  \nz.mem_2242_sv2v_reg ,\nz.mem_2241_sv2v_reg ,\nz.mem_2240_sv2v_reg ,
  \nz.mem_2239_sv2v_reg ,\nz.mem_2238_sv2v_reg ,\nz.mem_2237_sv2v_reg ,\nz.mem_2236_sv2v_reg ,
  \nz.mem_2235_sv2v_reg ,\nz.mem_2234_sv2v_reg ,\nz.mem_2233_sv2v_reg ,
  \nz.mem_2232_sv2v_reg ,\nz.mem_2231_sv2v_reg ,\nz.mem_2230_sv2v_reg ,\nz.mem_2229_sv2v_reg ,
  \nz.mem_2228_sv2v_reg ,\nz.mem_2227_sv2v_reg ,\nz.mem_2226_sv2v_reg ,
  \nz.mem_2225_sv2v_reg ,\nz.mem_2224_sv2v_reg ,\nz.mem_2223_sv2v_reg ,\nz.mem_2222_sv2v_reg ,
  \nz.mem_2221_sv2v_reg ,\nz.mem_2220_sv2v_reg ,\nz.mem_2219_sv2v_reg ,
  \nz.mem_2218_sv2v_reg ,\nz.mem_2217_sv2v_reg ,\nz.mem_2216_sv2v_reg ,\nz.mem_2215_sv2v_reg ,
  \nz.mem_2214_sv2v_reg ,\nz.mem_2213_sv2v_reg ,\nz.mem_2212_sv2v_reg ,
  \nz.mem_2211_sv2v_reg ,\nz.mem_2210_sv2v_reg ,\nz.mem_2209_sv2v_reg ,\nz.mem_2208_sv2v_reg ,
  \nz.mem_2207_sv2v_reg ,\nz.mem_2206_sv2v_reg ,\nz.mem_2205_sv2v_reg ,
  \nz.mem_2204_sv2v_reg ,\nz.mem_2203_sv2v_reg ,\nz.mem_2202_sv2v_reg ,\nz.mem_2201_sv2v_reg ,
  \nz.mem_2200_sv2v_reg ,\nz.mem_2199_sv2v_reg ,\nz.mem_2198_sv2v_reg ,
  \nz.mem_2197_sv2v_reg ,\nz.mem_2196_sv2v_reg ,\nz.mem_2195_sv2v_reg ,\nz.mem_2194_sv2v_reg ,
  \nz.mem_2193_sv2v_reg ,\nz.mem_2192_sv2v_reg ,\nz.mem_2191_sv2v_reg ,
  \nz.mem_2190_sv2v_reg ,\nz.mem_2189_sv2v_reg ,\nz.mem_2188_sv2v_reg ,\nz.mem_2187_sv2v_reg ,
  \nz.mem_2186_sv2v_reg ,\nz.mem_2185_sv2v_reg ,\nz.mem_2184_sv2v_reg ,
  \nz.mem_2183_sv2v_reg ,\nz.mem_2182_sv2v_reg ,\nz.mem_2181_sv2v_reg ,\nz.mem_2180_sv2v_reg ,
  \nz.mem_2179_sv2v_reg ,\nz.mem_2178_sv2v_reg ,\nz.mem_2177_sv2v_reg ,
  \nz.mem_2176_sv2v_reg ,\nz.mem_2175_sv2v_reg ,\nz.mem_2174_sv2v_reg ,\nz.mem_2173_sv2v_reg ,
  \nz.mem_2172_sv2v_reg ,\nz.mem_2171_sv2v_reg ,\nz.mem_2170_sv2v_reg ,
  \nz.mem_2169_sv2v_reg ,\nz.mem_2168_sv2v_reg ,\nz.mem_2167_sv2v_reg ,\nz.mem_2166_sv2v_reg ,
  \nz.mem_2165_sv2v_reg ,\nz.mem_2164_sv2v_reg ,\nz.mem_2163_sv2v_reg ,
  \nz.mem_2162_sv2v_reg ,\nz.mem_2161_sv2v_reg ,\nz.mem_2160_sv2v_reg ,
  \nz.mem_2159_sv2v_reg ,\nz.mem_2158_sv2v_reg ,\nz.mem_2157_sv2v_reg ,\nz.mem_2156_sv2v_reg ,
  \nz.mem_2155_sv2v_reg ,\nz.mem_2154_sv2v_reg ,\nz.mem_2153_sv2v_reg ,
  \nz.mem_2152_sv2v_reg ,\nz.mem_2151_sv2v_reg ,\nz.mem_2150_sv2v_reg ,\nz.mem_2149_sv2v_reg ,
  \nz.mem_2148_sv2v_reg ,\nz.mem_2147_sv2v_reg ,\nz.mem_2146_sv2v_reg ,
  \nz.mem_2145_sv2v_reg ,\nz.mem_2144_sv2v_reg ,\nz.mem_2143_sv2v_reg ,\nz.mem_2142_sv2v_reg ,
  \nz.mem_2141_sv2v_reg ,\nz.mem_2140_sv2v_reg ,\nz.mem_2139_sv2v_reg ,
  \nz.mem_2138_sv2v_reg ,\nz.mem_2137_sv2v_reg ,\nz.mem_2136_sv2v_reg ,\nz.mem_2135_sv2v_reg ,
  \nz.mem_2134_sv2v_reg ,\nz.mem_2133_sv2v_reg ,\nz.mem_2132_sv2v_reg ,
  \nz.mem_2131_sv2v_reg ,\nz.mem_2130_sv2v_reg ,\nz.mem_2129_sv2v_reg ,\nz.mem_2128_sv2v_reg ,
  \nz.mem_2127_sv2v_reg ,\nz.mem_2126_sv2v_reg ,\nz.mem_2125_sv2v_reg ,
  \nz.mem_2124_sv2v_reg ,\nz.mem_2123_sv2v_reg ,\nz.mem_2122_sv2v_reg ,\nz.mem_2121_sv2v_reg ,
  \nz.mem_2120_sv2v_reg ,\nz.mem_2119_sv2v_reg ,\nz.mem_2118_sv2v_reg ,
  \nz.mem_2117_sv2v_reg ,\nz.mem_2116_sv2v_reg ,\nz.mem_2115_sv2v_reg ,\nz.mem_2114_sv2v_reg ,
  \nz.mem_2113_sv2v_reg ,\nz.mem_2112_sv2v_reg ,\nz.mem_2111_sv2v_reg ,
  \nz.mem_2110_sv2v_reg ,\nz.mem_2109_sv2v_reg ,\nz.mem_2108_sv2v_reg ,\nz.mem_2107_sv2v_reg ,
  \nz.mem_2106_sv2v_reg ,\nz.mem_2105_sv2v_reg ,\nz.mem_2104_sv2v_reg ,
  \nz.mem_2103_sv2v_reg ,\nz.mem_2102_sv2v_reg ,\nz.mem_2101_sv2v_reg ,\nz.mem_2100_sv2v_reg ,
  \nz.mem_2099_sv2v_reg ,\nz.mem_2098_sv2v_reg ,\nz.mem_2097_sv2v_reg ,
  \nz.mem_2096_sv2v_reg ,\nz.mem_2095_sv2v_reg ,\nz.mem_2094_sv2v_reg ,\nz.mem_2093_sv2v_reg ,
  \nz.mem_2092_sv2v_reg ,\nz.mem_2091_sv2v_reg ,\nz.mem_2090_sv2v_reg ,
  \nz.mem_2089_sv2v_reg ,\nz.mem_2088_sv2v_reg ,\nz.mem_2087_sv2v_reg ,\nz.mem_2086_sv2v_reg ,
  \nz.mem_2085_sv2v_reg ,\nz.mem_2084_sv2v_reg ,\nz.mem_2083_sv2v_reg ,
  \nz.mem_2082_sv2v_reg ,\nz.mem_2081_sv2v_reg ,\nz.mem_2080_sv2v_reg ,
  \nz.mem_2079_sv2v_reg ,\nz.mem_2078_sv2v_reg ,\nz.mem_2077_sv2v_reg ,\nz.mem_2076_sv2v_reg ,
  \nz.mem_2075_sv2v_reg ,\nz.mem_2074_sv2v_reg ,\nz.mem_2073_sv2v_reg ,
  \nz.mem_2072_sv2v_reg ,\nz.mem_2071_sv2v_reg ,\nz.mem_2070_sv2v_reg ,\nz.mem_2069_sv2v_reg ,
  \nz.mem_2068_sv2v_reg ,\nz.mem_2067_sv2v_reg ,\nz.mem_2066_sv2v_reg ,
  \nz.mem_2065_sv2v_reg ,\nz.mem_2064_sv2v_reg ,\nz.mem_2063_sv2v_reg ,\nz.mem_2062_sv2v_reg ,
  \nz.mem_2061_sv2v_reg ,\nz.mem_2060_sv2v_reg ,\nz.mem_2059_sv2v_reg ,
  \nz.mem_2058_sv2v_reg ,\nz.mem_2057_sv2v_reg ,\nz.mem_2056_sv2v_reg ,\nz.mem_2055_sv2v_reg ,
  \nz.mem_2054_sv2v_reg ,\nz.mem_2053_sv2v_reg ,\nz.mem_2052_sv2v_reg ,
  \nz.mem_2051_sv2v_reg ,\nz.mem_2050_sv2v_reg ,\nz.mem_2049_sv2v_reg ,\nz.mem_2048_sv2v_reg ,
  \nz.mem_2047_sv2v_reg ,\nz.mem_2046_sv2v_reg ,\nz.mem_2045_sv2v_reg ,
  \nz.mem_2044_sv2v_reg ,\nz.mem_2043_sv2v_reg ,\nz.mem_2042_sv2v_reg ,\nz.mem_2041_sv2v_reg ,
  \nz.mem_2040_sv2v_reg ,\nz.mem_2039_sv2v_reg ,\nz.mem_2038_sv2v_reg ,
  \nz.mem_2037_sv2v_reg ,\nz.mem_2036_sv2v_reg ,\nz.mem_2035_sv2v_reg ,\nz.mem_2034_sv2v_reg ,
  \nz.mem_2033_sv2v_reg ,\nz.mem_2032_sv2v_reg ,\nz.mem_2031_sv2v_reg ,
  \nz.mem_2030_sv2v_reg ,\nz.mem_2029_sv2v_reg ,\nz.mem_2028_sv2v_reg ,\nz.mem_2027_sv2v_reg ,
  \nz.mem_2026_sv2v_reg ,\nz.mem_2025_sv2v_reg ,\nz.mem_2024_sv2v_reg ,
  \nz.mem_2023_sv2v_reg ,\nz.mem_2022_sv2v_reg ,\nz.mem_2021_sv2v_reg ,\nz.mem_2020_sv2v_reg ,
  \nz.mem_2019_sv2v_reg ,\nz.mem_2018_sv2v_reg ,\nz.mem_2017_sv2v_reg ,
  \nz.mem_2016_sv2v_reg ,\nz.mem_2015_sv2v_reg ,\nz.mem_2014_sv2v_reg ,\nz.mem_2013_sv2v_reg ,
  \nz.mem_2012_sv2v_reg ,\nz.mem_2011_sv2v_reg ,\nz.mem_2010_sv2v_reg ,
  \nz.mem_2009_sv2v_reg ,\nz.mem_2008_sv2v_reg ,\nz.mem_2007_sv2v_reg ,\nz.mem_2006_sv2v_reg ,
  \nz.mem_2005_sv2v_reg ,\nz.mem_2004_sv2v_reg ,\nz.mem_2003_sv2v_reg ,
  \nz.mem_2002_sv2v_reg ,\nz.mem_2001_sv2v_reg ,\nz.mem_2000_sv2v_reg ,
  \nz.mem_1999_sv2v_reg ,\nz.mem_1998_sv2v_reg ,\nz.mem_1997_sv2v_reg ,\nz.mem_1996_sv2v_reg ,
  \nz.mem_1995_sv2v_reg ,\nz.mem_1994_sv2v_reg ,\nz.mem_1993_sv2v_reg ,
  \nz.mem_1992_sv2v_reg ,\nz.mem_1991_sv2v_reg ,\nz.mem_1990_sv2v_reg ,\nz.mem_1989_sv2v_reg ,
  \nz.mem_1988_sv2v_reg ,\nz.mem_1987_sv2v_reg ,\nz.mem_1986_sv2v_reg ,
  \nz.mem_1985_sv2v_reg ,\nz.mem_1984_sv2v_reg ,\nz.mem_1983_sv2v_reg ,\nz.mem_1982_sv2v_reg ,
  \nz.mem_1981_sv2v_reg ,\nz.mem_1980_sv2v_reg ,\nz.mem_1979_sv2v_reg ,
  \nz.mem_1978_sv2v_reg ,\nz.mem_1977_sv2v_reg ,\nz.mem_1976_sv2v_reg ,\nz.mem_1975_sv2v_reg ,
  \nz.mem_1974_sv2v_reg ,\nz.mem_1973_sv2v_reg ,\nz.mem_1972_sv2v_reg ,
  \nz.mem_1971_sv2v_reg ,\nz.mem_1970_sv2v_reg ,\nz.mem_1969_sv2v_reg ,\nz.mem_1968_sv2v_reg ,
  \nz.mem_1967_sv2v_reg ,\nz.mem_1966_sv2v_reg ,\nz.mem_1965_sv2v_reg ,
  \nz.mem_1964_sv2v_reg ,\nz.mem_1963_sv2v_reg ,\nz.mem_1962_sv2v_reg ,\nz.mem_1961_sv2v_reg ,
  \nz.mem_1960_sv2v_reg ,\nz.mem_1959_sv2v_reg ,\nz.mem_1958_sv2v_reg ,
  \nz.mem_1957_sv2v_reg ,\nz.mem_1956_sv2v_reg ,\nz.mem_1955_sv2v_reg ,\nz.mem_1954_sv2v_reg ,
  \nz.mem_1953_sv2v_reg ,\nz.mem_1952_sv2v_reg ,\nz.mem_1951_sv2v_reg ,
  \nz.mem_1950_sv2v_reg ,\nz.mem_1949_sv2v_reg ,\nz.mem_1948_sv2v_reg ,\nz.mem_1947_sv2v_reg ,
  \nz.mem_1946_sv2v_reg ,\nz.mem_1945_sv2v_reg ,\nz.mem_1944_sv2v_reg ,
  \nz.mem_1943_sv2v_reg ,\nz.mem_1942_sv2v_reg ,\nz.mem_1941_sv2v_reg ,\nz.mem_1940_sv2v_reg ,
  \nz.mem_1939_sv2v_reg ,\nz.mem_1938_sv2v_reg ,\nz.mem_1937_sv2v_reg ,
  \nz.mem_1936_sv2v_reg ,\nz.mem_1935_sv2v_reg ,\nz.mem_1934_sv2v_reg ,\nz.mem_1933_sv2v_reg ,
  \nz.mem_1932_sv2v_reg ,\nz.mem_1931_sv2v_reg ,\nz.mem_1930_sv2v_reg ,
  \nz.mem_1929_sv2v_reg ,\nz.mem_1928_sv2v_reg ,\nz.mem_1927_sv2v_reg ,\nz.mem_1926_sv2v_reg ,
  \nz.mem_1925_sv2v_reg ,\nz.mem_1924_sv2v_reg ,\nz.mem_1923_sv2v_reg ,
  \nz.mem_1922_sv2v_reg ,\nz.mem_1921_sv2v_reg ,\nz.mem_1920_sv2v_reg ,
  \nz.mem_1919_sv2v_reg ,\nz.mem_1918_sv2v_reg ,\nz.mem_1917_sv2v_reg ,\nz.mem_1916_sv2v_reg ,
  \nz.mem_1915_sv2v_reg ,\nz.mem_1914_sv2v_reg ,\nz.mem_1913_sv2v_reg ,
  \nz.mem_1912_sv2v_reg ,\nz.mem_1911_sv2v_reg ,\nz.mem_1910_sv2v_reg ,\nz.mem_1909_sv2v_reg ,
  \nz.mem_1908_sv2v_reg ,\nz.mem_1907_sv2v_reg ,\nz.mem_1906_sv2v_reg ,
  \nz.mem_1905_sv2v_reg ,\nz.mem_1904_sv2v_reg ,\nz.mem_1903_sv2v_reg ,\nz.mem_1902_sv2v_reg ,
  \nz.mem_1901_sv2v_reg ,\nz.mem_1900_sv2v_reg ,\nz.mem_1899_sv2v_reg ,
  \nz.mem_1898_sv2v_reg ,\nz.mem_1897_sv2v_reg ,\nz.mem_1896_sv2v_reg ,\nz.mem_1895_sv2v_reg ,
  \nz.mem_1894_sv2v_reg ,\nz.mem_1893_sv2v_reg ,\nz.mem_1892_sv2v_reg ,
  \nz.mem_1891_sv2v_reg ,\nz.mem_1890_sv2v_reg ,\nz.mem_1889_sv2v_reg ,\nz.mem_1888_sv2v_reg ,
  \nz.mem_1887_sv2v_reg ,\nz.mem_1886_sv2v_reg ,\nz.mem_1885_sv2v_reg ,
  \nz.mem_1884_sv2v_reg ,\nz.mem_1883_sv2v_reg ,\nz.mem_1882_sv2v_reg ,\nz.mem_1881_sv2v_reg ,
  \nz.mem_1880_sv2v_reg ,\nz.mem_1879_sv2v_reg ,\nz.mem_1878_sv2v_reg ,
  \nz.mem_1877_sv2v_reg ,\nz.mem_1876_sv2v_reg ,\nz.mem_1875_sv2v_reg ,\nz.mem_1874_sv2v_reg ,
  \nz.mem_1873_sv2v_reg ,\nz.mem_1872_sv2v_reg ,\nz.mem_1871_sv2v_reg ,
  \nz.mem_1870_sv2v_reg ,\nz.mem_1869_sv2v_reg ,\nz.mem_1868_sv2v_reg ,\nz.mem_1867_sv2v_reg ,
  \nz.mem_1866_sv2v_reg ,\nz.mem_1865_sv2v_reg ,\nz.mem_1864_sv2v_reg ,
  \nz.mem_1863_sv2v_reg ,\nz.mem_1862_sv2v_reg ,\nz.mem_1861_sv2v_reg ,\nz.mem_1860_sv2v_reg ,
  \nz.mem_1859_sv2v_reg ,\nz.mem_1858_sv2v_reg ,\nz.mem_1857_sv2v_reg ,
  \nz.mem_1856_sv2v_reg ,\nz.mem_1855_sv2v_reg ,\nz.mem_1854_sv2v_reg ,\nz.mem_1853_sv2v_reg ,
  \nz.mem_1852_sv2v_reg ,\nz.mem_1851_sv2v_reg ,\nz.mem_1850_sv2v_reg ,
  \nz.mem_1849_sv2v_reg ,\nz.mem_1848_sv2v_reg ,\nz.mem_1847_sv2v_reg ,\nz.mem_1846_sv2v_reg ,
  \nz.mem_1845_sv2v_reg ,\nz.mem_1844_sv2v_reg ,\nz.mem_1843_sv2v_reg ,
  \nz.mem_1842_sv2v_reg ,\nz.mem_1841_sv2v_reg ,\nz.mem_1840_sv2v_reg ,
  \nz.mem_1839_sv2v_reg ,\nz.mem_1838_sv2v_reg ,\nz.mem_1837_sv2v_reg ,\nz.mem_1836_sv2v_reg ,
  \nz.mem_1835_sv2v_reg ,\nz.mem_1834_sv2v_reg ,\nz.mem_1833_sv2v_reg ,
  \nz.mem_1832_sv2v_reg ,\nz.mem_1831_sv2v_reg ,\nz.mem_1830_sv2v_reg ,\nz.mem_1829_sv2v_reg ,
  \nz.mem_1828_sv2v_reg ,\nz.mem_1827_sv2v_reg ,\nz.mem_1826_sv2v_reg ,
  \nz.mem_1825_sv2v_reg ,\nz.mem_1824_sv2v_reg ,\nz.mem_1823_sv2v_reg ,\nz.mem_1822_sv2v_reg ,
  \nz.mem_1821_sv2v_reg ,\nz.mem_1820_sv2v_reg ,\nz.mem_1819_sv2v_reg ,
  \nz.mem_1818_sv2v_reg ,\nz.mem_1817_sv2v_reg ,\nz.mem_1816_sv2v_reg ,\nz.mem_1815_sv2v_reg ,
  \nz.mem_1814_sv2v_reg ,\nz.mem_1813_sv2v_reg ,\nz.mem_1812_sv2v_reg ,
  \nz.mem_1811_sv2v_reg ,\nz.mem_1810_sv2v_reg ,\nz.mem_1809_sv2v_reg ,\nz.mem_1808_sv2v_reg ,
  \nz.mem_1807_sv2v_reg ,\nz.mem_1806_sv2v_reg ,\nz.mem_1805_sv2v_reg ,
  \nz.mem_1804_sv2v_reg ,\nz.mem_1803_sv2v_reg ,\nz.mem_1802_sv2v_reg ,\nz.mem_1801_sv2v_reg ,
  \nz.mem_1800_sv2v_reg ,\nz.mem_1799_sv2v_reg ,\nz.mem_1798_sv2v_reg ,
  \nz.mem_1797_sv2v_reg ,\nz.mem_1796_sv2v_reg ,\nz.mem_1795_sv2v_reg ,\nz.mem_1794_sv2v_reg ,
  \nz.mem_1793_sv2v_reg ,\nz.mem_1792_sv2v_reg ,\nz.mem_1791_sv2v_reg ,
  \nz.mem_1790_sv2v_reg ,\nz.mem_1789_sv2v_reg ,\nz.mem_1788_sv2v_reg ,\nz.mem_1787_sv2v_reg ,
  \nz.mem_1786_sv2v_reg ,\nz.mem_1785_sv2v_reg ,\nz.mem_1784_sv2v_reg ,
  \nz.mem_1783_sv2v_reg ,\nz.mem_1782_sv2v_reg ,\nz.mem_1781_sv2v_reg ,\nz.mem_1780_sv2v_reg ,
  \nz.mem_1779_sv2v_reg ,\nz.mem_1778_sv2v_reg ,\nz.mem_1777_sv2v_reg ,
  \nz.mem_1776_sv2v_reg ,\nz.mem_1775_sv2v_reg ,\nz.mem_1774_sv2v_reg ,\nz.mem_1773_sv2v_reg ,
  \nz.mem_1772_sv2v_reg ,\nz.mem_1771_sv2v_reg ,\nz.mem_1770_sv2v_reg ,
  \nz.mem_1769_sv2v_reg ,\nz.mem_1768_sv2v_reg ,\nz.mem_1767_sv2v_reg ,\nz.mem_1766_sv2v_reg ,
  \nz.mem_1765_sv2v_reg ,\nz.mem_1764_sv2v_reg ,\nz.mem_1763_sv2v_reg ,
  \nz.mem_1762_sv2v_reg ,\nz.mem_1761_sv2v_reg ,\nz.mem_1760_sv2v_reg ,
  \nz.mem_1759_sv2v_reg ,\nz.mem_1758_sv2v_reg ,\nz.mem_1757_sv2v_reg ,\nz.mem_1756_sv2v_reg ,
  \nz.mem_1755_sv2v_reg ,\nz.mem_1754_sv2v_reg ,\nz.mem_1753_sv2v_reg ,
  \nz.mem_1752_sv2v_reg ,\nz.mem_1751_sv2v_reg ,\nz.mem_1750_sv2v_reg ,\nz.mem_1749_sv2v_reg ,
  \nz.mem_1748_sv2v_reg ,\nz.mem_1747_sv2v_reg ,\nz.mem_1746_sv2v_reg ,
  \nz.mem_1745_sv2v_reg ,\nz.mem_1744_sv2v_reg ,\nz.mem_1743_sv2v_reg ,\nz.mem_1742_sv2v_reg ,
  \nz.mem_1741_sv2v_reg ,\nz.mem_1740_sv2v_reg ,\nz.mem_1739_sv2v_reg ,
  \nz.mem_1738_sv2v_reg ,\nz.mem_1737_sv2v_reg ,\nz.mem_1736_sv2v_reg ,\nz.mem_1735_sv2v_reg ,
  \nz.mem_1734_sv2v_reg ,\nz.mem_1733_sv2v_reg ,\nz.mem_1732_sv2v_reg ,
  \nz.mem_1731_sv2v_reg ,\nz.mem_1730_sv2v_reg ,\nz.mem_1729_sv2v_reg ,\nz.mem_1728_sv2v_reg ,
  \nz.mem_1727_sv2v_reg ,\nz.mem_1726_sv2v_reg ,\nz.mem_1725_sv2v_reg ,
  \nz.mem_1724_sv2v_reg ,\nz.mem_1723_sv2v_reg ,\nz.mem_1722_sv2v_reg ,\nz.mem_1721_sv2v_reg ,
  \nz.mem_1720_sv2v_reg ,\nz.mem_1719_sv2v_reg ,\nz.mem_1718_sv2v_reg ,
  \nz.mem_1717_sv2v_reg ,\nz.mem_1716_sv2v_reg ,\nz.mem_1715_sv2v_reg ,\nz.mem_1714_sv2v_reg ,
  \nz.mem_1713_sv2v_reg ,\nz.mem_1712_sv2v_reg ,\nz.mem_1711_sv2v_reg ,
  \nz.mem_1710_sv2v_reg ,\nz.mem_1709_sv2v_reg ,\nz.mem_1708_sv2v_reg ,\nz.mem_1707_sv2v_reg ,
  \nz.mem_1706_sv2v_reg ,\nz.mem_1705_sv2v_reg ,\nz.mem_1704_sv2v_reg ,
  \nz.mem_1703_sv2v_reg ,\nz.mem_1702_sv2v_reg ,\nz.mem_1701_sv2v_reg ,\nz.mem_1700_sv2v_reg ,
  \nz.mem_1699_sv2v_reg ,\nz.mem_1698_sv2v_reg ,\nz.mem_1697_sv2v_reg ,
  \nz.mem_1696_sv2v_reg ,\nz.mem_1695_sv2v_reg ,\nz.mem_1694_sv2v_reg ,\nz.mem_1693_sv2v_reg ,
  \nz.mem_1692_sv2v_reg ,\nz.mem_1691_sv2v_reg ,\nz.mem_1690_sv2v_reg ,
  \nz.mem_1689_sv2v_reg ,\nz.mem_1688_sv2v_reg ,\nz.mem_1687_sv2v_reg ,\nz.mem_1686_sv2v_reg ,
  \nz.mem_1685_sv2v_reg ,\nz.mem_1684_sv2v_reg ,\nz.mem_1683_sv2v_reg ,
  \nz.mem_1682_sv2v_reg ,\nz.mem_1681_sv2v_reg ,\nz.mem_1680_sv2v_reg ,
  \nz.mem_1679_sv2v_reg ,\nz.mem_1678_sv2v_reg ,\nz.mem_1677_sv2v_reg ,\nz.mem_1676_sv2v_reg ,
  \nz.mem_1675_sv2v_reg ,\nz.mem_1674_sv2v_reg ,\nz.mem_1673_sv2v_reg ,
  \nz.mem_1672_sv2v_reg ,\nz.mem_1671_sv2v_reg ,\nz.mem_1670_sv2v_reg ,\nz.mem_1669_sv2v_reg ,
  \nz.mem_1668_sv2v_reg ,\nz.mem_1667_sv2v_reg ,\nz.mem_1666_sv2v_reg ,
  \nz.mem_1665_sv2v_reg ,\nz.mem_1664_sv2v_reg ,\nz.mem_1663_sv2v_reg ,\nz.mem_1662_sv2v_reg ,
  \nz.mem_1661_sv2v_reg ,\nz.mem_1660_sv2v_reg ,\nz.mem_1659_sv2v_reg ,
  \nz.mem_1658_sv2v_reg ,\nz.mem_1657_sv2v_reg ,\nz.mem_1656_sv2v_reg ,\nz.mem_1655_sv2v_reg ,
  \nz.mem_1654_sv2v_reg ,\nz.mem_1653_sv2v_reg ,\nz.mem_1652_sv2v_reg ,
  \nz.mem_1651_sv2v_reg ,\nz.mem_1650_sv2v_reg ,\nz.mem_1649_sv2v_reg ,\nz.mem_1648_sv2v_reg ,
  \nz.mem_1647_sv2v_reg ,\nz.mem_1646_sv2v_reg ,\nz.mem_1645_sv2v_reg ,
  \nz.mem_1644_sv2v_reg ,\nz.mem_1643_sv2v_reg ,\nz.mem_1642_sv2v_reg ,\nz.mem_1641_sv2v_reg ,
  \nz.mem_1640_sv2v_reg ,\nz.mem_1639_sv2v_reg ,\nz.mem_1638_sv2v_reg ,
  \nz.mem_1637_sv2v_reg ,\nz.mem_1636_sv2v_reg ,\nz.mem_1635_sv2v_reg ,\nz.mem_1634_sv2v_reg ,
  \nz.mem_1633_sv2v_reg ,\nz.mem_1632_sv2v_reg ,\nz.mem_1631_sv2v_reg ,
  \nz.mem_1630_sv2v_reg ,\nz.mem_1629_sv2v_reg ,\nz.mem_1628_sv2v_reg ,\nz.mem_1627_sv2v_reg ,
  \nz.mem_1626_sv2v_reg ,\nz.mem_1625_sv2v_reg ,\nz.mem_1624_sv2v_reg ,
  \nz.mem_1623_sv2v_reg ,\nz.mem_1622_sv2v_reg ,\nz.mem_1621_sv2v_reg ,\nz.mem_1620_sv2v_reg ,
  \nz.mem_1619_sv2v_reg ,\nz.mem_1618_sv2v_reg ,\nz.mem_1617_sv2v_reg ,
  \nz.mem_1616_sv2v_reg ,\nz.mem_1615_sv2v_reg ,\nz.mem_1614_sv2v_reg ,\nz.mem_1613_sv2v_reg ,
  \nz.mem_1612_sv2v_reg ,\nz.mem_1611_sv2v_reg ,\nz.mem_1610_sv2v_reg ,
  \nz.mem_1609_sv2v_reg ,\nz.mem_1608_sv2v_reg ,\nz.mem_1607_sv2v_reg ,\nz.mem_1606_sv2v_reg ,
  \nz.mem_1605_sv2v_reg ,\nz.mem_1604_sv2v_reg ,\nz.mem_1603_sv2v_reg ,
  \nz.mem_1602_sv2v_reg ,\nz.mem_1601_sv2v_reg ,\nz.mem_1600_sv2v_reg ,
  \nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,\nz.mem_1596_sv2v_reg ,
  \nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,\nz.mem_1593_sv2v_reg ,
  \nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,\nz.mem_1589_sv2v_reg ,
  \nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,\nz.mem_1586_sv2v_reg ,
  \nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,\nz.mem_1582_sv2v_reg ,
  \nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,\nz.mem_1579_sv2v_reg ,
  \nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,\nz.mem_1575_sv2v_reg ,
  \nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,\nz.mem_1572_sv2v_reg ,
  \nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,\nz.mem_1569_sv2v_reg ,\nz.mem_1568_sv2v_reg ,
  \nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,\nz.mem_1565_sv2v_reg ,
  \nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,\nz.mem_1562_sv2v_reg ,\nz.mem_1561_sv2v_reg ,
  \nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,\nz.mem_1558_sv2v_reg ,
  \nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,\nz.mem_1555_sv2v_reg ,\nz.mem_1554_sv2v_reg ,
  \nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,\nz.mem_1551_sv2v_reg ,
  \nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,\nz.mem_1548_sv2v_reg ,\nz.mem_1547_sv2v_reg ,
  \nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,\nz.mem_1544_sv2v_reg ,
  \nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,\nz.mem_1541_sv2v_reg ,\nz.mem_1540_sv2v_reg ,
  \nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,\nz.mem_1537_sv2v_reg ,
  \nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,\nz.mem_1534_sv2v_reg ,\nz.mem_1533_sv2v_reg ,
  \nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,\nz.mem_1530_sv2v_reg ,
  \nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,\nz.mem_1527_sv2v_reg ,\nz.mem_1526_sv2v_reg ,
  \nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,\nz.mem_1523_sv2v_reg ,
  \nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,\nz.mem_1520_sv2v_reg ,
  \nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,\nz.mem_1516_sv2v_reg ,
  \nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,\nz.mem_1513_sv2v_reg ,
  \nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,\nz.mem_1509_sv2v_reg ,
  \nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,\nz.mem_1506_sv2v_reg ,
  \nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,\nz.mem_1502_sv2v_reg ,
  \nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,\nz.mem_1499_sv2v_reg ,
  \nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,\nz.mem_1495_sv2v_reg ,
  \nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,\nz.mem_1492_sv2v_reg ,
  \nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,\nz.mem_1489_sv2v_reg ,\nz.mem_1488_sv2v_reg ,
  \nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,\nz.mem_1485_sv2v_reg ,
  \nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,\nz.mem_1482_sv2v_reg ,\nz.mem_1481_sv2v_reg ,
  \nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,\nz.mem_1478_sv2v_reg ,
  \nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,\nz.mem_1475_sv2v_reg ,\nz.mem_1474_sv2v_reg ,
  \nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,\nz.mem_1471_sv2v_reg ,
  \nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,\nz.mem_1468_sv2v_reg ,\nz.mem_1467_sv2v_reg ,
  \nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,\nz.mem_1464_sv2v_reg ,
  \nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,\nz.mem_1461_sv2v_reg ,\nz.mem_1460_sv2v_reg ,
  \nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,\nz.mem_1457_sv2v_reg ,
  \nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,\nz.mem_1454_sv2v_reg ,\nz.mem_1453_sv2v_reg ,
  \nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,\nz.mem_1450_sv2v_reg ,
  \nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,\nz.mem_1447_sv2v_reg ,\nz.mem_1446_sv2v_reg ,
  \nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,\nz.mem_1443_sv2v_reg ,
  \nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,\nz.mem_1440_sv2v_reg ,
  \nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,\nz.mem_1436_sv2v_reg ,
  \nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,\nz.mem_1433_sv2v_reg ,
  \nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,\nz.mem_1429_sv2v_reg ,
  \nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,\nz.mem_1426_sv2v_reg ,
  \nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,\nz.mem_1422_sv2v_reg ,
  \nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,\nz.mem_1419_sv2v_reg ,
  \nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,\nz.mem_1415_sv2v_reg ,
  \nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,\nz.mem_1412_sv2v_reg ,
  \nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,\nz.mem_1409_sv2v_reg ,\nz.mem_1408_sv2v_reg ,
  \nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,\nz.mem_1405_sv2v_reg ,
  \nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,\nz.mem_1402_sv2v_reg ,\nz.mem_1401_sv2v_reg ,
  \nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,\nz.mem_1398_sv2v_reg ,
  \nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,\nz.mem_1395_sv2v_reg ,\nz.mem_1394_sv2v_reg ,
  \nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,\nz.mem_1391_sv2v_reg ,
  \nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,\nz.mem_1388_sv2v_reg ,\nz.mem_1387_sv2v_reg ,
  \nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,\nz.mem_1384_sv2v_reg ,
  \nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,\nz.mem_1381_sv2v_reg ,\nz.mem_1380_sv2v_reg ,
  \nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,\nz.mem_1377_sv2v_reg ,
  \nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,\nz.mem_1374_sv2v_reg ,\nz.mem_1373_sv2v_reg ,
  \nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,\nz.mem_1370_sv2v_reg ,
  \nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,\nz.mem_1367_sv2v_reg ,\nz.mem_1366_sv2v_reg ,
  \nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,\nz.mem_1363_sv2v_reg ,
  \nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,\nz.mem_1360_sv2v_reg ,
  \nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,\nz.mem_1356_sv2v_reg ,
  \nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,\nz.mem_1353_sv2v_reg ,
  \nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,\nz.mem_1349_sv2v_reg ,
  \nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,\nz.mem_1346_sv2v_reg ,
  \nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,\nz.mem_1342_sv2v_reg ,
  \nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,\nz.mem_1339_sv2v_reg ,
  \nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,\nz.mem_1335_sv2v_reg ,
  \nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,\nz.mem_1332_sv2v_reg ,
  \nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,\nz.mem_1329_sv2v_reg ,\nz.mem_1328_sv2v_reg ,
  \nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,\nz.mem_1325_sv2v_reg ,
  \nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,\nz.mem_1322_sv2v_reg ,\nz.mem_1321_sv2v_reg ,
  \nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,\nz.mem_1318_sv2v_reg ,
  \nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,\nz.mem_1315_sv2v_reg ,\nz.mem_1314_sv2v_reg ,
  \nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,\nz.mem_1311_sv2v_reg ,
  \nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,\nz.mem_1308_sv2v_reg ,\nz.mem_1307_sv2v_reg ,
  \nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,\nz.mem_1304_sv2v_reg ,
  \nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,\nz.mem_1301_sv2v_reg ,\nz.mem_1300_sv2v_reg ,
  \nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,\nz.mem_1297_sv2v_reg ,
  \nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,\nz.mem_1294_sv2v_reg ,\nz.mem_1293_sv2v_reg ,
  \nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,\nz.mem_1290_sv2v_reg ,
  \nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,\nz.mem_1287_sv2v_reg ,\nz.mem_1286_sv2v_reg ,
  \nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,\nz.mem_1283_sv2v_reg ,
  \nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,\nz.mem_1280_sv2v_reg ,
  \nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,\nz.mem_1276_sv2v_reg ,
  \nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,\nz.mem_1273_sv2v_reg ,
  \nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,\nz.mem_1269_sv2v_reg ,
  \nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,\nz.mem_1266_sv2v_reg ,
  \nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,\nz.mem_1262_sv2v_reg ,
  \nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,\nz.mem_1259_sv2v_reg ,
  \nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,\nz.mem_1255_sv2v_reg ,
  \nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,\nz.mem_1252_sv2v_reg ,
  \nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,\nz.mem_1249_sv2v_reg ,\nz.mem_1248_sv2v_reg ,
  \nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,\nz.mem_1245_sv2v_reg ,
  \nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,\nz.mem_1242_sv2v_reg ,\nz.mem_1241_sv2v_reg ,
  \nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,\nz.mem_1238_sv2v_reg ,
  \nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,\nz.mem_1235_sv2v_reg ,\nz.mem_1234_sv2v_reg ,
  \nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,\nz.mem_1231_sv2v_reg ,
  \nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,\nz.mem_1228_sv2v_reg ,\nz.mem_1227_sv2v_reg ,
  \nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,\nz.mem_1224_sv2v_reg ,
  \nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,\nz.mem_1221_sv2v_reg ,\nz.mem_1220_sv2v_reg ,
  \nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,\nz.mem_1217_sv2v_reg ,
  \nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,\nz.mem_1214_sv2v_reg ,\nz.mem_1213_sv2v_reg ,
  \nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,\nz.mem_1210_sv2v_reg ,
  \nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,\nz.mem_1207_sv2v_reg ,\nz.mem_1206_sv2v_reg ,
  \nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,\nz.mem_1203_sv2v_reg ,
  \nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,\nz.mem_1200_sv2v_reg ,
  \nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,\nz.mem_1196_sv2v_reg ,
  \nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,\nz.mem_1193_sv2v_reg ,
  \nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,\nz.mem_1189_sv2v_reg ,
  \nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,\nz.mem_1186_sv2v_reg ,
  \nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,\nz.mem_1182_sv2v_reg ,
  \nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,\nz.mem_1179_sv2v_reg ,
  \nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,\nz.mem_1175_sv2v_reg ,
  \nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,\nz.mem_1172_sv2v_reg ,
  \nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,\nz.mem_1169_sv2v_reg ,\nz.mem_1168_sv2v_reg ,
  \nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,\nz.mem_1165_sv2v_reg ,
  \nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,\nz.mem_1162_sv2v_reg ,\nz.mem_1161_sv2v_reg ,
  \nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,\nz.mem_1158_sv2v_reg ,
  \nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,\nz.mem_1155_sv2v_reg ,\nz.mem_1154_sv2v_reg ,
  \nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,\nz.mem_1151_sv2v_reg ,
  \nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,\nz.mem_1148_sv2v_reg ,\nz.mem_1147_sv2v_reg ,
  \nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,\nz.mem_1144_sv2v_reg ,
  \nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,\nz.mem_1141_sv2v_reg ,\nz.mem_1140_sv2v_reg ,
  \nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,\nz.mem_1137_sv2v_reg ,
  \nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,\nz.mem_1134_sv2v_reg ,\nz.mem_1133_sv2v_reg ,
  \nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,\nz.mem_1130_sv2v_reg ,
  \nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,\nz.mem_1127_sv2v_reg ,\nz.mem_1126_sv2v_reg ,
  \nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,\nz.mem_1123_sv2v_reg ,
  \nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,\nz.mem_1120_sv2v_reg ,
  \nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,\nz.mem_1116_sv2v_reg ,
  \nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,\nz.mem_1113_sv2v_reg ,
  \nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,\nz.mem_1109_sv2v_reg ,
  \nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,\nz.mem_1106_sv2v_reg ,
  \nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,\nz.mem_1102_sv2v_reg ,
  \nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,\nz.mem_1099_sv2v_reg ,
  \nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,\nz.mem_1095_sv2v_reg ,
  \nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,\nz.mem_1092_sv2v_reg ,
  \nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,\nz.mem_1089_sv2v_reg ,\nz.mem_1088_sv2v_reg ,
  \nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,\nz.mem_1085_sv2v_reg ,
  \nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,\nz.mem_1082_sv2v_reg ,\nz.mem_1081_sv2v_reg ,
  \nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,\nz.mem_1078_sv2v_reg ,
  \nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,\nz.mem_1075_sv2v_reg ,\nz.mem_1074_sv2v_reg ,
  \nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,\nz.mem_1071_sv2v_reg ,
  \nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,\nz.mem_1068_sv2v_reg ,\nz.mem_1067_sv2v_reg ,
  \nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,\nz.mem_1064_sv2v_reg ,
  \nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,\nz.mem_1061_sv2v_reg ,\nz.mem_1060_sv2v_reg ,
  \nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,\nz.mem_1057_sv2v_reg ,
  \nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,\nz.mem_1054_sv2v_reg ,\nz.mem_1053_sv2v_reg ,
  \nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,\nz.mem_1050_sv2v_reg ,
  \nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,\nz.mem_1047_sv2v_reg ,\nz.mem_1046_sv2v_reg ,
  \nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,\nz.mem_1043_sv2v_reg ,
  \nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,\nz.mem_1040_sv2v_reg ,
  \nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,\nz.mem_1036_sv2v_reg ,
  \nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,\nz.mem_1033_sv2v_reg ,
  \nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,\nz.mem_1029_sv2v_reg ,
  \nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,\nz.mem_1026_sv2v_reg ,
  \nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,\nz.mem_1022_sv2v_reg ,
  \nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,\nz.mem_1019_sv2v_reg ,
  \nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,\nz.mem_1015_sv2v_reg ,
  \nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,\nz.mem_1012_sv2v_reg ,
  \nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,\nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,
  \nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,\nz.mem_1005_sv2v_reg ,
  \nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,\nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,
  \nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,\nz.mem_998_sv2v_reg ,
  \nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,\nz.mem_994_sv2v_reg ,
  \nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,\nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,
  \nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,\nz.mem_987_sv2v_reg ,
  \nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,\nz.mem_983_sv2v_reg ,
  \nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,\nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,
  \nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,\nz.mem_976_sv2v_reg ,
  \nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,\nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,
  \nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,\nz.mem_969_sv2v_reg ,
  \nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,\nz.mem_965_sv2v_reg ,
  \nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,\nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,
  \nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,\nz.mem_958_sv2v_reg ,
  \nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,\nz.mem_954_sv2v_reg ,
  \nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,\nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,
  \nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,\nz.mem_947_sv2v_reg ,
  \nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,\nz.mem_943_sv2v_reg ,
  \nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,\nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,
  \nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,\nz.mem_936_sv2v_reg ,
  \nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,\nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,
  \nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,\nz.mem_929_sv2v_reg ,
  \nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,\nz.mem_925_sv2v_reg ,
  \nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,\nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,
  \nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,\nz.mem_918_sv2v_reg ,
  \nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,\nz.mem_914_sv2v_reg ,
  \nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,\nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,
  \nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,\nz.mem_907_sv2v_reg ,
  \nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,\nz.mem_903_sv2v_reg ,
  \nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,\nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,
  \nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,\nz.mem_896_sv2v_reg ,
  \nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,\nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,
  \nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,\nz.mem_889_sv2v_reg ,
  \nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,\nz.mem_885_sv2v_reg ,
  \nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,\nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,
  \nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,\nz.mem_878_sv2v_reg ,
  \nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,\nz.mem_874_sv2v_reg ,
  \nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,\nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,
  \nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,\nz.mem_867_sv2v_reg ,
  \nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,\nz.mem_863_sv2v_reg ,
  \nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,\nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,
  \nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,\nz.mem_856_sv2v_reg ,
  \nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,\nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,
  \nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,\nz.mem_849_sv2v_reg ,
  \nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,\nz.mem_845_sv2v_reg ,
  \nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,\nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,
  \nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,\nz.mem_838_sv2v_reg ,
  \nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,\nz.mem_834_sv2v_reg ,
  \nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,\nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,
  \nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,\nz.mem_827_sv2v_reg ,
  \nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,\nz.mem_823_sv2v_reg ,
  \nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,\nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,
  \nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,\nz.mem_816_sv2v_reg ,
  \nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,\nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,
  \nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,\nz.mem_809_sv2v_reg ,
  \nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,\nz.mem_805_sv2v_reg ,
  \nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,\nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,
  \nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,\nz.mem_798_sv2v_reg ,
  \nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,\nz.mem_794_sv2v_reg ,
  \nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,\nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,
  \nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,\nz.mem_787_sv2v_reg ,
  \nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,\nz.mem_783_sv2v_reg ,
  \nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,\nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,
  \nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,\nz.mem_776_sv2v_reg ,
  \nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,\nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,
  \nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,\nz.mem_769_sv2v_reg ,
  \nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,\nz.mem_765_sv2v_reg ,
  \nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,\nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,
  \nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,\nz.mem_758_sv2v_reg ,
  \nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,\nz.mem_754_sv2v_reg ,
  \nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,\nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,
  \nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,\nz.mem_747_sv2v_reg ,
  \nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,\nz.mem_743_sv2v_reg ,
  \nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,\nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,
  \nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,\nz.mem_736_sv2v_reg ,
  \nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,\nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,
  \nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,\nz.mem_729_sv2v_reg ,
  \nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,\nz.mem_725_sv2v_reg ,
  \nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,\nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,
  \nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,\nz.mem_718_sv2v_reg ,
  \nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,\nz.mem_714_sv2v_reg ,
  \nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,\nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,
  \nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,\nz.mem_707_sv2v_reg ,
  \nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,\nz.mem_703_sv2v_reg ,
  \nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,\nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,
  \nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,\nz.mem_696_sv2v_reg ,
  \nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,\nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,
  \nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,\nz.mem_689_sv2v_reg ,
  \nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,\nz.mem_685_sv2v_reg ,
  \nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,
  \nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,\nz.mem_678_sv2v_reg ,
  \nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,\nz.mem_674_sv2v_reg ,
  \nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,
  \nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,\nz.mem_667_sv2v_reg ,
  \nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,\nz.mem_663_sv2v_reg ,
  \nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,
  \nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,\nz.mem_656_sv2v_reg ,
  \nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,
  \nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,\nz.mem_649_sv2v_reg ,
  \nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,\nz.mem_645_sv2v_reg ,
  \nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,
  \nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,\nz.mem_638_sv2v_reg ,
  \nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,\nz.mem_634_sv2v_reg ,
  \nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,
  \nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,\nz.mem_627_sv2v_reg ,
  \nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,\nz.mem_623_sv2v_reg ,
  \nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,
  \nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,\nz.mem_616_sv2v_reg ,
  \nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,
  \nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,\nz.mem_609_sv2v_reg ,
  \nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,\nz.mem_605_sv2v_reg ,
  \nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,
  \nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,\nz.mem_598_sv2v_reg ,
  \nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,\nz.mem_594_sv2v_reg ,
  \nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,
  \nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,\nz.mem_587_sv2v_reg ,
  \nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,\nz.mem_583_sv2v_reg ,
  \nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,
  \nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,\nz.mem_576_sv2v_reg ,
  \nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,
  \nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,\nz.mem_569_sv2v_reg ,
  \nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,\nz.mem_565_sv2v_reg ,
  \nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,
  \nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,\nz.mem_558_sv2v_reg ,
  \nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,\nz.mem_554_sv2v_reg ,
  \nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,
  \nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,\nz.mem_547_sv2v_reg ,
  \nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,\nz.mem_543_sv2v_reg ,
  \nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,
  \nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,\nz.mem_536_sv2v_reg ,
  \nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,
  \nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,\nz.mem_529_sv2v_reg ,
  \nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,\nz.mem_525_sv2v_reg ,
  \nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,
  \nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,\nz.mem_518_sv2v_reg ,
  \nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,\nz.mem_514_sv2v_reg ,
  \nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,
  \nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,\nz.mem_507_sv2v_reg ,
  \nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,\nz.mem_503_sv2v_reg ,
  \nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,
  \nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,\nz.mem_496_sv2v_reg ,
  \nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,
  \nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,\nz.mem_489_sv2v_reg ,
  \nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,\nz.mem_485_sv2v_reg ,
  \nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,
  \nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,\nz.mem_478_sv2v_reg ,
  \nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,\nz.mem_474_sv2v_reg ,
  \nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,
  \nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,\nz.mem_467_sv2v_reg ,
  \nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,\nz.mem_463_sv2v_reg ,
  \nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,
  \nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,\nz.mem_456_sv2v_reg ,
  \nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,
  \nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,\nz.mem_449_sv2v_reg ,
  \nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,\nz.mem_445_sv2v_reg ,
  \nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,
  \nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,\nz.mem_438_sv2v_reg ,
  \nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,\nz.mem_434_sv2v_reg ,
  \nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,
  \nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,\nz.mem_427_sv2v_reg ,
  \nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,\nz.mem_423_sv2v_reg ,
  \nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,
  \nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,\nz.mem_416_sv2v_reg ,
  \nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,
  \nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,\nz.mem_409_sv2v_reg ,
  \nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,\nz.mem_405_sv2v_reg ,
  \nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,
  \nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,\nz.mem_398_sv2v_reg ,
  \nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,\nz.mem_394_sv2v_reg ,
  \nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,
  \nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,\nz.mem_387_sv2v_reg ,
  \nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,\nz.mem_383_sv2v_reg ,
  \nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,
  \nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,\nz.mem_376_sv2v_reg ,
  \nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,
  \nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,\nz.mem_369_sv2v_reg ,
  \nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,\nz.mem_365_sv2v_reg ,
  \nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,
  \nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,\nz.mem_358_sv2v_reg ,
  \nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,\nz.mem_354_sv2v_reg ,
  \nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,
  \nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,\nz.mem_347_sv2v_reg ,
  \nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,\nz.mem_343_sv2v_reg ,
  \nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,
  \nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,\nz.mem_336_sv2v_reg ,
  \nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,
  \nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,\nz.mem_329_sv2v_reg ,
  \nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,\nz.mem_325_sv2v_reg ,
  \nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,
  \nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,\nz.mem_318_sv2v_reg ,
  \nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,\nz.mem_314_sv2v_reg ,
  \nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,
  \nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,\nz.mem_307_sv2v_reg ,
  \nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,\nz.mem_303_sv2v_reg ,
  \nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,
  \nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,\nz.mem_296_sv2v_reg ,
  \nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,
  \nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,\nz.mem_289_sv2v_reg ,
  \nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,\nz.mem_285_sv2v_reg ,
  \nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,
  \nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,\nz.mem_278_sv2v_reg ,
  \nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,\nz.mem_274_sv2v_reg ,
  \nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,
  \nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,\nz.mem_267_sv2v_reg ,
  \nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,\nz.mem_263_sv2v_reg ,
  \nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,
  \nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,\nz.mem_256_sv2v_reg ,
  \nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,
  \nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,\nz.mem_249_sv2v_reg ,
  \nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,\nz.mem_245_sv2v_reg ,
  \nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,
  \nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,\nz.mem_238_sv2v_reg ,
  \nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,\nz.mem_234_sv2v_reg ,
  \nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,
  \nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,\nz.mem_227_sv2v_reg ,
  \nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,\nz.mem_223_sv2v_reg ,
  \nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,
  \nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,\nz.mem_216_sv2v_reg ,
  \nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,
  \nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,\nz.mem_209_sv2v_reg ,
  \nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,\nz.mem_205_sv2v_reg ,
  \nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,
  \nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,\nz.mem_198_sv2v_reg ,
  \nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,\nz.mem_194_sv2v_reg ,
  \nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,
  \nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,\nz.mem_187_sv2v_reg ,
  \nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,\nz.mem_183_sv2v_reg ,
  \nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,
  \nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,\nz.mem_176_sv2v_reg ,
  \nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,
  \nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,\nz.mem_169_sv2v_reg ,
  \nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,\nz.mem_165_sv2v_reg ,
  \nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,
  \nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,\nz.mem_158_sv2v_reg ,
  \nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,\nz.mem_154_sv2v_reg ,
  \nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,
  \nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,\nz.mem_147_sv2v_reg ,
  \nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,\nz.mem_143_sv2v_reg ,
  \nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,
  \nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,\nz.mem_136_sv2v_reg ,
  \nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,
  \nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,\nz.mem_129_sv2v_reg ,
  \nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,
  \nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,
  \nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,
  \nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,
  \nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [2559] = \nz.mem_2559_sv2v_reg ;
  assign \nz.mem [2558] = \nz.mem_2558_sv2v_reg ;
  assign \nz.mem [2557] = \nz.mem_2557_sv2v_reg ;
  assign \nz.mem [2556] = \nz.mem_2556_sv2v_reg ;
  assign \nz.mem [2555] = \nz.mem_2555_sv2v_reg ;
  assign \nz.mem [2554] = \nz.mem_2554_sv2v_reg ;
  assign \nz.mem [2553] = \nz.mem_2553_sv2v_reg ;
  assign \nz.mem [2552] = \nz.mem_2552_sv2v_reg ;
  assign \nz.mem [2551] = \nz.mem_2551_sv2v_reg ;
  assign \nz.mem [2550] = \nz.mem_2550_sv2v_reg ;
  assign \nz.mem [2549] = \nz.mem_2549_sv2v_reg ;
  assign \nz.mem [2548] = \nz.mem_2548_sv2v_reg ;
  assign \nz.mem [2547] = \nz.mem_2547_sv2v_reg ;
  assign \nz.mem [2546] = \nz.mem_2546_sv2v_reg ;
  assign \nz.mem [2545] = \nz.mem_2545_sv2v_reg ;
  assign \nz.mem [2544] = \nz.mem_2544_sv2v_reg ;
  assign \nz.mem [2543] = \nz.mem_2543_sv2v_reg ;
  assign \nz.mem [2542] = \nz.mem_2542_sv2v_reg ;
  assign \nz.mem [2541] = \nz.mem_2541_sv2v_reg ;
  assign \nz.mem [2540] = \nz.mem_2540_sv2v_reg ;
  assign \nz.mem [2539] = \nz.mem_2539_sv2v_reg ;
  assign \nz.mem [2538] = \nz.mem_2538_sv2v_reg ;
  assign \nz.mem [2537] = \nz.mem_2537_sv2v_reg ;
  assign \nz.mem [2536] = \nz.mem_2536_sv2v_reg ;
  assign \nz.mem [2535] = \nz.mem_2535_sv2v_reg ;
  assign \nz.mem [2534] = \nz.mem_2534_sv2v_reg ;
  assign \nz.mem [2533] = \nz.mem_2533_sv2v_reg ;
  assign \nz.mem [2532] = \nz.mem_2532_sv2v_reg ;
  assign \nz.mem [2531] = \nz.mem_2531_sv2v_reg ;
  assign \nz.mem [2530] = \nz.mem_2530_sv2v_reg ;
  assign \nz.mem [2529] = \nz.mem_2529_sv2v_reg ;
  assign \nz.mem [2528] = \nz.mem_2528_sv2v_reg ;
  assign \nz.mem [2527] = \nz.mem_2527_sv2v_reg ;
  assign \nz.mem [2526] = \nz.mem_2526_sv2v_reg ;
  assign \nz.mem [2525] = \nz.mem_2525_sv2v_reg ;
  assign \nz.mem [2524] = \nz.mem_2524_sv2v_reg ;
  assign \nz.mem [2523] = \nz.mem_2523_sv2v_reg ;
  assign \nz.mem [2522] = \nz.mem_2522_sv2v_reg ;
  assign \nz.mem [2521] = \nz.mem_2521_sv2v_reg ;
  assign \nz.mem [2520] = \nz.mem_2520_sv2v_reg ;
  assign \nz.mem [2519] = \nz.mem_2519_sv2v_reg ;
  assign \nz.mem [2518] = \nz.mem_2518_sv2v_reg ;
  assign \nz.mem [2517] = \nz.mem_2517_sv2v_reg ;
  assign \nz.mem [2516] = \nz.mem_2516_sv2v_reg ;
  assign \nz.mem [2515] = \nz.mem_2515_sv2v_reg ;
  assign \nz.mem [2514] = \nz.mem_2514_sv2v_reg ;
  assign \nz.mem [2513] = \nz.mem_2513_sv2v_reg ;
  assign \nz.mem [2512] = \nz.mem_2512_sv2v_reg ;
  assign \nz.mem [2511] = \nz.mem_2511_sv2v_reg ;
  assign \nz.mem [2510] = \nz.mem_2510_sv2v_reg ;
  assign \nz.mem [2509] = \nz.mem_2509_sv2v_reg ;
  assign \nz.mem [2508] = \nz.mem_2508_sv2v_reg ;
  assign \nz.mem [2507] = \nz.mem_2507_sv2v_reg ;
  assign \nz.mem [2506] = \nz.mem_2506_sv2v_reg ;
  assign \nz.mem [2505] = \nz.mem_2505_sv2v_reg ;
  assign \nz.mem [2504] = \nz.mem_2504_sv2v_reg ;
  assign \nz.mem [2503] = \nz.mem_2503_sv2v_reg ;
  assign \nz.mem [2502] = \nz.mem_2502_sv2v_reg ;
  assign \nz.mem [2501] = \nz.mem_2501_sv2v_reg ;
  assign \nz.mem [2500] = \nz.mem_2500_sv2v_reg ;
  assign \nz.mem [2499] = \nz.mem_2499_sv2v_reg ;
  assign \nz.mem [2498] = \nz.mem_2498_sv2v_reg ;
  assign \nz.mem [2497] = \nz.mem_2497_sv2v_reg ;
  assign \nz.mem [2496] = \nz.mem_2496_sv2v_reg ;
  assign \nz.mem [2495] = \nz.mem_2495_sv2v_reg ;
  assign \nz.mem [2494] = \nz.mem_2494_sv2v_reg ;
  assign \nz.mem [2493] = \nz.mem_2493_sv2v_reg ;
  assign \nz.mem [2492] = \nz.mem_2492_sv2v_reg ;
  assign \nz.mem [2491] = \nz.mem_2491_sv2v_reg ;
  assign \nz.mem [2490] = \nz.mem_2490_sv2v_reg ;
  assign \nz.mem [2489] = \nz.mem_2489_sv2v_reg ;
  assign \nz.mem [2488] = \nz.mem_2488_sv2v_reg ;
  assign \nz.mem [2487] = \nz.mem_2487_sv2v_reg ;
  assign \nz.mem [2486] = \nz.mem_2486_sv2v_reg ;
  assign \nz.mem [2485] = \nz.mem_2485_sv2v_reg ;
  assign \nz.mem [2484] = \nz.mem_2484_sv2v_reg ;
  assign \nz.mem [2483] = \nz.mem_2483_sv2v_reg ;
  assign \nz.mem [2482] = \nz.mem_2482_sv2v_reg ;
  assign \nz.mem [2481] = \nz.mem_2481_sv2v_reg ;
  assign \nz.mem [2480] = \nz.mem_2480_sv2v_reg ;
  assign \nz.mem [2479] = \nz.mem_2479_sv2v_reg ;
  assign \nz.mem [2478] = \nz.mem_2478_sv2v_reg ;
  assign \nz.mem [2477] = \nz.mem_2477_sv2v_reg ;
  assign \nz.mem [2476] = \nz.mem_2476_sv2v_reg ;
  assign \nz.mem [2475] = \nz.mem_2475_sv2v_reg ;
  assign \nz.mem [2474] = \nz.mem_2474_sv2v_reg ;
  assign \nz.mem [2473] = \nz.mem_2473_sv2v_reg ;
  assign \nz.mem [2472] = \nz.mem_2472_sv2v_reg ;
  assign \nz.mem [2471] = \nz.mem_2471_sv2v_reg ;
  assign \nz.mem [2470] = \nz.mem_2470_sv2v_reg ;
  assign \nz.mem [2469] = \nz.mem_2469_sv2v_reg ;
  assign \nz.mem [2468] = \nz.mem_2468_sv2v_reg ;
  assign \nz.mem [2467] = \nz.mem_2467_sv2v_reg ;
  assign \nz.mem [2466] = \nz.mem_2466_sv2v_reg ;
  assign \nz.mem [2465] = \nz.mem_2465_sv2v_reg ;
  assign \nz.mem [2464] = \nz.mem_2464_sv2v_reg ;
  assign \nz.mem [2463] = \nz.mem_2463_sv2v_reg ;
  assign \nz.mem [2462] = \nz.mem_2462_sv2v_reg ;
  assign \nz.mem [2461] = \nz.mem_2461_sv2v_reg ;
  assign \nz.mem [2460] = \nz.mem_2460_sv2v_reg ;
  assign \nz.mem [2459] = \nz.mem_2459_sv2v_reg ;
  assign \nz.mem [2458] = \nz.mem_2458_sv2v_reg ;
  assign \nz.mem [2457] = \nz.mem_2457_sv2v_reg ;
  assign \nz.mem [2456] = \nz.mem_2456_sv2v_reg ;
  assign \nz.mem [2455] = \nz.mem_2455_sv2v_reg ;
  assign \nz.mem [2454] = \nz.mem_2454_sv2v_reg ;
  assign \nz.mem [2453] = \nz.mem_2453_sv2v_reg ;
  assign \nz.mem [2452] = \nz.mem_2452_sv2v_reg ;
  assign \nz.mem [2451] = \nz.mem_2451_sv2v_reg ;
  assign \nz.mem [2450] = \nz.mem_2450_sv2v_reg ;
  assign \nz.mem [2449] = \nz.mem_2449_sv2v_reg ;
  assign \nz.mem [2448] = \nz.mem_2448_sv2v_reg ;
  assign \nz.mem [2447] = \nz.mem_2447_sv2v_reg ;
  assign \nz.mem [2446] = \nz.mem_2446_sv2v_reg ;
  assign \nz.mem [2445] = \nz.mem_2445_sv2v_reg ;
  assign \nz.mem [2444] = \nz.mem_2444_sv2v_reg ;
  assign \nz.mem [2443] = \nz.mem_2443_sv2v_reg ;
  assign \nz.mem [2442] = \nz.mem_2442_sv2v_reg ;
  assign \nz.mem [2441] = \nz.mem_2441_sv2v_reg ;
  assign \nz.mem [2440] = \nz.mem_2440_sv2v_reg ;
  assign \nz.mem [2439] = \nz.mem_2439_sv2v_reg ;
  assign \nz.mem [2438] = \nz.mem_2438_sv2v_reg ;
  assign \nz.mem [2437] = \nz.mem_2437_sv2v_reg ;
  assign \nz.mem [2436] = \nz.mem_2436_sv2v_reg ;
  assign \nz.mem [2435] = \nz.mem_2435_sv2v_reg ;
  assign \nz.mem [2434] = \nz.mem_2434_sv2v_reg ;
  assign \nz.mem [2433] = \nz.mem_2433_sv2v_reg ;
  assign \nz.mem [2432] = \nz.mem_2432_sv2v_reg ;
  assign \nz.mem [2431] = \nz.mem_2431_sv2v_reg ;
  assign \nz.mem [2430] = \nz.mem_2430_sv2v_reg ;
  assign \nz.mem [2429] = \nz.mem_2429_sv2v_reg ;
  assign \nz.mem [2428] = \nz.mem_2428_sv2v_reg ;
  assign \nz.mem [2427] = \nz.mem_2427_sv2v_reg ;
  assign \nz.mem [2426] = \nz.mem_2426_sv2v_reg ;
  assign \nz.mem [2425] = \nz.mem_2425_sv2v_reg ;
  assign \nz.mem [2424] = \nz.mem_2424_sv2v_reg ;
  assign \nz.mem [2423] = \nz.mem_2423_sv2v_reg ;
  assign \nz.mem [2422] = \nz.mem_2422_sv2v_reg ;
  assign \nz.mem [2421] = \nz.mem_2421_sv2v_reg ;
  assign \nz.mem [2420] = \nz.mem_2420_sv2v_reg ;
  assign \nz.mem [2419] = \nz.mem_2419_sv2v_reg ;
  assign \nz.mem [2418] = \nz.mem_2418_sv2v_reg ;
  assign \nz.mem [2417] = \nz.mem_2417_sv2v_reg ;
  assign \nz.mem [2416] = \nz.mem_2416_sv2v_reg ;
  assign \nz.mem [2415] = \nz.mem_2415_sv2v_reg ;
  assign \nz.mem [2414] = \nz.mem_2414_sv2v_reg ;
  assign \nz.mem [2413] = \nz.mem_2413_sv2v_reg ;
  assign \nz.mem [2412] = \nz.mem_2412_sv2v_reg ;
  assign \nz.mem [2411] = \nz.mem_2411_sv2v_reg ;
  assign \nz.mem [2410] = \nz.mem_2410_sv2v_reg ;
  assign \nz.mem [2409] = \nz.mem_2409_sv2v_reg ;
  assign \nz.mem [2408] = \nz.mem_2408_sv2v_reg ;
  assign \nz.mem [2407] = \nz.mem_2407_sv2v_reg ;
  assign \nz.mem [2406] = \nz.mem_2406_sv2v_reg ;
  assign \nz.mem [2405] = \nz.mem_2405_sv2v_reg ;
  assign \nz.mem [2404] = \nz.mem_2404_sv2v_reg ;
  assign \nz.mem [2403] = \nz.mem_2403_sv2v_reg ;
  assign \nz.mem [2402] = \nz.mem_2402_sv2v_reg ;
  assign \nz.mem [2401] = \nz.mem_2401_sv2v_reg ;
  assign \nz.mem [2400] = \nz.mem_2400_sv2v_reg ;
  assign \nz.mem [2399] = \nz.mem_2399_sv2v_reg ;
  assign \nz.mem [2398] = \nz.mem_2398_sv2v_reg ;
  assign \nz.mem [2397] = \nz.mem_2397_sv2v_reg ;
  assign \nz.mem [2396] = \nz.mem_2396_sv2v_reg ;
  assign \nz.mem [2395] = \nz.mem_2395_sv2v_reg ;
  assign \nz.mem [2394] = \nz.mem_2394_sv2v_reg ;
  assign \nz.mem [2393] = \nz.mem_2393_sv2v_reg ;
  assign \nz.mem [2392] = \nz.mem_2392_sv2v_reg ;
  assign \nz.mem [2391] = \nz.mem_2391_sv2v_reg ;
  assign \nz.mem [2390] = \nz.mem_2390_sv2v_reg ;
  assign \nz.mem [2389] = \nz.mem_2389_sv2v_reg ;
  assign \nz.mem [2388] = \nz.mem_2388_sv2v_reg ;
  assign \nz.mem [2387] = \nz.mem_2387_sv2v_reg ;
  assign \nz.mem [2386] = \nz.mem_2386_sv2v_reg ;
  assign \nz.mem [2385] = \nz.mem_2385_sv2v_reg ;
  assign \nz.mem [2384] = \nz.mem_2384_sv2v_reg ;
  assign \nz.mem [2383] = \nz.mem_2383_sv2v_reg ;
  assign \nz.mem [2382] = \nz.mem_2382_sv2v_reg ;
  assign \nz.mem [2381] = \nz.mem_2381_sv2v_reg ;
  assign \nz.mem [2380] = \nz.mem_2380_sv2v_reg ;
  assign \nz.mem [2379] = \nz.mem_2379_sv2v_reg ;
  assign \nz.mem [2378] = \nz.mem_2378_sv2v_reg ;
  assign \nz.mem [2377] = \nz.mem_2377_sv2v_reg ;
  assign \nz.mem [2376] = \nz.mem_2376_sv2v_reg ;
  assign \nz.mem [2375] = \nz.mem_2375_sv2v_reg ;
  assign \nz.mem [2374] = \nz.mem_2374_sv2v_reg ;
  assign \nz.mem [2373] = \nz.mem_2373_sv2v_reg ;
  assign \nz.mem [2372] = \nz.mem_2372_sv2v_reg ;
  assign \nz.mem [2371] = \nz.mem_2371_sv2v_reg ;
  assign \nz.mem [2370] = \nz.mem_2370_sv2v_reg ;
  assign \nz.mem [2369] = \nz.mem_2369_sv2v_reg ;
  assign \nz.mem [2368] = \nz.mem_2368_sv2v_reg ;
  assign \nz.mem [2367] = \nz.mem_2367_sv2v_reg ;
  assign \nz.mem [2366] = \nz.mem_2366_sv2v_reg ;
  assign \nz.mem [2365] = \nz.mem_2365_sv2v_reg ;
  assign \nz.mem [2364] = \nz.mem_2364_sv2v_reg ;
  assign \nz.mem [2363] = \nz.mem_2363_sv2v_reg ;
  assign \nz.mem [2362] = \nz.mem_2362_sv2v_reg ;
  assign \nz.mem [2361] = \nz.mem_2361_sv2v_reg ;
  assign \nz.mem [2360] = \nz.mem_2360_sv2v_reg ;
  assign \nz.mem [2359] = \nz.mem_2359_sv2v_reg ;
  assign \nz.mem [2358] = \nz.mem_2358_sv2v_reg ;
  assign \nz.mem [2357] = \nz.mem_2357_sv2v_reg ;
  assign \nz.mem [2356] = \nz.mem_2356_sv2v_reg ;
  assign \nz.mem [2355] = \nz.mem_2355_sv2v_reg ;
  assign \nz.mem [2354] = \nz.mem_2354_sv2v_reg ;
  assign \nz.mem [2353] = \nz.mem_2353_sv2v_reg ;
  assign \nz.mem [2352] = \nz.mem_2352_sv2v_reg ;
  assign \nz.mem [2351] = \nz.mem_2351_sv2v_reg ;
  assign \nz.mem [2350] = \nz.mem_2350_sv2v_reg ;
  assign \nz.mem [2349] = \nz.mem_2349_sv2v_reg ;
  assign \nz.mem [2348] = \nz.mem_2348_sv2v_reg ;
  assign \nz.mem [2347] = \nz.mem_2347_sv2v_reg ;
  assign \nz.mem [2346] = \nz.mem_2346_sv2v_reg ;
  assign \nz.mem [2345] = \nz.mem_2345_sv2v_reg ;
  assign \nz.mem [2344] = \nz.mem_2344_sv2v_reg ;
  assign \nz.mem [2343] = \nz.mem_2343_sv2v_reg ;
  assign \nz.mem [2342] = \nz.mem_2342_sv2v_reg ;
  assign \nz.mem [2341] = \nz.mem_2341_sv2v_reg ;
  assign \nz.mem [2340] = \nz.mem_2340_sv2v_reg ;
  assign \nz.mem [2339] = \nz.mem_2339_sv2v_reg ;
  assign \nz.mem [2338] = \nz.mem_2338_sv2v_reg ;
  assign \nz.mem [2337] = \nz.mem_2337_sv2v_reg ;
  assign \nz.mem [2336] = \nz.mem_2336_sv2v_reg ;
  assign \nz.mem [2335] = \nz.mem_2335_sv2v_reg ;
  assign \nz.mem [2334] = \nz.mem_2334_sv2v_reg ;
  assign \nz.mem [2333] = \nz.mem_2333_sv2v_reg ;
  assign \nz.mem [2332] = \nz.mem_2332_sv2v_reg ;
  assign \nz.mem [2331] = \nz.mem_2331_sv2v_reg ;
  assign \nz.mem [2330] = \nz.mem_2330_sv2v_reg ;
  assign \nz.mem [2329] = \nz.mem_2329_sv2v_reg ;
  assign \nz.mem [2328] = \nz.mem_2328_sv2v_reg ;
  assign \nz.mem [2327] = \nz.mem_2327_sv2v_reg ;
  assign \nz.mem [2326] = \nz.mem_2326_sv2v_reg ;
  assign \nz.mem [2325] = \nz.mem_2325_sv2v_reg ;
  assign \nz.mem [2324] = \nz.mem_2324_sv2v_reg ;
  assign \nz.mem [2323] = \nz.mem_2323_sv2v_reg ;
  assign \nz.mem [2322] = \nz.mem_2322_sv2v_reg ;
  assign \nz.mem [2321] = \nz.mem_2321_sv2v_reg ;
  assign \nz.mem [2320] = \nz.mem_2320_sv2v_reg ;
  assign \nz.mem [2319] = \nz.mem_2319_sv2v_reg ;
  assign \nz.mem [2318] = \nz.mem_2318_sv2v_reg ;
  assign \nz.mem [2317] = \nz.mem_2317_sv2v_reg ;
  assign \nz.mem [2316] = \nz.mem_2316_sv2v_reg ;
  assign \nz.mem [2315] = \nz.mem_2315_sv2v_reg ;
  assign \nz.mem [2314] = \nz.mem_2314_sv2v_reg ;
  assign \nz.mem [2313] = \nz.mem_2313_sv2v_reg ;
  assign \nz.mem [2312] = \nz.mem_2312_sv2v_reg ;
  assign \nz.mem [2311] = \nz.mem_2311_sv2v_reg ;
  assign \nz.mem [2310] = \nz.mem_2310_sv2v_reg ;
  assign \nz.mem [2309] = \nz.mem_2309_sv2v_reg ;
  assign \nz.mem [2308] = \nz.mem_2308_sv2v_reg ;
  assign \nz.mem [2307] = \nz.mem_2307_sv2v_reg ;
  assign \nz.mem [2306] = \nz.mem_2306_sv2v_reg ;
  assign \nz.mem [2305] = \nz.mem_2305_sv2v_reg ;
  assign \nz.mem [2304] = \nz.mem_2304_sv2v_reg ;
  assign \nz.mem [2303] = \nz.mem_2303_sv2v_reg ;
  assign \nz.mem [2302] = \nz.mem_2302_sv2v_reg ;
  assign \nz.mem [2301] = \nz.mem_2301_sv2v_reg ;
  assign \nz.mem [2300] = \nz.mem_2300_sv2v_reg ;
  assign \nz.mem [2299] = \nz.mem_2299_sv2v_reg ;
  assign \nz.mem [2298] = \nz.mem_2298_sv2v_reg ;
  assign \nz.mem [2297] = \nz.mem_2297_sv2v_reg ;
  assign \nz.mem [2296] = \nz.mem_2296_sv2v_reg ;
  assign \nz.mem [2295] = \nz.mem_2295_sv2v_reg ;
  assign \nz.mem [2294] = \nz.mem_2294_sv2v_reg ;
  assign \nz.mem [2293] = \nz.mem_2293_sv2v_reg ;
  assign \nz.mem [2292] = \nz.mem_2292_sv2v_reg ;
  assign \nz.mem [2291] = \nz.mem_2291_sv2v_reg ;
  assign \nz.mem [2290] = \nz.mem_2290_sv2v_reg ;
  assign \nz.mem [2289] = \nz.mem_2289_sv2v_reg ;
  assign \nz.mem [2288] = \nz.mem_2288_sv2v_reg ;
  assign \nz.mem [2287] = \nz.mem_2287_sv2v_reg ;
  assign \nz.mem [2286] = \nz.mem_2286_sv2v_reg ;
  assign \nz.mem [2285] = \nz.mem_2285_sv2v_reg ;
  assign \nz.mem [2284] = \nz.mem_2284_sv2v_reg ;
  assign \nz.mem [2283] = \nz.mem_2283_sv2v_reg ;
  assign \nz.mem [2282] = \nz.mem_2282_sv2v_reg ;
  assign \nz.mem [2281] = \nz.mem_2281_sv2v_reg ;
  assign \nz.mem [2280] = \nz.mem_2280_sv2v_reg ;
  assign \nz.mem [2279] = \nz.mem_2279_sv2v_reg ;
  assign \nz.mem [2278] = \nz.mem_2278_sv2v_reg ;
  assign \nz.mem [2277] = \nz.mem_2277_sv2v_reg ;
  assign \nz.mem [2276] = \nz.mem_2276_sv2v_reg ;
  assign \nz.mem [2275] = \nz.mem_2275_sv2v_reg ;
  assign \nz.mem [2274] = \nz.mem_2274_sv2v_reg ;
  assign \nz.mem [2273] = \nz.mem_2273_sv2v_reg ;
  assign \nz.mem [2272] = \nz.mem_2272_sv2v_reg ;
  assign \nz.mem [2271] = \nz.mem_2271_sv2v_reg ;
  assign \nz.mem [2270] = \nz.mem_2270_sv2v_reg ;
  assign \nz.mem [2269] = \nz.mem_2269_sv2v_reg ;
  assign \nz.mem [2268] = \nz.mem_2268_sv2v_reg ;
  assign \nz.mem [2267] = \nz.mem_2267_sv2v_reg ;
  assign \nz.mem [2266] = \nz.mem_2266_sv2v_reg ;
  assign \nz.mem [2265] = \nz.mem_2265_sv2v_reg ;
  assign \nz.mem [2264] = \nz.mem_2264_sv2v_reg ;
  assign \nz.mem [2263] = \nz.mem_2263_sv2v_reg ;
  assign \nz.mem [2262] = \nz.mem_2262_sv2v_reg ;
  assign \nz.mem [2261] = \nz.mem_2261_sv2v_reg ;
  assign \nz.mem [2260] = \nz.mem_2260_sv2v_reg ;
  assign \nz.mem [2259] = \nz.mem_2259_sv2v_reg ;
  assign \nz.mem [2258] = \nz.mem_2258_sv2v_reg ;
  assign \nz.mem [2257] = \nz.mem_2257_sv2v_reg ;
  assign \nz.mem [2256] = \nz.mem_2256_sv2v_reg ;
  assign \nz.mem [2255] = \nz.mem_2255_sv2v_reg ;
  assign \nz.mem [2254] = \nz.mem_2254_sv2v_reg ;
  assign \nz.mem [2253] = \nz.mem_2253_sv2v_reg ;
  assign \nz.mem [2252] = \nz.mem_2252_sv2v_reg ;
  assign \nz.mem [2251] = \nz.mem_2251_sv2v_reg ;
  assign \nz.mem [2250] = \nz.mem_2250_sv2v_reg ;
  assign \nz.mem [2249] = \nz.mem_2249_sv2v_reg ;
  assign \nz.mem [2248] = \nz.mem_2248_sv2v_reg ;
  assign \nz.mem [2247] = \nz.mem_2247_sv2v_reg ;
  assign \nz.mem [2246] = \nz.mem_2246_sv2v_reg ;
  assign \nz.mem [2245] = \nz.mem_2245_sv2v_reg ;
  assign \nz.mem [2244] = \nz.mem_2244_sv2v_reg ;
  assign \nz.mem [2243] = \nz.mem_2243_sv2v_reg ;
  assign \nz.mem [2242] = \nz.mem_2242_sv2v_reg ;
  assign \nz.mem [2241] = \nz.mem_2241_sv2v_reg ;
  assign \nz.mem [2240] = \nz.mem_2240_sv2v_reg ;
  assign \nz.mem [2239] = \nz.mem_2239_sv2v_reg ;
  assign \nz.mem [2238] = \nz.mem_2238_sv2v_reg ;
  assign \nz.mem [2237] = \nz.mem_2237_sv2v_reg ;
  assign \nz.mem [2236] = \nz.mem_2236_sv2v_reg ;
  assign \nz.mem [2235] = \nz.mem_2235_sv2v_reg ;
  assign \nz.mem [2234] = \nz.mem_2234_sv2v_reg ;
  assign \nz.mem [2233] = \nz.mem_2233_sv2v_reg ;
  assign \nz.mem [2232] = \nz.mem_2232_sv2v_reg ;
  assign \nz.mem [2231] = \nz.mem_2231_sv2v_reg ;
  assign \nz.mem [2230] = \nz.mem_2230_sv2v_reg ;
  assign \nz.mem [2229] = \nz.mem_2229_sv2v_reg ;
  assign \nz.mem [2228] = \nz.mem_2228_sv2v_reg ;
  assign \nz.mem [2227] = \nz.mem_2227_sv2v_reg ;
  assign \nz.mem [2226] = \nz.mem_2226_sv2v_reg ;
  assign \nz.mem [2225] = \nz.mem_2225_sv2v_reg ;
  assign \nz.mem [2224] = \nz.mem_2224_sv2v_reg ;
  assign \nz.mem [2223] = \nz.mem_2223_sv2v_reg ;
  assign \nz.mem [2222] = \nz.mem_2222_sv2v_reg ;
  assign \nz.mem [2221] = \nz.mem_2221_sv2v_reg ;
  assign \nz.mem [2220] = \nz.mem_2220_sv2v_reg ;
  assign \nz.mem [2219] = \nz.mem_2219_sv2v_reg ;
  assign \nz.mem [2218] = \nz.mem_2218_sv2v_reg ;
  assign \nz.mem [2217] = \nz.mem_2217_sv2v_reg ;
  assign \nz.mem [2216] = \nz.mem_2216_sv2v_reg ;
  assign \nz.mem [2215] = \nz.mem_2215_sv2v_reg ;
  assign \nz.mem [2214] = \nz.mem_2214_sv2v_reg ;
  assign \nz.mem [2213] = \nz.mem_2213_sv2v_reg ;
  assign \nz.mem [2212] = \nz.mem_2212_sv2v_reg ;
  assign \nz.mem [2211] = \nz.mem_2211_sv2v_reg ;
  assign \nz.mem [2210] = \nz.mem_2210_sv2v_reg ;
  assign \nz.mem [2209] = \nz.mem_2209_sv2v_reg ;
  assign \nz.mem [2208] = \nz.mem_2208_sv2v_reg ;
  assign \nz.mem [2207] = \nz.mem_2207_sv2v_reg ;
  assign \nz.mem [2206] = \nz.mem_2206_sv2v_reg ;
  assign \nz.mem [2205] = \nz.mem_2205_sv2v_reg ;
  assign \nz.mem [2204] = \nz.mem_2204_sv2v_reg ;
  assign \nz.mem [2203] = \nz.mem_2203_sv2v_reg ;
  assign \nz.mem [2202] = \nz.mem_2202_sv2v_reg ;
  assign \nz.mem [2201] = \nz.mem_2201_sv2v_reg ;
  assign \nz.mem [2200] = \nz.mem_2200_sv2v_reg ;
  assign \nz.mem [2199] = \nz.mem_2199_sv2v_reg ;
  assign \nz.mem [2198] = \nz.mem_2198_sv2v_reg ;
  assign \nz.mem [2197] = \nz.mem_2197_sv2v_reg ;
  assign \nz.mem [2196] = \nz.mem_2196_sv2v_reg ;
  assign \nz.mem [2195] = \nz.mem_2195_sv2v_reg ;
  assign \nz.mem [2194] = \nz.mem_2194_sv2v_reg ;
  assign \nz.mem [2193] = \nz.mem_2193_sv2v_reg ;
  assign \nz.mem [2192] = \nz.mem_2192_sv2v_reg ;
  assign \nz.mem [2191] = \nz.mem_2191_sv2v_reg ;
  assign \nz.mem [2190] = \nz.mem_2190_sv2v_reg ;
  assign \nz.mem [2189] = \nz.mem_2189_sv2v_reg ;
  assign \nz.mem [2188] = \nz.mem_2188_sv2v_reg ;
  assign \nz.mem [2187] = \nz.mem_2187_sv2v_reg ;
  assign \nz.mem [2186] = \nz.mem_2186_sv2v_reg ;
  assign \nz.mem [2185] = \nz.mem_2185_sv2v_reg ;
  assign \nz.mem [2184] = \nz.mem_2184_sv2v_reg ;
  assign \nz.mem [2183] = \nz.mem_2183_sv2v_reg ;
  assign \nz.mem [2182] = \nz.mem_2182_sv2v_reg ;
  assign \nz.mem [2181] = \nz.mem_2181_sv2v_reg ;
  assign \nz.mem [2180] = \nz.mem_2180_sv2v_reg ;
  assign \nz.mem [2179] = \nz.mem_2179_sv2v_reg ;
  assign \nz.mem [2178] = \nz.mem_2178_sv2v_reg ;
  assign \nz.mem [2177] = \nz.mem_2177_sv2v_reg ;
  assign \nz.mem [2176] = \nz.mem_2176_sv2v_reg ;
  assign \nz.mem [2175] = \nz.mem_2175_sv2v_reg ;
  assign \nz.mem [2174] = \nz.mem_2174_sv2v_reg ;
  assign \nz.mem [2173] = \nz.mem_2173_sv2v_reg ;
  assign \nz.mem [2172] = \nz.mem_2172_sv2v_reg ;
  assign \nz.mem [2171] = \nz.mem_2171_sv2v_reg ;
  assign \nz.mem [2170] = \nz.mem_2170_sv2v_reg ;
  assign \nz.mem [2169] = \nz.mem_2169_sv2v_reg ;
  assign \nz.mem [2168] = \nz.mem_2168_sv2v_reg ;
  assign \nz.mem [2167] = \nz.mem_2167_sv2v_reg ;
  assign \nz.mem [2166] = \nz.mem_2166_sv2v_reg ;
  assign \nz.mem [2165] = \nz.mem_2165_sv2v_reg ;
  assign \nz.mem [2164] = \nz.mem_2164_sv2v_reg ;
  assign \nz.mem [2163] = \nz.mem_2163_sv2v_reg ;
  assign \nz.mem [2162] = \nz.mem_2162_sv2v_reg ;
  assign \nz.mem [2161] = \nz.mem_2161_sv2v_reg ;
  assign \nz.mem [2160] = \nz.mem_2160_sv2v_reg ;
  assign \nz.mem [2159] = \nz.mem_2159_sv2v_reg ;
  assign \nz.mem [2158] = \nz.mem_2158_sv2v_reg ;
  assign \nz.mem [2157] = \nz.mem_2157_sv2v_reg ;
  assign \nz.mem [2156] = \nz.mem_2156_sv2v_reg ;
  assign \nz.mem [2155] = \nz.mem_2155_sv2v_reg ;
  assign \nz.mem [2154] = \nz.mem_2154_sv2v_reg ;
  assign \nz.mem [2153] = \nz.mem_2153_sv2v_reg ;
  assign \nz.mem [2152] = \nz.mem_2152_sv2v_reg ;
  assign \nz.mem [2151] = \nz.mem_2151_sv2v_reg ;
  assign \nz.mem [2150] = \nz.mem_2150_sv2v_reg ;
  assign \nz.mem [2149] = \nz.mem_2149_sv2v_reg ;
  assign \nz.mem [2148] = \nz.mem_2148_sv2v_reg ;
  assign \nz.mem [2147] = \nz.mem_2147_sv2v_reg ;
  assign \nz.mem [2146] = \nz.mem_2146_sv2v_reg ;
  assign \nz.mem [2145] = \nz.mem_2145_sv2v_reg ;
  assign \nz.mem [2144] = \nz.mem_2144_sv2v_reg ;
  assign \nz.mem [2143] = \nz.mem_2143_sv2v_reg ;
  assign \nz.mem [2142] = \nz.mem_2142_sv2v_reg ;
  assign \nz.mem [2141] = \nz.mem_2141_sv2v_reg ;
  assign \nz.mem [2140] = \nz.mem_2140_sv2v_reg ;
  assign \nz.mem [2139] = \nz.mem_2139_sv2v_reg ;
  assign \nz.mem [2138] = \nz.mem_2138_sv2v_reg ;
  assign \nz.mem [2137] = \nz.mem_2137_sv2v_reg ;
  assign \nz.mem [2136] = \nz.mem_2136_sv2v_reg ;
  assign \nz.mem [2135] = \nz.mem_2135_sv2v_reg ;
  assign \nz.mem [2134] = \nz.mem_2134_sv2v_reg ;
  assign \nz.mem [2133] = \nz.mem_2133_sv2v_reg ;
  assign \nz.mem [2132] = \nz.mem_2132_sv2v_reg ;
  assign \nz.mem [2131] = \nz.mem_2131_sv2v_reg ;
  assign \nz.mem [2130] = \nz.mem_2130_sv2v_reg ;
  assign \nz.mem [2129] = \nz.mem_2129_sv2v_reg ;
  assign \nz.mem [2128] = \nz.mem_2128_sv2v_reg ;
  assign \nz.mem [2127] = \nz.mem_2127_sv2v_reg ;
  assign \nz.mem [2126] = \nz.mem_2126_sv2v_reg ;
  assign \nz.mem [2125] = \nz.mem_2125_sv2v_reg ;
  assign \nz.mem [2124] = \nz.mem_2124_sv2v_reg ;
  assign \nz.mem [2123] = \nz.mem_2123_sv2v_reg ;
  assign \nz.mem [2122] = \nz.mem_2122_sv2v_reg ;
  assign \nz.mem [2121] = \nz.mem_2121_sv2v_reg ;
  assign \nz.mem [2120] = \nz.mem_2120_sv2v_reg ;
  assign \nz.mem [2119] = \nz.mem_2119_sv2v_reg ;
  assign \nz.mem [2118] = \nz.mem_2118_sv2v_reg ;
  assign \nz.mem [2117] = \nz.mem_2117_sv2v_reg ;
  assign \nz.mem [2116] = \nz.mem_2116_sv2v_reg ;
  assign \nz.mem [2115] = \nz.mem_2115_sv2v_reg ;
  assign \nz.mem [2114] = \nz.mem_2114_sv2v_reg ;
  assign \nz.mem [2113] = \nz.mem_2113_sv2v_reg ;
  assign \nz.mem [2112] = \nz.mem_2112_sv2v_reg ;
  assign \nz.mem [2111] = \nz.mem_2111_sv2v_reg ;
  assign \nz.mem [2110] = \nz.mem_2110_sv2v_reg ;
  assign \nz.mem [2109] = \nz.mem_2109_sv2v_reg ;
  assign \nz.mem [2108] = \nz.mem_2108_sv2v_reg ;
  assign \nz.mem [2107] = \nz.mem_2107_sv2v_reg ;
  assign \nz.mem [2106] = \nz.mem_2106_sv2v_reg ;
  assign \nz.mem [2105] = \nz.mem_2105_sv2v_reg ;
  assign \nz.mem [2104] = \nz.mem_2104_sv2v_reg ;
  assign \nz.mem [2103] = \nz.mem_2103_sv2v_reg ;
  assign \nz.mem [2102] = \nz.mem_2102_sv2v_reg ;
  assign \nz.mem [2101] = \nz.mem_2101_sv2v_reg ;
  assign \nz.mem [2100] = \nz.mem_2100_sv2v_reg ;
  assign \nz.mem [2099] = \nz.mem_2099_sv2v_reg ;
  assign \nz.mem [2098] = \nz.mem_2098_sv2v_reg ;
  assign \nz.mem [2097] = \nz.mem_2097_sv2v_reg ;
  assign \nz.mem [2096] = \nz.mem_2096_sv2v_reg ;
  assign \nz.mem [2095] = \nz.mem_2095_sv2v_reg ;
  assign \nz.mem [2094] = \nz.mem_2094_sv2v_reg ;
  assign \nz.mem [2093] = \nz.mem_2093_sv2v_reg ;
  assign \nz.mem [2092] = \nz.mem_2092_sv2v_reg ;
  assign \nz.mem [2091] = \nz.mem_2091_sv2v_reg ;
  assign \nz.mem [2090] = \nz.mem_2090_sv2v_reg ;
  assign \nz.mem [2089] = \nz.mem_2089_sv2v_reg ;
  assign \nz.mem [2088] = \nz.mem_2088_sv2v_reg ;
  assign \nz.mem [2087] = \nz.mem_2087_sv2v_reg ;
  assign \nz.mem [2086] = \nz.mem_2086_sv2v_reg ;
  assign \nz.mem [2085] = \nz.mem_2085_sv2v_reg ;
  assign \nz.mem [2084] = \nz.mem_2084_sv2v_reg ;
  assign \nz.mem [2083] = \nz.mem_2083_sv2v_reg ;
  assign \nz.mem [2082] = \nz.mem_2082_sv2v_reg ;
  assign \nz.mem [2081] = \nz.mem_2081_sv2v_reg ;
  assign \nz.mem [2080] = \nz.mem_2080_sv2v_reg ;
  assign \nz.mem [2079] = \nz.mem_2079_sv2v_reg ;
  assign \nz.mem [2078] = \nz.mem_2078_sv2v_reg ;
  assign \nz.mem [2077] = \nz.mem_2077_sv2v_reg ;
  assign \nz.mem [2076] = \nz.mem_2076_sv2v_reg ;
  assign \nz.mem [2075] = \nz.mem_2075_sv2v_reg ;
  assign \nz.mem [2074] = \nz.mem_2074_sv2v_reg ;
  assign \nz.mem [2073] = \nz.mem_2073_sv2v_reg ;
  assign \nz.mem [2072] = \nz.mem_2072_sv2v_reg ;
  assign \nz.mem [2071] = \nz.mem_2071_sv2v_reg ;
  assign \nz.mem [2070] = \nz.mem_2070_sv2v_reg ;
  assign \nz.mem [2069] = \nz.mem_2069_sv2v_reg ;
  assign \nz.mem [2068] = \nz.mem_2068_sv2v_reg ;
  assign \nz.mem [2067] = \nz.mem_2067_sv2v_reg ;
  assign \nz.mem [2066] = \nz.mem_2066_sv2v_reg ;
  assign \nz.mem [2065] = \nz.mem_2065_sv2v_reg ;
  assign \nz.mem [2064] = \nz.mem_2064_sv2v_reg ;
  assign \nz.mem [2063] = \nz.mem_2063_sv2v_reg ;
  assign \nz.mem [2062] = \nz.mem_2062_sv2v_reg ;
  assign \nz.mem [2061] = \nz.mem_2061_sv2v_reg ;
  assign \nz.mem [2060] = \nz.mem_2060_sv2v_reg ;
  assign \nz.mem [2059] = \nz.mem_2059_sv2v_reg ;
  assign \nz.mem [2058] = \nz.mem_2058_sv2v_reg ;
  assign \nz.mem [2057] = \nz.mem_2057_sv2v_reg ;
  assign \nz.mem [2056] = \nz.mem_2056_sv2v_reg ;
  assign \nz.mem [2055] = \nz.mem_2055_sv2v_reg ;
  assign \nz.mem [2054] = \nz.mem_2054_sv2v_reg ;
  assign \nz.mem [2053] = \nz.mem_2053_sv2v_reg ;
  assign \nz.mem [2052] = \nz.mem_2052_sv2v_reg ;
  assign \nz.mem [2051] = \nz.mem_2051_sv2v_reg ;
  assign \nz.mem [2050] = \nz.mem_2050_sv2v_reg ;
  assign \nz.mem [2049] = \nz.mem_2049_sv2v_reg ;
  assign \nz.mem [2048] = \nz.mem_2048_sv2v_reg ;
  assign \nz.mem [2047] = \nz.mem_2047_sv2v_reg ;
  assign \nz.mem [2046] = \nz.mem_2046_sv2v_reg ;
  assign \nz.mem [2045] = \nz.mem_2045_sv2v_reg ;
  assign \nz.mem [2044] = \nz.mem_2044_sv2v_reg ;
  assign \nz.mem [2043] = \nz.mem_2043_sv2v_reg ;
  assign \nz.mem [2042] = \nz.mem_2042_sv2v_reg ;
  assign \nz.mem [2041] = \nz.mem_2041_sv2v_reg ;
  assign \nz.mem [2040] = \nz.mem_2040_sv2v_reg ;
  assign \nz.mem [2039] = \nz.mem_2039_sv2v_reg ;
  assign \nz.mem [2038] = \nz.mem_2038_sv2v_reg ;
  assign \nz.mem [2037] = \nz.mem_2037_sv2v_reg ;
  assign \nz.mem [2036] = \nz.mem_2036_sv2v_reg ;
  assign \nz.mem [2035] = \nz.mem_2035_sv2v_reg ;
  assign \nz.mem [2034] = \nz.mem_2034_sv2v_reg ;
  assign \nz.mem [2033] = \nz.mem_2033_sv2v_reg ;
  assign \nz.mem [2032] = \nz.mem_2032_sv2v_reg ;
  assign \nz.mem [2031] = \nz.mem_2031_sv2v_reg ;
  assign \nz.mem [2030] = \nz.mem_2030_sv2v_reg ;
  assign \nz.mem [2029] = \nz.mem_2029_sv2v_reg ;
  assign \nz.mem [2028] = \nz.mem_2028_sv2v_reg ;
  assign \nz.mem [2027] = \nz.mem_2027_sv2v_reg ;
  assign \nz.mem [2026] = \nz.mem_2026_sv2v_reg ;
  assign \nz.mem [2025] = \nz.mem_2025_sv2v_reg ;
  assign \nz.mem [2024] = \nz.mem_2024_sv2v_reg ;
  assign \nz.mem [2023] = \nz.mem_2023_sv2v_reg ;
  assign \nz.mem [2022] = \nz.mem_2022_sv2v_reg ;
  assign \nz.mem [2021] = \nz.mem_2021_sv2v_reg ;
  assign \nz.mem [2020] = \nz.mem_2020_sv2v_reg ;
  assign \nz.mem [2019] = \nz.mem_2019_sv2v_reg ;
  assign \nz.mem [2018] = \nz.mem_2018_sv2v_reg ;
  assign \nz.mem [2017] = \nz.mem_2017_sv2v_reg ;
  assign \nz.mem [2016] = \nz.mem_2016_sv2v_reg ;
  assign \nz.mem [2015] = \nz.mem_2015_sv2v_reg ;
  assign \nz.mem [2014] = \nz.mem_2014_sv2v_reg ;
  assign \nz.mem [2013] = \nz.mem_2013_sv2v_reg ;
  assign \nz.mem [2012] = \nz.mem_2012_sv2v_reg ;
  assign \nz.mem [2011] = \nz.mem_2011_sv2v_reg ;
  assign \nz.mem [2010] = \nz.mem_2010_sv2v_reg ;
  assign \nz.mem [2009] = \nz.mem_2009_sv2v_reg ;
  assign \nz.mem [2008] = \nz.mem_2008_sv2v_reg ;
  assign \nz.mem [2007] = \nz.mem_2007_sv2v_reg ;
  assign \nz.mem [2006] = \nz.mem_2006_sv2v_reg ;
  assign \nz.mem [2005] = \nz.mem_2005_sv2v_reg ;
  assign \nz.mem [2004] = \nz.mem_2004_sv2v_reg ;
  assign \nz.mem [2003] = \nz.mem_2003_sv2v_reg ;
  assign \nz.mem [2002] = \nz.mem_2002_sv2v_reg ;
  assign \nz.mem [2001] = \nz.mem_2001_sv2v_reg ;
  assign \nz.mem [2000] = \nz.mem_2000_sv2v_reg ;
  assign \nz.mem [1999] = \nz.mem_1999_sv2v_reg ;
  assign \nz.mem [1998] = \nz.mem_1998_sv2v_reg ;
  assign \nz.mem [1997] = \nz.mem_1997_sv2v_reg ;
  assign \nz.mem [1996] = \nz.mem_1996_sv2v_reg ;
  assign \nz.mem [1995] = \nz.mem_1995_sv2v_reg ;
  assign \nz.mem [1994] = \nz.mem_1994_sv2v_reg ;
  assign \nz.mem [1993] = \nz.mem_1993_sv2v_reg ;
  assign \nz.mem [1992] = \nz.mem_1992_sv2v_reg ;
  assign \nz.mem [1991] = \nz.mem_1991_sv2v_reg ;
  assign \nz.mem [1990] = \nz.mem_1990_sv2v_reg ;
  assign \nz.mem [1989] = \nz.mem_1989_sv2v_reg ;
  assign \nz.mem [1988] = \nz.mem_1988_sv2v_reg ;
  assign \nz.mem [1987] = \nz.mem_1987_sv2v_reg ;
  assign \nz.mem [1986] = \nz.mem_1986_sv2v_reg ;
  assign \nz.mem [1985] = \nz.mem_1985_sv2v_reg ;
  assign \nz.mem [1984] = \nz.mem_1984_sv2v_reg ;
  assign \nz.mem [1983] = \nz.mem_1983_sv2v_reg ;
  assign \nz.mem [1982] = \nz.mem_1982_sv2v_reg ;
  assign \nz.mem [1981] = \nz.mem_1981_sv2v_reg ;
  assign \nz.mem [1980] = \nz.mem_1980_sv2v_reg ;
  assign \nz.mem [1979] = \nz.mem_1979_sv2v_reg ;
  assign \nz.mem [1978] = \nz.mem_1978_sv2v_reg ;
  assign \nz.mem [1977] = \nz.mem_1977_sv2v_reg ;
  assign \nz.mem [1976] = \nz.mem_1976_sv2v_reg ;
  assign \nz.mem [1975] = \nz.mem_1975_sv2v_reg ;
  assign \nz.mem [1974] = \nz.mem_1974_sv2v_reg ;
  assign \nz.mem [1973] = \nz.mem_1973_sv2v_reg ;
  assign \nz.mem [1972] = \nz.mem_1972_sv2v_reg ;
  assign \nz.mem [1971] = \nz.mem_1971_sv2v_reg ;
  assign \nz.mem [1970] = \nz.mem_1970_sv2v_reg ;
  assign \nz.mem [1969] = \nz.mem_1969_sv2v_reg ;
  assign \nz.mem [1968] = \nz.mem_1968_sv2v_reg ;
  assign \nz.mem [1967] = \nz.mem_1967_sv2v_reg ;
  assign \nz.mem [1966] = \nz.mem_1966_sv2v_reg ;
  assign \nz.mem [1965] = \nz.mem_1965_sv2v_reg ;
  assign \nz.mem [1964] = \nz.mem_1964_sv2v_reg ;
  assign \nz.mem [1963] = \nz.mem_1963_sv2v_reg ;
  assign \nz.mem [1962] = \nz.mem_1962_sv2v_reg ;
  assign \nz.mem [1961] = \nz.mem_1961_sv2v_reg ;
  assign \nz.mem [1960] = \nz.mem_1960_sv2v_reg ;
  assign \nz.mem [1959] = \nz.mem_1959_sv2v_reg ;
  assign \nz.mem [1958] = \nz.mem_1958_sv2v_reg ;
  assign \nz.mem [1957] = \nz.mem_1957_sv2v_reg ;
  assign \nz.mem [1956] = \nz.mem_1956_sv2v_reg ;
  assign \nz.mem [1955] = \nz.mem_1955_sv2v_reg ;
  assign \nz.mem [1954] = \nz.mem_1954_sv2v_reg ;
  assign \nz.mem [1953] = \nz.mem_1953_sv2v_reg ;
  assign \nz.mem [1952] = \nz.mem_1952_sv2v_reg ;
  assign \nz.mem [1951] = \nz.mem_1951_sv2v_reg ;
  assign \nz.mem [1950] = \nz.mem_1950_sv2v_reg ;
  assign \nz.mem [1949] = \nz.mem_1949_sv2v_reg ;
  assign \nz.mem [1948] = \nz.mem_1948_sv2v_reg ;
  assign \nz.mem [1947] = \nz.mem_1947_sv2v_reg ;
  assign \nz.mem [1946] = \nz.mem_1946_sv2v_reg ;
  assign \nz.mem [1945] = \nz.mem_1945_sv2v_reg ;
  assign \nz.mem [1944] = \nz.mem_1944_sv2v_reg ;
  assign \nz.mem [1943] = \nz.mem_1943_sv2v_reg ;
  assign \nz.mem [1942] = \nz.mem_1942_sv2v_reg ;
  assign \nz.mem [1941] = \nz.mem_1941_sv2v_reg ;
  assign \nz.mem [1940] = \nz.mem_1940_sv2v_reg ;
  assign \nz.mem [1939] = \nz.mem_1939_sv2v_reg ;
  assign \nz.mem [1938] = \nz.mem_1938_sv2v_reg ;
  assign \nz.mem [1937] = \nz.mem_1937_sv2v_reg ;
  assign \nz.mem [1936] = \nz.mem_1936_sv2v_reg ;
  assign \nz.mem [1935] = \nz.mem_1935_sv2v_reg ;
  assign \nz.mem [1934] = \nz.mem_1934_sv2v_reg ;
  assign \nz.mem [1933] = \nz.mem_1933_sv2v_reg ;
  assign \nz.mem [1932] = \nz.mem_1932_sv2v_reg ;
  assign \nz.mem [1931] = \nz.mem_1931_sv2v_reg ;
  assign \nz.mem [1930] = \nz.mem_1930_sv2v_reg ;
  assign \nz.mem [1929] = \nz.mem_1929_sv2v_reg ;
  assign \nz.mem [1928] = \nz.mem_1928_sv2v_reg ;
  assign \nz.mem [1927] = \nz.mem_1927_sv2v_reg ;
  assign \nz.mem [1926] = \nz.mem_1926_sv2v_reg ;
  assign \nz.mem [1925] = \nz.mem_1925_sv2v_reg ;
  assign \nz.mem [1924] = \nz.mem_1924_sv2v_reg ;
  assign \nz.mem [1923] = \nz.mem_1923_sv2v_reg ;
  assign \nz.mem [1922] = \nz.mem_1922_sv2v_reg ;
  assign \nz.mem [1921] = \nz.mem_1921_sv2v_reg ;
  assign \nz.mem [1920] = \nz.mem_1920_sv2v_reg ;
  assign \nz.mem [1919] = \nz.mem_1919_sv2v_reg ;
  assign \nz.mem [1918] = \nz.mem_1918_sv2v_reg ;
  assign \nz.mem [1917] = \nz.mem_1917_sv2v_reg ;
  assign \nz.mem [1916] = \nz.mem_1916_sv2v_reg ;
  assign \nz.mem [1915] = \nz.mem_1915_sv2v_reg ;
  assign \nz.mem [1914] = \nz.mem_1914_sv2v_reg ;
  assign \nz.mem [1913] = \nz.mem_1913_sv2v_reg ;
  assign \nz.mem [1912] = \nz.mem_1912_sv2v_reg ;
  assign \nz.mem [1911] = \nz.mem_1911_sv2v_reg ;
  assign \nz.mem [1910] = \nz.mem_1910_sv2v_reg ;
  assign \nz.mem [1909] = \nz.mem_1909_sv2v_reg ;
  assign \nz.mem [1908] = \nz.mem_1908_sv2v_reg ;
  assign \nz.mem [1907] = \nz.mem_1907_sv2v_reg ;
  assign \nz.mem [1906] = \nz.mem_1906_sv2v_reg ;
  assign \nz.mem [1905] = \nz.mem_1905_sv2v_reg ;
  assign \nz.mem [1904] = \nz.mem_1904_sv2v_reg ;
  assign \nz.mem [1903] = \nz.mem_1903_sv2v_reg ;
  assign \nz.mem [1902] = \nz.mem_1902_sv2v_reg ;
  assign \nz.mem [1901] = \nz.mem_1901_sv2v_reg ;
  assign \nz.mem [1900] = \nz.mem_1900_sv2v_reg ;
  assign \nz.mem [1899] = \nz.mem_1899_sv2v_reg ;
  assign \nz.mem [1898] = \nz.mem_1898_sv2v_reg ;
  assign \nz.mem [1897] = \nz.mem_1897_sv2v_reg ;
  assign \nz.mem [1896] = \nz.mem_1896_sv2v_reg ;
  assign \nz.mem [1895] = \nz.mem_1895_sv2v_reg ;
  assign \nz.mem [1894] = \nz.mem_1894_sv2v_reg ;
  assign \nz.mem [1893] = \nz.mem_1893_sv2v_reg ;
  assign \nz.mem [1892] = \nz.mem_1892_sv2v_reg ;
  assign \nz.mem [1891] = \nz.mem_1891_sv2v_reg ;
  assign \nz.mem [1890] = \nz.mem_1890_sv2v_reg ;
  assign \nz.mem [1889] = \nz.mem_1889_sv2v_reg ;
  assign \nz.mem [1888] = \nz.mem_1888_sv2v_reg ;
  assign \nz.mem [1887] = \nz.mem_1887_sv2v_reg ;
  assign \nz.mem [1886] = \nz.mem_1886_sv2v_reg ;
  assign \nz.mem [1885] = \nz.mem_1885_sv2v_reg ;
  assign \nz.mem [1884] = \nz.mem_1884_sv2v_reg ;
  assign \nz.mem [1883] = \nz.mem_1883_sv2v_reg ;
  assign \nz.mem [1882] = \nz.mem_1882_sv2v_reg ;
  assign \nz.mem [1881] = \nz.mem_1881_sv2v_reg ;
  assign \nz.mem [1880] = \nz.mem_1880_sv2v_reg ;
  assign \nz.mem [1879] = \nz.mem_1879_sv2v_reg ;
  assign \nz.mem [1878] = \nz.mem_1878_sv2v_reg ;
  assign \nz.mem [1877] = \nz.mem_1877_sv2v_reg ;
  assign \nz.mem [1876] = \nz.mem_1876_sv2v_reg ;
  assign \nz.mem [1875] = \nz.mem_1875_sv2v_reg ;
  assign \nz.mem [1874] = \nz.mem_1874_sv2v_reg ;
  assign \nz.mem [1873] = \nz.mem_1873_sv2v_reg ;
  assign \nz.mem [1872] = \nz.mem_1872_sv2v_reg ;
  assign \nz.mem [1871] = \nz.mem_1871_sv2v_reg ;
  assign \nz.mem [1870] = \nz.mem_1870_sv2v_reg ;
  assign \nz.mem [1869] = \nz.mem_1869_sv2v_reg ;
  assign \nz.mem [1868] = \nz.mem_1868_sv2v_reg ;
  assign \nz.mem [1867] = \nz.mem_1867_sv2v_reg ;
  assign \nz.mem [1866] = \nz.mem_1866_sv2v_reg ;
  assign \nz.mem [1865] = \nz.mem_1865_sv2v_reg ;
  assign \nz.mem [1864] = \nz.mem_1864_sv2v_reg ;
  assign \nz.mem [1863] = \nz.mem_1863_sv2v_reg ;
  assign \nz.mem [1862] = \nz.mem_1862_sv2v_reg ;
  assign \nz.mem [1861] = \nz.mem_1861_sv2v_reg ;
  assign \nz.mem [1860] = \nz.mem_1860_sv2v_reg ;
  assign \nz.mem [1859] = \nz.mem_1859_sv2v_reg ;
  assign \nz.mem [1858] = \nz.mem_1858_sv2v_reg ;
  assign \nz.mem [1857] = \nz.mem_1857_sv2v_reg ;
  assign \nz.mem [1856] = \nz.mem_1856_sv2v_reg ;
  assign \nz.mem [1855] = \nz.mem_1855_sv2v_reg ;
  assign \nz.mem [1854] = \nz.mem_1854_sv2v_reg ;
  assign \nz.mem [1853] = \nz.mem_1853_sv2v_reg ;
  assign \nz.mem [1852] = \nz.mem_1852_sv2v_reg ;
  assign \nz.mem [1851] = \nz.mem_1851_sv2v_reg ;
  assign \nz.mem [1850] = \nz.mem_1850_sv2v_reg ;
  assign \nz.mem [1849] = \nz.mem_1849_sv2v_reg ;
  assign \nz.mem [1848] = \nz.mem_1848_sv2v_reg ;
  assign \nz.mem [1847] = \nz.mem_1847_sv2v_reg ;
  assign \nz.mem [1846] = \nz.mem_1846_sv2v_reg ;
  assign \nz.mem [1845] = \nz.mem_1845_sv2v_reg ;
  assign \nz.mem [1844] = \nz.mem_1844_sv2v_reg ;
  assign \nz.mem [1843] = \nz.mem_1843_sv2v_reg ;
  assign \nz.mem [1842] = \nz.mem_1842_sv2v_reg ;
  assign \nz.mem [1841] = \nz.mem_1841_sv2v_reg ;
  assign \nz.mem [1840] = \nz.mem_1840_sv2v_reg ;
  assign \nz.mem [1839] = \nz.mem_1839_sv2v_reg ;
  assign \nz.mem [1838] = \nz.mem_1838_sv2v_reg ;
  assign \nz.mem [1837] = \nz.mem_1837_sv2v_reg ;
  assign \nz.mem [1836] = \nz.mem_1836_sv2v_reg ;
  assign \nz.mem [1835] = \nz.mem_1835_sv2v_reg ;
  assign \nz.mem [1834] = \nz.mem_1834_sv2v_reg ;
  assign \nz.mem [1833] = \nz.mem_1833_sv2v_reg ;
  assign \nz.mem [1832] = \nz.mem_1832_sv2v_reg ;
  assign \nz.mem [1831] = \nz.mem_1831_sv2v_reg ;
  assign \nz.mem [1830] = \nz.mem_1830_sv2v_reg ;
  assign \nz.mem [1829] = \nz.mem_1829_sv2v_reg ;
  assign \nz.mem [1828] = \nz.mem_1828_sv2v_reg ;
  assign \nz.mem [1827] = \nz.mem_1827_sv2v_reg ;
  assign \nz.mem [1826] = \nz.mem_1826_sv2v_reg ;
  assign \nz.mem [1825] = \nz.mem_1825_sv2v_reg ;
  assign \nz.mem [1824] = \nz.mem_1824_sv2v_reg ;
  assign \nz.mem [1823] = \nz.mem_1823_sv2v_reg ;
  assign \nz.mem [1822] = \nz.mem_1822_sv2v_reg ;
  assign \nz.mem [1821] = \nz.mem_1821_sv2v_reg ;
  assign \nz.mem [1820] = \nz.mem_1820_sv2v_reg ;
  assign \nz.mem [1819] = \nz.mem_1819_sv2v_reg ;
  assign \nz.mem [1818] = \nz.mem_1818_sv2v_reg ;
  assign \nz.mem [1817] = \nz.mem_1817_sv2v_reg ;
  assign \nz.mem [1816] = \nz.mem_1816_sv2v_reg ;
  assign \nz.mem [1815] = \nz.mem_1815_sv2v_reg ;
  assign \nz.mem [1814] = \nz.mem_1814_sv2v_reg ;
  assign \nz.mem [1813] = \nz.mem_1813_sv2v_reg ;
  assign \nz.mem [1812] = \nz.mem_1812_sv2v_reg ;
  assign \nz.mem [1811] = \nz.mem_1811_sv2v_reg ;
  assign \nz.mem [1810] = \nz.mem_1810_sv2v_reg ;
  assign \nz.mem [1809] = \nz.mem_1809_sv2v_reg ;
  assign \nz.mem [1808] = \nz.mem_1808_sv2v_reg ;
  assign \nz.mem [1807] = \nz.mem_1807_sv2v_reg ;
  assign \nz.mem [1806] = \nz.mem_1806_sv2v_reg ;
  assign \nz.mem [1805] = \nz.mem_1805_sv2v_reg ;
  assign \nz.mem [1804] = \nz.mem_1804_sv2v_reg ;
  assign \nz.mem [1803] = \nz.mem_1803_sv2v_reg ;
  assign \nz.mem [1802] = \nz.mem_1802_sv2v_reg ;
  assign \nz.mem [1801] = \nz.mem_1801_sv2v_reg ;
  assign \nz.mem [1800] = \nz.mem_1800_sv2v_reg ;
  assign \nz.mem [1799] = \nz.mem_1799_sv2v_reg ;
  assign \nz.mem [1798] = \nz.mem_1798_sv2v_reg ;
  assign \nz.mem [1797] = \nz.mem_1797_sv2v_reg ;
  assign \nz.mem [1796] = \nz.mem_1796_sv2v_reg ;
  assign \nz.mem [1795] = \nz.mem_1795_sv2v_reg ;
  assign \nz.mem [1794] = \nz.mem_1794_sv2v_reg ;
  assign \nz.mem [1793] = \nz.mem_1793_sv2v_reg ;
  assign \nz.mem [1792] = \nz.mem_1792_sv2v_reg ;
  assign \nz.mem [1791] = \nz.mem_1791_sv2v_reg ;
  assign \nz.mem [1790] = \nz.mem_1790_sv2v_reg ;
  assign \nz.mem [1789] = \nz.mem_1789_sv2v_reg ;
  assign \nz.mem [1788] = \nz.mem_1788_sv2v_reg ;
  assign \nz.mem [1787] = \nz.mem_1787_sv2v_reg ;
  assign \nz.mem [1786] = \nz.mem_1786_sv2v_reg ;
  assign \nz.mem [1785] = \nz.mem_1785_sv2v_reg ;
  assign \nz.mem [1784] = \nz.mem_1784_sv2v_reg ;
  assign \nz.mem [1783] = \nz.mem_1783_sv2v_reg ;
  assign \nz.mem [1782] = \nz.mem_1782_sv2v_reg ;
  assign \nz.mem [1781] = \nz.mem_1781_sv2v_reg ;
  assign \nz.mem [1780] = \nz.mem_1780_sv2v_reg ;
  assign \nz.mem [1779] = \nz.mem_1779_sv2v_reg ;
  assign \nz.mem [1778] = \nz.mem_1778_sv2v_reg ;
  assign \nz.mem [1777] = \nz.mem_1777_sv2v_reg ;
  assign \nz.mem [1776] = \nz.mem_1776_sv2v_reg ;
  assign \nz.mem [1775] = \nz.mem_1775_sv2v_reg ;
  assign \nz.mem [1774] = \nz.mem_1774_sv2v_reg ;
  assign \nz.mem [1773] = \nz.mem_1773_sv2v_reg ;
  assign \nz.mem [1772] = \nz.mem_1772_sv2v_reg ;
  assign \nz.mem [1771] = \nz.mem_1771_sv2v_reg ;
  assign \nz.mem [1770] = \nz.mem_1770_sv2v_reg ;
  assign \nz.mem [1769] = \nz.mem_1769_sv2v_reg ;
  assign \nz.mem [1768] = \nz.mem_1768_sv2v_reg ;
  assign \nz.mem [1767] = \nz.mem_1767_sv2v_reg ;
  assign \nz.mem [1766] = \nz.mem_1766_sv2v_reg ;
  assign \nz.mem [1765] = \nz.mem_1765_sv2v_reg ;
  assign \nz.mem [1764] = \nz.mem_1764_sv2v_reg ;
  assign \nz.mem [1763] = \nz.mem_1763_sv2v_reg ;
  assign \nz.mem [1762] = \nz.mem_1762_sv2v_reg ;
  assign \nz.mem [1761] = \nz.mem_1761_sv2v_reg ;
  assign \nz.mem [1760] = \nz.mem_1760_sv2v_reg ;
  assign \nz.mem [1759] = \nz.mem_1759_sv2v_reg ;
  assign \nz.mem [1758] = \nz.mem_1758_sv2v_reg ;
  assign \nz.mem [1757] = \nz.mem_1757_sv2v_reg ;
  assign \nz.mem [1756] = \nz.mem_1756_sv2v_reg ;
  assign \nz.mem [1755] = \nz.mem_1755_sv2v_reg ;
  assign \nz.mem [1754] = \nz.mem_1754_sv2v_reg ;
  assign \nz.mem [1753] = \nz.mem_1753_sv2v_reg ;
  assign \nz.mem [1752] = \nz.mem_1752_sv2v_reg ;
  assign \nz.mem [1751] = \nz.mem_1751_sv2v_reg ;
  assign \nz.mem [1750] = \nz.mem_1750_sv2v_reg ;
  assign \nz.mem [1749] = \nz.mem_1749_sv2v_reg ;
  assign \nz.mem [1748] = \nz.mem_1748_sv2v_reg ;
  assign \nz.mem [1747] = \nz.mem_1747_sv2v_reg ;
  assign \nz.mem [1746] = \nz.mem_1746_sv2v_reg ;
  assign \nz.mem [1745] = \nz.mem_1745_sv2v_reg ;
  assign \nz.mem [1744] = \nz.mem_1744_sv2v_reg ;
  assign \nz.mem [1743] = \nz.mem_1743_sv2v_reg ;
  assign \nz.mem [1742] = \nz.mem_1742_sv2v_reg ;
  assign \nz.mem [1741] = \nz.mem_1741_sv2v_reg ;
  assign \nz.mem [1740] = \nz.mem_1740_sv2v_reg ;
  assign \nz.mem [1739] = \nz.mem_1739_sv2v_reg ;
  assign \nz.mem [1738] = \nz.mem_1738_sv2v_reg ;
  assign \nz.mem [1737] = \nz.mem_1737_sv2v_reg ;
  assign \nz.mem [1736] = \nz.mem_1736_sv2v_reg ;
  assign \nz.mem [1735] = \nz.mem_1735_sv2v_reg ;
  assign \nz.mem [1734] = \nz.mem_1734_sv2v_reg ;
  assign \nz.mem [1733] = \nz.mem_1733_sv2v_reg ;
  assign \nz.mem [1732] = \nz.mem_1732_sv2v_reg ;
  assign \nz.mem [1731] = \nz.mem_1731_sv2v_reg ;
  assign \nz.mem [1730] = \nz.mem_1730_sv2v_reg ;
  assign \nz.mem [1729] = \nz.mem_1729_sv2v_reg ;
  assign \nz.mem [1728] = \nz.mem_1728_sv2v_reg ;
  assign \nz.mem [1727] = \nz.mem_1727_sv2v_reg ;
  assign \nz.mem [1726] = \nz.mem_1726_sv2v_reg ;
  assign \nz.mem [1725] = \nz.mem_1725_sv2v_reg ;
  assign \nz.mem [1724] = \nz.mem_1724_sv2v_reg ;
  assign \nz.mem [1723] = \nz.mem_1723_sv2v_reg ;
  assign \nz.mem [1722] = \nz.mem_1722_sv2v_reg ;
  assign \nz.mem [1721] = \nz.mem_1721_sv2v_reg ;
  assign \nz.mem [1720] = \nz.mem_1720_sv2v_reg ;
  assign \nz.mem [1719] = \nz.mem_1719_sv2v_reg ;
  assign \nz.mem [1718] = \nz.mem_1718_sv2v_reg ;
  assign \nz.mem [1717] = \nz.mem_1717_sv2v_reg ;
  assign \nz.mem [1716] = \nz.mem_1716_sv2v_reg ;
  assign \nz.mem [1715] = \nz.mem_1715_sv2v_reg ;
  assign \nz.mem [1714] = \nz.mem_1714_sv2v_reg ;
  assign \nz.mem [1713] = \nz.mem_1713_sv2v_reg ;
  assign \nz.mem [1712] = \nz.mem_1712_sv2v_reg ;
  assign \nz.mem [1711] = \nz.mem_1711_sv2v_reg ;
  assign \nz.mem [1710] = \nz.mem_1710_sv2v_reg ;
  assign \nz.mem [1709] = \nz.mem_1709_sv2v_reg ;
  assign \nz.mem [1708] = \nz.mem_1708_sv2v_reg ;
  assign \nz.mem [1707] = \nz.mem_1707_sv2v_reg ;
  assign \nz.mem [1706] = \nz.mem_1706_sv2v_reg ;
  assign \nz.mem [1705] = \nz.mem_1705_sv2v_reg ;
  assign \nz.mem [1704] = \nz.mem_1704_sv2v_reg ;
  assign \nz.mem [1703] = \nz.mem_1703_sv2v_reg ;
  assign \nz.mem [1702] = \nz.mem_1702_sv2v_reg ;
  assign \nz.mem [1701] = \nz.mem_1701_sv2v_reg ;
  assign \nz.mem [1700] = \nz.mem_1700_sv2v_reg ;
  assign \nz.mem [1699] = \nz.mem_1699_sv2v_reg ;
  assign \nz.mem [1698] = \nz.mem_1698_sv2v_reg ;
  assign \nz.mem [1697] = \nz.mem_1697_sv2v_reg ;
  assign \nz.mem [1696] = \nz.mem_1696_sv2v_reg ;
  assign \nz.mem [1695] = \nz.mem_1695_sv2v_reg ;
  assign \nz.mem [1694] = \nz.mem_1694_sv2v_reg ;
  assign \nz.mem [1693] = \nz.mem_1693_sv2v_reg ;
  assign \nz.mem [1692] = \nz.mem_1692_sv2v_reg ;
  assign \nz.mem [1691] = \nz.mem_1691_sv2v_reg ;
  assign \nz.mem [1690] = \nz.mem_1690_sv2v_reg ;
  assign \nz.mem [1689] = \nz.mem_1689_sv2v_reg ;
  assign \nz.mem [1688] = \nz.mem_1688_sv2v_reg ;
  assign \nz.mem [1687] = \nz.mem_1687_sv2v_reg ;
  assign \nz.mem [1686] = \nz.mem_1686_sv2v_reg ;
  assign \nz.mem [1685] = \nz.mem_1685_sv2v_reg ;
  assign \nz.mem [1684] = \nz.mem_1684_sv2v_reg ;
  assign \nz.mem [1683] = \nz.mem_1683_sv2v_reg ;
  assign \nz.mem [1682] = \nz.mem_1682_sv2v_reg ;
  assign \nz.mem [1681] = \nz.mem_1681_sv2v_reg ;
  assign \nz.mem [1680] = \nz.mem_1680_sv2v_reg ;
  assign \nz.mem [1679] = \nz.mem_1679_sv2v_reg ;
  assign \nz.mem [1678] = \nz.mem_1678_sv2v_reg ;
  assign \nz.mem [1677] = \nz.mem_1677_sv2v_reg ;
  assign \nz.mem [1676] = \nz.mem_1676_sv2v_reg ;
  assign \nz.mem [1675] = \nz.mem_1675_sv2v_reg ;
  assign \nz.mem [1674] = \nz.mem_1674_sv2v_reg ;
  assign \nz.mem [1673] = \nz.mem_1673_sv2v_reg ;
  assign \nz.mem [1672] = \nz.mem_1672_sv2v_reg ;
  assign \nz.mem [1671] = \nz.mem_1671_sv2v_reg ;
  assign \nz.mem [1670] = \nz.mem_1670_sv2v_reg ;
  assign \nz.mem [1669] = \nz.mem_1669_sv2v_reg ;
  assign \nz.mem [1668] = \nz.mem_1668_sv2v_reg ;
  assign \nz.mem [1667] = \nz.mem_1667_sv2v_reg ;
  assign \nz.mem [1666] = \nz.mem_1666_sv2v_reg ;
  assign \nz.mem [1665] = \nz.mem_1665_sv2v_reg ;
  assign \nz.mem [1664] = \nz.mem_1664_sv2v_reg ;
  assign \nz.mem [1663] = \nz.mem_1663_sv2v_reg ;
  assign \nz.mem [1662] = \nz.mem_1662_sv2v_reg ;
  assign \nz.mem [1661] = \nz.mem_1661_sv2v_reg ;
  assign \nz.mem [1660] = \nz.mem_1660_sv2v_reg ;
  assign \nz.mem [1659] = \nz.mem_1659_sv2v_reg ;
  assign \nz.mem [1658] = \nz.mem_1658_sv2v_reg ;
  assign \nz.mem [1657] = \nz.mem_1657_sv2v_reg ;
  assign \nz.mem [1656] = \nz.mem_1656_sv2v_reg ;
  assign \nz.mem [1655] = \nz.mem_1655_sv2v_reg ;
  assign \nz.mem [1654] = \nz.mem_1654_sv2v_reg ;
  assign \nz.mem [1653] = \nz.mem_1653_sv2v_reg ;
  assign \nz.mem [1652] = \nz.mem_1652_sv2v_reg ;
  assign \nz.mem [1651] = \nz.mem_1651_sv2v_reg ;
  assign \nz.mem [1650] = \nz.mem_1650_sv2v_reg ;
  assign \nz.mem [1649] = \nz.mem_1649_sv2v_reg ;
  assign \nz.mem [1648] = \nz.mem_1648_sv2v_reg ;
  assign \nz.mem [1647] = \nz.mem_1647_sv2v_reg ;
  assign \nz.mem [1646] = \nz.mem_1646_sv2v_reg ;
  assign \nz.mem [1645] = \nz.mem_1645_sv2v_reg ;
  assign \nz.mem [1644] = \nz.mem_1644_sv2v_reg ;
  assign \nz.mem [1643] = \nz.mem_1643_sv2v_reg ;
  assign \nz.mem [1642] = \nz.mem_1642_sv2v_reg ;
  assign \nz.mem [1641] = \nz.mem_1641_sv2v_reg ;
  assign \nz.mem [1640] = \nz.mem_1640_sv2v_reg ;
  assign \nz.mem [1639] = \nz.mem_1639_sv2v_reg ;
  assign \nz.mem [1638] = \nz.mem_1638_sv2v_reg ;
  assign \nz.mem [1637] = \nz.mem_1637_sv2v_reg ;
  assign \nz.mem [1636] = \nz.mem_1636_sv2v_reg ;
  assign \nz.mem [1635] = \nz.mem_1635_sv2v_reg ;
  assign \nz.mem [1634] = \nz.mem_1634_sv2v_reg ;
  assign \nz.mem [1633] = \nz.mem_1633_sv2v_reg ;
  assign \nz.mem [1632] = \nz.mem_1632_sv2v_reg ;
  assign \nz.mem [1631] = \nz.mem_1631_sv2v_reg ;
  assign \nz.mem [1630] = \nz.mem_1630_sv2v_reg ;
  assign \nz.mem [1629] = \nz.mem_1629_sv2v_reg ;
  assign \nz.mem [1628] = \nz.mem_1628_sv2v_reg ;
  assign \nz.mem [1627] = \nz.mem_1627_sv2v_reg ;
  assign \nz.mem [1626] = \nz.mem_1626_sv2v_reg ;
  assign \nz.mem [1625] = \nz.mem_1625_sv2v_reg ;
  assign \nz.mem [1624] = \nz.mem_1624_sv2v_reg ;
  assign \nz.mem [1623] = \nz.mem_1623_sv2v_reg ;
  assign \nz.mem [1622] = \nz.mem_1622_sv2v_reg ;
  assign \nz.mem [1621] = \nz.mem_1621_sv2v_reg ;
  assign \nz.mem [1620] = \nz.mem_1620_sv2v_reg ;
  assign \nz.mem [1619] = \nz.mem_1619_sv2v_reg ;
  assign \nz.mem [1618] = \nz.mem_1618_sv2v_reg ;
  assign \nz.mem [1617] = \nz.mem_1617_sv2v_reg ;
  assign \nz.mem [1616] = \nz.mem_1616_sv2v_reg ;
  assign \nz.mem [1615] = \nz.mem_1615_sv2v_reg ;
  assign \nz.mem [1614] = \nz.mem_1614_sv2v_reg ;
  assign \nz.mem [1613] = \nz.mem_1613_sv2v_reg ;
  assign \nz.mem [1612] = \nz.mem_1612_sv2v_reg ;
  assign \nz.mem [1611] = \nz.mem_1611_sv2v_reg ;
  assign \nz.mem [1610] = \nz.mem_1610_sv2v_reg ;
  assign \nz.mem [1609] = \nz.mem_1609_sv2v_reg ;
  assign \nz.mem [1608] = \nz.mem_1608_sv2v_reg ;
  assign \nz.mem [1607] = \nz.mem_1607_sv2v_reg ;
  assign \nz.mem [1606] = \nz.mem_1606_sv2v_reg ;
  assign \nz.mem [1605] = \nz.mem_1605_sv2v_reg ;
  assign \nz.mem [1604] = \nz.mem_1604_sv2v_reg ;
  assign \nz.mem [1603] = \nz.mem_1603_sv2v_reg ;
  assign \nz.mem [1602] = \nz.mem_1602_sv2v_reg ;
  assign \nz.mem [1601] = \nz.mem_1601_sv2v_reg ;
  assign \nz.mem [1600] = \nz.mem_1600_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [39] = (N115)? \nz.mem [39] : 
                             (N117)? \nz.mem [79] : 
                             (N119)? \nz.mem [119] : 
                             (N121)? \nz.mem [159] : 
                             (N123)? \nz.mem [199] : 
                             (N125)? \nz.mem [239] : 
                             (N127)? \nz.mem [279] : 
                             (N129)? \nz.mem [319] : 
                             (N131)? \nz.mem [359] : 
                             (N133)? \nz.mem [399] : 
                             (N135)? \nz.mem [439] : 
                             (N137)? \nz.mem [479] : 
                             (N139)? \nz.mem [519] : 
                             (N141)? \nz.mem [559] : 
                             (N143)? \nz.mem [599] : 
                             (N145)? \nz.mem [639] : 
                             (N147)? \nz.mem [679] : 
                             (N149)? \nz.mem [719] : 
                             (N151)? \nz.mem [759] : 
                             (N153)? \nz.mem [799] : 
                             (N155)? \nz.mem [839] : 
                             (N157)? \nz.mem [879] : 
                             (N159)? \nz.mem [919] : 
                             (N161)? \nz.mem [959] : 
                             (N163)? \nz.mem [999] : 
                             (N165)? \nz.mem [1039] : 
                             (N167)? \nz.mem [1079] : 
                             (N169)? \nz.mem [1119] : 
                             (N171)? \nz.mem [1159] : 
                             (N173)? \nz.mem [1199] : 
                             (N175)? \nz.mem [1239] : 
                             (N177)? \nz.mem [1279] : 
                             (N116)? \nz.mem [1319] : 
                             (N118)? \nz.mem [1359] : 
                             (N120)? \nz.mem [1399] : 
                             (N122)? \nz.mem [1439] : 
                             (N124)? \nz.mem [1479] : 
                             (N126)? \nz.mem [1519] : 
                             (N128)? \nz.mem [1559] : 
                             (N130)? \nz.mem [1599] : 
                             (N132)? \nz.mem [1639] : 
                             (N134)? \nz.mem [1679] : 
                             (N136)? \nz.mem [1719] : 
                             (N138)? \nz.mem [1759] : 
                             (N140)? \nz.mem [1799] : 
                             (N142)? \nz.mem [1839] : 
                             (N144)? \nz.mem [1879] : 
                             (N146)? \nz.mem [1919] : 
                             (N148)? \nz.mem [1959] : 
                             (N150)? \nz.mem [1999] : 
                             (N152)? \nz.mem [2039] : 
                             (N154)? \nz.mem [2079] : 
                             (N156)? \nz.mem [2119] : 
                             (N158)? \nz.mem [2159] : 
                             (N160)? \nz.mem [2199] : 
                             (N162)? \nz.mem [2239] : 
                             (N164)? \nz.mem [2279] : 
                             (N166)? \nz.mem [2319] : 
                             (N168)? \nz.mem [2359] : 
                             (N170)? \nz.mem [2399] : 
                             (N172)? \nz.mem [2439] : 
                             (N174)? \nz.mem [2479] : 
                             (N176)? \nz.mem [2519] : 
                             (N178)? \nz.mem [2559] : 1'b0;
  assign \nz.data_out [38] = (N115)? \nz.mem [38] : 
                             (N117)? \nz.mem [78] : 
                             (N119)? \nz.mem [118] : 
                             (N121)? \nz.mem [158] : 
                             (N123)? \nz.mem [198] : 
                             (N125)? \nz.mem [238] : 
                             (N127)? \nz.mem [278] : 
                             (N129)? \nz.mem [318] : 
                             (N131)? \nz.mem [358] : 
                             (N133)? \nz.mem [398] : 
                             (N135)? \nz.mem [438] : 
                             (N137)? \nz.mem [478] : 
                             (N139)? \nz.mem [518] : 
                             (N141)? \nz.mem [558] : 
                             (N143)? \nz.mem [598] : 
                             (N145)? \nz.mem [638] : 
                             (N147)? \nz.mem [678] : 
                             (N149)? \nz.mem [718] : 
                             (N151)? \nz.mem [758] : 
                             (N153)? \nz.mem [798] : 
                             (N155)? \nz.mem [838] : 
                             (N157)? \nz.mem [878] : 
                             (N159)? \nz.mem [918] : 
                             (N161)? \nz.mem [958] : 
                             (N163)? \nz.mem [998] : 
                             (N165)? \nz.mem [1038] : 
                             (N167)? \nz.mem [1078] : 
                             (N169)? \nz.mem [1118] : 
                             (N171)? \nz.mem [1158] : 
                             (N173)? \nz.mem [1198] : 
                             (N175)? \nz.mem [1238] : 
                             (N177)? \nz.mem [1278] : 
                             (N116)? \nz.mem [1318] : 
                             (N118)? \nz.mem [1358] : 
                             (N120)? \nz.mem [1398] : 
                             (N122)? \nz.mem [1438] : 
                             (N124)? \nz.mem [1478] : 
                             (N126)? \nz.mem [1518] : 
                             (N128)? \nz.mem [1558] : 
                             (N130)? \nz.mem [1598] : 
                             (N132)? \nz.mem [1638] : 
                             (N134)? \nz.mem [1678] : 
                             (N136)? \nz.mem [1718] : 
                             (N138)? \nz.mem [1758] : 
                             (N140)? \nz.mem [1798] : 
                             (N142)? \nz.mem [1838] : 
                             (N144)? \nz.mem [1878] : 
                             (N146)? \nz.mem [1918] : 
                             (N148)? \nz.mem [1958] : 
                             (N150)? \nz.mem [1998] : 
                             (N152)? \nz.mem [2038] : 
                             (N154)? \nz.mem [2078] : 
                             (N156)? \nz.mem [2118] : 
                             (N158)? \nz.mem [2158] : 
                             (N160)? \nz.mem [2198] : 
                             (N162)? \nz.mem [2238] : 
                             (N164)? \nz.mem [2278] : 
                             (N166)? \nz.mem [2318] : 
                             (N168)? \nz.mem [2358] : 
                             (N170)? \nz.mem [2398] : 
                             (N172)? \nz.mem [2438] : 
                             (N174)? \nz.mem [2478] : 
                             (N176)? \nz.mem [2518] : 
                             (N178)? \nz.mem [2558] : 1'b0;
  assign \nz.data_out [37] = (N115)? \nz.mem [37] : 
                             (N117)? \nz.mem [77] : 
                             (N119)? \nz.mem [117] : 
                             (N121)? \nz.mem [157] : 
                             (N123)? \nz.mem [197] : 
                             (N125)? \nz.mem [237] : 
                             (N127)? \nz.mem [277] : 
                             (N129)? \nz.mem [317] : 
                             (N131)? \nz.mem [357] : 
                             (N133)? \nz.mem [397] : 
                             (N135)? \nz.mem [437] : 
                             (N137)? \nz.mem [477] : 
                             (N139)? \nz.mem [517] : 
                             (N141)? \nz.mem [557] : 
                             (N143)? \nz.mem [597] : 
                             (N145)? \nz.mem [637] : 
                             (N147)? \nz.mem [677] : 
                             (N149)? \nz.mem [717] : 
                             (N151)? \nz.mem [757] : 
                             (N153)? \nz.mem [797] : 
                             (N155)? \nz.mem [837] : 
                             (N157)? \nz.mem [877] : 
                             (N159)? \nz.mem [917] : 
                             (N161)? \nz.mem [957] : 
                             (N163)? \nz.mem [997] : 
                             (N165)? \nz.mem [1037] : 
                             (N167)? \nz.mem [1077] : 
                             (N169)? \nz.mem [1117] : 
                             (N171)? \nz.mem [1157] : 
                             (N173)? \nz.mem [1197] : 
                             (N175)? \nz.mem [1237] : 
                             (N177)? \nz.mem [1277] : 
                             (N116)? \nz.mem [1317] : 
                             (N118)? \nz.mem [1357] : 
                             (N120)? \nz.mem [1397] : 
                             (N122)? \nz.mem [1437] : 
                             (N124)? \nz.mem [1477] : 
                             (N126)? \nz.mem [1517] : 
                             (N128)? \nz.mem [1557] : 
                             (N130)? \nz.mem [1597] : 
                             (N132)? \nz.mem [1637] : 
                             (N134)? \nz.mem [1677] : 
                             (N136)? \nz.mem [1717] : 
                             (N138)? \nz.mem [1757] : 
                             (N140)? \nz.mem [1797] : 
                             (N142)? \nz.mem [1837] : 
                             (N144)? \nz.mem [1877] : 
                             (N146)? \nz.mem [1917] : 
                             (N148)? \nz.mem [1957] : 
                             (N150)? \nz.mem [1997] : 
                             (N152)? \nz.mem [2037] : 
                             (N154)? \nz.mem [2077] : 
                             (N156)? \nz.mem [2117] : 
                             (N158)? \nz.mem [2157] : 
                             (N160)? \nz.mem [2197] : 
                             (N162)? \nz.mem [2237] : 
                             (N164)? \nz.mem [2277] : 
                             (N166)? \nz.mem [2317] : 
                             (N168)? \nz.mem [2357] : 
                             (N170)? \nz.mem [2397] : 
                             (N172)? \nz.mem [2437] : 
                             (N174)? \nz.mem [2477] : 
                             (N176)? \nz.mem [2517] : 
                             (N178)? \nz.mem [2557] : 1'b0;
  assign \nz.data_out [36] = (N115)? \nz.mem [36] : 
                             (N117)? \nz.mem [76] : 
                             (N119)? \nz.mem [116] : 
                             (N121)? \nz.mem [156] : 
                             (N123)? \nz.mem [196] : 
                             (N125)? \nz.mem [236] : 
                             (N127)? \nz.mem [276] : 
                             (N129)? \nz.mem [316] : 
                             (N131)? \nz.mem [356] : 
                             (N133)? \nz.mem [396] : 
                             (N135)? \nz.mem [436] : 
                             (N137)? \nz.mem [476] : 
                             (N139)? \nz.mem [516] : 
                             (N141)? \nz.mem [556] : 
                             (N143)? \nz.mem [596] : 
                             (N145)? \nz.mem [636] : 
                             (N147)? \nz.mem [676] : 
                             (N149)? \nz.mem [716] : 
                             (N151)? \nz.mem [756] : 
                             (N153)? \nz.mem [796] : 
                             (N155)? \nz.mem [836] : 
                             (N157)? \nz.mem [876] : 
                             (N159)? \nz.mem [916] : 
                             (N161)? \nz.mem [956] : 
                             (N163)? \nz.mem [996] : 
                             (N165)? \nz.mem [1036] : 
                             (N167)? \nz.mem [1076] : 
                             (N169)? \nz.mem [1116] : 
                             (N171)? \nz.mem [1156] : 
                             (N173)? \nz.mem [1196] : 
                             (N175)? \nz.mem [1236] : 
                             (N177)? \nz.mem [1276] : 
                             (N116)? \nz.mem [1316] : 
                             (N118)? \nz.mem [1356] : 
                             (N120)? \nz.mem [1396] : 
                             (N122)? \nz.mem [1436] : 
                             (N124)? \nz.mem [1476] : 
                             (N126)? \nz.mem [1516] : 
                             (N128)? \nz.mem [1556] : 
                             (N130)? \nz.mem [1596] : 
                             (N132)? \nz.mem [1636] : 
                             (N134)? \nz.mem [1676] : 
                             (N136)? \nz.mem [1716] : 
                             (N138)? \nz.mem [1756] : 
                             (N140)? \nz.mem [1796] : 
                             (N142)? \nz.mem [1836] : 
                             (N144)? \nz.mem [1876] : 
                             (N146)? \nz.mem [1916] : 
                             (N148)? \nz.mem [1956] : 
                             (N150)? \nz.mem [1996] : 
                             (N152)? \nz.mem [2036] : 
                             (N154)? \nz.mem [2076] : 
                             (N156)? \nz.mem [2116] : 
                             (N158)? \nz.mem [2156] : 
                             (N160)? \nz.mem [2196] : 
                             (N162)? \nz.mem [2236] : 
                             (N164)? \nz.mem [2276] : 
                             (N166)? \nz.mem [2316] : 
                             (N168)? \nz.mem [2356] : 
                             (N170)? \nz.mem [2396] : 
                             (N172)? \nz.mem [2436] : 
                             (N174)? \nz.mem [2476] : 
                             (N176)? \nz.mem [2516] : 
                             (N178)? \nz.mem [2556] : 1'b0;
  assign \nz.data_out [35] = (N115)? \nz.mem [35] : 
                             (N117)? \nz.mem [75] : 
                             (N119)? \nz.mem [115] : 
                             (N121)? \nz.mem [155] : 
                             (N123)? \nz.mem [195] : 
                             (N125)? \nz.mem [235] : 
                             (N127)? \nz.mem [275] : 
                             (N129)? \nz.mem [315] : 
                             (N131)? \nz.mem [355] : 
                             (N133)? \nz.mem [395] : 
                             (N135)? \nz.mem [435] : 
                             (N137)? \nz.mem [475] : 
                             (N139)? \nz.mem [515] : 
                             (N141)? \nz.mem [555] : 
                             (N143)? \nz.mem [595] : 
                             (N145)? \nz.mem [635] : 
                             (N147)? \nz.mem [675] : 
                             (N149)? \nz.mem [715] : 
                             (N151)? \nz.mem [755] : 
                             (N153)? \nz.mem [795] : 
                             (N155)? \nz.mem [835] : 
                             (N157)? \nz.mem [875] : 
                             (N159)? \nz.mem [915] : 
                             (N161)? \nz.mem [955] : 
                             (N163)? \nz.mem [995] : 
                             (N165)? \nz.mem [1035] : 
                             (N167)? \nz.mem [1075] : 
                             (N169)? \nz.mem [1115] : 
                             (N171)? \nz.mem [1155] : 
                             (N173)? \nz.mem [1195] : 
                             (N175)? \nz.mem [1235] : 
                             (N177)? \nz.mem [1275] : 
                             (N116)? \nz.mem [1315] : 
                             (N118)? \nz.mem [1355] : 
                             (N120)? \nz.mem [1395] : 
                             (N122)? \nz.mem [1435] : 
                             (N124)? \nz.mem [1475] : 
                             (N126)? \nz.mem [1515] : 
                             (N128)? \nz.mem [1555] : 
                             (N130)? \nz.mem [1595] : 
                             (N132)? \nz.mem [1635] : 
                             (N134)? \nz.mem [1675] : 
                             (N136)? \nz.mem [1715] : 
                             (N138)? \nz.mem [1755] : 
                             (N140)? \nz.mem [1795] : 
                             (N142)? \nz.mem [1835] : 
                             (N144)? \nz.mem [1875] : 
                             (N146)? \nz.mem [1915] : 
                             (N148)? \nz.mem [1955] : 
                             (N150)? \nz.mem [1995] : 
                             (N152)? \nz.mem [2035] : 
                             (N154)? \nz.mem [2075] : 
                             (N156)? \nz.mem [2115] : 
                             (N158)? \nz.mem [2155] : 
                             (N160)? \nz.mem [2195] : 
                             (N162)? \nz.mem [2235] : 
                             (N164)? \nz.mem [2275] : 
                             (N166)? \nz.mem [2315] : 
                             (N168)? \nz.mem [2355] : 
                             (N170)? \nz.mem [2395] : 
                             (N172)? \nz.mem [2435] : 
                             (N174)? \nz.mem [2475] : 
                             (N176)? \nz.mem [2515] : 
                             (N178)? \nz.mem [2555] : 1'b0;
  assign \nz.data_out [34] = (N115)? \nz.mem [34] : 
                             (N117)? \nz.mem [74] : 
                             (N119)? \nz.mem [114] : 
                             (N121)? \nz.mem [154] : 
                             (N123)? \nz.mem [194] : 
                             (N125)? \nz.mem [234] : 
                             (N127)? \nz.mem [274] : 
                             (N129)? \nz.mem [314] : 
                             (N131)? \nz.mem [354] : 
                             (N133)? \nz.mem [394] : 
                             (N135)? \nz.mem [434] : 
                             (N137)? \nz.mem [474] : 
                             (N139)? \nz.mem [514] : 
                             (N141)? \nz.mem [554] : 
                             (N143)? \nz.mem [594] : 
                             (N145)? \nz.mem [634] : 
                             (N147)? \nz.mem [674] : 
                             (N149)? \nz.mem [714] : 
                             (N151)? \nz.mem [754] : 
                             (N153)? \nz.mem [794] : 
                             (N155)? \nz.mem [834] : 
                             (N157)? \nz.mem [874] : 
                             (N159)? \nz.mem [914] : 
                             (N161)? \nz.mem [954] : 
                             (N163)? \nz.mem [994] : 
                             (N165)? \nz.mem [1034] : 
                             (N167)? \nz.mem [1074] : 
                             (N169)? \nz.mem [1114] : 
                             (N171)? \nz.mem [1154] : 
                             (N173)? \nz.mem [1194] : 
                             (N175)? \nz.mem [1234] : 
                             (N177)? \nz.mem [1274] : 
                             (N116)? \nz.mem [1314] : 
                             (N118)? \nz.mem [1354] : 
                             (N120)? \nz.mem [1394] : 
                             (N122)? \nz.mem [1434] : 
                             (N124)? \nz.mem [1474] : 
                             (N126)? \nz.mem [1514] : 
                             (N128)? \nz.mem [1554] : 
                             (N130)? \nz.mem [1594] : 
                             (N132)? \nz.mem [1634] : 
                             (N134)? \nz.mem [1674] : 
                             (N136)? \nz.mem [1714] : 
                             (N138)? \nz.mem [1754] : 
                             (N140)? \nz.mem [1794] : 
                             (N142)? \nz.mem [1834] : 
                             (N144)? \nz.mem [1874] : 
                             (N146)? \nz.mem [1914] : 
                             (N148)? \nz.mem [1954] : 
                             (N150)? \nz.mem [1994] : 
                             (N152)? \nz.mem [2034] : 
                             (N154)? \nz.mem [2074] : 
                             (N156)? \nz.mem [2114] : 
                             (N158)? \nz.mem [2154] : 
                             (N160)? \nz.mem [2194] : 
                             (N162)? \nz.mem [2234] : 
                             (N164)? \nz.mem [2274] : 
                             (N166)? \nz.mem [2314] : 
                             (N168)? \nz.mem [2354] : 
                             (N170)? \nz.mem [2394] : 
                             (N172)? \nz.mem [2434] : 
                             (N174)? \nz.mem [2474] : 
                             (N176)? \nz.mem [2514] : 
                             (N178)? \nz.mem [2554] : 1'b0;
  assign \nz.data_out [33] = (N115)? \nz.mem [33] : 
                             (N117)? \nz.mem [73] : 
                             (N119)? \nz.mem [113] : 
                             (N121)? \nz.mem [153] : 
                             (N123)? \nz.mem [193] : 
                             (N125)? \nz.mem [233] : 
                             (N127)? \nz.mem [273] : 
                             (N129)? \nz.mem [313] : 
                             (N131)? \nz.mem [353] : 
                             (N133)? \nz.mem [393] : 
                             (N135)? \nz.mem [433] : 
                             (N137)? \nz.mem [473] : 
                             (N139)? \nz.mem [513] : 
                             (N141)? \nz.mem [553] : 
                             (N143)? \nz.mem [593] : 
                             (N145)? \nz.mem [633] : 
                             (N147)? \nz.mem [673] : 
                             (N149)? \nz.mem [713] : 
                             (N151)? \nz.mem [753] : 
                             (N153)? \nz.mem [793] : 
                             (N155)? \nz.mem [833] : 
                             (N157)? \nz.mem [873] : 
                             (N159)? \nz.mem [913] : 
                             (N161)? \nz.mem [953] : 
                             (N163)? \nz.mem [993] : 
                             (N165)? \nz.mem [1033] : 
                             (N167)? \nz.mem [1073] : 
                             (N169)? \nz.mem [1113] : 
                             (N171)? \nz.mem [1153] : 
                             (N173)? \nz.mem [1193] : 
                             (N175)? \nz.mem [1233] : 
                             (N177)? \nz.mem [1273] : 
                             (N116)? \nz.mem [1313] : 
                             (N118)? \nz.mem [1353] : 
                             (N120)? \nz.mem [1393] : 
                             (N122)? \nz.mem [1433] : 
                             (N124)? \nz.mem [1473] : 
                             (N126)? \nz.mem [1513] : 
                             (N128)? \nz.mem [1553] : 
                             (N130)? \nz.mem [1593] : 
                             (N132)? \nz.mem [1633] : 
                             (N134)? \nz.mem [1673] : 
                             (N136)? \nz.mem [1713] : 
                             (N138)? \nz.mem [1753] : 
                             (N140)? \nz.mem [1793] : 
                             (N142)? \nz.mem [1833] : 
                             (N144)? \nz.mem [1873] : 
                             (N146)? \nz.mem [1913] : 
                             (N148)? \nz.mem [1953] : 
                             (N150)? \nz.mem [1993] : 
                             (N152)? \nz.mem [2033] : 
                             (N154)? \nz.mem [2073] : 
                             (N156)? \nz.mem [2113] : 
                             (N158)? \nz.mem [2153] : 
                             (N160)? \nz.mem [2193] : 
                             (N162)? \nz.mem [2233] : 
                             (N164)? \nz.mem [2273] : 
                             (N166)? \nz.mem [2313] : 
                             (N168)? \nz.mem [2353] : 
                             (N170)? \nz.mem [2393] : 
                             (N172)? \nz.mem [2433] : 
                             (N174)? \nz.mem [2473] : 
                             (N176)? \nz.mem [2513] : 
                             (N178)? \nz.mem [2553] : 1'b0;
  assign \nz.data_out [32] = (N115)? \nz.mem [32] : 
                             (N117)? \nz.mem [72] : 
                             (N119)? \nz.mem [112] : 
                             (N121)? \nz.mem [152] : 
                             (N123)? \nz.mem [192] : 
                             (N125)? \nz.mem [232] : 
                             (N127)? \nz.mem [272] : 
                             (N129)? \nz.mem [312] : 
                             (N131)? \nz.mem [352] : 
                             (N133)? \nz.mem [392] : 
                             (N135)? \nz.mem [432] : 
                             (N137)? \nz.mem [472] : 
                             (N139)? \nz.mem [512] : 
                             (N141)? \nz.mem [552] : 
                             (N143)? \nz.mem [592] : 
                             (N145)? \nz.mem [632] : 
                             (N147)? \nz.mem [672] : 
                             (N149)? \nz.mem [712] : 
                             (N151)? \nz.mem [752] : 
                             (N153)? \nz.mem [792] : 
                             (N155)? \nz.mem [832] : 
                             (N157)? \nz.mem [872] : 
                             (N159)? \nz.mem [912] : 
                             (N161)? \nz.mem [952] : 
                             (N163)? \nz.mem [992] : 
                             (N165)? \nz.mem [1032] : 
                             (N167)? \nz.mem [1072] : 
                             (N169)? \nz.mem [1112] : 
                             (N171)? \nz.mem [1152] : 
                             (N173)? \nz.mem [1192] : 
                             (N175)? \nz.mem [1232] : 
                             (N177)? \nz.mem [1272] : 
                             (N116)? \nz.mem [1312] : 
                             (N118)? \nz.mem [1352] : 
                             (N120)? \nz.mem [1392] : 
                             (N122)? \nz.mem [1432] : 
                             (N124)? \nz.mem [1472] : 
                             (N126)? \nz.mem [1512] : 
                             (N128)? \nz.mem [1552] : 
                             (N130)? \nz.mem [1592] : 
                             (N132)? \nz.mem [1632] : 
                             (N134)? \nz.mem [1672] : 
                             (N136)? \nz.mem [1712] : 
                             (N138)? \nz.mem [1752] : 
                             (N140)? \nz.mem [1792] : 
                             (N142)? \nz.mem [1832] : 
                             (N144)? \nz.mem [1872] : 
                             (N146)? \nz.mem [1912] : 
                             (N148)? \nz.mem [1952] : 
                             (N150)? \nz.mem [1992] : 
                             (N152)? \nz.mem [2032] : 
                             (N154)? \nz.mem [2072] : 
                             (N156)? \nz.mem [2112] : 
                             (N158)? \nz.mem [2152] : 
                             (N160)? \nz.mem [2192] : 
                             (N162)? \nz.mem [2232] : 
                             (N164)? \nz.mem [2272] : 
                             (N166)? \nz.mem [2312] : 
                             (N168)? \nz.mem [2352] : 
                             (N170)? \nz.mem [2392] : 
                             (N172)? \nz.mem [2432] : 
                             (N174)? \nz.mem [2472] : 
                             (N176)? \nz.mem [2512] : 
                             (N178)? \nz.mem [2552] : 1'b0;
  assign \nz.data_out [31] = (N115)? \nz.mem [31] : 
                             (N117)? \nz.mem [71] : 
                             (N119)? \nz.mem [111] : 
                             (N121)? \nz.mem [151] : 
                             (N123)? \nz.mem [191] : 
                             (N125)? \nz.mem [231] : 
                             (N127)? \nz.mem [271] : 
                             (N129)? \nz.mem [311] : 
                             (N131)? \nz.mem [351] : 
                             (N133)? \nz.mem [391] : 
                             (N135)? \nz.mem [431] : 
                             (N137)? \nz.mem [471] : 
                             (N139)? \nz.mem [511] : 
                             (N141)? \nz.mem [551] : 
                             (N143)? \nz.mem [591] : 
                             (N145)? \nz.mem [631] : 
                             (N147)? \nz.mem [671] : 
                             (N149)? \nz.mem [711] : 
                             (N151)? \nz.mem [751] : 
                             (N153)? \nz.mem [791] : 
                             (N155)? \nz.mem [831] : 
                             (N157)? \nz.mem [871] : 
                             (N159)? \nz.mem [911] : 
                             (N161)? \nz.mem [951] : 
                             (N163)? \nz.mem [991] : 
                             (N165)? \nz.mem [1031] : 
                             (N167)? \nz.mem [1071] : 
                             (N169)? \nz.mem [1111] : 
                             (N171)? \nz.mem [1151] : 
                             (N173)? \nz.mem [1191] : 
                             (N175)? \nz.mem [1231] : 
                             (N177)? \nz.mem [1271] : 
                             (N116)? \nz.mem [1311] : 
                             (N118)? \nz.mem [1351] : 
                             (N120)? \nz.mem [1391] : 
                             (N122)? \nz.mem [1431] : 
                             (N124)? \nz.mem [1471] : 
                             (N126)? \nz.mem [1511] : 
                             (N128)? \nz.mem [1551] : 
                             (N130)? \nz.mem [1591] : 
                             (N132)? \nz.mem [1631] : 
                             (N134)? \nz.mem [1671] : 
                             (N136)? \nz.mem [1711] : 
                             (N138)? \nz.mem [1751] : 
                             (N140)? \nz.mem [1791] : 
                             (N142)? \nz.mem [1831] : 
                             (N144)? \nz.mem [1871] : 
                             (N146)? \nz.mem [1911] : 
                             (N148)? \nz.mem [1951] : 
                             (N150)? \nz.mem [1991] : 
                             (N152)? \nz.mem [2031] : 
                             (N154)? \nz.mem [2071] : 
                             (N156)? \nz.mem [2111] : 
                             (N158)? \nz.mem [2151] : 
                             (N160)? \nz.mem [2191] : 
                             (N162)? \nz.mem [2231] : 
                             (N164)? \nz.mem [2271] : 
                             (N166)? \nz.mem [2311] : 
                             (N168)? \nz.mem [2351] : 
                             (N170)? \nz.mem [2391] : 
                             (N172)? \nz.mem [2431] : 
                             (N174)? \nz.mem [2471] : 
                             (N176)? \nz.mem [2511] : 
                             (N178)? \nz.mem [2551] : 1'b0;
  assign \nz.data_out [30] = (N115)? \nz.mem [30] : 
                             (N117)? \nz.mem [70] : 
                             (N119)? \nz.mem [110] : 
                             (N121)? \nz.mem [150] : 
                             (N123)? \nz.mem [190] : 
                             (N125)? \nz.mem [230] : 
                             (N127)? \nz.mem [270] : 
                             (N129)? \nz.mem [310] : 
                             (N131)? \nz.mem [350] : 
                             (N133)? \nz.mem [390] : 
                             (N135)? \nz.mem [430] : 
                             (N137)? \nz.mem [470] : 
                             (N139)? \nz.mem [510] : 
                             (N141)? \nz.mem [550] : 
                             (N143)? \nz.mem [590] : 
                             (N145)? \nz.mem [630] : 
                             (N147)? \nz.mem [670] : 
                             (N149)? \nz.mem [710] : 
                             (N151)? \nz.mem [750] : 
                             (N153)? \nz.mem [790] : 
                             (N155)? \nz.mem [830] : 
                             (N157)? \nz.mem [870] : 
                             (N159)? \nz.mem [910] : 
                             (N161)? \nz.mem [950] : 
                             (N163)? \nz.mem [990] : 
                             (N165)? \nz.mem [1030] : 
                             (N167)? \nz.mem [1070] : 
                             (N169)? \nz.mem [1110] : 
                             (N171)? \nz.mem [1150] : 
                             (N173)? \nz.mem [1190] : 
                             (N175)? \nz.mem [1230] : 
                             (N177)? \nz.mem [1270] : 
                             (N116)? \nz.mem [1310] : 
                             (N118)? \nz.mem [1350] : 
                             (N120)? \nz.mem [1390] : 
                             (N122)? \nz.mem [1430] : 
                             (N124)? \nz.mem [1470] : 
                             (N126)? \nz.mem [1510] : 
                             (N128)? \nz.mem [1550] : 
                             (N130)? \nz.mem [1590] : 
                             (N132)? \nz.mem [1630] : 
                             (N134)? \nz.mem [1670] : 
                             (N136)? \nz.mem [1710] : 
                             (N138)? \nz.mem [1750] : 
                             (N140)? \nz.mem [1790] : 
                             (N142)? \nz.mem [1830] : 
                             (N144)? \nz.mem [1870] : 
                             (N146)? \nz.mem [1910] : 
                             (N148)? \nz.mem [1950] : 
                             (N150)? \nz.mem [1990] : 
                             (N152)? \nz.mem [2030] : 
                             (N154)? \nz.mem [2070] : 
                             (N156)? \nz.mem [2110] : 
                             (N158)? \nz.mem [2150] : 
                             (N160)? \nz.mem [2190] : 
                             (N162)? \nz.mem [2230] : 
                             (N164)? \nz.mem [2270] : 
                             (N166)? \nz.mem [2310] : 
                             (N168)? \nz.mem [2350] : 
                             (N170)? \nz.mem [2390] : 
                             (N172)? \nz.mem [2430] : 
                             (N174)? \nz.mem [2470] : 
                             (N176)? \nz.mem [2510] : 
                             (N178)? \nz.mem [2550] : 1'b0;
  assign \nz.data_out [29] = (N115)? \nz.mem [29] : 
                             (N117)? \nz.mem [69] : 
                             (N119)? \nz.mem [109] : 
                             (N121)? \nz.mem [149] : 
                             (N123)? \nz.mem [189] : 
                             (N125)? \nz.mem [229] : 
                             (N127)? \nz.mem [269] : 
                             (N129)? \nz.mem [309] : 
                             (N131)? \nz.mem [349] : 
                             (N133)? \nz.mem [389] : 
                             (N135)? \nz.mem [429] : 
                             (N137)? \nz.mem [469] : 
                             (N139)? \nz.mem [509] : 
                             (N141)? \nz.mem [549] : 
                             (N143)? \nz.mem [589] : 
                             (N145)? \nz.mem [629] : 
                             (N147)? \nz.mem [669] : 
                             (N149)? \nz.mem [709] : 
                             (N151)? \nz.mem [749] : 
                             (N153)? \nz.mem [789] : 
                             (N155)? \nz.mem [829] : 
                             (N157)? \nz.mem [869] : 
                             (N159)? \nz.mem [909] : 
                             (N161)? \nz.mem [949] : 
                             (N163)? \nz.mem [989] : 
                             (N165)? \nz.mem [1029] : 
                             (N167)? \nz.mem [1069] : 
                             (N169)? \nz.mem [1109] : 
                             (N171)? \nz.mem [1149] : 
                             (N173)? \nz.mem [1189] : 
                             (N175)? \nz.mem [1229] : 
                             (N177)? \nz.mem [1269] : 
                             (N116)? \nz.mem [1309] : 
                             (N118)? \nz.mem [1349] : 
                             (N120)? \nz.mem [1389] : 
                             (N122)? \nz.mem [1429] : 
                             (N124)? \nz.mem [1469] : 
                             (N126)? \nz.mem [1509] : 
                             (N128)? \nz.mem [1549] : 
                             (N130)? \nz.mem [1589] : 
                             (N132)? \nz.mem [1629] : 
                             (N134)? \nz.mem [1669] : 
                             (N136)? \nz.mem [1709] : 
                             (N138)? \nz.mem [1749] : 
                             (N140)? \nz.mem [1789] : 
                             (N142)? \nz.mem [1829] : 
                             (N144)? \nz.mem [1869] : 
                             (N146)? \nz.mem [1909] : 
                             (N148)? \nz.mem [1949] : 
                             (N150)? \nz.mem [1989] : 
                             (N152)? \nz.mem [2029] : 
                             (N154)? \nz.mem [2069] : 
                             (N156)? \nz.mem [2109] : 
                             (N158)? \nz.mem [2149] : 
                             (N160)? \nz.mem [2189] : 
                             (N162)? \nz.mem [2229] : 
                             (N164)? \nz.mem [2269] : 
                             (N166)? \nz.mem [2309] : 
                             (N168)? \nz.mem [2349] : 
                             (N170)? \nz.mem [2389] : 
                             (N172)? \nz.mem [2429] : 
                             (N174)? \nz.mem [2469] : 
                             (N176)? \nz.mem [2509] : 
                             (N178)? \nz.mem [2549] : 1'b0;
  assign \nz.data_out [28] = (N115)? \nz.mem [28] : 
                             (N117)? \nz.mem [68] : 
                             (N119)? \nz.mem [108] : 
                             (N121)? \nz.mem [148] : 
                             (N123)? \nz.mem [188] : 
                             (N125)? \nz.mem [228] : 
                             (N127)? \nz.mem [268] : 
                             (N129)? \nz.mem [308] : 
                             (N131)? \nz.mem [348] : 
                             (N133)? \nz.mem [388] : 
                             (N135)? \nz.mem [428] : 
                             (N137)? \nz.mem [468] : 
                             (N139)? \nz.mem [508] : 
                             (N141)? \nz.mem [548] : 
                             (N143)? \nz.mem [588] : 
                             (N145)? \nz.mem [628] : 
                             (N147)? \nz.mem [668] : 
                             (N149)? \nz.mem [708] : 
                             (N151)? \nz.mem [748] : 
                             (N153)? \nz.mem [788] : 
                             (N155)? \nz.mem [828] : 
                             (N157)? \nz.mem [868] : 
                             (N159)? \nz.mem [908] : 
                             (N161)? \nz.mem [948] : 
                             (N163)? \nz.mem [988] : 
                             (N165)? \nz.mem [1028] : 
                             (N167)? \nz.mem [1068] : 
                             (N169)? \nz.mem [1108] : 
                             (N171)? \nz.mem [1148] : 
                             (N173)? \nz.mem [1188] : 
                             (N175)? \nz.mem [1228] : 
                             (N177)? \nz.mem [1268] : 
                             (N116)? \nz.mem [1308] : 
                             (N118)? \nz.mem [1348] : 
                             (N120)? \nz.mem [1388] : 
                             (N122)? \nz.mem [1428] : 
                             (N124)? \nz.mem [1468] : 
                             (N126)? \nz.mem [1508] : 
                             (N128)? \nz.mem [1548] : 
                             (N130)? \nz.mem [1588] : 
                             (N132)? \nz.mem [1628] : 
                             (N134)? \nz.mem [1668] : 
                             (N136)? \nz.mem [1708] : 
                             (N138)? \nz.mem [1748] : 
                             (N140)? \nz.mem [1788] : 
                             (N142)? \nz.mem [1828] : 
                             (N144)? \nz.mem [1868] : 
                             (N146)? \nz.mem [1908] : 
                             (N148)? \nz.mem [1948] : 
                             (N150)? \nz.mem [1988] : 
                             (N152)? \nz.mem [2028] : 
                             (N154)? \nz.mem [2068] : 
                             (N156)? \nz.mem [2108] : 
                             (N158)? \nz.mem [2148] : 
                             (N160)? \nz.mem [2188] : 
                             (N162)? \nz.mem [2228] : 
                             (N164)? \nz.mem [2268] : 
                             (N166)? \nz.mem [2308] : 
                             (N168)? \nz.mem [2348] : 
                             (N170)? \nz.mem [2388] : 
                             (N172)? \nz.mem [2428] : 
                             (N174)? \nz.mem [2468] : 
                             (N176)? \nz.mem [2508] : 
                             (N178)? \nz.mem [2548] : 1'b0;
  assign \nz.data_out [27] = (N115)? \nz.mem [27] : 
                             (N117)? \nz.mem [67] : 
                             (N119)? \nz.mem [107] : 
                             (N121)? \nz.mem [147] : 
                             (N123)? \nz.mem [187] : 
                             (N125)? \nz.mem [227] : 
                             (N127)? \nz.mem [267] : 
                             (N129)? \nz.mem [307] : 
                             (N131)? \nz.mem [347] : 
                             (N133)? \nz.mem [387] : 
                             (N135)? \nz.mem [427] : 
                             (N137)? \nz.mem [467] : 
                             (N139)? \nz.mem [507] : 
                             (N141)? \nz.mem [547] : 
                             (N143)? \nz.mem [587] : 
                             (N145)? \nz.mem [627] : 
                             (N147)? \nz.mem [667] : 
                             (N149)? \nz.mem [707] : 
                             (N151)? \nz.mem [747] : 
                             (N153)? \nz.mem [787] : 
                             (N155)? \nz.mem [827] : 
                             (N157)? \nz.mem [867] : 
                             (N159)? \nz.mem [907] : 
                             (N161)? \nz.mem [947] : 
                             (N163)? \nz.mem [987] : 
                             (N165)? \nz.mem [1027] : 
                             (N167)? \nz.mem [1067] : 
                             (N169)? \nz.mem [1107] : 
                             (N171)? \nz.mem [1147] : 
                             (N173)? \nz.mem [1187] : 
                             (N175)? \nz.mem [1227] : 
                             (N177)? \nz.mem [1267] : 
                             (N116)? \nz.mem [1307] : 
                             (N118)? \nz.mem [1347] : 
                             (N120)? \nz.mem [1387] : 
                             (N122)? \nz.mem [1427] : 
                             (N124)? \nz.mem [1467] : 
                             (N126)? \nz.mem [1507] : 
                             (N128)? \nz.mem [1547] : 
                             (N130)? \nz.mem [1587] : 
                             (N132)? \nz.mem [1627] : 
                             (N134)? \nz.mem [1667] : 
                             (N136)? \nz.mem [1707] : 
                             (N138)? \nz.mem [1747] : 
                             (N140)? \nz.mem [1787] : 
                             (N142)? \nz.mem [1827] : 
                             (N144)? \nz.mem [1867] : 
                             (N146)? \nz.mem [1907] : 
                             (N148)? \nz.mem [1947] : 
                             (N150)? \nz.mem [1987] : 
                             (N152)? \nz.mem [2027] : 
                             (N154)? \nz.mem [2067] : 
                             (N156)? \nz.mem [2107] : 
                             (N158)? \nz.mem [2147] : 
                             (N160)? \nz.mem [2187] : 
                             (N162)? \nz.mem [2227] : 
                             (N164)? \nz.mem [2267] : 
                             (N166)? \nz.mem [2307] : 
                             (N168)? \nz.mem [2347] : 
                             (N170)? \nz.mem [2387] : 
                             (N172)? \nz.mem [2427] : 
                             (N174)? \nz.mem [2467] : 
                             (N176)? \nz.mem [2507] : 
                             (N178)? \nz.mem [2547] : 1'b0;
  assign \nz.data_out [26] = (N115)? \nz.mem [26] : 
                             (N117)? \nz.mem [66] : 
                             (N119)? \nz.mem [106] : 
                             (N121)? \nz.mem [146] : 
                             (N123)? \nz.mem [186] : 
                             (N125)? \nz.mem [226] : 
                             (N127)? \nz.mem [266] : 
                             (N129)? \nz.mem [306] : 
                             (N131)? \nz.mem [346] : 
                             (N133)? \nz.mem [386] : 
                             (N135)? \nz.mem [426] : 
                             (N137)? \nz.mem [466] : 
                             (N139)? \nz.mem [506] : 
                             (N141)? \nz.mem [546] : 
                             (N143)? \nz.mem [586] : 
                             (N145)? \nz.mem [626] : 
                             (N147)? \nz.mem [666] : 
                             (N149)? \nz.mem [706] : 
                             (N151)? \nz.mem [746] : 
                             (N153)? \nz.mem [786] : 
                             (N155)? \nz.mem [826] : 
                             (N157)? \nz.mem [866] : 
                             (N159)? \nz.mem [906] : 
                             (N161)? \nz.mem [946] : 
                             (N163)? \nz.mem [986] : 
                             (N165)? \nz.mem [1026] : 
                             (N167)? \nz.mem [1066] : 
                             (N169)? \nz.mem [1106] : 
                             (N171)? \nz.mem [1146] : 
                             (N173)? \nz.mem [1186] : 
                             (N175)? \nz.mem [1226] : 
                             (N177)? \nz.mem [1266] : 
                             (N116)? \nz.mem [1306] : 
                             (N118)? \nz.mem [1346] : 
                             (N120)? \nz.mem [1386] : 
                             (N122)? \nz.mem [1426] : 
                             (N124)? \nz.mem [1466] : 
                             (N126)? \nz.mem [1506] : 
                             (N128)? \nz.mem [1546] : 
                             (N130)? \nz.mem [1586] : 
                             (N132)? \nz.mem [1626] : 
                             (N134)? \nz.mem [1666] : 
                             (N136)? \nz.mem [1706] : 
                             (N138)? \nz.mem [1746] : 
                             (N140)? \nz.mem [1786] : 
                             (N142)? \nz.mem [1826] : 
                             (N144)? \nz.mem [1866] : 
                             (N146)? \nz.mem [1906] : 
                             (N148)? \nz.mem [1946] : 
                             (N150)? \nz.mem [1986] : 
                             (N152)? \nz.mem [2026] : 
                             (N154)? \nz.mem [2066] : 
                             (N156)? \nz.mem [2106] : 
                             (N158)? \nz.mem [2146] : 
                             (N160)? \nz.mem [2186] : 
                             (N162)? \nz.mem [2226] : 
                             (N164)? \nz.mem [2266] : 
                             (N166)? \nz.mem [2306] : 
                             (N168)? \nz.mem [2346] : 
                             (N170)? \nz.mem [2386] : 
                             (N172)? \nz.mem [2426] : 
                             (N174)? \nz.mem [2466] : 
                             (N176)? \nz.mem [2506] : 
                             (N178)? \nz.mem [2546] : 1'b0;
  assign \nz.data_out [25] = (N115)? \nz.mem [25] : 
                             (N117)? \nz.mem [65] : 
                             (N119)? \nz.mem [105] : 
                             (N121)? \nz.mem [145] : 
                             (N123)? \nz.mem [185] : 
                             (N125)? \nz.mem [225] : 
                             (N127)? \nz.mem [265] : 
                             (N129)? \nz.mem [305] : 
                             (N131)? \nz.mem [345] : 
                             (N133)? \nz.mem [385] : 
                             (N135)? \nz.mem [425] : 
                             (N137)? \nz.mem [465] : 
                             (N139)? \nz.mem [505] : 
                             (N141)? \nz.mem [545] : 
                             (N143)? \nz.mem [585] : 
                             (N145)? \nz.mem [625] : 
                             (N147)? \nz.mem [665] : 
                             (N149)? \nz.mem [705] : 
                             (N151)? \nz.mem [745] : 
                             (N153)? \nz.mem [785] : 
                             (N155)? \nz.mem [825] : 
                             (N157)? \nz.mem [865] : 
                             (N159)? \nz.mem [905] : 
                             (N161)? \nz.mem [945] : 
                             (N163)? \nz.mem [985] : 
                             (N165)? \nz.mem [1025] : 
                             (N167)? \nz.mem [1065] : 
                             (N169)? \nz.mem [1105] : 
                             (N171)? \nz.mem [1145] : 
                             (N173)? \nz.mem [1185] : 
                             (N175)? \nz.mem [1225] : 
                             (N177)? \nz.mem [1265] : 
                             (N116)? \nz.mem [1305] : 
                             (N118)? \nz.mem [1345] : 
                             (N120)? \nz.mem [1385] : 
                             (N122)? \nz.mem [1425] : 
                             (N124)? \nz.mem [1465] : 
                             (N126)? \nz.mem [1505] : 
                             (N128)? \nz.mem [1545] : 
                             (N130)? \nz.mem [1585] : 
                             (N132)? \nz.mem [1625] : 
                             (N134)? \nz.mem [1665] : 
                             (N136)? \nz.mem [1705] : 
                             (N138)? \nz.mem [1745] : 
                             (N140)? \nz.mem [1785] : 
                             (N142)? \nz.mem [1825] : 
                             (N144)? \nz.mem [1865] : 
                             (N146)? \nz.mem [1905] : 
                             (N148)? \nz.mem [1945] : 
                             (N150)? \nz.mem [1985] : 
                             (N152)? \nz.mem [2025] : 
                             (N154)? \nz.mem [2065] : 
                             (N156)? \nz.mem [2105] : 
                             (N158)? \nz.mem [2145] : 
                             (N160)? \nz.mem [2185] : 
                             (N162)? \nz.mem [2225] : 
                             (N164)? \nz.mem [2265] : 
                             (N166)? \nz.mem [2305] : 
                             (N168)? \nz.mem [2345] : 
                             (N170)? \nz.mem [2385] : 
                             (N172)? \nz.mem [2425] : 
                             (N174)? \nz.mem [2465] : 
                             (N176)? \nz.mem [2505] : 
                             (N178)? \nz.mem [2545] : 1'b0;
  assign \nz.data_out [24] = (N115)? \nz.mem [24] : 
                             (N117)? \nz.mem [64] : 
                             (N119)? \nz.mem [104] : 
                             (N121)? \nz.mem [144] : 
                             (N123)? \nz.mem [184] : 
                             (N125)? \nz.mem [224] : 
                             (N127)? \nz.mem [264] : 
                             (N129)? \nz.mem [304] : 
                             (N131)? \nz.mem [344] : 
                             (N133)? \nz.mem [384] : 
                             (N135)? \nz.mem [424] : 
                             (N137)? \nz.mem [464] : 
                             (N139)? \nz.mem [504] : 
                             (N141)? \nz.mem [544] : 
                             (N143)? \nz.mem [584] : 
                             (N145)? \nz.mem [624] : 
                             (N147)? \nz.mem [664] : 
                             (N149)? \nz.mem [704] : 
                             (N151)? \nz.mem [744] : 
                             (N153)? \nz.mem [784] : 
                             (N155)? \nz.mem [824] : 
                             (N157)? \nz.mem [864] : 
                             (N159)? \nz.mem [904] : 
                             (N161)? \nz.mem [944] : 
                             (N163)? \nz.mem [984] : 
                             (N165)? \nz.mem [1024] : 
                             (N167)? \nz.mem [1064] : 
                             (N169)? \nz.mem [1104] : 
                             (N171)? \nz.mem [1144] : 
                             (N173)? \nz.mem [1184] : 
                             (N175)? \nz.mem [1224] : 
                             (N177)? \nz.mem [1264] : 
                             (N116)? \nz.mem [1304] : 
                             (N118)? \nz.mem [1344] : 
                             (N120)? \nz.mem [1384] : 
                             (N122)? \nz.mem [1424] : 
                             (N124)? \nz.mem [1464] : 
                             (N126)? \nz.mem [1504] : 
                             (N128)? \nz.mem [1544] : 
                             (N130)? \nz.mem [1584] : 
                             (N132)? \nz.mem [1624] : 
                             (N134)? \nz.mem [1664] : 
                             (N136)? \nz.mem [1704] : 
                             (N138)? \nz.mem [1744] : 
                             (N140)? \nz.mem [1784] : 
                             (N142)? \nz.mem [1824] : 
                             (N144)? \nz.mem [1864] : 
                             (N146)? \nz.mem [1904] : 
                             (N148)? \nz.mem [1944] : 
                             (N150)? \nz.mem [1984] : 
                             (N152)? \nz.mem [2024] : 
                             (N154)? \nz.mem [2064] : 
                             (N156)? \nz.mem [2104] : 
                             (N158)? \nz.mem [2144] : 
                             (N160)? \nz.mem [2184] : 
                             (N162)? \nz.mem [2224] : 
                             (N164)? \nz.mem [2264] : 
                             (N166)? \nz.mem [2304] : 
                             (N168)? \nz.mem [2344] : 
                             (N170)? \nz.mem [2384] : 
                             (N172)? \nz.mem [2424] : 
                             (N174)? \nz.mem [2464] : 
                             (N176)? \nz.mem [2504] : 
                             (N178)? \nz.mem [2544] : 1'b0;
  assign \nz.data_out [23] = (N115)? \nz.mem [23] : 
                             (N117)? \nz.mem [63] : 
                             (N119)? \nz.mem [103] : 
                             (N121)? \nz.mem [143] : 
                             (N123)? \nz.mem [183] : 
                             (N125)? \nz.mem [223] : 
                             (N127)? \nz.mem [263] : 
                             (N129)? \nz.mem [303] : 
                             (N131)? \nz.mem [343] : 
                             (N133)? \nz.mem [383] : 
                             (N135)? \nz.mem [423] : 
                             (N137)? \nz.mem [463] : 
                             (N139)? \nz.mem [503] : 
                             (N141)? \nz.mem [543] : 
                             (N143)? \nz.mem [583] : 
                             (N145)? \nz.mem [623] : 
                             (N147)? \nz.mem [663] : 
                             (N149)? \nz.mem [703] : 
                             (N151)? \nz.mem [743] : 
                             (N153)? \nz.mem [783] : 
                             (N155)? \nz.mem [823] : 
                             (N157)? \nz.mem [863] : 
                             (N159)? \nz.mem [903] : 
                             (N161)? \nz.mem [943] : 
                             (N163)? \nz.mem [983] : 
                             (N165)? \nz.mem [1023] : 
                             (N167)? \nz.mem [1063] : 
                             (N169)? \nz.mem [1103] : 
                             (N171)? \nz.mem [1143] : 
                             (N173)? \nz.mem [1183] : 
                             (N175)? \nz.mem [1223] : 
                             (N177)? \nz.mem [1263] : 
                             (N116)? \nz.mem [1303] : 
                             (N118)? \nz.mem [1343] : 
                             (N120)? \nz.mem [1383] : 
                             (N122)? \nz.mem [1423] : 
                             (N124)? \nz.mem [1463] : 
                             (N126)? \nz.mem [1503] : 
                             (N128)? \nz.mem [1543] : 
                             (N130)? \nz.mem [1583] : 
                             (N132)? \nz.mem [1623] : 
                             (N134)? \nz.mem [1663] : 
                             (N136)? \nz.mem [1703] : 
                             (N138)? \nz.mem [1743] : 
                             (N140)? \nz.mem [1783] : 
                             (N142)? \nz.mem [1823] : 
                             (N144)? \nz.mem [1863] : 
                             (N146)? \nz.mem [1903] : 
                             (N148)? \nz.mem [1943] : 
                             (N150)? \nz.mem [1983] : 
                             (N152)? \nz.mem [2023] : 
                             (N154)? \nz.mem [2063] : 
                             (N156)? \nz.mem [2103] : 
                             (N158)? \nz.mem [2143] : 
                             (N160)? \nz.mem [2183] : 
                             (N162)? \nz.mem [2223] : 
                             (N164)? \nz.mem [2263] : 
                             (N166)? \nz.mem [2303] : 
                             (N168)? \nz.mem [2343] : 
                             (N170)? \nz.mem [2383] : 
                             (N172)? \nz.mem [2423] : 
                             (N174)? \nz.mem [2463] : 
                             (N176)? \nz.mem [2503] : 
                             (N178)? \nz.mem [2543] : 1'b0;
  assign \nz.data_out [22] = (N115)? \nz.mem [22] : 
                             (N117)? \nz.mem [62] : 
                             (N119)? \nz.mem [102] : 
                             (N121)? \nz.mem [142] : 
                             (N123)? \nz.mem [182] : 
                             (N125)? \nz.mem [222] : 
                             (N127)? \nz.mem [262] : 
                             (N129)? \nz.mem [302] : 
                             (N131)? \nz.mem [342] : 
                             (N133)? \nz.mem [382] : 
                             (N135)? \nz.mem [422] : 
                             (N137)? \nz.mem [462] : 
                             (N139)? \nz.mem [502] : 
                             (N141)? \nz.mem [542] : 
                             (N143)? \nz.mem [582] : 
                             (N145)? \nz.mem [622] : 
                             (N147)? \nz.mem [662] : 
                             (N149)? \nz.mem [702] : 
                             (N151)? \nz.mem [742] : 
                             (N153)? \nz.mem [782] : 
                             (N155)? \nz.mem [822] : 
                             (N157)? \nz.mem [862] : 
                             (N159)? \nz.mem [902] : 
                             (N161)? \nz.mem [942] : 
                             (N163)? \nz.mem [982] : 
                             (N165)? \nz.mem [1022] : 
                             (N167)? \nz.mem [1062] : 
                             (N169)? \nz.mem [1102] : 
                             (N171)? \nz.mem [1142] : 
                             (N173)? \nz.mem [1182] : 
                             (N175)? \nz.mem [1222] : 
                             (N177)? \nz.mem [1262] : 
                             (N116)? \nz.mem [1302] : 
                             (N118)? \nz.mem [1342] : 
                             (N120)? \nz.mem [1382] : 
                             (N122)? \nz.mem [1422] : 
                             (N124)? \nz.mem [1462] : 
                             (N126)? \nz.mem [1502] : 
                             (N128)? \nz.mem [1542] : 
                             (N130)? \nz.mem [1582] : 
                             (N132)? \nz.mem [1622] : 
                             (N134)? \nz.mem [1662] : 
                             (N136)? \nz.mem [1702] : 
                             (N138)? \nz.mem [1742] : 
                             (N140)? \nz.mem [1782] : 
                             (N142)? \nz.mem [1822] : 
                             (N144)? \nz.mem [1862] : 
                             (N146)? \nz.mem [1902] : 
                             (N148)? \nz.mem [1942] : 
                             (N150)? \nz.mem [1982] : 
                             (N152)? \nz.mem [2022] : 
                             (N154)? \nz.mem [2062] : 
                             (N156)? \nz.mem [2102] : 
                             (N158)? \nz.mem [2142] : 
                             (N160)? \nz.mem [2182] : 
                             (N162)? \nz.mem [2222] : 
                             (N164)? \nz.mem [2262] : 
                             (N166)? \nz.mem [2302] : 
                             (N168)? \nz.mem [2342] : 
                             (N170)? \nz.mem [2382] : 
                             (N172)? \nz.mem [2422] : 
                             (N174)? \nz.mem [2462] : 
                             (N176)? \nz.mem [2502] : 
                             (N178)? \nz.mem [2542] : 1'b0;
  assign \nz.data_out [21] = (N115)? \nz.mem [21] : 
                             (N117)? \nz.mem [61] : 
                             (N119)? \nz.mem [101] : 
                             (N121)? \nz.mem [141] : 
                             (N123)? \nz.mem [181] : 
                             (N125)? \nz.mem [221] : 
                             (N127)? \nz.mem [261] : 
                             (N129)? \nz.mem [301] : 
                             (N131)? \nz.mem [341] : 
                             (N133)? \nz.mem [381] : 
                             (N135)? \nz.mem [421] : 
                             (N137)? \nz.mem [461] : 
                             (N139)? \nz.mem [501] : 
                             (N141)? \nz.mem [541] : 
                             (N143)? \nz.mem [581] : 
                             (N145)? \nz.mem [621] : 
                             (N147)? \nz.mem [661] : 
                             (N149)? \nz.mem [701] : 
                             (N151)? \nz.mem [741] : 
                             (N153)? \nz.mem [781] : 
                             (N155)? \nz.mem [821] : 
                             (N157)? \nz.mem [861] : 
                             (N159)? \nz.mem [901] : 
                             (N161)? \nz.mem [941] : 
                             (N163)? \nz.mem [981] : 
                             (N165)? \nz.mem [1021] : 
                             (N167)? \nz.mem [1061] : 
                             (N169)? \nz.mem [1101] : 
                             (N171)? \nz.mem [1141] : 
                             (N173)? \nz.mem [1181] : 
                             (N175)? \nz.mem [1221] : 
                             (N177)? \nz.mem [1261] : 
                             (N116)? \nz.mem [1301] : 
                             (N118)? \nz.mem [1341] : 
                             (N120)? \nz.mem [1381] : 
                             (N122)? \nz.mem [1421] : 
                             (N124)? \nz.mem [1461] : 
                             (N126)? \nz.mem [1501] : 
                             (N128)? \nz.mem [1541] : 
                             (N130)? \nz.mem [1581] : 
                             (N132)? \nz.mem [1621] : 
                             (N134)? \nz.mem [1661] : 
                             (N136)? \nz.mem [1701] : 
                             (N138)? \nz.mem [1741] : 
                             (N140)? \nz.mem [1781] : 
                             (N142)? \nz.mem [1821] : 
                             (N144)? \nz.mem [1861] : 
                             (N146)? \nz.mem [1901] : 
                             (N148)? \nz.mem [1941] : 
                             (N150)? \nz.mem [1981] : 
                             (N152)? \nz.mem [2021] : 
                             (N154)? \nz.mem [2061] : 
                             (N156)? \nz.mem [2101] : 
                             (N158)? \nz.mem [2141] : 
                             (N160)? \nz.mem [2181] : 
                             (N162)? \nz.mem [2221] : 
                             (N164)? \nz.mem [2261] : 
                             (N166)? \nz.mem [2301] : 
                             (N168)? \nz.mem [2341] : 
                             (N170)? \nz.mem [2381] : 
                             (N172)? \nz.mem [2421] : 
                             (N174)? \nz.mem [2461] : 
                             (N176)? \nz.mem [2501] : 
                             (N178)? \nz.mem [2541] : 1'b0;
  assign \nz.data_out [20] = (N115)? \nz.mem [20] : 
                             (N117)? \nz.mem [60] : 
                             (N119)? \nz.mem [100] : 
                             (N121)? \nz.mem [140] : 
                             (N123)? \nz.mem [180] : 
                             (N125)? \nz.mem [220] : 
                             (N127)? \nz.mem [260] : 
                             (N129)? \nz.mem [300] : 
                             (N131)? \nz.mem [340] : 
                             (N133)? \nz.mem [380] : 
                             (N135)? \nz.mem [420] : 
                             (N137)? \nz.mem [460] : 
                             (N139)? \nz.mem [500] : 
                             (N141)? \nz.mem [540] : 
                             (N143)? \nz.mem [580] : 
                             (N145)? \nz.mem [620] : 
                             (N147)? \nz.mem [660] : 
                             (N149)? \nz.mem [700] : 
                             (N151)? \nz.mem [740] : 
                             (N153)? \nz.mem [780] : 
                             (N155)? \nz.mem [820] : 
                             (N157)? \nz.mem [860] : 
                             (N159)? \nz.mem [900] : 
                             (N161)? \nz.mem [940] : 
                             (N163)? \nz.mem [980] : 
                             (N165)? \nz.mem [1020] : 
                             (N167)? \nz.mem [1060] : 
                             (N169)? \nz.mem [1100] : 
                             (N171)? \nz.mem [1140] : 
                             (N173)? \nz.mem [1180] : 
                             (N175)? \nz.mem [1220] : 
                             (N177)? \nz.mem [1260] : 
                             (N116)? \nz.mem [1300] : 
                             (N118)? \nz.mem [1340] : 
                             (N120)? \nz.mem [1380] : 
                             (N122)? \nz.mem [1420] : 
                             (N124)? \nz.mem [1460] : 
                             (N126)? \nz.mem [1500] : 
                             (N128)? \nz.mem [1540] : 
                             (N130)? \nz.mem [1580] : 
                             (N132)? \nz.mem [1620] : 
                             (N134)? \nz.mem [1660] : 
                             (N136)? \nz.mem [1700] : 
                             (N138)? \nz.mem [1740] : 
                             (N140)? \nz.mem [1780] : 
                             (N142)? \nz.mem [1820] : 
                             (N144)? \nz.mem [1860] : 
                             (N146)? \nz.mem [1900] : 
                             (N148)? \nz.mem [1940] : 
                             (N150)? \nz.mem [1980] : 
                             (N152)? \nz.mem [2020] : 
                             (N154)? \nz.mem [2060] : 
                             (N156)? \nz.mem [2100] : 
                             (N158)? \nz.mem [2140] : 
                             (N160)? \nz.mem [2180] : 
                             (N162)? \nz.mem [2220] : 
                             (N164)? \nz.mem [2260] : 
                             (N166)? \nz.mem [2300] : 
                             (N168)? \nz.mem [2340] : 
                             (N170)? \nz.mem [2380] : 
                             (N172)? \nz.mem [2420] : 
                             (N174)? \nz.mem [2460] : 
                             (N176)? \nz.mem [2500] : 
                             (N178)? \nz.mem [2540] : 1'b0;
  assign \nz.data_out [19] = (N115)? \nz.mem [19] : 
                             (N117)? \nz.mem [59] : 
                             (N119)? \nz.mem [99] : 
                             (N121)? \nz.mem [139] : 
                             (N123)? \nz.mem [179] : 
                             (N125)? \nz.mem [219] : 
                             (N127)? \nz.mem [259] : 
                             (N129)? \nz.mem [299] : 
                             (N131)? \nz.mem [339] : 
                             (N133)? \nz.mem [379] : 
                             (N135)? \nz.mem [419] : 
                             (N137)? \nz.mem [459] : 
                             (N139)? \nz.mem [499] : 
                             (N141)? \nz.mem [539] : 
                             (N143)? \nz.mem [579] : 
                             (N145)? \nz.mem [619] : 
                             (N147)? \nz.mem [659] : 
                             (N149)? \nz.mem [699] : 
                             (N151)? \nz.mem [739] : 
                             (N153)? \nz.mem [779] : 
                             (N155)? \nz.mem [819] : 
                             (N157)? \nz.mem [859] : 
                             (N159)? \nz.mem [899] : 
                             (N161)? \nz.mem [939] : 
                             (N163)? \nz.mem [979] : 
                             (N165)? \nz.mem [1019] : 
                             (N167)? \nz.mem [1059] : 
                             (N169)? \nz.mem [1099] : 
                             (N171)? \nz.mem [1139] : 
                             (N173)? \nz.mem [1179] : 
                             (N175)? \nz.mem [1219] : 
                             (N177)? \nz.mem [1259] : 
                             (N116)? \nz.mem [1299] : 
                             (N118)? \nz.mem [1339] : 
                             (N120)? \nz.mem [1379] : 
                             (N122)? \nz.mem [1419] : 
                             (N124)? \nz.mem [1459] : 
                             (N126)? \nz.mem [1499] : 
                             (N128)? \nz.mem [1539] : 
                             (N130)? \nz.mem [1579] : 
                             (N132)? \nz.mem [1619] : 
                             (N134)? \nz.mem [1659] : 
                             (N136)? \nz.mem [1699] : 
                             (N138)? \nz.mem [1739] : 
                             (N140)? \nz.mem [1779] : 
                             (N142)? \nz.mem [1819] : 
                             (N144)? \nz.mem [1859] : 
                             (N146)? \nz.mem [1899] : 
                             (N148)? \nz.mem [1939] : 
                             (N150)? \nz.mem [1979] : 
                             (N152)? \nz.mem [2019] : 
                             (N154)? \nz.mem [2059] : 
                             (N156)? \nz.mem [2099] : 
                             (N158)? \nz.mem [2139] : 
                             (N160)? \nz.mem [2179] : 
                             (N162)? \nz.mem [2219] : 
                             (N164)? \nz.mem [2259] : 
                             (N166)? \nz.mem [2299] : 
                             (N168)? \nz.mem [2339] : 
                             (N170)? \nz.mem [2379] : 
                             (N172)? \nz.mem [2419] : 
                             (N174)? \nz.mem [2459] : 
                             (N176)? \nz.mem [2499] : 
                             (N178)? \nz.mem [2539] : 1'b0;
  assign \nz.data_out [18] = (N115)? \nz.mem [18] : 
                             (N117)? \nz.mem [58] : 
                             (N119)? \nz.mem [98] : 
                             (N121)? \nz.mem [138] : 
                             (N123)? \nz.mem [178] : 
                             (N125)? \nz.mem [218] : 
                             (N127)? \nz.mem [258] : 
                             (N129)? \nz.mem [298] : 
                             (N131)? \nz.mem [338] : 
                             (N133)? \nz.mem [378] : 
                             (N135)? \nz.mem [418] : 
                             (N137)? \nz.mem [458] : 
                             (N139)? \nz.mem [498] : 
                             (N141)? \nz.mem [538] : 
                             (N143)? \nz.mem [578] : 
                             (N145)? \nz.mem [618] : 
                             (N147)? \nz.mem [658] : 
                             (N149)? \nz.mem [698] : 
                             (N151)? \nz.mem [738] : 
                             (N153)? \nz.mem [778] : 
                             (N155)? \nz.mem [818] : 
                             (N157)? \nz.mem [858] : 
                             (N159)? \nz.mem [898] : 
                             (N161)? \nz.mem [938] : 
                             (N163)? \nz.mem [978] : 
                             (N165)? \nz.mem [1018] : 
                             (N167)? \nz.mem [1058] : 
                             (N169)? \nz.mem [1098] : 
                             (N171)? \nz.mem [1138] : 
                             (N173)? \nz.mem [1178] : 
                             (N175)? \nz.mem [1218] : 
                             (N177)? \nz.mem [1258] : 
                             (N116)? \nz.mem [1298] : 
                             (N118)? \nz.mem [1338] : 
                             (N120)? \nz.mem [1378] : 
                             (N122)? \nz.mem [1418] : 
                             (N124)? \nz.mem [1458] : 
                             (N126)? \nz.mem [1498] : 
                             (N128)? \nz.mem [1538] : 
                             (N130)? \nz.mem [1578] : 
                             (N132)? \nz.mem [1618] : 
                             (N134)? \nz.mem [1658] : 
                             (N136)? \nz.mem [1698] : 
                             (N138)? \nz.mem [1738] : 
                             (N140)? \nz.mem [1778] : 
                             (N142)? \nz.mem [1818] : 
                             (N144)? \nz.mem [1858] : 
                             (N146)? \nz.mem [1898] : 
                             (N148)? \nz.mem [1938] : 
                             (N150)? \nz.mem [1978] : 
                             (N152)? \nz.mem [2018] : 
                             (N154)? \nz.mem [2058] : 
                             (N156)? \nz.mem [2098] : 
                             (N158)? \nz.mem [2138] : 
                             (N160)? \nz.mem [2178] : 
                             (N162)? \nz.mem [2218] : 
                             (N164)? \nz.mem [2258] : 
                             (N166)? \nz.mem [2298] : 
                             (N168)? \nz.mem [2338] : 
                             (N170)? \nz.mem [2378] : 
                             (N172)? \nz.mem [2418] : 
                             (N174)? \nz.mem [2458] : 
                             (N176)? \nz.mem [2498] : 
                             (N178)? \nz.mem [2538] : 1'b0;
  assign \nz.data_out [17] = (N115)? \nz.mem [17] : 
                             (N117)? \nz.mem [57] : 
                             (N119)? \nz.mem [97] : 
                             (N121)? \nz.mem [137] : 
                             (N123)? \nz.mem [177] : 
                             (N125)? \nz.mem [217] : 
                             (N127)? \nz.mem [257] : 
                             (N129)? \nz.mem [297] : 
                             (N131)? \nz.mem [337] : 
                             (N133)? \nz.mem [377] : 
                             (N135)? \nz.mem [417] : 
                             (N137)? \nz.mem [457] : 
                             (N139)? \nz.mem [497] : 
                             (N141)? \nz.mem [537] : 
                             (N143)? \nz.mem [577] : 
                             (N145)? \nz.mem [617] : 
                             (N147)? \nz.mem [657] : 
                             (N149)? \nz.mem [697] : 
                             (N151)? \nz.mem [737] : 
                             (N153)? \nz.mem [777] : 
                             (N155)? \nz.mem [817] : 
                             (N157)? \nz.mem [857] : 
                             (N159)? \nz.mem [897] : 
                             (N161)? \nz.mem [937] : 
                             (N163)? \nz.mem [977] : 
                             (N165)? \nz.mem [1017] : 
                             (N167)? \nz.mem [1057] : 
                             (N169)? \nz.mem [1097] : 
                             (N171)? \nz.mem [1137] : 
                             (N173)? \nz.mem [1177] : 
                             (N175)? \nz.mem [1217] : 
                             (N177)? \nz.mem [1257] : 
                             (N116)? \nz.mem [1297] : 
                             (N118)? \nz.mem [1337] : 
                             (N120)? \nz.mem [1377] : 
                             (N122)? \nz.mem [1417] : 
                             (N124)? \nz.mem [1457] : 
                             (N126)? \nz.mem [1497] : 
                             (N128)? \nz.mem [1537] : 
                             (N130)? \nz.mem [1577] : 
                             (N132)? \nz.mem [1617] : 
                             (N134)? \nz.mem [1657] : 
                             (N136)? \nz.mem [1697] : 
                             (N138)? \nz.mem [1737] : 
                             (N140)? \nz.mem [1777] : 
                             (N142)? \nz.mem [1817] : 
                             (N144)? \nz.mem [1857] : 
                             (N146)? \nz.mem [1897] : 
                             (N148)? \nz.mem [1937] : 
                             (N150)? \nz.mem [1977] : 
                             (N152)? \nz.mem [2017] : 
                             (N154)? \nz.mem [2057] : 
                             (N156)? \nz.mem [2097] : 
                             (N158)? \nz.mem [2137] : 
                             (N160)? \nz.mem [2177] : 
                             (N162)? \nz.mem [2217] : 
                             (N164)? \nz.mem [2257] : 
                             (N166)? \nz.mem [2297] : 
                             (N168)? \nz.mem [2337] : 
                             (N170)? \nz.mem [2377] : 
                             (N172)? \nz.mem [2417] : 
                             (N174)? \nz.mem [2457] : 
                             (N176)? \nz.mem [2497] : 
                             (N178)? \nz.mem [2537] : 1'b0;
  assign \nz.data_out [16] = (N115)? \nz.mem [16] : 
                             (N117)? \nz.mem [56] : 
                             (N119)? \nz.mem [96] : 
                             (N121)? \nz.mem [136] : 
                             (N123)? \nz.mem [176] : 
                             (N125)? \nz.mem [216] : 
                             (N127)? \nz.mem [256] : 
                             (N129)? \nz.mem [296] : 
                             (N131)? \nz.mem [336] : 
                             (N133)? \nz.mem [376] : 
                             (N135)? \nz.mem [416] : 
                             (N137)? \nz.mem [456] : 
                             (N139)? \nz.mem [496] : 
                             (N141)? \nz.mem [536] : 
                             (N143)? \nz.mem [576] : 
                             (N145)? \nz.mem [616] : 
                             (N147)? \nz.mem [656] : 
                             (N149)? \nz.mem [696] : 
                             (N151)? \nz.mem [736] : 
                             (N153)? \nz.mem [776] : 
                             (N155)? \nz.mem [816] : 
                             (N157)? \nz.mem [856] : 
                             (N159)? \nz.mem [896] : 
                             (N161)? \nz.mem [936] : 
                             (N163)? \nz.mem [976] : 
                             (N165)? \nz.mem [1016] : 
                             (N167)? \nz.mem [1056] : 
                             (N169)? \nz.mem [1096] : 
                             (N171)? \nz.mem [1136] : 
                             (N173)? \nz.mem [1176] : 
                             (N175)? \nz.mem [1216] : 
                             (N177)? \nz.mem [1256] : 
                             (N116)? \nz.mem [1296] : 
                             (N118)? \nz.mem [1336] : 
                             (N120)? \nz.mem [1376] : 
                             (N122)? \nz.mem [1416] : 
                             (N124)? \nz.mem [1456] : 
                             (N126)? \nz.mem [1496] : 
                             (N128)? \nz.mem [1536] : 
                             (N130)? \nz.mem [1576] : 
                             (N132)? \nz.mem [1616] : 
                             (N134)? \nz.mem [1656] : 
                             (N136)? \nz.mem [1696] : 
                             (N138)? \nz.mem [1736] : 
                             (N140)? \nz.mem [1776] : 
                             (N142)? \nz.mem [1816] : 
                             (N144)? \nz.mem [1856] : 
                             (N146)? \nz.mem [1896] : 
                             (N148)? \nz.mem [1936] : 
                             (N150)? \nz.mem [1976] : 
                             (N152)? \nz.mem [2016] : 
                             (N154)? \nz.mem [2056] : 
                             (N156)? \nz.mem [2096] : 
                             (N158)? \nz.mem [2136] : 
                             (N160)? \nz.mem [2176] : 
                             (N162)? \nz.mem [2216] : 
                             (N164)? \nz.mem [2256] : 
                             (N166)? \nz.mem [2296] : 
                             (N168)? \nz.mem [2336] : 
                             (N170)? \nz.mem [2376] : 
                             (N172)? \nz.mem [2416] : 
                             (N174)? \nz.mem [2456] : 
                             (N176)? \nz.mem [2496] : 
                             (N178)? \nz.mem [2536] : 1'b0;
  assign \nz.data_out [15] = (N115)? \nz.mem [15] : 
                             (N117)? \nz.mem [55] : 
                             (N119)? \nz.mem [95] : 
                             (N121)? \nz.mem [135] : 
                             (N123)? \nz.mem [175] : 
                             (N125)? \nz.mem [215] : 
                             (N127)? \nz.mem [255] : 
                             (N129)? \nz.mem [295] : 
                             (N131)? \nz.mem [335] : 
                             (N133)? \nz.mem [375] : 
                             (N135)? \nz.mem [415] : 
                             (N137)? \nz.mem [455] : 
                             (N139)? \nz.mem [495] : 
                             (N141)? \nz.mem [535] : 
                             (N143)? \nz.mem [575] : 
                             (N145)? \nz.mem [615] : 
                             (N147)? \nz.mem [655] : 
                             (N149)? \nz.mem [695] : 
                             (N151)? \nz.mem [735] : 
                             (N153)? \nz.mem [775] : 
                             (N155)? \nz.mem [815] : 
                             (N157)? \nz.mem [855] : 
                             (N159)? \nz.mem [895] : 
                             (N161)? \nz.mem [935] : 
                             (N163)? \nz.mem [975] : 
                             (N165)? \nz.mem [1015] : 
                             (N167)? \nz.mem [1055] : 
                             (N169)? \nz.mem [1095] : 
                             (N171)? \nz.mem [1135] : 
                             (N173)? \nz.mem [1175] : 
                             (N175)? \nz.mem [1215] : 
                             (N177)? \nz.mem [1255] : 
                             (N116)? \nz.mem [1295] : 
                             (N118)? \nz.mem [1335] : 
                             (N120)? \nz.mem [1375] : 
                             (N122)? \nz.mem [1415] : 
                             (N124)? \nz.mem [1455] : 
                             (N126)? \nz.mem [1495] : 
                             (N128)? \nz.mem [1535] : 
                             (N130)? \nz.mem [1575] : 
                             (N132)? \nz.mem [1615] : 
                             (N134)? \nz.mem [1655] : 
                             (N136)? \nz.mem [1695] : 
                             (N138)? \nz.mem [1735] : 
                             (N140)? \nz.mem [1775] : 
                             (N142)? \nz.mem [1815] : 
                             (N144)? \nz.mem [1855] : 
                             (N146)? \nz.mem [1895] : 
                             (N148)? \nz.mem [1935] : 
                             (N150)? \nz.mem [1975] : 
                             (N152)? \nz.mem [2015] : 
                             (N154)? \nz.mem [2055] : 
                             (N156)? \nz.mem [2095] : 
                             (N158)? \nz.mem [2135] : 
                             (N160)? \nz.mem [2175] : 
                             (N162)? \nz.mem [2215] : 
                             (N164)? \nz.mem [2255] : 
                             (N166)? \nz.mem [2295] : 
                             (N168)? \nz.mem [2335] : 
                             (N170)? \nz.mem [2375] : 
                             (N172)? \nz.mem [2415] : 
                             (N174)? \nz.mem [2455] : 
                             (N176)? \nz.mem [2495] : 
                             (N178)? \nz.mem [2535] : 1'b0;
  assign \nz.data_out [14] = (N115)? \nz.mem [14] : 
                             (N117)? \nz.mem [54] : 
                             (N119)? \nz.mem [94] : 
                             (N121)? \nz.mem [134] : 
                             (N123)? \nz.mem [174] : 
                             (N125)? \nz.mem [214] : 
                             (N127)? \nz.mem [254] : 
                             (N129)? \nz.mem [294] : 
                             (N131)? \nz.mem [334] : 
                             (N133)? \nz.mem [374] : 
                             (N135)? \nz.mem [414] : 
                             (N137)? \nz.mem [454] : 
                             (N139)? \nz.mem [494] : 
                             (N141)? \nz.mem [534] : 
                             (N143)? \nz.mem [574] : 
                             (N145)? \nz.mem [614] : 
                             (N147)? \nz.mem [654] : 
                             (N149)? \nz.mem [694] : 
                             (N151)? \nz.mem [734] : 
                             (N153)? \nz.mem [774] : 
                             (N155)? \nz.mem [814] : 
                             (N157)? \nz.mem [854] : 
                             (N159)? \nz.mem [894] : 
                             (N161)? \nz.mem [934] : 
                             (N163)? \nz.mem [974] : 
                             (N165)? \nz.mem [1014] : 
                             (N167)? \nz.mem [1054] : 
                             (N169)? \nz.mem [1094] : 
                             (N171)? \nz.mem [1134] : 
                             (N173)? \nz.mem [1174] : 
                             (N175)? \nz.mem [1214] : 
                             (N177)? \nz.mem [1254] : 
                             (N116)? \nz.mem [1294] : 
                             (N118)? \nz.mem [1334] : 
                             (N120)? \nz.mem [1374] : 
                             (N122)? \nz.mem [1414] : 
                             (N124)? \nz.mem [1454] : 
                             (N126)? \nz.mem [1494] : 
                             (N128)? \nz.mem [1534] : 
                             (N130)? \nz.mem [1574] : 
                             (N132)? \nz.mem [1614] : 
                             (N134)? \nz.mem [1654] : 
                             (N136)? \nz.mem [1694] : 
                             (N138)? \nz.mem [1734] : 
                             (N140)? \nz.mem [1774] : 
                             (N142)? \nz.mem [1814] : 
                             (N144)? \nz.mem [1854] : 
                             (N146)? \nz.mem [1894] : 
                             (N148)? \nz.mem [1934] : 
                             (N150)? \nz.mem [1974] : 
                             (N152)? \nz.mem [2014] : 
                             (N154)? \nz.mem [2054] : 
                             (N156)? \nz.mem [2094] : 
                             (N158)? \nz.mem [2134] : 
                             (N160)? \nz.mem [2174] : 
                             (N162)? \nz.mem [2214] : 
                             (N164)? \nz.mem [2254] : 
                             (N166)? \nz.mem [2294] : 
                             (N168)? \nz.mem [2334] : 
                             (N170)? \nz.mem [2374] : 
                             (N172)? \nz.mem [2414] : 
                             (N174)? \nz.mem [2454] : 
                             (N176)? \nz.mem [2494] : 
                             (N178)? \nz.mem [2534] : 1'b0;
  assign \nz.data_out [13] = (N115)? \nz.mem [13] : 
                             (N117)? \nz.mem [53] : 
                             (N119)? \nz.mem [93] : 
                             (N121)? \nz.mem [133] : 
                             (N123)? \nz.mem [173] : 
                             (N125)? \nz.mem [213] : 
                             (N127)? \nz.mem [253] : 
                             (N129)? \nz.mem [293] : 
                             (N131)? \nz.mem [333] : 
                             (N133)? \nz.mem [373] : 
                             (N135)? \nz.mem [413] : 
                             (N137)? \nz.mem [453] : 
                             (N139)? \nz.mem [493] : 
                             (N141)? \nz.mem [533] : 
                             (N143)? \nz.mem [573] : 
                             (N145)? \nz.mem [613] : 
                             (N147)? \nz.mem [653] : 
                             (N149)? \nz.mem [693] : 
                             (N151)? \nz.mem [733] : 
                             (N153)? \nz.mem [773] : 
                             (N155)? \nz.mem [813] : 
                             (N157)? \nz.mem [853] : 
                             (N159)? \nz.mem [893] : 
                             (N161)? \nz.mem [933] : 
                             (N163)? \nz.mem [973] : 
                             (N165)? \nz.mem [1013] : 
                             (N167)? \nz.mem [1053] : 
                             (N169)? \nz.mem [1093] : 
                             (N171)? \nz.mem [1133] : 
                             (N173)? \nz.mem [1173] : 
                             (N175)? \nz.mem [1213] : 
                             (N177)? \nz.mem [1253] : 
                             (N116)? \nz.mem [1293] : 
                             (N118)? \nz.mem [1333] : 
                             (N120)? \nz.mem [1373] : 
                             (N122)? \nz.mem [1413] : 
                             (N124)? \nz.mem [1453] : 
                             (N126)? \nz.mem [1493] : 
                             (N128)? \nz.mem [1533] : 
                             (N130)? \nz.mem [1573] : 
                             (N132)? \nz.mem [1613] : 
                             (N134)? \nz.mem [1653] : 
                             (N136)? \nz.mem [1693] : 
                             (N138)? \nz.mem [1733] : 
                             (N140)? \nz.mem [1773] : 
                             (N142)? \nz.mem [1813] : 
                             (N144)? \nz.mem [1853] : 
                             (N146)? \nz.mem [1893] : 
                             (N148)? \nz.mem [1933] : 
                             (N150)? \nz.mem [1973] : 
                             (N152)? \nz.mem [2013] : 
                             (N154)? \nz.mem [2053] : 
                             (N156)? \nz.mem [2093] : 
                             (N158)? \nz.mem [2133] : 
                             (N160)? \nz.mem [2173] : 
                             (N162)? \nz.mem [2213] : 
                             (N164)? \nz.mem [2253] : 
                             (N166)? \nz.mem [2293] : 
                             (N168)? \nz.mem [2333] : 
                             (N170)? \nz.mem [2373] : 
                             (N172)? \nz.mem [2413] : 
                             (N174)? \nz.mem [2453] : 
                             (N176)? \nz.mem [2493] : 
                             (N178)? \nz.mem [2533] : 1'b0;
  assign \nz.data_out [12] = (N115)? \nz.mem [12] : 
                             (N117)? \nz.mem [52] : 
                             (N119)? \nz.mem [92] : 
                             (N121)? \nz.mem [132] : 
                             (N123)? \nz.mem [172] : 
                             (N125)? \nz.mem [212] : 
                             (N127)? \nz.mem [252] : 
                             (N129)? \nz.mem [292] : 
                             (N131)? \nz.mem [332] : 
                             (N133)? \nz.mem [372] : 
                             (N135)? \nz.mem [412] : 
                             (N137)? \nz.mem [452] : 
                             (N139)? \nz.mem [492] : 
                             (N141)? \nz.mem [532] : 
                             (N143)? \nz.mem [572] : 
                             (N145)? \nz.mem [612] : 
                             (N147)? \nz.mem [652] : 
                             (N149)? \nz.mem [692] : 
                             (N151)? \nz.mem [732] : 
                             (N153)? \nz.mem [772] : 
                             (N155)? \nz.mem [812] : 
                             (N157)? \nz.mem [852] : 
                             (N159)? \nz.mem [892] : 
                             (N161)? \nz.mem [932] : 
                             (N163)? \nz.mem [972] : 
                             (N165)? \nz.mem [1012] : 
                             (N167)? \nz.mem [1052] : 
                             (N169)? \nz.mem [1092] : 
                             (N171)? \nz.mem [1132] : 
                             (N173)? \nz.mem [1172] : 
                             (N175)? \nz.mem [1212] : 
                             (N177)? \nz.mem [1252] : 
                             (N116)? \nz.mem [1292] : 
                             (N118)? \nz.mem [1332] : 
                             (N120)? \nz.mem [1372] : 
                             (N122)? \nz.mem [1412] : 
                             (N124)? \nz.mem [1452] : 
                             (N126)? \nz.mem [1492] : 
                             (N128)? \nz.mem [1532] : 
                             (N130)? \nz.mem [1572] : 
                             (N132)? \nz.mem [1612] : 
                             (N134)? \nz.mem [1652] : 
                             (N136)? \nz.mem [1692] : 
                             (N138)? \nz.mem [1732] : 
                             (N140)? \nz.mem [1772] : 
                             (N142)? \nz.mem [1812] : 
                             (N144)? \nz.mem [1852] : 
                             (N146)? \nz.mem [1892] : 
                             (N148)? \nz.mem [1932] : 
                             (N150)? \nz.mem [1972] : 
                             (N152)? \nz.mem [2012] : 
                             (N154)? \nz.mem [2052] : 
                             (N156)? \nz.mem [2092] : 
                             (N158)? \nz.mem [2132] : 
                             (N160)? \nz.mem [2172] : 
                             (N162)? \nz.mem [2212] : 
                             (N164)? \nz.mem [2252] : 
                             (N166)? \nz.mem [2292] : 
                             (N168)? \nz.mem [2332] : 
                             (N170)? \nz.mem [2372] : 
                             (N172)? \nz.mem [2412] : 
                             (N174)? \nz.mem [2452] : 
                             (N176)? \nz.mem [2492] : 
                             (N178)? \nz.mem [2532] : 1'b0;
  assign \nz.data_out [11] = (N115)? \nz.mem [11] : 
                             (N117)? \nz.mem [51] : 
                             (N119)? \nz.mem [91] : 
                             (N121)? \nz.mem [131] : 
                             (N123)? \nz.mem [171] : 
                             (N125)? \nz.mem [211] : 
                             (N127)? \nz.mem [251] : 
                             (N129)? \nz.mem [291] : 
                             (N131)? \nz.mem [331] : 
                             (N133)? \nz.mem [371] : 
                             (N135)? \nz.mem [411] : 
                             (N137)? \nz.mem [451] : 
                             (N139)? \nz.mem [491] : 
                             (N141)? \nz.mem [531] : 
                             (N143)? \nz.mem [571] : 
                             (N145)? \nz.mem [611] : 
                             (N147)? \nz.mem [651] : 
                             (N149)? \nz.mem [691] : 
                             (N151)? \nz.mem [731] : 
                             (N153)? \nz.mem [771] : 
                             (N155)? \nz.mem [811] : 
                             (N157)? \nz.mem [851] : 
                             (N159)? \nz.mem [891] : 
                             (N161)? \nz.mem [931] : 
                             (N163)? \nz.mem [971] : 
                             (N165)? \nz.mem [1011] : 
                             (N167)? \nz.mem [1051] : 
                             (N169)? \nz.mem [1091] : 
                             (N171)? \nz.mem [1131] : 
                             (N173)? \nz.mem [1171] : 
                             (N175)? \nz.mem [1211] : 
                             (N177)? \nz.mem [1251] : 
                             (N116)? \nz.mem [1291] : 
                             (N118)? \nz.mem [1331] : 
                             (N120)? \nz.mem [1371] : 
                             (N122)? \nz.mem [1411] : 
                             (N124)? \nz.mem [1451] : 
                             (N126)? \nz.mem [1491] : 
                             (N128)? \nz.mem [1531] : 
                             (N130)? \nz.mem [1571] : 
                             (N132)? \nz.mem [1611] : 
                             (N134)? \nz.mem [1651] : 
                             (N136)? \nz.mem [1691] : 
                             (N138)? \nz.mem [1731] : 
                             (N140)? \nz.mem [1771] : 
                             (N142)? \nz.mem [1811] : 
                             (N144)? \nz.mem [1851] : 
                             (N146)? \nz.mem [1891] : 
                             (N148)? \nz.mem [1931] : 
                             (N150)? \nz.mem [1971] : 
                             (N152)? \nz.mem [2011] : 
                             (N154)? \nz.mem [2051] : 
                             (N156)? \nz.mem [2091] : 
                             (N158)? \nz.mem [2131] : 
                             (N160)? \nz.mem [2171] : 
                             (N162)? \nz.mem [2211] : 
                             (N164)? \nz.mem [2251] : 
                             (N166)? \nz.mem [2291] : 
                             (N168)? \nz.mem [2331] : 
                             (N170)? \nz.mem [2371] : 
                             (N172)? \nz.mem [2411] : 
                             (N174)? \nz.mem [2451] : 
                             (N176)? \nz.mem [2491] : 
                             (N178)? \nz.mem [2531] : 1'b0;
  assign \nz.data_out [10] = (N115)? \nz.mem [10] : 
                             (N117)? \nz.mem [50] : 
                             (N119)? \nz.mem [90] : 
                             (N121)? \nz.mem [130] : 
                             (N123)? \nz.mem [170] : 
                             (N125)? \nz.mem [210] : 
                             (N127)? \nz.mem [250] : 
                             (N129)? \nz.mem [290] : 
                             (N131)? \nz.mem [330] : 
                             (N133)? \nz.mem [370] : 
                             (N135)? \nz.mem [410] : 
                             (N137)? \nz.mem [450] : 
                             (N139)? \nz.mem [490] : 
                             (N141)? \nz.mem [530] : 
                             (N143)? \nz.mem [570] : 
                             (N145)? \nz.mem [610] : 
                             (N147)? \nz.mem [650] : 
                             (N149)? \nz.mem [690] : 
                             (N151)? \nz.mem [730] : 
                             (N153)? \nz.mem [770] : 
                             (N155)? \nz.mem [810] : 
                             (N157)? \nz.mem [850] : 
                             (N159)? \nz.mem [890] : 
                             (N161)? \nz.mem [930] : 
                             (N163)? \nz.mem [970] : 
                             (N165)? \nz.mem [1010] : 
                             (N167)? \nz.mem [1050] : 
                             (N169)? \nz.mem [1090] : 
                             (N171)? \nz.mem [1130] : 
                             (N173)? \nz.mem [1170] : 
                             (N175)? \nz.mem [1210] : 
                             (N177)? \nz.mem [1250] : 
                             (N116)? \nz.mem [1290] : 
                             (N118)? \nz.mem [1330] : 
                             (N120)? \nz.mem [1370] : 
                             (N122)? \nz.mem [1410] : 
                             (N124)? \nz.mem [1450] : 
                             (N126)? \nz.mem [1490] : 
                             (N128)? \nz.mem [1530] : 
                             (N130)? \nz.mem [1570] : 
                             (N132)? \nz.mem [1610] : 
                             (N134)? \nz.mem [1650] : 
                             (N136)? \nz.mem [1690] : 
                             (N138)? \nz.mem [1730] : 
                             (N140)? \nz.mem [1770] : 
                             (N142)? \nz.mem [1810] : 
                             (N144)? \nz.mem [1850] : 
                             (N146)? \nz.mem [1890] : 
                             (N148)? \nz.mem [1930] : 
                             (N150)? \nz.mem [1970] : 
                             (N152)? \nz.mem [2010] : 
                             (N154)? \nz.mem [2050] : 
                             (N156)? \nz.mem [2090] : 
                             (N158)? \nz.mem [2130] : 
                             (N160)? \nz.mem [2170] : 
                             (N162)? \nz.mem [2210] : 
                             (N164)? \nz.mem [2250] : 
                             (N166)? \nz.mem [2290] : 
                             (N168)? \nz.mem [2330] : 
                             (N170)? \nz.mem [2370] : 
                             (N172)? \nz.mem [2410] : 
                             (N174)? \nz.mem [2450] : 
                             (N176)? \nz.mem [2490] : 
                             (N178)? \nz.mem [2530] : 1'b0;
  assign \nz.data_out [9] = (N115)? \nz.mem [9] : 
                            (N117)? \nz.mem [49] : 
                            (N119)? \nz.mem [89] : 
                            (N121)? \nz.mem [129] : 
                            (N123)? \nz.mem [169] : 
                            (N125)? \nz.mem [209] : 
                            (N127)? \nz.mem [249] : 
                            (N129)? \nz.mem [289] : 
                            (N131)? \nz.mem [329] : 
                            (N133)? \nz.mem [369] : 
                            (N135)? \nz.mem [409] : 
                            (N137)? \nz.mem [449] : 
                            (N139)? \nz.mem [489] : 
                            (N141)? \nz.mem [529] : 
                            (N143)? \nz.mem [569] : 
                            (N145)? \nz.mem [609] : 
                            (N147)? \nz.mem [649] : 
                            (N149)? \nz.mem [689] : 
                            (N151)? \nz.mem [729] : 
                            (N153)? \nz.mem [769] : 
                            (N155)? \nz.mem [809] : 
                            (N157)? \nz.mem [849] : 
                            (N159)? \nz.mem [889] : 
                            (N161)? \nz.mem [929] : 
                            (N163)? \nz.mem [969] : 
                            (N165)? \nz.mem [1009] : 
                            (N167)? \nz.mem [1049] : 
                            (N169)? \nz.mem [1089] : 
                            (N171)? \nz.mem [1129] : 
                            (N173)? \nz.mem [1169] : 
                            (N175)? \nz.mem [1209] : 
                            (N177)? \nz.mem [1249] : 
                            (N116)? \nz.mem [1289] : 
                            (N118)? \nz.mem [1329] : 
                            (N120)? \nz.mem [1369] : 
                            (N122)? \nz.mem [1409] : 
                            (N124)? \nz.mem [1449] : 
                            (N126)? \nz.mem [1489] : 
                            (N128)? \nz.mem [1529] : 
                            (N130)? \nz.mem [1569] : 
                            (N132)? \nz.mem [1609] : 
                            (N134)? \nz.mem [1649] : 
                            (N136)? \nz.mem [1689] : 
                            (N138)? \nz.mem [1729] : 
                            (N140)? \nz.mem [1769] : 
                            (N142)? \nz.mem [1809] : 
                            (N144)? \nz.mem [1849] : 
                            (N146)? \nz.mem [1889] : 
                            (N148)? \nz.mem [1929] : 
                            (N150)? \nz.mem [1969] : 
                            (N152)? \nz.mem [2009] : 
                            (N154)? \nz.mem [2049] : 
                            (N156)? \nz.mem [2089] : 
                            (N158)? \nz.mem [2129] : 
                            (N160)? \nz.mem [2169] : 
                            (N162)? \nz.mem [2209] : 
                            (N164)? \nz.mem [2249] : 
                            (N166)? \nz.mem [2289] : 
                            (N168)? \nz.mem [2329] : 
                            (N170)? \nz.mem [2369] : 
                            (N172)? \nz.mem [2409] : 
                            (N174)? \nz.mem [2449] : 
                            (N176)? \nz.mem [2489] : 
                            (N178)? \nz.mem [2529] : 1'b0;
  assign \nz.data_out [8] = (N115)? \nz.mem [8] : 
                            (N117)? \nz.mem [48] : 
                            (N119)? \nz.mem [88] : 
                            (N121)? \nz.mem [128] : 
                            (N123)? \nz.mem [168] : 
                            (N125)? \nz.mem [208] : 
                            (N127)? \nz.mem [248] : 
                            (N129)? \nz.mem [288] : 
                            (N131)? \nz.mem [328] : 
                            (N133)? \nz.mem [368] : 
                            (N135)? \nz.mem [408] : 
                            (N137)? \nz.mem [448] : 
                            (N139)? \nz.mem [488] : 
                            (N141)? \nz.mem [528] : 
                            (N143)? \nz.mem [568] : 
                            (N145)? \nz.mem [608] : 
                            (N147)? \nz.mem [648] : 
                            (N149)? \nz.mem [688] : 
                            (N151)? \nz.mem [728] : 
                            (N153)? \nz.mem [768] : 
                            (N155)? \nz.mem [808] : 
                            (N157)? \nz.mem [848] : 
                            (N159)? \nz.mem [888] : 
                            (N161)? \nz.mem [928] : 
                            (N163)? \nz.mem [968] : 
                            (N165)? \nz.mem [1008] : 
                            (N167)? \nz.mem [1048] : 
                            (N169)? \nz.mem [1088] : 
                            (N171)? \nz.mem [1128] : 
                            (N173)? \nz.mem [1168] : 
                            (N175)? \nz.mem [1208] : 
                            (N177)? \nz.mem [1248] : 
                            (N116)? \nz.mem [1288] : 
                            (N118)? \nz.mem [1328] : 
                            (N120)? \nz.mem [1368] : 
                            (N122)? \nz.mem [1408] : 
                            (N124)? \nz.mem [1448] : 
                            (N126)? \nz.mem [1488] : 
                            (N128)? \nz.mem [1528] : 
                            (N130)? \nz.mem [1568] : 
                            (N132)? \nz.mem [1608] : 
                            (N134)? \nz.mem [1648] : 
                            (N136)? \nz.mem [1688] : 
                            (N138)? \nz.mem [1728] : 
                            (N140)? \nz.mem [1768] : 
                            (N142)? \nz.mem [1808] : 
                            (N144)? \nz.mem [1848] : 
                            (N146)? \nz.mem [1888] : 
                            (N148)? \nz.mem [1928] : 
                            (N150)? \nz.mem [1968] : 
                            (N152)? \nz.mem [2008] : 
                            (N154)? \nz.mem [2048] : 
                            (N156)? \nz.mem [2088] : 
                            (N158)? \nz.mem [2128] : 
                            (N160)? \nz.mem [2168] : 
                            (N162)? \nz.mem [2208] : 
                            (N164)? \nz.mem [2248] : 
                            (N166)? \nz.mem [2288] : 
                            (N168)? \nz.mem [2328] : 
                            (N170)? \nz.mem [2368] : 
                            (N172)? \nz.mem [2408] : 
                            (N174)? \nz.mem [2448] : 
                            (N176)? \nz.mem [2488] : 
                            (N178)? \nz.mem [2528] : 1'b0;
  assign \nz.data_out [7] = (N115)? \nz.mem [7] : 
                            (N117)? \nz.mem [47] : 
                            (N119)? \nz.mem [87] : 
                            (N121)? \nz.mem [127] : 
                            (N123)? \nz.mem [167] : 
                            (N125)? \nz.mem [207] : 
                            (N127)? \nz.mem [247] : 
                            (N129)? \nz.mem [287] : 
                            (N131)? \nz.mem [327] : 
                            (N133)? \nz.mem [367] : 
                            (N135)? \nz.mem [407] : 
                            (N137)? \nz.mem [447] : 
                            (N139)? \nz.mem [487] : 
                            (N141)? \nz.mem [527] : 
                            (N143)? \nz.mem [567] : 
                            (N145)? \nz.mem [607] : 
                            (N147)? \nz.mem [647] : 
                            (N149)? \nz.mem [687] : 
                            (N151)? \nz.mem [727] : 
                            (N153)? \nz.mem [767] : 
                            (N155)? \nz.mem [807] : 
                            (N157)? \nz.mem [847] : 
                            (N159)? \nz.mem [887] : 
                            (N161)? \nz.mem [927] : 
                            (N163)? \nz.mem [967] : 
                            (N165)? \nz.mem [1007] : 
                            (N167)? \nz.mem [1047] : 
                            (N169)? \nz.mem [1087] : 
                            (N171)? \nz.mem [1127] : 
                            (N173)? \nz.mem [1167] : 
                            (N175)? \nz.mem [1207] : 
                            (N177)? \nz.mem [1247] : 
                            (N116)? \nz.mem [1287] : 
                            (N118)? \nz.mem [1327] : 
                            (N120)? \nz.mem [1367] : 
                            (N122)? \nz.mem [1407] : 
                            (N124)? \nz.mem [1447] : 
                            (N126)? \nz.mem [1487] : 
                            (N128)? \nz.mem [1527] : 
                            (N130)? \nz.mem [1567] : 
                            (N132)? \nz.mem [1607] : 
                            (N134)? \nz.mem [1647] : 
                            (N136)? \nz.mem [1687] : 
                            (N138)? \nz.mem [1727] : 
                            (N140)? \nz.mem [1767] : 
                            (N142)? \nz.mem [1807] : 
                            (N144)? \nz.mem [1847] : 
                            (N146)? \nz.mem [1887] : 
                            (N148)? \nz.mem [1927] : 
                            (N150)? \nz.mem [1967] : 
                            (N152)? \nz.mem [2007] : 
                            (N154)? \nz.mem [2047] : 
                            (N156)? \nz.mem [2087] : 
                            (N158)? \nz.mem [2127] : 
                            (N160)? \nz.mem [2167] : 
                            (N162)? \nz.mem [2207] : 
                            (N164)? \nz.mem [2247] : 
                            (N166)? \nz.mem [2287] : 
                            (N168)? \nz.mem [2327] : 
                            (N170)? \nz.mem [2367] : 
                            (N172)? \nz.mem [2407] : 
                            (N174)? \nz.mem [2447] : 
                            (N176)? \nz.mem [2487] : 
                            (N178)? \nz.mem [2527] : 1'b0;
  assign \nz.data_out [6] = (N115)? \nz.mem [6] : 
                            (N117)? \nz.mem [46] : 
                            (N119)? \nz.mem [86] : 
                            (N121)? \nz.mem [126] : 
                            (N123)? \nz.mem [166] : 
                            (N125)? \nz.mem [206] : 
                            (N127)? \nz.mem [246] : 
                            (N129)? \nz.mem [286] : 
                            (N131)? \nz.mem [326] : 
                            (N133)? \nz.mem [366] : 
                            (N135)? \nz.mem [406] : 
                            (N137)? \nz.mem [446] : 
                            (N139)? \nz.mem [486] : 
                            (N141)? \nz.mem [526] : 
                            (N143)? \nz.mem [566] : 
                            (N145)? \nz.mem [606] : 
                            (N147)? \nz.mem [646] : 
                            (N149)? \nz.mem [686] : 
                            (N151)? \nz.mem [726] : 
                            (N153)? \nz.mem [766] : 
                            (N155)? \nz.mem [806] : 
                            (N157)? \nz.mem [846] : 
                            (N159)? \nz.mem [886] : 
                            (N161)? \nz.mem [926] : 
                            (N163)? \nz.mem [966] : 
                            (N165)? \nz.mem [1006] : 
                            (N167)? \nz.mem [1046] : 
                            (N169)? \nz.mem [1086] : 
                            (N171)? \nz.mem [1126] : 
                            (N173)? \nz.mem [1166] : 
                            (N175)? \nz.mem [1206] : 
                            (N177)? \nz.mem [1246] : 
                            (N116)? \nz.mem [1286] : 
                            (N118)? \nz.mem [1326] : 
                            (N120)? \nz.mem [1366] : 
                            (N122)? \nz.mem [1406] : 
                            (N124)? \nz.mem [1446] : 
                            (N126)? \nz.mem [1486] : 
                            (N128)? \nz.mem [1526] : 
                            (N130)? \nz.mem [1566] : 
                            (N132)? \nz.mem [1606] : 
                            (N134)? \nz.mem [1646] : 
                            (N136)? \nz.mem [1686] : 
                            (N138)? \nz.mem [1726] : 
                            (N140)? \nz.mem [1766] : 
                            (N142)? \nz.mem [1806] : 
                            (N144)? \nz.mem [1846] : 
                            (N146)? \nz.mem [1886] : 
                            (N148)? \nz.mem [1926] : 
                            (N150)? \nz.mem [1966] : 
                            (N152)? \nz.mem [2006] : 
                            (N154)? \nz.mem [2046] : 
                            (N156)? \nz.mem [2086] : 
                            (N158)? \nz.mem [2126] : 
                            (N160)? \nz.mem [2166] : 
                            (N162)? \nz.mem [2206] : 
                            (N164)? \nz.mem [2246] : 
                            (N166)? \nz.mem [2286] : 
                            (N168)? \nz.mem [2326] : 
                            (N170)? \nz.mem [2366] : 
                            (N172)? \nz.mem [2406] : 
                            (N174)? \nz.mem [2446] : 
                            (N176)? \nz.mem [2486] : 
                            (N178)? \nz.mem [2526] : 1'b0;
  assign \nz.data_out [5] = (N115)? \nz.mem [5] : 
                            (N117)? \nz.mem [45] : 
                            (N119)? \nz.mem [85] : 
                            (N121)? \nz.mem [125] : 
                            (N123)? \nz.mem [165] : 
                            (N125)? \nz.mem [205] : 
                            (N127)? \nz.mem [245] : 
                            (N129)? \nz.mem [285] : 
                            (N131)? \nz.mem [325] : 
                            (N133)? \nz.mem [365] : 
                            (N135)? \nz.mem [405] : 
                            (N137)? \nz.mem [445] : 
                            (N139)? \nz.mem [485] : 
                            (N141)? \nz.mem [525] : 
                            (N143)? \nz.mem [565] : 
                            (N145)? \nz.mem [605] : 
                            (N147)? \nz.mem [645] : 
                            (N149)? \nz.mem [685] : 
                            (N151)? \nz.mem [725] : 
                            (N153)? \nz.mem [765] : 
                            (N155)? \nz.mem [805] : 
                            (N157)? \nz.mem [845] : 
                            (N159)? \nz.mem [885] : 
                            (N161)? \nz.mem [925] : 
                            (N163)? \nz.mem [965] : 
                            (N165)? \nz.mem [1005] : 
                            (N167)? \nz.mem [1045] : 
                            (N169)? \nz.mem [1085] : 
                            (N171)? \nz.mem [1125] : 
                            (N173)? \nz.mem [1165] : 
                            (N175)? \nz.mem [1205] : 
                            (N177)? \nz.mem [1245] : 
                            (N116)? \nz.mem [1285] : 
                            (N118)? \nz.mem [1325] : 
                            (N120)? \nz.mem [1365] : 
                            (N122)? \nz.mem [1405] : 
                            (N124)? \nz.mem [1445] : 
                            (N126)? \nz.mem [1485] : 
                            (N128)? \nz.mem [1525] : 
                            (N130)? \nz.mem [1565] : 
                            (N132)? \nz.mem [1605] : 
                            (N134)? \nz.mem [1645] : 
                            (N136)? \nz.mem [1685] : 
                            (N138)? \nz.mem [1725] : 
                            (N140)? \nz.mem [1765] : 
                            (N142)? \nz.mem [1805] : 
                            (N144)? \nz.mem [1845] : 
                            (N146)? \nz.mem [1885] : 
                            (N148)? \nz.mem [1925] : 
                            (N150)? \nz.mem [1965] : 
                            (N152)? \nz.mem [2005] : 
                            (N154)? \nz.mem [2045] : 
                            (N156)? \nz.mem [2085] : 
                            (N158)? \nz.mem [2125] : 
                            (N160)? \nz.mem [2165] : 
                            (N162)? \nz.mem [2205] : 
                            (N164)? \nz.mem [2245] : 
                            (N166)? \nz.mem [2285] : 
                            (N168)? \nz.mem [2325] : 
                            (N170)? \nz.mem [2365] : 
                            (N172)? \nz.mem [2405] : 
                            (N174)? \nz.mem [2445] : 
                            (N176)? \nz.mem [2485] : 
                            (N178)? \nz.mem [2525] : 1'b0;
  assign \nz.data_out [4] = (N115)? \nz.mem [4] : 
                            (N117)? \nz.mem [44] : 
                            (N119)? \nz.mem [84] : 
                            (N121)? \nz.mem [124] : 
                            (N123)? \nz.mem [164] : 
                            (N125)? \nz.mem [204] : 
                            (N127)? \nz.mem [244] : 
                            (N129)? \nz.mem [284] : 
                            (N131)? \nz.mem [324] : 
                            (N133)? \nz.mem [364] : 
                            (N135)? \nz.mem [404] : 
                            (N137)? \nz.mem [444] : 
                            (N139)? \nz.mem [484] : 
                            (N141)? \nz.mem [524] : 
                            (N143)? \nz.mem [564] : 
                            (N145)? \nz.mem [604] : 
                            (N147)? \nz.mem [644] : 
                            (N149)? \nz.mem [684] : 
                            (N151)? \nz.mem [724] : 
                            (N153)? \nz.mem [764] : 
                            (N155)? \nz.mem [804] : 
                            (N157)? \nz.mem [844] : 
                            (N159)? \nz.mem [884] : 
                            (N161)? \nz.mem [924] : 
                            (N163)? \nz.mem [964] : 
                            (N165)? \nz.mem [1004] : 
                            (N167)? \nz.mem [1044] : 
                            (N169)? \nz.mem [1084] : 
                            (N171)? \nz.mem [1124] : 
                            (N173)? \nz.mem [1164] : 
                            (N175)? \nz.mem [1204] : 
                            (N177)? \nz.mem [1244] : 
                            (N116)? \nz.mem [1284] : 
                            (N118)? \nz.mem [1324] : 
                            (N120)? \nz.mem [1364] : 
                            (N122)? \nz.mem [1404] : 
                            (N124)? \nz.mem [1444] : 
                            (N126)? \nz.mem [1484] : 
                            (N128)? \nz.mem [1524] : 
                            (N130)? \nz.mem [1564] : 
                            (N132)? \nz.mem [1604] : 
                            (N134)? \nz.mem [1644] : 
                            (N136)? \nz.mem [1684] : 
                            (N138)? \nz.mem [1724] : 
                            (N140)? \nz.mem [1764] : 
                            (N142)? \nz.mem [1804] : 
                            (N144)? \nz.mem [1844] : 
                            (N146)? \nz.mem [1884] : 
                            (N148)? \nz.mem [1924] : 
                            (N150)? \nz.mem [1964] : 
                            (N152)? \nz.mem [2004] : 
                            (N154)? \nz.mem [2044] : 
                            (N156)? \nz.mem [2084] : 
                            (N158)? \nz.mem [2124] : 
                            (N160)? \nz.mem [2164] : 
                            (N162)? \nz.mem [2204] : 
                            (N164)? \nz.mem [2244] : 
                            (N166)? \nz.mem [2284] : 
                            (N168)? \nz.mem [2324] : 
                            (N170)? \nz.mem [2364] : 
                            (N172)? \nz.mem [2404] : 
                            (N174)? \nz.mem [2444] : 
                            (N176)? \nz.mem [2484] : 
                            (N178)? \nz.mem [2524] : 1'b0;
  assign \nz.data_out [3] = (N115)? \nz.mem [3] : 
                            (N117)? \nz.mem [43] : 
                            (N119)? \nz.mem [83] : 
                            (N121)? \nz.mem [123] : 
                            (N123)? \nz.mem [163] : 
                            (N125)? \nz.mem [203] : 
                            (N127)? \nz.mem [243] : 
                            (N129)? \nz.mem [283] : 
                            (N131)? \nz.mem [323] : 
                            (N133)? \nz.mem [363] : 
                            (N135)? \nz.mem [403] : 
                            (N137)? \nz.mem [443] : 
                            (N139)? \nz.mem [483] : 
                            (N141)? \nz.mem [523] : 
                            (N143)? \nz.mem [563] : 
                            (N145)? \nz.mem [603] : 
                            (N147)? \nz.mem [643] : 
                            (N149)? \nz.mem [683] : 
                            (N151)? \nz.mem [723] : 
                            (N153)? \nz.mem [763] : 
                            (N155)? \nz.mem [803] : 
                            (N157)? \nz.mem [843] : 
                            (N159)? \nz.mem [883] : 
                            (N161)? \nz.mem [923] : 
                            (N163)? \nz.mem [963] : 
                            (N165)? \nz.mem [1003] : 
                            (N167)? \nz.mem [1043] : 
                            (N169)? \nz.mem [1083] : 
                            (N171)? \nz.mem [1123] : 
                            (N173)? \nz.mem [1163] : 
                            (N175)? \nz.mem [1203] : 
                            (N177)? \nz.mem [1243] : 
                            (N116)? \nz.mem [1283] : 
                            (N118)? \nz.mem [1323] : 
                            (N120)? \nz.mem [1363] : 
                            (N122)? \nz.mem [1403] : 
                            (N124)? \nz.mem [1443] : 
                            (N126)? \nz.mem [1483] : 
                            (N128)? \nz.mem [1523] : 
                            (N130)? \nz.mem [1563] : 
                            (N132)? \nz.mem [1603] : 
                            (N134)? \nz.mem [1643] : 
                            (N136)? \nz.mem [1683] : 
                            (N138)? \nz.mem [1723] : 
                            (N140)? \nz.mem [1763] : 
                            (N142)? \nz.mem [1803] : 
                            (N144)? \nz.mem [1843] : 
                            (N146)? \nz.mem [1883] : 
                            (N148)? \nz.mem [1923] : 
                            (N150)? \nz.mem [1963] : 
                            (N152)? \nz.mem [2003] : 
                            (N154)? \nz.mem [2043] : 
                            (N156)? \nz.mem [2083] : 
                            (N158)? \nz.mem [2123] : 
                            (N160)? \nz.mem [2163] : 
                            (N162)? \nz.mem [2203] : 
                            (N164)? \nz.mem [2243] : 
                            (N166)? \nz.mem [2283] : 
                            (N168)? \nz.mem [2323] : 
                            (N170)? \nz.mem [2363] : 
                            (N172)? \nz.mem [2403] : 
                            (N174)? \nz.mem [2443] : 
                            (N176)? \nz.mem [2483] : 
                            (N178)? \nz.mem [2523] : 1'b0;
  assign \nz.data_out [2] = (N115)? \nz.mem [2] : 
                            (N117)? \nz.mem [42] : 
                            (N119)? \nz.mem [82] : 
                            (N121)? \nz.mem [122] : 
                            (N123)? \nz.mem [162] : 
                            (N125)? \nz.mem [202] : 
                            (N127)? \nz.mem [242] : 
                            (N129)? \nz.mem [282] : 
                            (N131)? \nz.mem [322] : 
                            (N133)? \nz.mem [362] : 
                            (N135)? \nz.mem [402] : 
                            (N137)? \nz.mem [442] : 
                            (N139)? \nz.mem [482] : 
                            (N141)? \nz.mem [522] : 
                            (N143)? \nz.mem [562] : 
                            (N145)? \nz.mem [602] : 
                            (N147)? \nz.mem [642] : 
                            (N149)? \nz.mem [682] : 
                            (N151)? \nz.mem [722] : 
                            (N153)? \nz.mem [762] : 
                            (N155)? \nz.mem [802] : 
                            (N157)? \nz.mem [842] : 
                            (N159)? \nz.mem [882] : 
                            (N161)? \nz.mem [922] : 
                            (N163)? \nz.mem [962] : 
                            (N165)? \nz.mem [1002] : 
                            (N167)? \nz.mem [1042] : 
                            (N169)? \nz.mem [1082] : 
                            (N171)? \nz.mem [1122] : 
                            (N173)? \nz.mem [1162] : 
                            (N175)? \nz.mem [1202] : 
                            (N177)? \nz.mem [1242] : 
                            (N116)? \nz.mem [1282] : 
                            (N118)? \nz.mem [1322] : 
                            (N120)? \nz.mem [1362] : 
                            (N122)? \nz.mem [1402] : 
                            (N124)? \nz.mem [1442] : 
                            (N126)? \nz.mem [1482] : 
                            (N128)? \nz.mem [1522] : 
                            (N130)? \nz.mem [1562] : 
                            (N132)? \nz.mem [1602] : 
                            (N134)? \nz.mem [1642] : 
                            (N136)? \nz.mem [1682] : 
                            (N138)? \nz.mem [1722] : 
                            (N140)? \nz.mem [1762] : 
                            (N142)? \nz.mem [1802] : 
                            (N144)? \nz.mem [1842] : 
                            (N146)? \nz.mem [1882] : 
                            (N148)? \nz.mem [1922] : 
                            (N150)? \nz.mem [1962] : 
                            (N152)? \nz.mem [2002] : 
                            (N154)? \nz.mem [2042] : 
                            (N156)? \nz.mem [2082] : 
                            (N158)? \nz.mem [2122] : 
                            (N160)? \nz.mem [2162] : 
                            (N162)? \nz.mem [2202] : 
                            (N164)? \nz.mem [2242] : 
                            (N166)? \nz.mem [2282] : 
                            (N168)? \nz.mem [2322] : 
                            (N170)? \nz.mem [2362] : 
                            (N172)? \nz.mem [2402] : 
                            (N174)? \nz.mem [2442] : 
                            (N176)? \nz.mem [2482] : 
                            (N178)? \nz.mem [2522] : 1'b0;
  assign \nz.data_out [1] = (N115)? \nz.mem [1] : 
                            (N117)? \nz.mem [41] : 
                            (N119)? \nz.mem [81] : 
                            (N121)? \nz.mem [121] : 
                            (N123)? \nz.mem [161] : 
                            (N125)? \nz.mem [201] : 
                            (N127)? \nz.mem [241] : 
                            (N129)? \nz.mem [281] : 
                            (N131)? \nz.mem [321] : 
                            (N133)? \nz.mem [361] : 
                            (N135)? \nz.mem [401] : 
                            (N137)? \nz.mem [441] : 
                            (N139)? \nz.mem [481] : 
                            (N141)? \nz.mem [521] : 
                            (N143)? \nz.mem [561] : 
                            (N145)? \nz.mem [601] : 
                            (N147)? \nz.mem [641] : 
                            (N149)? \nz.mem [681] : 
                            (N151)? \nz.mem [721] : 
                            (N153)? \nz.mem [761] : 
                            (N155)? \nz.mem [801] : 
                            (N157)? \nz.mem [841] : 
                            (N159)? \nz.mem [881] : 
                            (N161)? \nz.mem [921] : 
                            (N163)? \nz.mem [961] : 
                            (N165)? \nz.mem [1001] : 
                            (N167)? \nz.mem [1041] : 
                            (N169)? \nz.mem [1081] : 
                            (N171)? \nz.mem [1121] : 
                            (N173)? \nz.mem [1161] : 
                            (N175)? \nz.mem [1201] : 
                            (N177)? \nz.mem [1241] : 
                            (N116)? \nz.mem [1281] : 
                            (N118)? \nz.mem [1321] : 
                            (N120)? \nz.mem [1361] : 
                            (N122)? \nz.mem [1401] : 
                            (N124)? \nz.mem [1441] : 
                            (N126)? \nz.mem [1481] : 
                            (N128)? \nz.mem [1521] : 
                            (N130)? \nz.mem [1561] : 
                            (N132)? \nz.mem [1601] : 
                            (N134)? \nz.mem [1641] : 
                            (N136)? \nz.mem [1681] : 
                            (N138)? \nz.mem [1721] : 
                            (N140)? \nz.mem [1761] : 
                            (N142)? \nz.mem [1801] : 
                            (N144)? \nz.mem [1841] : 
                            (N146)? \nz.mem [1881] : 
                            (N148)? \nz.mem [1921] : 
                            (N150)? \nz.mem [1961] : 
                            (N152)? \nz.mem [2001] : 
                            (N154)? \nz.mem [2041] : 
                            (N156)? \nz.mem [2081] : 
                            (N158)? \nz.mem [2121] : 
                            (N160)? \nz.mem [2161] : 
                            (N162)? \nz.mem [2201] : 
                            (N164)? \nz.mem [2241] : 
                            (N166)? \nz.mem [2281] : 
                            (N168)? \nz.mem [2321] : 
                            (N170)? \nz.mem [2361] : 
                            (N172)? \nz.mem [2401] : 
                            (N174)? \nz.mem [2441] : 
                            (N176)? \nz.mem [2481] : 
                            (N178)? \nz.mem [2521] : 1'b0;
  assign \nz.data_out [0] = (N115)? \nz.mem [0] : 
                            (N117)? \nz.mem [40] : 
                            (N119)? \nz.mem [80] : 
                            (N121)? \nz.mem [120] : 
                            (N123)? \nz.mem [160] : 
                            (N125)? \nz.mem [200] : 
                            (N127)? \nz.mem [240] : 
                            (N129)? \nz.mem [280] : 
                            (N131)? \nz.mem [320] : 
                            (N133)? \nz.mem [360] : 
                            (N135)? \nz.mem [400] : 
                            (N137)? \nz.mem [440] : 
                            (N139)? \nz.mem [480] : 
                            (N141)? \nz.mem [520] : 
                            (N143)? \nz.mem [560] : 
                            (N145)? \nz.mem [600] : 
                            (N147)? \nz.mem [640] : 
                            (N149)? \nz.mem [680] : 
                            (N151)? \nz.mem [720] : 
                            (N153)? \nz.mem [760] : 
                            (N155)? \nz.mem [800] : 
                            (N157)? \nz.mem [840] : 
                            (N159)? \nz.mem [880] : 
                            (N161)? \nz.mem [920] : 
                            (N163)? \nz.mem [960] : 
                            (N165)? \nz.mem [1000] : 
                            (N167)? \nz.mem [1040] : 
                            (N169)? \nz.mem [1080] : 
                            (N171)? \nz.mem [1120] : 
                            (N173)? \nz.mem [1160] : 
                            (N175)? \nz.mem [1200] : 
                            (N177)? \nz.mem [1240] : 
                            (N116)? \nz.mem [1280] : 
                            (N118)? \nz.mem [1320] : 
                            (N120)? \nz.mem [1360] : 
                            (N122)? \nz.mem [1400] : 
                            (N124)? \nz.mem [1440] : 
                            (N126)? \nz.mem [1480] : 
                            (N128)? \nz.mem [1520] : 
                            (N130)? \nz.mem [1560] : 
                            (N132)? \nz.mem [1600] : 
                            (N134)? \nz.mem [1640] : 
                            (N136)? \nz.mem [1680] : 
                            (N138)? \nz.mem [1720] : 
                            (N140)? \nz.mem [1760] : 
                            (N142)? \nz.mem [1800] : 
                            (N144)? \nz.mem [1840] : 
                            (N146)? \nz.mem [1880] : 
                            (N148)? \nz.mem [1920] : 
                            (N150)? \nz.mem [1960] : 
                            (N152)? \nz.mem [2000] : 
                            (N154)? \nz.mem [2040] : 
                            (N156)? \nz.mem [2080] : 
                            (N158)? \nz.mem [2120] : 
                            (N160)? \nz.mem [2160] : 
                            (N162)? \nz.mem [2200] : 
                            (N164)? \nz.mem [2240] : 
                            (N166)? \nz.mem [2280] : 
                            (N168)? \nz.mem [2320] : 
                            (N170)? \nz.mem [2360] : 
                            (N172)? \nz.mem [2400] : 
                            (N174)? \nz.mem [2440] : 
                            (N176)? \nz.mem [2480] : 
                            (N178)? \nz.mem [2520] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p40
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N5811 = addr_i[5] & N5869;
  assign N5812 = addr_i[5] & N5870;
  assign N5813 = addr_i[5] & N5871;
  assign N5814 = addr_i[2] & N5881;
  assign N5815 = addr_i[2] & N5882;
  assign N5816 = addr_i[2] & N5883;
  assign N415 = N5811 & N5814;
  assign N414 = N5811 & N5815;
  assign N413 = N5811 & N5816;
  assign N412 = N5811 & N5888;
  assign N411 = N5811 & N5831;
  assign N410 = N5811 & N5832;
  assign N409 = N5811 & N5833;
  assign N408 = N5811 & N5834;
  assign N407 = N5812 & N5814;
  assign N406 = N5812 & N5815;
  assign N405 = N5812 & N5816;
  assign N404 = N5812 & N5888;
  assign N403 = N5812 & N5831;
  assign N402 = N5812 & N5832;
  assign N401 = N5812 & N5833;
  assign N400 = N5812 & N5834;
  assign N399 = N5813 & N5814;
  assign N398 = N5813 & N5815;
  assign N397 = N5813 & N5816;
  assign N396 = N5813 & N5888;
  assign N395 = N5813 & N5831;
  assign N394 = N5813 & N5832;
  assign N393 = N5813 & N5833;
  assign N392 = N5813 & N5834;
  assign N391 = N5876 & N5814;
  assign N390 = N5876 & N5815;
  assign N389 = N5876 & N5816;
  assign N388 = N5826 & N5814;
  assign N387 = N5826 & N5815;
  assign N386 = N5826 & N5816;
  assign N385 = N5827 & N5814;
  assign N384 = N5827 & N5815;
  assign N383 = N5827 & N5816;
  assign N382 = N5828 & N5814;
  assign N381 = N5828 & N5815;
  assign N380 = N5828 & N5816;
  assign N379 = N5829 & N5814;
  assign N378 = N5829 & N5815;
  assign N377 = N5829 & N5816;
  assign N884 = N5835 & N5888;
  assign N883 = N5836 & N5888;
  assign N882 = N5837 & N5888;
  assign N881 = N5876 & N5838;
  assign N880 = N5876 & N5839;
  assign N879 = N5876 & N5840;
  assign N878 = N5876 & N5831;
  assign N877 = N5876 & N5832;
  assign N876 = N5876 & N5833;
  assign N875 = N5876 & N5834;
  assign N874 = N5826 & N5888;
  assign N873 = N5827 & N5888;
  assign N872 = N5828 & N5888;
  assign N871 = N5829 & N5888;
  assign N5817 = N5825 & N5869;
  assign N5818 = N5825 & N5870;
  assign N5819 = N5825 & N5871;
  assign N5820 = N5825 & N5872;
  assign N5821 = N5830 & N5881;
  assign N5822 = N5830 & N5882;
  assign N5823 = N5830 & N5883;
  assign N5824 = N5830 & N5884;
  assign N1127 = N5835 & N5821;
  assign N1126 = N5835 & N5822;
  assign N1125 = N5835 & N5823;
  assign N1124 = N5835 & N5824;
  assign N1123 = N5836 & N5821;
  assign N1122 = N5836 & N5822;
  assign N1121 = N5836 & N5823;
  assign N1120 = N5836 & N5824;
  assign N1119 = N5837 & N5821;
  assign N1118 = N5837 & N5822;
  assign N1117 = N5837 & N5823;
  assign N1116 = N5837 & N5824;
  assign N1115 = N5859 & N5821;
  assign N1114 = N5859 & N5822;
  assign N1113 = N5859 & N5823;
  assign N1112 = N5859 & N5824;
  assign N1111 = N5817 & N5838;
  assign N1110 = N5817 & N5839;
  assign N1109 = N5817 & N5840;
  assign N1108 = N5817 & N5864;
  assign N1107 = N5817 & N5821;
  assign N1106 = N5817 & N5822;
  assign N1105 = N5817 & N5823;
  assign N1104 = N5817 & N5824;
  assign N1103 = N5818 & N5838;
  assign N1102 = N5818 & N5839;
  assign N1101 = N5818 & N5840;
  assign N1100 = N5818 & N5864;
  assign N1099 = N5818 & N5821;
  assign N1098 = N5818 & N5822;
  assign N1097 = N5818 & N5823;
  assign N1096 = N5818 & N5824;
  assign N1095 = N5819 & N5838;
  assign N1094 = N5819 & N5839;
  assign N1093 = N5819 & N5840;
  assign N1092 = N5819 & N5864;
  assign N1091 = N5819 & N5821;
  assign N1090 = N5819 & N5822;
  assign N1089 = N5819 & N5823;
  assign N1088 = N5819 & N5824;
  assign N1087 = N5820 & N5838;
  assign N1086 = N5820 & N5839;
  assign N1085 = N5820 & N5840;
  assign N1084 = N5820 & N5864;
  assign N1083 = N5820 & N5821;
  assign N1082 = N5820 & N5822;
  assign N1081 = N5820 & N5823;
  assign N1080 = N5820 & N5824;
  assign N5825 = ~addr_i[5];
  assign N5826 = N5825 & N5869;
  assign N5827 = N5825 & N5870;
  assign N5828 = N5825 & N5871;
  assign N5829 = N5825 & N5872;
  assign N5830 = ~addr_i[2];
  assign N5831 = N5830 & N5881;
  assign N5832 = N5830 & N5882;
  assign N5833 = N5830 & N5883;
  assign N5834 = N5830 & N5884;
  assign N1240 = N5835 & N5831;
  assign N1239 = N5835 & N5832;
  assign N1238 = N5835 & N5833;
  assign N1237 = N5835 & N5834;
  assign N1236 = N5836 & N5831;
  assign N1235 = N5836 & N5832;
  assign N1234 = N5836 & N5833;
  assign N1233 = N5836 & N5834;
  assign N1232 = N5837 & N5831;
  assign N1231 = N5837 & N5832;
  assign N1230 = N5837 & N5833;
  assign N1229 = N5837 & N5834;
  assign N1228 = N5859 & N5831;
  assign N1227 = N5859 & N5832;
  assign N1226 = N5859 & N5833;
  assign N1225 = N5859 & N5834;
  assign N1224 = N5826 & N5838;
  assign N1223 = N5826 & N5839;
  assign N1222 = N5826 & N5840;
  assign N1221 = N5826 & N5864;
  assign N1220 = N5826 & N5831;
  assign N1219 = N5826 & N5832;
  assign N1218 = N5826 & N5833;
  assign N1217 = N5826 & N5834;
  assign N1216 = N5827 & N5838;
  assign N1215 = N5827 & N5839;
  assign N1214 = N5827 & N5840;
  assign N1213 = N5827 & N5864;
  assign N1212 = N5827 & N5831;
  assign N1211 = N5827 & N5832;
  assign N1210 = N5827 & N5833;
  assign N1209 = N5827 & N5834;
  assign N1208 = N5828 & N5838;
  assign N1207 = N5828 & N5839;
  assign N1206 = N5828 & N5840;
  assign N1205 = N5828 & N5864;
  assign N1204 = N5828 & N5831;
  assign N1203 = N5828 & N5832;
  assign N1202 = N5828 & N5833;
  assign N1201 = N5828 & N5834;
  assign N1200 = N5829 & N5838;
  assign N1199 = N5829 & N5839;
  assign N1198 = N5829 & N5840;
  assign N1197 = N5829 & N5864;
  assign N1196 = N5829 & N5831;
  assign N1195 = N5829 & N5832;
  assign N1194 = N5829 & N5833;
  assign N1193 = N5829 & N5834;
  assign N5835 = addr_i[5] & N5869;
  assign N5836 = addr_i[5] & N5870;
  assign N5837 = addr_i[5] & N5871;
  assign N5838 = addr_i[2] & N5881;
  assign N5839 = addr_i[2] & N5882;
  assign N5840 = addr_i[2] & N5883;
  assign N1344 = N5835 & N5838;
  assign N1343 = N5835 & N5839;
  assign N1342 = N5835 & N5840;
  assign N1341 = N5835 & N5864;
  assign N1340 = N5835 & N5889;
  assign N1339 = N5835 & N5890;
  assign N1338 = N5835 & N5891;
  assign N1337 = N5835 & N5892;
  assign N1336 = N5836 & N5838;
  assign N1335 = N5836 & N5839;
  assign N1334 = N5836 & N5840;
  assign N1333 = N5836 & N5864;
  assign N1332 = N5836 & N5889;
  assign N1331 = N5836 & N5890;
  assign N1330 = N5836 & N5891;
  assign N1329 = N5836 & N5892;
  assign N1328 = N5837 & N5838;
  assign N1327 = N5837 & N5839;
  assign N1326 = N5837 & N5840;
  assign N1325 = N5837 & N5864;
  assign N1324 = N5837 & N5889;
  assign N1323 = N5837 & N5890;
  assign N1322 = N5837 & N5891;
  assign N1321 = N5837 & N5892;
  assign N1320 = N5859 & N5838;
  assign N1319 = N5859 & N5839;
  assign N1318 = N5859 & N5840;
  assign N1317 = N5877 & N5838;
  assign N1316 = N5877 & N5839;
  assign N1315 = N5877 & N5840;
  assign N1314 = N5878 & N5838;
  assign N1313 = N5878 & N5839;
  assign N1312 = N5878 & N5840;
  assign N1311 = N5879 & N5838;
  assign N1310 = N5879 & N5839;
  assign N1309 = N5879 & N5840;
  assign N1308 = N5880 & N5838;
  assign N1307 = N5880 & N5839;
  assign N1306 = N5880 & N5840;
  assign N1748 = N5841 & N5864;
  assign N1747 = N5842 & N5864;
  assign N1746 = N5843 & N5864;
  assign N1745 = N5859 & N5844;
  assign N1744 = N5859 & N5845;
  assign N1743 = N5859 & N5846;
  assign N1742 = N5859 & N5889;
  assign N1741 = N5859 & N5890;
  assign N1740 = N5859 & N5891;
  assign N1739 = N5859 & N5892;
  assign N1738 = N5877 & N5864;
  assign N1737 = N5878 & N5864;
  assign N1736 = N5879 & N5864;
  assign N1735 = N5880 & N5864;
  assign N2040 = N5841 & N5889;
  assign N2039 = N5841 & N5890;
  assign N2038 = N5841 & N5891;
  assign N2037 = N5841 & N5892;
  assign N2036 = N5842 & N5889;
  assign N2035 = N5842 & N5890;
  assign N2034 = N5842 & N5891;
  assign N2033 = N5842 & N5892;
  assign N2032 = N5843 & N5889;
  assign N2031 = N5843 & N5890;
  assign N2030 = N5843 & N5891;
  assign N2029 = N5843 & N5892;
  assign N2028 = N5849 & N5889;
  assign N2027 = N5849 & N5890;
  assign N2026 = N5849 & N5891;
  assign N2025 = N5849 & N5892;
  assign N2024 = N5877 & N5844;
  assign N2023 = N5877 & N5845;
  assign N2022 = N5877 & N5846;
  assign N2021 = N5877 & N5854;
  assign N2020 = N5878 & N5844;
  assign N2019 = N5878 & N5845;
  assign N2018 = N5878 & N5846;
  assign N2017 = N5878 & N5854;
  assign N2016 = N5879 & N5844;
  assign N2015 = N5879 & N5845;
  assign N2014 = N5879 & N5846;
  assign N2013 = N5879 & N5854;
  assign N2012 = N5880 & N5844;
  assign N2011 = N5880 & N5845;
  assign N2010 = N5880 & N5846;
  assign N2009 = N5880 & N5854;
  assign N5841 = addr_i[5] & N5869;
  assign N5842 = addr_i[5] & N5870;
  assign N5843 = addr_i[5] & N5871;
  assign N5844 = addr_i[2] & N5881;
  assign N5845 = addr_i[2] & N5882;
  assign N5846 = addr_i[2] & N5883;
  assign N2209 = N5841 & N5844;
  assign N2208 = N5841 & N5845;
  assign N2207 = N5841 & N5846;
  assign N2206 = N5841 & N5854;
  assign N2205 = N5841 & N5865;
  assign N2204 = N5841 & N5866;
  assign N2203 = N5841 & N5867;
  assign N2202 = N5841 & N5868;
  assign N2201 = N5842 & N5844;
  assign N2200 = N5842 & N5845;
  assign N2199 = N5842 & N5846;
  assign N2198 = N5842 & N5854;
  assign N2197 = N5842 & N5865;
  assign N2196 = N5842 & N5866;
  assign N2195 = N5842 & N5867;
  assign N2194 = N5842 & N5868;
  assign N2193 = N5843 & N5844;
  assign N2192 = N5843 & N5845;
  assign N2191 = N5843 & N5846;
  assign N2190 = N5843 & N5854;
  assign N2189 = N5843 & N5865;
  assign N2188 = N5843 & N5866;
  assign N2187 = N5843 & N5867;
  assign N2186 = N5843 & N5868;
  assign N2185 = N5849 & N5844;
  assign N2184 = N5849 & N5845;
  assign N2183 = N5849 & N5846;
  assign N2182 = N5860 & N5844;
  assign N2181 = N5860 & N5845;
  assign N2180 = N5860 & N5846;
  assign N2179 = N5861 & N5844;
  assign N2178 = N5861 & N5845;
  assign N2177 = N5861 & N5846;
  assign N2176 = N5862 & N5844;
  assign N2175 = N5862 & N5845;
  assign N2174 = N5862 & N5846;
  assign N2173 = N5863 & N5844;
  assign N2172 = N5863 & N5845;
  assign N2171 = N5863 & N5846;
  assign N2542 = N5849 & N5865;
  assign N2541 = N5849 & N5866;
  assign N2540 = N5849 & N5867;
  assign N2539 = N5849 & N5868;
  assign N2538 = N5860 & N5854;
  assign N2537 = N5861 & N5854;
  assign N2536 = N5862 & N5854;
  assign N2535 = N5863 & N5854;
  assign N5847 = addr_i[5] & N5872;
  assign N5848 = addr_i[2] & N5884;
  assign N2817 = N5873 & N5848;
  assign N2816 = N5874 & N5848;
  assign N2815 = N5875 & N5848;
  assign N2814 = N5847 & N5885;
  assign N2813 = N5847 & N5886;
  assign N2812 = N5847 & N5887;
  assign N2811 = N5847 & N5848;
  assign N2810 = N5847 & N5865;
  assign N2809 = N5847 & N5866;
  assign N2808 = N5847 & N5867;
  assign N2807 = N5847 & N5868;
  assign N2806 = N5860 & N5848;
  assign N2805 = N5861 & N5848;
  assign N2804 = N5862 & N5848;
  assign N2803 = N5863 & N5848;
  assign N5849 = addr_i[5] & N5872;
  assign N5850 = N5825 & N5869;
  assign N5851 = N5825 & N5870;
  assign N5852 = N5825 & N5871;
  assign N5853 = N5825 & N5872;
  assign N5854 = addr_i[2] & N5884;
  assign N5855 = N5830 & N5881;
  assign N5856 = N5830 & N5882;
  assign N5857 = N5830 & N5883;
  assign N5858 = N5830 & N5884;
  assign N2937 = N5873 & N5854;
  assign N2936 = N5873 & N5855;
  assign N2935 = N5873 & N5856;
  assign N2934 = N5873 & N5857;
  assign N2933 = N5873 & N5858;
  assign N2932 = N5874 & N5854;
  assign N2931 = N5874 & N5855;
  assign N2930 = N5874 & N5856;
  assign N2929 = N5874 & N5857;
  assign N2928 = N5874 & N5858;
  assign N2927 = N5875 & N5854;
  assign N2926 = N5875 & N5855;
  assign N2925 = N5875 & N5856;
  assign N2924 = N5875 & N5857;
  assign N2923 = N5875 & N5858;
  assign N2922 = N5849 & N5885;
  assign N2921 = N5849 & N5886;
  assign N2920 = N5849 & N5887;
  assign N2919 = N5849 & N5854;
  assign N2918 = N5849 & N5855;
  assign N2917 = N5849 & N5856;
  assign N2916 = N5849 & N5857;
  assign N2915 = N5849 & N5858;
  assign N2914 = N5850 & N5885;
  assign N2913 = N5850 & N5886;
  assign N2912 = N5850 & N5887;
  assign N2911 = N5850 & N5854;
  assign N2910 = N5850 & N5855;
  assign N2909 = N5850 & N5856;
  assign N2908 = N5850 & N5857;
  assign N2907 = N5850 & N5858;
  assign N2906 = N5851 & N5885;
  assign N2905 = N5851 & N5886;
  assign N2904 = N5851 & N5887;
  assign N2903 = N5851 & N5854;
  assign N2902 = N5851 & N5855;
  assign N2901 = N5851 & N5856;
  assign N2900 = N5851 & N5857;
  assign N2899 = N5851 & N5858;
  assign N2898 = N5852 & N5885;
  assign N2897 = N5852 & N5886;
  assign N2896 = N5852 & N5887;
  assign N2895 = N5852 & N5854;
  assign N2894 = N5852 & N5855;
  assign N2893 = N5852 & N5856;
  assign N2892 = N5852 & N5857;
  assign N2891 = N5852 & N5858;
  assign N2890 = N5853 & N5885;
  assign N2889 = N5853 & N5886;
  assign N2888 = N5853 & N5887;
  assign N2887 = N5853 & N5854;
  assign N2886 = N5853 & N5855;
  assign N2885 = N5853 & N5856;
  assign N2884 = N5853 & N5857;
  assign N2883 = N5853 & N5858;
  assign N5859 = addr_i[5] & N5872;
  assign N5860 = N5825 & N5869;
  assign N5861 = N5825 & N5870;
  assign N5862 = N5825 & N5871;
  assign N5863 = N5825 & N5872;
  assign N5864 = addr_i[2] & N5884;
  assign N5865 = N5830 & N5881;
  assign N5866 = N5830 & N5882;
  assign N5867 = N5830 & N5883;
  assign N5868 = N5830 & N5884;
  assign N3057 = N5873 & N5864;
  assign N3056 = N5873 & N5865;
  assign N3055 = N5873 & N5866;
  assign N3054 = N5873 & N5867;
  assign N3053 = N5873 & N5868;
  assign N3052 = N5874 & N5864;
  assign N3051 = N5874 & N5865;
  assign N3050 = N5874 & N5866;
  assign N3049 = N5874 & N5867;
  assign N3048 = N5874 & N5868;
  assign N3047 = N5875 & N5864;
  assign N3046 = N5875 & N5865;
  assign N3045 = N5875 & N5866;
  assign N3044 = N5875 & N5867;
  assign N3043 = N5875 & N5868;
  assign N3042 = N5859 & N5885;
  assign N3041 = N5859 & N5886;
  assign N3040 = N5859 & N5887;
  assign N3039 = N5859 & N5864;
  assign N3038 = N5859 & N5865;
  assign N3037 = N5859 & N5866;
  assign N3036 = N5859 & N5867;
  assign N3035 = N5859 & N5868;
  assign N3034 = N5860 & N5885;
  assign N3033 = N5860 & N5886;
  assign N3032 = N5860 & N5887;
  assign N3031 = N5860 & N5864;
  assign N3030 = N5860 & N5865;
  assign N3029 = N5860 & N5866;
  assign N3028 = N5860 & N5867;
  assign N3027 = N5860 & N5868;
  assign N3026 = N5861 & N5885;
  assign N3025 = N5861 & N5886;
  assign N3024 = N5861 & N5887;
  assign N3023 = N5861 & N5864;
  assign N3022 = N5861 & N5865;
  assign N3021 = N5861 & N5866;
  assign N3020 = N5861 & N5867;
  assign N3019 = N5861 & N5868;
  assign N3018 = N5862 & N5885;
  assign N3017 = N5862 & N5886;
  assign N3016 = N5862 & N5887;
  assign N3015 = N5862 & N5864;
  assign N3014 = N5862 & N5865;
  assign N3013 = N5862 & N5866;
  assign N3012 = N5862 & N5867;
  assign N3011 = N5862 & N5868;
  assign N3010 = N5863 & N5885;
  assign N3009 = N5863 & N5886;
  assign N3008 = N5863 & N5887;
  assign N3007 = N5863 & N5864;
  assign N3006 = N5863 & N5865;
  assign N3005 = N5863 & N5866;
  assign N3004 = N5863 & N5867;
  assign N3003 = N5863 & N5868;
  assign N5869 = addr_i[3] & addr_i[4];
  assign N5870 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N5871 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N5872 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N5873 = addr_i[5] & N5869;
  assign N5874 = addr_i[5] & N5870;
  assign N5875 = addr_i[5] & N5871;
  assign N5876 = addr_i[5] & N5872;
  assign N5877 = N5825 & N5869;
  assign N5878 = N5825 & N5870;
  assign N5879 = N5825 & N5871;
  assign N5880 = N5825 & N5872;
  assign N5881 = addr_i[0] & addr_i[1];
  assign N5882 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N5883 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N5884 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N5885 = addr_i[2] & N5881;
  assign N5886 = addr_i[2] & N5882;
  assign N5887 = addr_i[2] & N5883;
  assign N5888 = addr_i[2] & N5884;
  assign N5889 = N5830 & N5881;
  assign N5890 = N5830 & N5882;
  assign N5891 = N5830 & N5883;
  assign N5892 = N5830 & N5884;
  assign N3186 = N5873 & N5885;
  assign N3185 = N5873 & N5886;
  assign N3184 = N5873 & N5887;
  assign N3183 = N5873 & N5888;
  assign N3182 = N5873 & N5889;
  assign N3181 = N5873 & N5890;
  assign N3180 = N5873 & N5891;
  assign N3179 = N5873 & N5892;
  assign N3178 = N5874 & N5885;
  assign N3177 = N5874 & N5886;
  assign N3176 = N5874 & N5887;
  assign N3175 = N5874 & N5888;
  assign N3174 = N5874 & N5889;
  assign N3173 = N5874 & N5890;
  assign N3172 = N5874 & N5891;
  assign N3171 = N5874 & N5892;
  assign N3170 = N5875 & N5885;
  assign N3169 = N5875 & N5886;
  assign N3168 = N5875 & N5887;
  assign N3167 = N5875 & N5888;
  assign N3166 = N5875 & N5889;
  assign N3165 = N5875 & N5890;
  assign N3164 = N5875 & N5891;
  assign N3163 = N5875 & N5892;
  assign N3162 = N5876 & N5885;
  assign N3161 = N5876 & N5886;
  assign N3160 = N5876 & N5887;
  assign N3159 = N5876 & N5888;
  assign N3158 = N5876 & N5889;
  assign N3157 = N5876 & N5890;
  assign N3156 = N5876 & N5891;
  assign N3155 = N5876 & N5892;
  assign N3154 = N5877 & N5885;
  assign N3153 = N5877 & N5886;
  assign N3152 = N5877 & N5887;
  assign N3151 = N5877 & N5888;
  assign N3150 = N5877 & N5889;
  assign N3149 = N5877 & N5890;
  assign N3148 = N5877 & N5891;
  assign N3147 = N5877 & N5892;
  assign N3146 = N5878 & N5885;
  assign N3145 = N5878 & N5886;
  assign N3144 = N5878 & N5887;
  assign N3143 = N5878 & N5888;
  assign N3142 = N5878 & N5889;
  assign N3141 = N5878 & N5890;
  assign N3140 = N5878 & N5891;
  assign N3139 = N5878 & N5892;
  assign N3138 = N5879 & N5885;
  assign N3137 = N5879 & N5886;
  assign N3136 = N5879 & N5887;
  assign N3135 = N5879 & N5888;
  assign N3134 = N5879 & N5889;
  assign N3133 = N5879 & N5890;
  assign N3132 = N5879 & N5891;
  assign N3131 = N5879 & N5892;
  assign N3130 = N5880 & N5885;
  assign N3129 = N5880 & N5886;
  assign N3128 = N5880 & N5887;
  assign N3127 = N5880 & N5888;
  assign N3126 = N5880 & N5889;
  assign N3125 = N5880 & N5890;
  assign N3124 = N5880 & N5891;
  assign N3123 = N5880 & N5892;
  assign { N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182 } = (N8)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N181)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247 } = (N9)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N246)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312 } = (N10)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N311)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416 } = (N11)? { N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N3159, N878, N877, N876, N875, N388, N387, N386, N874, N1220, N1219, N1218, N1217, N385, N384, N383, N873, N1212, N1211, N1210, N1209, N382, N381, N380, N872, N1204, N1203, N1202, N1201, N379, N378, N377, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N376)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481 } = (N12)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N480)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546 } = (N13)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N545)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611 } = (N14)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N610)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676 } = (N15)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N675)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = w_mask_i[7];
  assign { N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741 } = (N16)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N740)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_mask_i[8];
  assign { N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806 } = (N17)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N805)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N17 = w_mask_i[9];
  assign { N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885 } = (N18)? { N1344, N1343, N1342, N884, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N883, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N882, N1232, N1231, N1230, N1229, N881, N880, N879, N3159, N878, N877, N876, N875, N1224, N1223, N1222, N874, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N873, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N872, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N871, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N870)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N18 = w_mask_i[10];
  assign { N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950 } = (N19)? { N1344, N1343, N1342, N1341, N1127, N1126, N1125, N1124, N1336, N1335, N1334, N1333, N1123, N1122, N1121, N1120, N1328, N1327, N1326, N1325, N1119, N1118, N1117, N1116, N1320, N1319, N1318, N3039, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                            (N949)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = w_mask_i[11];
  assign { N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015 } = (N20)? { N1344, N1343, N1342, N1341, N1127, N1126, N1125, N1124, N1336, N1335, N1334, N1333, N1123, N1122, N1121, N1120, N1328, N1327, N1326, N1325, N1119, N1118, N1117, N1116, N1320, N1319, N1318, N3039, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1014)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = w_mask_i[12];
  assign { N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128 } = (N21)? { N1344, N1343, N1342, N1341, N1127, N1126, N1125, N1124, N1336, N1335, N1334, N1333, N1123, N1122, N1121, N1120, N1328, N1327, N1326, N1325, N1119, N1118, N1117, N1116, N1320, N1319, N1318, N3039, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1079)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N21 = w_mask_i[13];
  assign { N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241 } = (N22)? { N1344, N1343, N1342, N1341, N1240, N1239, N1238, N1237, N1336, N1335, N1334, N1333, N1236, N1235, N1234, N1233, N1328, N1327, N1326, N1325, N1232, N1231, N1230, N1229, N1320, N1319, N1318, N3039, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1192)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = w_mask_i[14];
  assign { N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345 } = (N23)? { N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N3039, N1742, N1741, N1740, N1739, N1317, N1316, N1315, N1738, N3150, N3149, N3148, N3147, N1314, N1313, N1312, N1737, N3142, N3141, N3140, N3139, N1311, N1310, N1309, N1736, N3134, N3133, N3132, N3131, N1308, N1307, N1306, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1305)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N23 = w_mask_i[15];
  assign { N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410 } = (N24)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1409)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N24 = w_mask_i[16];
  assign { N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475 } = (N25)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1474)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = w_mask_i[17];
  assign { N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540 } = (N26)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1539)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = w_mask_i[18];
  assign { N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605 } = (N27)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1604)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N27 = w_mask_i[19];
  assign { N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670 } = (N28)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1669)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N28 = w_mask_i[20];
  assign { N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749 } = (N29)? { N2209, N2208, N2207, N1748, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N1747, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N1746, N2032, N2031, N2030, N2029, N1745, N1744, N1743, N3039, N1742, N1741, N1740, N1739, N2024, N2023, N2022, N1738, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N1737, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N1736, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N1735, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1734)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N29 = w_mask_i[21];
  assign { N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814 } = (N30)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1813)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = w_mask_i[22];
  assign { N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879 } = (N31)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1878)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N31 = w_mask_i[23];
  assign { N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944 } = (N32)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1943)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = w_mask_i[24];
  assign { N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041 } = (N33)? { N2209, N2208, N2207, N2206, N2040, N2039, N2038, N2037, N2201, N2200, N2199, N2198, N2036, N2035, N2034, N2033, N2193, N2192, N2191, N2190, N2032, N2031, N2030, N2029, N2185, N2184, N2183, N2919, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N3150, N3149, N3148, N3147, N2020, N2019, N2018, N2017, N3142, N3141, N3140, N3139, N2016, N2015, N2014, N2013, N3134, N3133, N3132, N3131, N2012, N2011, N2010, N2009, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2008)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = w_mask_i[25];
  assign { N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106 } = (N34)? { N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2919, N2542, N2541, N2540, N2539, N2182, N2181, N2180, N2538, N3030, N3029, N3028, N3027, N2179, N2178, N2177, N2537, N3022, N3021, N3020, N3019, N2176, N2175, N2174, N2536, N3014, N3013, N3012, N3011, N2173, N2172, N2171, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2105)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N34 = w_mask_i[26];
  assign { N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210 } = (N35)? { N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2919, N2542, N2541, N2540, N2539, N2182, N2181, N2180, N2538, N3030, N3029, N3028, N3027, N2179, N2178, N2177, N2537, N3022, N3021, N3020, N3019, N2176, N2175, N2174, N2536, N3014, N3013, N3012, N3011, N2173, N2172, N2171, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2170)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N35 = w_mask_i[27];
  assign { N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275 } = (N36)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2274)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N36 = w_mask_i[28];
  assign { N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340 } = (N37)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2339)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N37 = w_mask_i[29];
  assign { N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405 } = (N38)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2404)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N38 = w_mask_i[30];
  assign { N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470 } = (N39)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2469)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N39 = w_mask_i[31];
  assign { N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543 } = (N40)? { N3186, N3185, N3184, N2937, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2932, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2927, N3046, N3045, N3044, N3043, N2922, N2921, N2920, N2919, N2542, N2541, N2540, N2539, N3034, N3033, N3032, N2538, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2537, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2536, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2535, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = w_mask_i[32];
  assign { N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608 } = (N41)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2607)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N41 = w_mask_i[33];
  assign { N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673 } = (N42)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2672)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = w_mask_i[34];
  assign { N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738 } = (N43)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2737)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N43 = w_mask_i[35];
  assign { N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818 } = (N44)? { N3186, N3185, N3184, N2817, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N2816, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N2815, N3046, N3045, N3044, N3043, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N3034, N3033, N3032, N2806, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N2805, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N2804, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N2803, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2802)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N44 = w_mask_i[36];
  assign { N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938 } = (N45)? { N3186, N3185, N3184, N2937, N2936, N2935, N2934, N2933, N3178, N3177, N3176, N2932, N2931, N2930, N2929, N2928, N3170, N3169, N3168, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2882)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N45 = w_mask_i[37];
  assign { N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058 } = (N46)? { N3186, N3185, N3184, N3057, N3056, N3055, N3054, N3053, N3178, N3177, N3176, N3052, N3051, N3050, N3049, N3048, N3170, N3169, N3168, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3002)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N46 = w_mask_i[38];
  assign { N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187 } = (N47)? { N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3122)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N47 = w_mask_i[39];
  assign { N5810, N5809, N5808, N5807, N5806, N5805, N5804, N5803, N5802, N5801, N5800, N5799, N5798, N5797, N5796, N5795, N5794, N5793, N5792, N5791, N5790, N5789, N5788, N5787, N5786, N5785, N5784, N5783, N5782, N5781, N5780, N5779, N5778, N5777, N5776, N5775, N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, N5755, N5754, N5753, N5752, N5751, N5750, N5749, N5748, N5747, N5746, N5745, N5744, N5743, N5742, N5741, N5740, N5739, N5738, N5737, N5736, N5735, N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721, N5720, N5719, N5718, N5717, N5716, N5715, N5714, N5713, N5712, N5711, N5710, N5709, N5708, N5707, N5706, N5705, N5704, N5703, N5702, N5701, N5700, N5699, N5698, N5697, N5696, N5695, N5694, N5693, N5692, N5691, N5690, N5689, N5688, N5687, N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, N5676, N5675, N5674, N5673, N5672, N5671, N5670, N5669, N5668, N5667, N5666, N5665, N5664, N5663, N5662, N5661, N5660, N5659, N5658, N5657, N5656, N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642, N5641, N5640, N5639, N5638, N5637, N5636, N5635, N5634, N5633, N5632, N5631, N5630, N5629, N5628, N5627, N5626, N5625, N5624, N5623, N5622, N5621, N5620, N5619, N5618, N5617, N5616, N5615, N5614, N5613, N5612, N5611, N5610, N5609, N5608, N5607, N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5587, N5586, N5585, N5584, N5583, N5582, N5581, N5580, N5579, N5578, N5577, N5576, N5575, N5574, N5573, N5572, N5571, N5570, N5569, N5568, N5567, N5566, N5565, N5564, N5563, N5562, N5561, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553, N5552, N5551, N5550, N5549, N5548, N5547, N5546, N5545, N5544, N5543, N5542, N5541, N5540, N5539, N5538, N5537, N5536, N5535, N5534, N5533, N5532, N5531, N5530, N5529, N5528, N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, N5507, N5506, N5505, N5504, N5503, N5502, N5501, N5500, N5499, N5498, N5497, N5496, N5495, N5494, N5493, N5492, N5491, N5490, N5489, N5488, N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474, N5473, N5472, N5471, N5470, N5469, N5468, N5467, N5466, N5465, N5464, N5463, N5462, N5461, N5460, N5459, N5458, N5457, N5456, N5455, N5454, N5453, N5452, N5451, N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442, N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, N5418, N5417, N5416, N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385, N5384, N5383, N5382, N5381, N5380, N5379, N5378, N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368, N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321, N5320, N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306, N5305, N5304, N5303, N5302, N5301, N5300, N5299, N5298, N5297, N5296, N5295, N5294, N5293, N5292, N5291, N5290, N5289, N5288, N5287, N5286, N5285, N5284, N5283, N5282, N5281, N5280, N5279, N5278, N5277, N5276, N5275, N5274, N5273, N5272, N5271, N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, N5250, N5249, N5248, N5247, N5246, N5245, N5244, N5243, N5242, N5241, N5240, N5239, N5238, N5237, N5236, N5235, N5234, N5233, N5232, N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217, N5216, N5215, N5214, N5213, N5212, N5211, N5210, N5209, N5208, N5207, N5206, N5205, N5204, N5203, N5202, N5201, N5200, N5199, N5198, N5197, N5196, N5195, N5194, N5193, N5192, N5191, N5190, N5189, N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, N5168, N5167, N5166, N5165, N5164, N5163, N5162, N5161, N5160, N5159, N5158, N5157, N5156, N5155, N5154, N5153, N5152, N5151, N5150, N5149, N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135, N5134, N5133, N5132, N5131, N5130, N5129, N5128, N5127, N5126, N5125, N5124, N5123, N5122, N5121, N5120, N5119, N5118, N5117, N5116, N5115, N5114, N5113, N5112, N5111, N5110, N5109, N5108, N5107, N5106, N5105, N5104, N5103, N5102, N5101, N5100, N5099, N5098, N5097, N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487, N4486, N4485, N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421, N4420, N4419, N4418, N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342, N4341, N4340, N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207, N4206, N4205, N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074, N4073, N4072, N4071, N4070, N4069, N4068, N4067, N4066, N4065, N4064, N4063, N4062, N4061, N4060, N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991, N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926, N3925, N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861, N3860, N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251 } = (N48)? { N3250, N3121, N3001, N2881, N2801, N2736, N2671, N2606, N2533, N2468, N2403, N2338, N2273, N2169, N2104, N2007, N1942, N1877, N1812, N1733, N1668, N1603, N1538, N1473, N1408, N1304, N1191, N1078, N1013, N948, N869, N804, N739, N674, N609, N544, N479, N375, N310, N245, N3249, N3120, N3000, N2880, N2800, N2735, N2670, N2605, N2532, N2467, N2402, N2337, N2272, N2168, N2103, N2006, N1941, N1876, N1811, N1732, N1667, N1602, N1537, N1472, N1407, N1303, N1190, N1077, N1012, N947, N868, N803, N738, N673, N608, N543, N478, N374, N309, N244, N3248, N3119, N2999, N2879, N2799, N2734, N2669, N2604, N2531, N2466, N2401, N2336, N2271, N2167, N2102, N2005, N1940, N1875, N1810, N1731, N1666, N1601, N1536, N1471, N1406, N1302, N1189, N1076, N1011, N946, N867, N802, N737, N672, N607, N542, N477, N373, N308, N243, N3247, N3118, N2998, N2878, N2798, N2733, N2668, N2603, N2530, N2465, N2400, N2335, N2270, N2166, N2101, N2004, N1939, N1874, N1809, N1730, N1665, N1600, N1535, N1470, N1405, N1301, N1188, N1075, N1010, N945, N866, N801, N736, N671, N606, N541, N476, N372, N307, N242, N3246, N3117, N2997, N2877, N2797, N2732, N2667, N2602, N2529, N2464, N2399, N2334, N2269, N2165, N2100, N2003, N1938, N1873, N1808, N1729, N1664, N1599, N1534, N1469, N1404, N1300, N1187, N1074, N1009, N944, N865, N800, N735, N670, N605, N540, N475, N371, N306, N241, N3245, N3116, N2996, N2876, N2796, N2731, N2666, N2601, N2528, N2463, N2398, N2333, N2268, N2164, N2099, N2002, N1937, N1872, N1807, N1728, N1663, N1598, N1533, N1468, N1403, N1299, N1186, N1073, N1008, N943, N864, N799, N734, N669, N604, N539, N474, N370, N305, N240, N3244, N3115, N2995, N2875, N2795, N2730, N2665, N2600, N2527, N2462, N2397, N2332, N2267, N2163, N2098, N2001, N1936, N1871, N1806, N1727, N1662, N1597, N1532, N1467, N1402, N1298, N1185, N1072, N1007, N942, N863, N798, N733, N668, N603, N538, N473, N369, N304, N239, N3243, N3114, N2994, N2874, N2794, N2729, N2664, N2599, N2526, N2461, N2396, N2331, N2266, N2162, N2097, N2000, N1935, N1870, N1805, N1726, N1661, N1596, N1531, N1466, N1401, N1297, N1184, N1071, N1006, N941, N862, N797, N732, N667, N602, N537, N472, N368, N303, N238, N3242, N3113, N2993, N2873, N2793, N2728, N2663, N2598, N2525, N2460, N2395, N2330, N2265, N2161, N2096, N1999, N1934, N1869, N1804, N1725, N1660, N1595, N1530, N1465, N1400, N1296, N1183, N1070, N1005, N940, N861, N796, N731, N666, N601, N536, N471, N367, N302, N237, N3241, N3112, N2992, N2872, N2792, N2727, N2662, N2597, N2524, N2459, N2394, N2329, N2264, N2160, N2095, N1998, N1933, N1868, N1803, N1724, N1659, N1594, N1529, N1464, N1399, N1295, N1182, N1069, N1004, N939, N860, N795, N730, N665, N600, N535, N470, N366, N301, N236, N3240, N3111, N2991, N2871, N2791, N2726, N2661, N2596, N2523, N2458, N2393, N2328, N2263, N2159, N2094, N1997, N1932, N1867, N1802, N1723, N1658, N1593, N1528, N1463, N1398, N1294, N1181, N1068, N1003, N938, N859, N794, N729, N664, N599, N534, N469, N365, N300, N235, N3239, N3110, N2990, N2870, N2790, N2725, N2660, N2595, N2522, N2457, N2392, N2327, N2262, N2158, N2093, N1996, N1931, N1866, N1801, N1722, N1657, N1592, N1527, N1462, N1397, N1293, N1180, N1067, N1002, N937, N858, N793, N728, N663, N598, N533, N468, N364, N299, N234, N3238, N3109, N2989, N2869, N2789, N2724, N2659, N2594, N2521, N2456, N2391, N2326, N2261, N2157, N2092, N1995, N1930, N1865, N1800, N1721, N1656, N1591, N1526, N1461, N1396, N1292, N1179, N1066, N1001, N936, N857, N792, N727, N662, N597, N532, N467, N363, N298, N233, N3237, N3108, N2988, N2868, N2788, N2723, N2658, N2593, N2520, N2455, N2390, N2325, N2260, N2156, N2091, N1994, N1929, N1864, N1799, N1720, N1655, N1590, N1525, N1460, N1395, N1291, N1178, N1065, N1000, N935, N856, N791, N726, N661, N596, N531, N466, N362, N297, N232, N3236, N3107, N2987, N2867, N2787, N2722, N2657, N2592, N2519, N2454, N2389, N2324, N2259, N2155, N2090, N1993, N1928, N1863, N1798, N1719, N1654, N1589, N1524, N1459, N1394, N1290, N1177, N1064, N999, N934, N855, N790, N725, N660, N595, N530, N465, N361, N296, N231, N3235, N3106, N2986, N2866, N2786, N2721, N2656, N2591, N2518, N2453, N2388, N2323, N2258, N2154, N2089, N1992, N1927, N1862, N1797, N1718, N1653, N1588, N1523, N1458, N1393, N1289, N1176, N1063, N998, N933, N854, N789, N724, N659, N594, N529, N464, N360, N295, N230, N3234, N3105, N2985, N2865, N2785, N2720, N2655, N2590, N2517, N2452, N2387, N2322, N2257, N2153, N2088, N1991, N1926, N1861, N1796, N1717, N1652, N1587, N1522, N1457, N1392, N1288, N1175, N1062, N997, N932, N853, N788, N723, N658, N593, N528, N463, N359, N294, N229, N3233, N3104, N2984, N2864, N2784, N2719, N2654, N2589, N2516, N2451, N2386, N2321, N2256, N2152, N2087, N1990, N1925, N1860, N1795, N1716, N1651, N1586, N1521, N1456, N1391, N1287, N1174, N1061, N996, N931, N852, N787, N722, N657, N592, N527, N462, N358, N293, N228, N3232, N3103, N2983, N2863, N2783, N2718, N2653, N2588, N2515, N2450, N2385, N2320, N2255, N2151, N2086, N1989, N1924, N1859, N1794, N1715, N1650, N1585, N1520, N1455, N1390, N1286, N1173, N1060, N995, N930, N851, N786, N721, N656, N591, N526, N461, N357, N292, N227, N3231, N3102, N2982, N2862, N2782, N2717, N2652, N2587, N2514, N2449, N2384, N2319, N2254, N2150, N2085, N1988, N1923, N1858, N1793, N1714, N1649, N1584, N1519, N1454, N1389, N1285, N1172, N1059, N994, N929, N850, N785, N720, N655, N590, N525, N460, N356, N291, N226, N3230, N3101, N2981, N2861, N2781, N2716, N2651, N2586, N2513, N2448, N2383, N2318, N2253, N2149, N2084, N1987, N1922, N1857, N1792, N1713, N1648, N1583, N1518, N1453, N1388, N1284, N1171, N1058, N993, N928, N849, N784, N719, N654, N589, N524, N459, N355, N290, N225, N3229, N3100, N2980, N2860, N2780, N2715, N2650, N2585, N2512, N2447, N2382, N2317, N2252, N2148, N2083, N1986, N1921, N1856, N1791, N1712, N1647, N1582, N1517, N1452, N1387, N1283, N1170, N1057, N992, N927, N848, N783, N718, N653, N588, N523, N458, N354, N289, N224, N3228, N3099, N2979, N2859, N2779, N2714, N2649, N2584, N2511, N2446, N2381, N2316, N2251, N2147, N2082, N1985, N1920, N1855, N1790, N1711, N1646, N1581, N1516, N1451, N1386, N1282, N1169, N1056, N991, N926, N847, N782, N717, N652, N587, N522, N457, N353, N288, N223, N3227, N3098, N2978, N2858, N2778, N2713, N2648, N2583, N2510, N2445, N2380, N2315, N2250, N2146, N2081, N1984, N1919, N1854, N1789, N1710, N1645, N1580, N1515, N1450, N1385, N1281, N1168, N1055, N990, N925, N846, N781, N716, N651, N586, N521, N456, N352, N287, N222, N3226, N3097, N2977, N2857, N2777, N2712, N2647, N2582, N2509, N2444, N2379, N2314, N2249, N2145, N2080, N1983, N1918, N1853, N1788, N1709, N1644, N1579, N1514, N1449, N1384, N1280, N1167, N1054, N989, N924, N845, N780, N715, N650, N585, N520, N455, N351, N286, N221, N3225, N3096, N2976, N2856, N2776, N2711, N2646, N2581, N2508, N2443, N2378, N2313, N2248, N2144, N2079, N1982, N1917, N1852, N1787, N1708, N1643, N1578, N1513, N1448, N1383, N1279, N1166, N1053, N988, N923, N844, N779, N714, N649, N584, N519, N454, N350, N285, N220, N3224, N3095, N2975, N2855, N2775, N2710, N2645, N2580, N2507, N2442, N2377, N2312, N2247, N2143, N2078, N1981, N1916, N1851, N1786, N1707, N1642, N1577, N1512, N1447, N1382, N1278, N1165, N1052, N987, N922, N843, N778, N713, N648, N583, N518, N453, N349, N284, N219, N3223, N3094, N2974, N2854, N2774, N2709, N2644, N2579, N2506, N2441, N2376, N2311, N2246, N2142, N2077, N1980, N1915, N1850, N1785, N1706, N1641, N1576, N1511, N1446, N1381, N1277, N1164, N1051, N986, N921, N842, N777, N712, N647, N582, N517, N452, N348, N283, N218, N3222, N3093, N2973, N2853, N2773, N2708, N2643, N2578, N2505, N2440, N2375, N2310, N2245, N2141, N2076, N1979, N1914, N1849, N1784, N1705, N1640, N1575, N1510, N1445, N1380, N1276, N1163, N1050, N985, N920, N841, N776, N711, N646, N581, N516, N451, N347, N282, N217, N3221, N3092, N2972, N2852, N2772, N2707, N2642, N2577, N2504, N2439, N2374, N2309, N2244, N2140, N2075, N1978, N1913, N1848, N1783, N1704, N1639, N1574, N1509, N1444, N1379, N1275, N1162, N1049, N984, N919, N840, N775, N710, N645, N580, N515, N450, N346, N281, N216, N3220, N3091, N2971, N2851, N2771, N2706, N2641, N2576, N2503, N2438, N2373, N2308, N2243, N2139, N2074, N1977, N1912, N1847, N1782, N1703, N1638, N1573, N1508, N1443, N1378, N1274, N1161, N1048, N983, N918, N839, N774, N709, N644, N579, N514, N449, N345, N280, N215, N3219, N3090, N2970, N2850, N2770, N2705, N2640, N2575, N2502, N2437, N2372, N2307, N2242, N2138, N2073, N1976, N1911, N1846, N1781, N1702, N1637, N1572, N1507, N1442, N1377, N1273, N1160, N1047, N982, N917, N838, N773, N708, N643, N578, N513, N448, N344, N279, N214, N3218, N3089, N2969, N2849, N2769, N2704, N2639, N2574, N2501, N2436, N2371, N2306, N2241, N2137, N2072, N1975, N1910, N1845, N1780, N1701, N1636, N1571, N1506, N1441, N1376, N1272, N1159, N1046, N981, N916, N837, N772, N707, N642, N577, N512, N447, N343, N278, N213, N3217, N3088, N2968, N2848, N2768, N2703, N2638, N2573, N2500, N2435, N2370, N2305, N2240, N2136, N2071, N1974, N1909, N1844, N1779, N1700, N1635, N1570, N1505, N1440, N1375, N1271, N1158, N1045, N980, N915, N836, N771, N706, N641, N576, N511, N446, N342, N277, N212, N3216, N3087, N2967, N2847, N2767, N2702, N2637, N2572, N2499, N2434, N2369, N2304, N2239, N2135, N2070, N1973, N1908, N1843, N1778, N1699, N1634, N1569, N1504, N1439, N1374, N1270, N1157, N1044, N979, N914, N835, N770, N705, N640, N575, N510, N445, N341, N276, N211, N3215, N3086, N2966, N2846, N2766, N2701, N2636, N2571, N2498, N2433, N2368, N2303, N2238, N2134, N2069, N1972, N1907, N1842, N1777, N1698, N1633, N1568, N1503, N1438, N1373, N1269, N1156, N1043, N978, N913, N834, N769, N704, N639, N574, N509, N444, N340, N275, N210, N3214, N3085, N2965, N2845, N2765, N2700, N2635, N2570, N2497, N2432, N2367, N2302, N2237, N2133, N2068, N1971, N1906, N1841, N1776, N1697, N1632, N1567, N1502, N1437, N1372, N1268, N1155, N1042, N977, N912, N833, N768, N703, N638, N573, N508, N443, N339, N274, N209, N3213, N3084, N2964, N2844, N2764, N2699, N2634, N2569, N2496, N2431, N2366, N2301, N2236, N2132, N2067, N1970, N1905, N1840, N1775, N1696, N1631, N1566, N1501, N1436, N1371, N1267, N1154, N1041, N976, N911, N832, N767, N702, N637, N572, N507, N442, N338, N273, N208, N3212, N3083, N2963, N2843, N2763, N2698, N2633, N2568, N2495, N2430, N2365, N2300, N2235, N2131, N2066, N1969, N1904, N1839, N1774, N1695, N1630, N1565, N1500, N1435, N1370, N1266, N1153, N1040, N975, N910, N831, N766, N701, N636, N571, N506, N441, N337, N272, N207, N3211, N3082, N2962, N2842, N2762, N2697, N2632, N2567, N2494, N2429, N2364, N2299, N2234, N2130, N2065, N1968, N1903, N1838, N1773, N1694, N1629, N1564, N1499, N1434, N1369, N1265, N1152, N1039, N974, N909, N830, N765, N700, N635, N570, N505, N440, N336, N271, N206, N3210, N3081, N2961, N2841, N2761, N2696, N2631, N2566, N2493, N2428, N2363, N2298, N2233, N2129, N2064, N1967, N1902, N1837, N1772, N1693, N1628, N1563, N1498, N1433, N1368, N1264, N1151, N1038, N973, N908, N829, N764, N699, N634, N569, N504, N439, N335, N270, N205, N3209, N3080, N2960, N2840, N2760, N2695, N2630, N2565, N2492, N2427, N2362, N2297, N2232, N2128, N2063, N1966, N1901, N1836, N1771, N1692, N1627, N1562, N1497, N1432, N1367, N1263, N1150, N1037, N972, N907, N828, N763, N698, N633, N568, N503, N438, N334, N269, N204, N3208, N3079, N2959, N2839, N2759, N2694, N2629, N2564, N2491, N2426, N2361, N2296, N2231, N2127, N2062, N1965, N1900, N1835, N1770, N1691, N1626, N1561, N1496, N1431, N1366, N1262, N1149, N1036, N971, N906, N827, N762, N697, N632, N567, N502, N437, N333, N268, N203, N3207, N3078, N2958, N2838, N2758, N2693, N2628, N2563, N2490, N2425, N2360, N2295, N2230, N2126, N2061, N1964, N1899, N1834, N1769, N1690, N1625, N1560, N1495, N1430, N1365, N1261, N1148, N1035, N970, N905, N826, N761, N696, N631, N566, N501, N436, N332, N267, N202, N3206, N3077, N2957, N2837, N2757, N2692, N2627, N2562, N2489, N2424, N2359, N2294, N2229, N2125, N2060, N1963, N1898, N1833, N1768, N1689, N1624, N1559, N1494, N1429, N1364, N1260, N1147, N1034, N969, N904, N825, N760, N695, N630, N565, N500, N435, N331, N266, N201, N3205, N3076, N2956, N2836, N2756, N2691, N2626, N2561, N2488, N2423, N2358, N2293, N2228, N2124, N2059, N1962, N1897, N1832, N1767, N1688, N1623, N1558, N1493, N1428, N1363, N1259, N1146, N1033, N968, N903, N824, N759, N694, N629, N564, N499, N434, N330, N265, N200, N3204, N3075, N2955, N2835, N2755, N2690, N2625, N2560, N2487, N2422, N2357, N2292, N2227, N2123, N2058, N1961, N1896, N1831, N1766, N1687, N1622, N1557, N1492, N1427, N1362, N1258, N1145, N1032, N967, N902, N823, N758, N693, N628, N563, N498, N433, N329, N264, N199, N3203, N3074, N2954, N2834, N2754, N2689, N2624, N2559, N2486, N2421, N2356, N2291, N2226, N2122, N2057, N1960, N1895, N1830, N1765, N1686, N1621, N1556, N1491, N1426, N1361, N1257, N1144, N1031, N966, N901, N822, N757, N692, N627, N562, N497, N432, N328, N263, N198, N3202, N3073, N2953, N2833, N2753, N2688, N2623, N2558, N2485, N2420, N2355, N2290, N2225, N2121, N2056, N1959, N1894, N1829, N1764, N1685, N1620, N1555, N1490, N1425, N1360, N1256, N1143, N1030, N965, N900, N821, N756, N691, N626, N561, N496, N431, N327, N262, N197, N3201, N3072, N2952, N2832, N2752, N2687, N2622, N2557, N2484, N2419, N2354, N2289, N2224, N2120, N2055, N1958, N1893, N1828, N1763, N1684, N1619, N1554, N1489, N1424, N1359, N1255, N1142, N1029, N964, N899, N820, N755, N690, N625, N560, N495, N430, N326, N261, N196, N3200, N3071, N2951, N2831, N2751, N2686, N2621, N2556, N2483, N2418, N2353, N2288, N2223, N2119, N2054, N1957, N1892, N1827, N1762, N1683, N1618, N1553, N1488, N1423, N1358, N1254, N1141, N1028, N963, N898, N819, N754, N689, N624, N559, N494, N429, N325, N260, N195, N3199, N3070, N2950, N2830, N2750, N2685, N2620, N2555, N2482, N2417, N2352, N2287, N2222, N2118, N2053, N1956, N1891, N1826, N1761, N1682, N1617, N1552, N1487, N1422, N1357, N1253, N1140, N1027, N962, N897, N818, N753, N688, N623, N558, N493, N428, N324, N259, N194, N3198, N3069, N2949, N2829, N2749, N2684, N2619, N2554, N2481, N2416, N2351, N2286, N2221, N2117, N2052, N1955, N1890, N1825, N1760, N1681, N1616, N1551, N1486, N1421, N1356, N1252, N1139, N1026, N961, N896, N817, N752, N687, N622, N557, N492, N427, N323, N258, N193, N3197, N3068, N2948, N2828, N2748, N2683, N2618, N2553, N2480, N2415, N2350, N2285, N2220, N2116, N2051, N1954, N1889, N1824, N1759, N1680, N1615, N1550, N1485, N1420, N1355, N1251, N1138, N1025, N960, N895, N816, N751, N686, N621, N556, N491, N426, N322, N257, N192, N3196, N3067, N2947, N2827, N2747, N2682, N2617, N2552, N2479, N2414, N2349, N2284, N2219, N2115, N2050, N1953, N1888, N1823, N1758, N1679, N1614, N1549, N1484, N1419, N1354, N1250, N1137, N1024, N959, N894, N815, N750, N685, N620, N555, N490, N425, N321, N256, N191, N3195, N3066, N2946, N2826, N2746, N2681, N2616, N2551, N2478, N2413, N2348, N2283, N2218, N2114, N2049, N1952, N1887, N1822, N1757, N1678, N1613, N1548, N1483, N1418, N1353, N1249, N1136, N1023, N958, N893, N814, N749, N684, N619, N554, N489, N424, N320, N255, N190, N3194, N3065, N2945, N2825, N2745, N2680, N2615, N2550, N2477, N2412, N2347, N2282, N2217, N2113, N2048, N1951, N1886, N1821, N1756, N1677, N1612, N1547, N1482, N1417, N1352, N1248, N1135, N1022, N957, N892, N813, N748, N683, N618, N553, N488, N423, N319, N254, N189, N3193, N3064, N2944, N2824, N2744, N2679, N2614, N2549, N2476, N2411, N2346, N2281, N2216, N2112, N2047, N1950, N1885, N1820, N1755, N1676, N1611, N1546, N1481, N1416, N1351, N1247, N1134, N1021, N956, N891, N812, N747, N682, N617, N552, N487, N422, N318, N253, N188, N3192, N3063, N2943, N2823, N2743, N2678, N2613, N2548, N2475, N2410, N2345, N2280, N2215, N2111, N2046, N1949, N1884, N1819, N1754, N1675, N1610, N1545, N1480, N1415, N1350, N1246, N1133, N1020, N955, N890, N811, N746, N681, N616, N551, N486, N421, N317, N252, N187, N3191, N3062, N2942, N2822, N2742, N2677, N2612, N2547, N2474, N2409, N2344, N2279, N2214, N2110, N2045, N1948, N1883, N1818, N1753, N1674, N1609, N1544, N1479, N1414, N1349, N1245, N1132, N1019, N954, N889, N810, N745, N680, N615, N550, N485, N420, N316, N251, N186, N3190, N3061, N2941, N2821, N2741, N2676, N2611, N2546, N2473, N2408, N2343, N2278, N2213, N2109, N2044, N1947, N1882, N1817, N1752, N1673, N1608, N1543, N1478, N1413, N1348, N1244, N1131, N1018, N953, N888, N809, N744, N679, N614, N549, N484, N419, N315, N250, N185, N3189, N3060, N2940, N2820, N2740, N2675, N2610, N2545, N2472, N2407, N2342, N2277, N2212, N2108, N2043, N1946, N1881, N1816, N1751, N1672, N1607, N1542, N1477, N1412, N1347, N1243, N1130, N1017, N952, N887, N808, N743, N678, N613, N548, N483, N418, N314, N249, N184, N3188, N3059, N2939, N2819, N2739, N2674, N2609, N2544, N2471, N2406, N2341, N2276, N2211, N2107, N2042, N1945, N1880, N1815, N1750, N1671, N1606, N1541, N1476, N1411, N1346, N1242, N1129, N1016, N951, N886, N807, N742, N677, N612, N547, N482, N417, N313, N248, N183, N3187, N3058, N2938, N2818, N2738, N2673, N2608, N2543, N2470, N2405, N2340, N2275, N2210, N2106, N2041, N1944, N1879, N1814, N1749, N1670, N1605, N1540, N1475, N1410, N1345, N1241, N1128, N1015, N950, N885, N806, N741, N676, N611, N546, N481, N416, N312, N247, N182 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N180)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N48 = N179;
  assign \nz.read_en  = v_i & N5893;
  assign N5893 = ~w_i;
  assign N49 = ~\nz.addr_r [0];
  assign N50 = ~\nz.addr_r [1];
  assign N51 = N49 & N50;
  assign N52 = N49 & \nz.addr_r [1];
  assign N53 = \nz.addr_r [0] & N50;
  assign N54 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N55 = ~\nz.addr_r [2];
  assign N56 = N51 & N55;
  assign N57 = N51 & \nz.addr_r [2];
  assign N58 = N53 & N55;
  assign N59 = N53 & \nz.addr_r [2];
  assign N60 = N52 & N55;
  assign N61 = N52 & \nz.addr_r [2];
  assign N62 = N54 & N55;
  assign N63 = N54 & \nz.addr_r [2];
  assign N64 = ~\nz.addr_r [3];
  assign N65 = N56 & N64;
  assign N66 = N56 & \nz.addr_r [3];
  assign N67 = N58 & N64;
  assign N68 = N58 & \nz.addr_r [3];
  assign N69 = N60 & N64;
  assign N70 = N60 & \nz.addr_r [3];
  assign N71 = N62 & N64;
  assign N72 = N62 & \nz.addr_r [3];
  assign N73 = N57 & N64;
  assign N74 = N57 & \nz.addr_r [3];
  assign N75 = N59 & N64;
  assign N76 = N59 & \nz.addr_r [3];
  assign N77 = N61 & N64;
  assign N78 = N61 & \nz.addr_r [3];
  assign N79 = N63 & N64;
  assign N80 = N63 & \nz.addr_r [3];
  assign N81 = ~\nz.addr_r [4];
  assign N82 = N65 & N81;
  assign N83 = N65 & \nz.addr_r [4];
  assign N84 = N67 & N81;
  assign N85 = N67 & \nz.addr_r [4];
  assign N86 = N69 & N81;
  assign N87 = N69 & \nz.addr_r [4];
  assign N88 = N71 & N81;
  assign N89 = N71 & \nz.addr_r [4];
  assign N90 = N73 & N81;
  assign N91 = N73 & \nz.addr_r [4];
  assign N92 = N75 & N81;
  assign N93 = N75 & \nz.addr_r [4];
  assign N94 = N77 & N81;
  assign N95 = N77 & \nz.addr_r [4];
  assign N96 = N79 & N81;
  assign N97 = N79 & \nz.addr_r [4];
  assign N98 = N66 & N81;
  assign N99 = N66 & \nz.addr_r [4];
  assign N100 = N68 & N81;
  assign N101 = N68 & \nz.addr_r [4];
  assign N102 = N70 & N81;
  assign N103 = N70 & \nz.addr_r [4];
  assign N104 = N72 & N81;
  assign N105 = N72 & \nz.addr_r [4];
  assign N106 = N74 & N81;
  assign N107 = N74 & \nz.addr_r [4];
  assign N108 = N76 & N81;
  assign N109 = N76 & \nz.addr_r [4];
  assign N110 = N78 & N81;
  assign N111 = N78 & \nz.addr_r [4];
  assign N112 = N80 & N81;
  assign N113 = N80 & \nz.addr_r [4];
  assign N114 = ~\nz.addr_r [5];
  assign N115 = N82 & N114;
  assign N116 = N82 & \nz.addr_r [5];
  assign N117 = N84 & N114;
  assign N118 = N84 & \nz.addr_r [5];
  assign N119 = N86 & N114;
  assign N120 = N86 & \nz.addr_r [5];
  assign N121 = N88 & N114;
  assign N122 = N88 & \nz.addr_r [5];
  assign N123 = N90 & N114;
  assign N124 = N90 & \nz.addr_r [5];
  assign N125 = N92 & N114;
  assign N126 = N92 & \nz.addr_r [5];
  assign N127 = N94 & N114;
  assign N128 = N94 & \nz.addr_r [5];
  assign N129 = N96 & N114;
  assign N130 = N96 & \nz.addr_r [5];
  assign N131 = N98 & N114;
  assign N132 = N98 & \nz.addr_r [5];
  assign N133 = N100 & N114;
  assign N134 = N100 & \nz.addr_r [5];
  assign N135 = N102 & N114;
  assign N136 = N102 & \nz.addr_r [5];
  assign N137 = N104 & N114;
  assign N138 = N104 & \nz.addr_r [5];
  assign N139 = N106 & N114;
  assign N140 = N106 & \nz.addr_r [5];
  assign N141 = N108 & N114;
  assign N142 = N108 & \nz.addr_r [5];
  assign N143 = N110 & N114;
  assign N144 = N110 & \nz.addr_r [5];
  assign N145 = N112 & N114;
  assign N146 = N112 & \nz.addr_r [5];
  assign N147 = N83 & N114;
  assign N148 = N83 & \nz.addr_r [5];
  assign N149 = N85 & N114;
  assign N150 = N85 & \nz.addr_r [5];
  assign N151 = N87 & N114;
  assign N152 = N87 & \nz.addr_r [5];
  assign N153 = N89 & N114;
  assign N154 = N89 & \nz.addr_r [5];
  assign N155 = N91 & N114;
  assign N156 = N91 & \nz.addr_r [5];
  assign N157 = N93 & N114;
  assign N158 = N93 & \nz.addr_r [5];
  assign N159 = N95 & N114;
  assign N160 = N95 & \nz.addr_r [5];
  assign N161 = N97 & N114;
  assign N162 = N97 & \nz.addr_r [5];
  assign N163 = N99 & N114;
  assign N164 = N99 & \nz.addr_r [5];
  assign N165 = N101 & N114;
  assign N166 = N101 & \nz.addr_r [5];
  assign N167 = N103 & N114;
  assign N168 = N103 & \nz.addr_r [5];
  assign N169 = N105 & N114;
  assign N170 = N105 & \nz.addr_r [5];
  assign N171 = N107 & N114;
  assign N172 = N107 & \nz.addr_r [5];
  assign N173 = N109 & N114;
  assign N174 = N109 & \nz.addr_r [5];
  assign N175 = N111 & N114;
  assign N176 = N111 & \nz.addr_r [5];
  assign N177 = N113 & N114;
  assign N178 = N113 & \nz.addr_r [5];
  assign N179 = v_i & w_i;
  assign N180 = ~N179;
  assign N181 = ~w_mask_i[0];
  assign N246 = ~w_mask_i[1];
  assign N311 = ~w_mask_i[2];
  assign N376 = ~w_mask_i[3];
  assign N480 = ~w_mask_i[4];
  assign N545 = ~w_mask_i[5];
  assign N610 = ~w_mask_i[6];
  assign N675 = ~w_mask_i[7];
  assign N740 = ~w_mask_i[8];
  assign N805 = ~w_mask_i[9];
  assign N870 = ~w_mask_i[10];
  assign N949 = ~w_mask_i[11];
  assign N1014 = ~w_mask_i[12];
  assign N1079 = ~w_mask_i[13];
  assign N1192 = ~w_mask_i[14];
  assign N1305 = ~w_mask_i[15];
  assign N1409 = ~w_mask_i[16];
  assign N1474 = ~w_mask_i[17];
  assign N1539 = ~w_mask_i[18];
  assign N1604 = ~w_mask_i[19];
  assign N1669 = ~w_mask_i[20];
  assign N1734 = ~w_mask_i[21];
  assign N1813 = ~w_mask_i[22];
  assign N1878 = ~w_mask_i[23];
  assign N1943 = ~w_mask_i[24];
  assign N2008 = ~w_mask_i[25];
  assign N2105 = ~w_mask_i[26];
  assign N2170 = ~w_mask_i[27];
  assign N2274 = ~w_mask_i[28];
  assign N2339 = ~w_mask_i[29];
  assign N2404 = ~w_mask_i[30];
  assign N2469 = ~w_mask_i[31];
  assign N2534 = ~w_mask_i[32];
  assign N2607 = ~w_mask_i[33];
  assign N2672 = ~w_mask_i[34];
  assign N2737 = ~w_mask_i[35];
  assign N2802 = ~w_mask_i[36];
  assign N2882 = ~w_mask_i[37];
  assign N3002 = ~w_mask_i[38];
  assign N3122 = ~w_mask_i[39];

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N5810) begin
      \nz.mem_2559_sv2v_reg  <= data_i[39];
    end 
    if(N5809) begin
      \nz.mem_2558_sv2v_reg  <= data_i[38];
    end 
    if(N5808) begin
      \nz.mem_2557_sv2v_reg  <= data_i[37];
    end 
    if(N5807) begin
      \nz.mem_2556_sv2v_reg  <= data_i[36];
    end 
    if(N5806) begin
      \nz.mem_2555_sv2v_reg  <= data_i[35];
    end 
    if(N5805) begin
      \nz.mem_2554_sv2v_reg  <= data_i[34];
    end 
    if(N5804) begin
      \nz.mem_2553_sv2v_reg  <= data_i[33];
    end 
    if(N5803) begin
      \nz.mem_2552_sv2v_reg  <= data_i[32];
    end 
    if(N5802) begin
      \nz.mem_2551_sv2v_reg  <= data_i[31];
    end 
    if(N5801) begin
      \nz.mem_2550_sv2v_reg  <= data_i[30];
    end 
    if(N5800) begin
      \nz.mem_2549_sv2v_reg  <= data_i[29];
    end 
    if(N5799) begin
      \nz.mem_2548_sv2v_reg  <= data_i[28];
    end 
    if(N5798) begin
      \nz.mem_2547_sv2v_reg  <= data_i[27];
    end 
    if(N5797) begin
      \nz.mem_2546_sv2v_reg  <= data_i[26];
    end 
    if(N5796) begin
      \nz.mem_2545_sv2v_reg  <= data_i[25];
    end 
    if(N5795) begin
      \nz.mem_2544_sv2v_reg  <= data_i[24];
    end 
    if(N5794) begin
      \nz.mem_2543_sv2v_reg  <= data_i[23];
    end 
    if(N5793) begin
      \nz.mem_2542_sv2v_reg  <= data_i[22];
    end 
    if(N5792) begin
      \nz.mem_2541_sv2v_reg  <= data_i[21];
    end 
    if(N5791) begin
      \nz.mem_2540_sv2v_reg  <= data_i[20];
    end 
    if(N5790) begin
      \nz.mem_2539_sv2v_reg  <= data_i[19];
    end 
    if(N5789) begin
      \nz.mem_2538_sv2v_reg  <= data_i[18];
    end 
    if(N5788) begin
      \nz.mem_2537_sv2v_reg  <= data_i[17];
    end 
    if(N5787) begin
      \nz.mem_2536_sv2v_reg  <= data_i[16];
    end 
    if(N5786) begin
      \nz.mem_2535_sv2v_reg  <= data_i[15];
    end 
    if(N5785) begin
      \nz.mem_2534_sv2v_reg  <= data_i[14];
    end 
    if(N5784) begin
      \nz.mem_2533_sv2v_reg  <= data_i[13];
    end 
    if(N5783) begin
      \nz.mem_2532_sv2v_reg  <= data_i[12];
    end 
    if(N5782) begin
      \nz.mem_2531_sv2v_reg  <= data_i[11];
    end 
    if(N5781) begin
      \nz.mem_2530_sv2v_reg  <= data_i[10];
    end 
    if(N5780) begin
      \nz.mem_2529_sv2v_reg  <= data_i[9];
    end 
    if(N5779) begin
      \nz.mem_2528_sv2v_reg  <= data_i[8];
    end 
    if(N5778) begin
      \nz.mem_2527_sv2v_reg  <= data_i[7];
    end 
    if(N5777) begin
      \nz.mem_2526_sv2v_reg  <= data_i[6];
    end 
    if(N5776) begin
      \nz.mem_2525_sv2v_reg  <= data_i[5];
    end 
    if(N5775) begin
      \nz.mem_2524_sv2v_reg  <= data_i[4];
    end 
    if(N5774) begin
      \nz.mem_2523_sv2v_reg  <= data_i[3];
    end 
    if(N5773) begin
      \nz.mem_2522_sv2v_reg  <= data_i[2];
    end 
    if(N5772) begin
      \nz.mem_2521_sv2v_reg  <= data_i[1];
    end 
    if(N5771) begin
      \nz.mem_2520_sv2v_reg  <= data_i[0];
    end 
    if(N5770) begin
      \nz.mem_2519_sv2v_reg  <= data_i[39];
    end 
    if(N5769) begin
      \nz.mem_2518_sv2v_reg  <= data_i[38];
    end 
    if(N5768) begin
      \nz.mem_2517_sv2v_reg  <= data_i[37];
    end 
    if(N5767) begin
      \nz.mem_2516_sv2v_reg  <= data_i[36];
    end 
    if(N5766) begin
      \nz.mem_2515_sv2v_reg  <= data_i[35];
    end 
    if(N5765) begin
      \nz.mem_2514_sv2v_reg  <= data_i[34];
    end 
    if(N5764) begin
      \nz.mem_2513_sv2v_reg  <= data_i[33];
    end 
    if(N5763) begin
      \nz.mem_2512_sv2v_reg  <= data_i[32];
    end 
    if(N5762) begin
      \nz.mem_2511_sv2v_reg  <= data_i[31];
    end 
    if(N5761) begin
      \nz.mem_2510_sv2v_reg  <= data_i[30];
    end 
    if(N5760) begin
      \nz.mem_2509_sv2v_reg  <= data_i[29];
    end 
    if(N5759) begin
      \nz.mem_2508_sv2v_reg  <= data_i[28];
    end 
    if(N5758) begin
      \nz.mem_2507_sv2v_reg  <= data_i[27];
    end 
    if(N5757) begin
      \nz.mem_2506_sv2v_reg  <= data_i[26];
    end 
    if(N5756) begin
      \nz.mem_2505_sv2v_reg  <= data_i[25];
    end 
    if(N5755) begin
      \nz.mem_2504_sv2v_reg  <= data_i[24];
    end 
    if(N5754) begin
      \nz.mem_2503_sv2v_reg  <= data_i[23];
    end 
    if(N5753) begin
      \nz.mem_2502_sv2v_reg  <= data_i[22];
    end 
    if(N5752) begin
      \nz.mem_2501_sv2v_reg  <= data_i[21];
    end 
    if(N5751) begin
      \nz.mem_2500_sv2v_reg  <= data_i[20];
    end 
    if(N5750) begin
      \nz.mem_2499_sv2v_reg  <= data_i[19];
    end 
    if(N5749) begin
      \nz.mem_2498_sv2v_reg  <= data_i[18];
    end 
    if(N5748) begin
      \nz.mem_2497_sv2v_reg  <= data_i[17];
    end 
    if(N5747) begin
      \nz.mem_2496_sv2v_reg  <= data_i[16];
    end 
    if(N5746) begin
      \nz.mem_2495_sv2v_reg  <= data_i[15];
    end 
    if(N5745) begin
      \nz.mem_2494_sv2v_reg  <= data_i[14];
    end 
    if(N5744) begin
      \nz.mem_2493_sv2v_reg  <= data_i[13];
    end 
    if(N5743) begin
      \nz.mem_2492_sv2v_reg  <= data_i[12];
    end 
    if(N5742) begin
      \nz.mem_2491_sv2v_reg  <= data_i[11];
    end 
    if(N5741) begin
      \nz.mem_2490_sv2v_reg  <= data_i[10];
    end 
    if(N5740) begin
      \nz.mem_2489_sv2v_reg  <= data_i[9];
    end 
    if(N5739) begin
      \nz.mem_2488_sv2v_reg  <= data_i[8];
    end 
    if(N5738) begin
      \nz.mem_2487_sv2v_reg  <= data_i[7];
    end 
    if(N5737) begin
      \nz.mem_2486_sv2v_reg  <= data_i[6];
    end 
    if(N5736) begin
      \nz.mem_2485_sv2v_reg  <= data_i[5];
    end 
    if(N5735) begin
      \nz.mem_2484_sv2v_reg  <= data_i[4];
    end 
    if(N5734) begin
      \nz.mem_2483_sv2v_reg  <= data_i[3];
    end 
    if(N5733) begin
      \nz.mem_2482_sv2v_reg  <= data_i[2];
    end 
    if(N5732) begin
      \nz.mem_2481_sv2v_reg  <= data_i[1];
    end 
    if(N5731) begin
      \nz.mem_2480_sv2v_reg  <= data_i[0];
    end 
    if(N5730) begin
      \nz.mem_2479_sv2v_reg  <= data_i[39];
    end 
    if(N5729) begin
      \nz.mem_2478_sv2v_reg  <= data_i[38];
    end 
    if(N5728) begin
      \nz.mem_2477_sv2v_reg  <= data_i[37];
    end 
    if(N5727) begin
      \nz.mem_2476_sv2v_reg  <= data_i[36];
    end 
    if(N5726) begin
      \nz.mem_2475_sv2v_reg  <= data_i[35];
    end 
    if(N5725) begin
      \nz.mem_2474_sv2v_reg  <= data_i[34];
    end 
    if(N5724) begin
      \nz.mem_2473_sv2v_reg  <= data_i[33];
    end 
    if(N5723) begin
      \nz.mem_2472_sv2v_reg  <= data_i[32];
    end 
    if(N5722) begin
      \nz.mem_2471_sv2v_reg  <= data_i[31];
    end 
    if(N5721) begin
      \nz.mem_2470_sv2v_reg  <= data_i[30];
    end 
    if(N5720) begin
      \nz.mem_2469_sv2v_reg  <= data_i[29];
    end 
    if(N5719) begin
      \nz.mem_2468_sv2v_reg  <= data_i[28];
    end 
    if(N5718) begin
      \nz.mem_2467_sv2v_reg  <= data_i[27];
    end 
    if(N5717) begin
      \nz.mem_2466_sv2v_reg  <= data_i[26];
    end 
    if(N5716) begin
      \nz.mem_2465_sv2v_reg  <= data_i[25];
    end 
    if(N5715) begin
      \nz.mem_2464_sv2v_reg  <= data_i[24];
    end 
    if(N5714) begin
      \nz.mem_2463_sv2v_reg  <= data_i[23];
    end 
    if(N5713) begin
      \nz.mem_2462_sv2v_reg  <= data_i[22];
    end 
    if(N5712) begin
      \nz.mem_2461_sv2v_reg  <= data_i[21];
    end 
    if(N5711) begin
      \nz.mem_2460_sv2v_reg  <= data_i[20];
    end 
    if(N5710) begin
      \nz.mem_2459_sv2v_reg  <= data_i[19];
    end 
    if(N5709) begin
      \nz.mem_2458_sv2v_reg  <= data_i[18];
    end 
    if(N5708) begin
      \nz.mem_2457_sv2v_reg  <= data_i[17];
    end 
    if(N5707) begin
      \nz.mem_2456_sv2v_reg  <= data_i[16];
    end 
    if(N5706) begin
      \nz.mem_2455_sv2v_reg  <= data_i[15];
    end 
    if(N5705) begin
      \nz.mem_2454_sv2v_reg  <= data_i[14];
    end 
    if(N5704) begin
      \nz.mem_2453_sv2v_reg  <= data_i[13];
    end 
    if(N5703) begin
      \nz.mem_2452_sv2v_reg  <= data_i[12];
    end 
    if(N5702) begin
      \nz.mem_2451_sv2v_reg  <= data_i[11];
    end 
    if(N5701) begin
      \nz.mem_2450_sv2v_reg  <= data_i[10];
    end 
    if(N5700) begin
      \nz.mem_2449_sv2v_reg  <= data_i[9];
    end 
    if(N5699) begin
      \nz.mem_2448_sv2v_reg  <= data_i[8];
    end 
    if(N5698) begin
      \nz.mem_2447_sv2v_reg  <= data_i[7];
    end 
    if(N5697) begin
      \nz.mem_2446_sv2v_reg  <= data_i[6];
    end 
    if(N5696) begin
      \nz.mem_2445_sv2v_reg  <= data_i[5];
    end 
    if(N5695) begin
      \nz.mem_2444_sv2v_reg  <= data_i[4];
    end 
    if(N5694) begin
      \nz.mem_2443_sv2v_reg  <= data_i[3];
    end 
    if(N5693) begin
      \nz.mem_2442_sv2v_reg  <= data_i[2];
    end 
    if(N5692) begin
      \nz.mem_2441_sv2v_reg  <= data_i[1];
    end 
    if(N5691) begin
      \nz.mem_2440_sv2v_reg  <= data_i[0];
    end 
    if(N5690) begin
      \nz.mem_2439_sv2v_reg  <= data_i[39];
    end 
    if(N5689) begin
      \nz.mem_2438_sv2v_reg  <= data_i[38];
    end 
    if(N5688) begin
      \nz.mem_2437_sv2v_reg  <= data_i[37];
    end 
    if(N5687) begin
      \nz.mem_2436_sv2v_reg  <= data_i[36];
    end 
    if(N5686) begin
      \nz.mem_2435_sv2v_reg  <= data_i[35];
    end 
    if(N5685) begin
      \nz.mem_2434_sv2v_reg  <= data_i[34];
    end 
    if(N5684) begin
      \nz.mem_2433_sv2v_reg  <= data_i[33];
    end 
    if(N5683) begin
      \nz.mem_2432_sv2v_reg  <= data_i[32];
    end 
    if(N5682) begin
      \nz.mem_2431_sv2v_reg  <= data_i[31];
    end 
    if(N5681) begin
      \nz.mem_2430_sv2v_reg  <= data_i[30];
    end 
    if(N5680) begin
      \nz.mem_2429_sv2v_reg  <= data_i[29];
    end 
    if(N5679) begin
      \nz.mem_2428_sv2v_reg  <= data_i[28];
    end 
    if(N5678) begin
      \nz.mem_2427_sv2v_reg  <= data_i[27];
    end 
    if(N5677) begin
      \nz.mem_2426_sv2v_reg  <= data_i[26];
    end 
    if(N5676) begin
      \nz.mem_2425_sv2v_reg  <= data_i[25];
    end 
    if(N5675) begin
      \nz.mem_2424_sv2v_reg  <= data_i[24];
    end 
    if(N5674) begin
      \nz.mem_2423_sv2v_reg  <= data_i[23];
    end 
    if(N5673) begin
      \nz.mem_2422_sv2v_reg  <= data_i[22];
    end 
    if(N5672) begin
      \nz.mem_2421_sv2v_reg  <= data_i[21];
    end 
    if(N5671) begin
      \nz.mem_2420_sv2v_reg  <= data_i[20];
    end 
    if(N5670) begin
      \nz.mem_2419_sv2v_reg  <= data_i[19];
    end 
    if(N5669) begin
      \nz.mem_2418_sv2v_reg  <= data_i[18];
    end 
    if(N5668) begin
      \nz.mem_2417_sv2v_reg  <= data_i[17];
    end 
    if(N5667) begin
      \nz.mem_2416_sv2v_reg  <= data_i[16];
    end 
    if(N5666) begin
      \nz.mem_2415_sv2v_reg  <= data_i[15];
    end 
    if(N5665) begin
      \nz.mem_2414_sv2v_reg  <= data_i[14];
    end 
    if(N5664) begin
      \nz.mem_2413_sv2v_reg  <= data_i[13];
    end 
    if(N5663) begin
      \nz.mem_2412_sv2v_reg  <= data_i[12];
    end 
    if(N5662) begin
      \nz.mem_2411_sv2v_reg  <= data_i[11];
    end 
    if(N5661) begin
      \nz.mem_2410_sv2v_reg  <= data_i[10];
    end 
    if(N5660) begin
      \nz.mem_2409_sv2v_reg  <= data_i[9];
    end 
    if(N5659) begin
      \nz.mem_2408_sv2v_reg  <= data_i[8];
    end 
    if(N5658) begin
      \nz.mem_2407_sv2v_reg  <= data_i[7];
    end 
    if(N5657) begin
      \nz.mem_2406_sv2v_reg  <= data_i[6];
    end 
    if(N5656) begin
      \nz.mem_2405_sv2v_reg  <= data_i[5];
    end 
    if(N5655) begin
      \nz.mem_2404_sv2v_reg  <= data_i[4];
    end 
    if(N5654) begin
      \nz.mem_2403_sv2v_reg  <= data_i[3];
    end 
    if(N5653) begin
      \nz.mem_2402_sv2v_reg  <= data_i[2];
    end 
    if(N5652) begin
      \nz.mem_2401_sv2v_reg  <= data_i[1];
    end 
    if(N5651) begin
      \nz.mem_2400_sv2v_reg  <= data_i[0];
    end 
    if(N5650) begin
      \nz.mem_2399_sv2v_reg  <= data_i[39];
    end 
    if(N5649) begin
      \nz.mem_2398_sv2v_reg  <= data_i[38];
    end 
    if(N5648) begin
      \nz.mem_2397_sv2v_reg  <= data_i[37];
    end 
    if(N5647) begin
      \nz.mem_2396_sv2v_reg  <= data_i[36];
    end 
    if(N5646) begin
      \nz.mem_2395_sv2v_reg  <= data_i[35];
    end 
    if(N5645) begin
      \nz.mem_2394_sv2v_reg  <= data_i[34];
    end 
    if(N5644) begin
      \nz.mem_2393_sv2v_reg  <= data_i[33];
    end 
    if(N5643) begin
      \nz.mem_2392_sv2v_reg  <= data_i[32];
    end 
    if(N5642) begin
      \nz.mem_2391_sv2v_reg  <= data_i[31];
    end 
    if(N5641) begin
      \nz.mem_2390_sv2v_reg  <= data_i[30];
    end 
    if(N5640) begin
      \nz.mem_2389_sv2v_reg  <= data_i[29];
    end 
    if(N5639) begin
      \nz.mem_2388_sv2v_reg  <= data_i[28];
    end 
    if(N5638) begin
      \nz.mem_2387_sv2v_reg  <= data_i[27];
    end 
    if(N5637) begin
      \nz.mem_2386_sv2v_reg  <= data_i[26];
    end 
    if(N5636) begin
      \nz.mem_2385_sv2v_reg  <= data_i[25];
    end 
    if(N5635) begin
      \nz.mem_2384_sv2v_reg  <= data_i[24];
    end 
    if(N5634) begin
      \nz.mem_2383_sv2v_reg  <= data_i[23];
    end 
    if(N5633) begin
      \nz.mem_2382_sv2v_reg  <= data_i[22];
    end 
    if(N5632) begin
      \nz.mem_2381_sv2v_reg  <= data_i[21];
    end 
    if(N5631) begin
      \nz.mem_2380_sv2v_reg  <= data_i[20];
    end 
    if(N5630) begin
      \nz.mem_2379_sv2v_reg  <= data_i[19];
    end 
    if(N5629) begin
      \nz.mem_2378_sv2v_reg  <= data_i[18];
    end 
    if(N5628) begin
      \nz.mem_2377_sv2v_reg  <= data_i[17];
    end 
    if(N5627) begin
      \nz.mem_2376_sv2v_reg  <= data_i[16];
    end 
    if(N5626) begin
      \nz.mem_2375_sv2v_reg  <= data_i[15];
    end 
    if(N5625) begin
      \nz.mem_2374_sv2v_reg  <= data_i[14];
    end 
    if(N5624) begin
      \nz.mem_2373_sv2v_reg  <= data_i[13];
    end 
    if(N5623) begin
      \nz.mem_2372_sv2v_reg  <= data_i[12];
    end 
    if(N5622) begin
      \nz.mem_2371_sv2v_reg  <= data_i[11];
    end 
    if(N5621) begin
      \nz.mem_2370_sv2v_reg  <= data_i[10];
    end 
    if(N5620) begin
      \nz.mem_2369_sv2v_reg  <= data_i[9];
    end 
    if(N5619) begin
      \nz.mem_2368_sv2v_reg  <= data_i[8];
    end 
    if(N5618) begin
      \nz.mem_2367_sv2v_reg  <= data_i[7];
    end 
    if(N5617) begin
      \nz.mem_2366_sv2v_reg  <= data_i[6];
    end 
    if(N5616) begin
      \nz.mem_2365_sv2v_reg  <= data_i[5];
    end 
    if(N5615) begin
      \nz.mem_2364_sv2v_reg  <= data_i[4];
    end 
    if(N5614) begin
      \nz.mem_2363_sv2v_reg  <= data_i[3];
    end 
    if(N5613) begin
      \nz.mem_2362_sv2v_reg  <= data_i[2];
    end 
    if(N5612) begin
      \nz.mem_2361_sv2v_reg  <= data_i[1];
    end 
    if(N5611) begin
      \nz.mem_2360_sv2v_reg  <= data_i[0];
    end 
    if(N5610) begin
      \nz.mem_2359_sv2v_reg  <= data_i[39];
    end 
    if(N5609) begin
      \nz.mem_2358_sv2v_reg  <= data_i[38];
    end 
    if(N5608) begin
      \nz.mem_2357_sv2v_reg  <= data_i[37];
    end 
    if(N5607) begin
      \nz.mem_2356_sv2v_reg  <= data_i[36];
    end 
    if(N5606) begin
      \nz.mem_2355_sv2v_reg  <= data_i[35];
    end 
    if(N5605) begin
      \nz.mem_2354_sv2v_reg  <= data_i[34];
    end 
    if(N5604) begin
      \nz.mem_2353_sv2v_reg  <= data_i[33];
    end 
    if(N5603) begin
      \nz.mem_2352_sv2v_reg  <= data_i[32];
    end 
    if(N5602) begin
      \nz.mem_2351_sv2v_reg  <= data_i[31];
    end 
    if(N5601) begin
      \nz.mem_2350_sv2v_reg  <= data_i[30];
    end 
    if(N5600) begin
      \nz.mem_2349_sv2v_reg  <= data_i[29];
    end 
    if(N5599) begin
      \nz.mem_2348_sv2v_reg  <= data_i[28];
    end 
    if(N5598) begin
      \nz.mem_2347_sv2v_reg  <= data_i[27];
    end 
    if(N5597) begin
      \nz.mem_2346_sv2v_reg  <= data_i[26];
    end 
    if(N5596) begin
      \nz.mem_2345_sv2v_reg  <= data_i[25];
    end 
    if(N5595) begin
      \nz.mem_2344_sv2v_reg  <= data_i[24];
    end 
    if(N5594) begin
      \nz.mem_2343_sv2v_reg  <= data_i[23];
    end 
    if(N5593) begin
      \nz.mem_2342_sv2v_reg  <= data_i[22];
    end 
    if(N5592) begin
      \nz.mem_2341_sv2v_reg  <= data_i[21];
    end 
    if(N5591) begin
      \nz.mem_2340_sv2v_reg  <= data_i[20];
    end 
    if(N5590) begin
      \nz.mem_2339_sv2v_reg  <= data_i[19];
    end 
    if(N5589) begin
      \nz.mem_2338_sv2v_reg  <= data_i[18];
    end 
    if(N5588) begin
      \nz.mem_2337_sv2v_reg  <= data_i[17];
    end 
    if(N5587) begin
      \nz.mem_2336_sv2v_reg  <= data_i[16];
    end 
    if(N5586) begin
      \nz.mem_2335_sv2v_reg  <= data_i[15];
    end 
    if(N5585) begin
      \nz.mem_2334_sv2v_reg  <= data_i[14];
    end 
    if(N5584) begin
      \nz.mem_2333_sv2v_reg  <= data_i[13];
    end 
    if(N5583) begin
      \nz.mem_2332_sv2v_reg  <= data_i[12];
    end 
    if(N5582) begin
      \nz.mem_2331_sv2v_reg  <= data_i[11];
    end 
    if(N5581) begin
      \nz.mem_2330_sv2v_reg  <= data_i[10];
    end 
    if(N5580) begin
      \nz.mem_2329_sv2v_reg  <= data_i[9];
    end 
    if(N5579) begin
      \nz.mem_2328_sv2v_reg  <= data_i[8];
    end 
    if(N5578) begin
      \nz.mem_2327_sv2v_reg  <= data_i[7];
    end 
    if(N5577) begin
      \nz.mem_2326_sv2v_reg  <= data_i[6];
    end 
    if(N5576) begin
      \nz.mem_2325_sv2v_reg  <= data_i[5];
    end 
    if(N5575) begin
      \nz.mem_2324_sv2v_reg  <= data_i[4];
    end 
    if(N5574) begin
      \nz.mem_2323_sv2v_reg  <= data_i[3];
    end 
    if(N5573) begin
      \nz.mem_2322_sv2v_reg  <= data_i[2];
    end 
    if(N5572) begin
      \nz.mem_2321_sv2v_reg  <= data_i[1];
    end 
    if(N5571) begin
      \nz.mem_2320_sv2v_reg  <= data_i[0];
    end 
    if(N5570) begin
      \nz.mem_2319_sv2v_reg  <= data_i[39];
    end 
    if(N5569) begin
      \nz.mem_2318_sv2v_reg  <= data_i[38];
    end 
    if(N5568) begin
      \nz.mem_2317_sv2v_reg  <= data_i[37];
    end 
    if(N5567) begin
      \nz.mem_2316_sv2v_reg  <= data_i[36];
    end 
    if(N5566) begin
      \nz.mem_2315_sv2v_reg  <= data_i[35];
    end 
    if(N5565) begin
      \nz.mem_2314_sv2v_reg  <= data_i[34];
    end 
    if(N5564) begin
      \nz.mem_2313_sv2v_reg  <= data_i[33];
    end 
    if(N5563) begin
      \nz.mem_2312_sv2v_reg  <= data_i[32];
    end 
    if(N5562) begin
      \nz.mem_2311_sv2v_reg  <= data_i[31];
    end 
    if(N5561) begin
      \nz.mem_2310_sv2v_reg  <= data_i[30];
    end 
    if(N5560) begin
      \nz.mem_2309_sv2v_reg  <= data_i[29];
    end 
    if(N5559) begin
      \nz.mem_2308_sv2v_reg  <= data_i[28];
    end 
    if(N5558) begin
      \nz.mem_2307_sv2v_reg  <= data_i[27];
    end 
    if(N5557) begin
      \nz.mem_2306_sv2v_reg  <= data_i[26];
    end 
    if(N5556) begin
      \nz.mem_2305_sv2v_reg  <= data_i[25];
    end 
    if(N5555) begin
      \nz.mem_2304_sv2v_reg  <= data_i[24];
    end 
    if(N5554) begin
      \nz.mem_2303_sv2v_reg  <= data_i[23];
    end 
    if(N5553) begin
      \nz.mem_2302_sv2v_reg  <= data_i[22];
    end 
    if(N5552) begin
      \nz.mem_2301_sv2v_reg  <= data_i[21];
    end 
    if(N5551) begin
      \nz.mem_2300_sv2v_reg  <= data_i[20];
    end 
    if(N5550) begin
      \nz.mem_2299_sv2v_reg  <= data_i[19];
    end 
    if(N5549) begin
      \nz.mem_2298_sv2v_reg  <= data_i[18];
    end 
    if(N5548) begin
      \nz.mem_2297_sv2v_reg  <= data_i[17];
    end 
    if(N5547) begin
      \nz.mem_2296_sv2v_reg  <= data_i[16];
    end 
    if(N5546) begin
      \nz.mem_2295_sv2v_reg  <= data_i[15];
    end 
    if(N5545) begin
      \nz.mem_2294_sv2v_reg  <= data_i[14];
    end 
    if(N5544) begin
      \nz.mem_2293_sv2v_reg  <= data_i[13];
    end 
    if(N5543) begin
      \nz.mem_2292_sv2v_reg  <= data_i[12];
    end 
    if(N5542) begin
      \nz.mem_2291_sv2v_reg  <= data_i[11];
    end 
    if(N5541) begin
      \nz.mem_2290_sv2v_reg  <= data_i[10];
    end 
    if(N5540) begin
      \nz.mem_2289_sv2v_reg  <= data_i[9];
    end 
    if(N5539) begin
      \nz.mem_2288_sv2v_reg  <= data_i[8];
    end 
    if(N5538) begin
      \nz.mem_2287_sv2v_reg  <= data_i[7];
    end 
    if(N5537) begin
      \nz.mem_2286_sv2v_reg  <= data_i[6];
    end 
    if(N5536) begin
      \nz.mem_2285_sv2v_reg  <= data_i[5];
    end 
    if(N5535) begin
      \nz.mem_2284_sv2v_reg  <= data_i[4];
    end 
    if(N5534) begin
      \nz.mem_2283_sv2v_reg  <= data_i[3];
    end 
    if(N5533) begin
      \nz.mem_2282_sv2v_reg  <= data_i[2];
    end 
    if(N5532) begin
      \nz.mem_2281_sv2v_reg  <= data_i[1];
    end 
    if(N5531) begin
      \nz.mem_2280_sv2v_reg  <= data_i[0];
    end 
    if(N5530) begin
      \nz.mem_2279_sv2v_reg  <= data_i[39];
    end 
    if(N5529) begin
      \nz.mem_2278_sv2v_reg  <= data_i[38];
    end 
    if(N5528) begin
      \nz.mem_2277_sv2v_reg  <= data_i[37];
    end 
    if(N5527) begin
      \nz.mem_2276_sv2v_reg  <= data_i[36];
    end 
    if(N5526) begin
      \nz.mem_2275_sv2v_reg  <= data_i[35];
    end 
    if(N5525) begin
      \nz.mem_2274_sv2v_reg  <= data_i[34];
    end 
    if(N5524) begin
      \nz.mem_2273_sv2v_reg  <= data_i[33];
    end 
    if(N5523) begin
      \nz.mem_2272_sv2v_reg  <= data_i[32];
    end 
    if(N5522) begin
      \nz.mem_2271_sv2v_reg  <= data_i[31];
    end 
    if(N5521) begin
      \nz.mem_2270_sv2v_reg  <= data_i[30];
    end 
    if(N5520) begin
      \nz.mem_2269_sv2v_reg  <= data_i[29];
    end 
    if(N5519) begin
      \nz.mem_2268_sv2v_reg  <= data_i[28];
    end 
    if(N5518) begin
      \nz.mem_2267_sv2v_reg  <= data_i[27];
    end 
    if(N5517) begin
      \nz.mem_2266_sv2v_reg  <= data_i[26];
    end 
    if(N5516) begin
      \nz.mem_2265_sv2v_reg  <= data_i[25];
    end 
    if(N5515) begin
      \nz.mem_2264_sv2v_reg  <= data_i[24];
    end 
    if(N5514) begin
      \nz.mem_2263_sv2v_reg  <= data_i[23];
    end 
    if(N5513) begin
      \nz.mem_2262_sv2v_reg  <= data_i[22];
    end 
    if(N5512) begin
      \nz.mem_2261_sv2v_reg  <= data_i[21];
    end 
    if(N5511) begin
      \nz.mem_2260_sv2v_reg  <= data_i[20];
    end 
    if(N5510) begin
      \nz.mem_2259_sv2v_reg  <= data_i[19];
    end 
    if(N5509) begin
      \nz.mem_2258_sv2v_reg  <= data_i[18];
    end 
    if(N5508) begin
      \nz.mem_2257_sv2v_reg  <= data_i[17];
    end 
    if(N5507) begin
      \nz.mem_2256_sv2v_reg  <= data_i[16];
    end 
    if(N5506) begin
      \nz.mem_2255_sv2v_reg  <= data_i[15];
    end 
    if(N5505) begin
      \nz.mem_2254_sv2v_reg  <= data_i[14];
    end 
    if(N5504) begin
      \nz.mem_2253_sv2v_reg  <= data_i[13];
    end 
    if(N5503) begin
      \nz.mem_2252_sv2v_reg  <= data_i[12];
    end 
    if(N5502) begin
      \nz.mem_2251_sv2v_reg  <= data_i[11];
    end 
    if(N5501) begin
      \nz.mem_2250_sv2v_reg  <= data_i[10];
    end 
    if(N5500) begin
      \nz.mem_2249_sv2v_reg  <= data_i[9];
    end 
    if(N5499) begin
      \nz.mem_2248_sv2v_reg  <= data_i[8];
    end 
    if(N5498) begin
      \nz.mem_2247_sv2v_reg  <= data_i[7];
    end 
    if(N5497) begin
      \nz.mem_2246_sv2v_reg  <= data_i[6];
    end 
    if(N5496) begin
      \nz.mem_2245_sv2v_reg  <= data_i[5];
    end 
    if(N5495) begin
      \nz.mem_2244_sv2v_reg  <= data_i[4];
    end 
    if(N5494) begin
      \nz.mem_2243_sv2v_reg  <= data_i[3];
    end 
    if(N5493) begin
      \nz.mem_2242_sv2v_reg  <= data_i[2];
    end 
    if(N5492) begin
      \nz.mem_2241_sv2v_reg  <= data_i[1];
    end 
    if(N5491) begin
      \nz.mem_2240_sv2v_reg  <= data_i[0];
    end 
    if(N5490) begin
      \nz.mem_2239_sv2v_reg  <= data_i[39];
    end 
    if(N5489) begin
      \nz.mem_2238_sv2v_reg  <= data_i[38];
    end 
    if(N5488) begin
      \nz.mem_2237_sv2v_reg  <= data_i[37];
    end 
    if(N5487) begin
      \nz.mem_2236_sv2v_reg  <= data_i[36];
    end 
    if(N5486) begin
      \nz.mem_2235_sv2v_reg  <= data_i[35];
    end 
    if(N5485) begin
      \nz.mem_2234_sv2v_reg  <= data_i[34];
    end 
    if(N5484) begin
      \nz.mem_2233_sv2v_reg  <= data_i[33];
    end 
    if(N5483) begin
      \nz.mem_2232_sv2v_reg  <= data_i[32];
    end 
    if(N5482) begin
      \nz.mem_2231_sv2v_reg  <= data_i[31];
    end 
    if(N5481) begin
      \nz.mem_2230_sv2v_reg  <= data_i[30];
    end 
    if(N5480) begin
      \nz.mem_2229_sv2v_reg  <= data_i[29];
    end 
    if(N5479) begin
      \nz.mem_2228_sv2v_reg  <= data_i[28];
    end 
    if(N5478) begin
      \nz.mem_2227_sv2v_reg  <= data_i[27];
    end 
    if(N5477) begin
      \nz.mem_2226_sv2v_reg  <= data_i[26];
    end 
    if(N5476) begin
      \nz.mem_2225_sv2v_reg  <= data_i[25];
    end 
    if(N5475) begin
      \nz.mem_2224_sv2v_reg  <= data_i[24];
    end 
    if(N5474) begin
      \nz.mem_2223_sv2v_reg  <= data_i[23];
    end 
    if(N5473) begin
      \nz.mem_2222_sv2v_reg  <= data_i[22];
    end 
    if(N5472) begin
      \nz.mem_2221_sv2v_reg  <= data_i[21];
    end 
    if(N5471) begin
      \nz.mem_2220_sv2v_reg  <= data_i[20];
    end 
    if(N5470) begin
      \nz.mem_2219_sv2v_reg  <= data_i[19];
    end 
    if(N5469) begin
      \nz.mem_2218_sv2v_reg  <= data_i[18];
    end 
    if(N5468) begin
      \nz.mem_2217_sv2v_reg  <= data_i[17];
    end 
    if(N5467) begin
      \nz.mem_2216_sv2v_reg  <= data_i[16];
    end 
    if(N5466) begin
      \nz.mem_2215_sv2v_reg  <= data_i[15];
    end 
    if(N5465) begin
      \nz.mem_2214_sv2v_reg  <= data_i[14];
    end 
    if(N5464) begin
      \nz.mem_2213_sv2v_reg  <= data_i[13];
    end 
    if(N5463) begin
      \nz.mem_2212_sv2v_reg  <= data_i[12];
    end 
    if(N5462) begin
      \nz.mem_2211_sv2v_reg  <= data_i[11];
    end 
    if(N5461) begin
      \nz.mem_2210_sv2v_reg  <= data_i[10];
    end 
    if(N5460) begin
      \nz.mem_2209_sv2v_reg  <= data_i[9];
    end 
    if(N5459) begin
      \nz.mem_2208_sv2v_reg  <= data_i[8];
    end 
    if(N5458) begin
      \nz.mem_2207_sv2v_reg  <= data_i[7];
    end 
    if(N5457) begin
      \nz.mem_2206_sv2v_reg  <= data_i[6];
    end 
    if(N5456) begin
      \nz.mem_2205_sv2v_reg  <= data_i[5];
    end 
    if(N5455) begin
      \nz.mem_2204_sv2v_reg  <= data_i[4];
    end 
    if(N5454) begin
      \nz.mem_2203_sv2v_reg  <= data_i[3];
    end 
    if(N5453) begin
      \nz.mem_2202_sv2v_reg  <= data_i[2];
    end 
    if(N5452) begin
      \nz.mem_2201_sv2v_reg  <= data_i[1];
    end 
    if(N5451) begin
      \nz.mem_2200_sv2v_reg  <= data_i[0];
    end 
    if(N5450) begin
      \nz.mem_2199_sv2v_reg  <= data_i[39];
    end 
    if(N5449) begin
      \nz.mem_2198_sv2v_reg  <= data_i[38];
    end 
    if(N5448) begin
      \nz.mem_2197_sv2v_reg  <= data_i[37];
    end 
    if(N5447) begin
      \nz.mem_2196_sv2v_reg  <= data_i[36];
    end 
    if(N5446) begin
      \nz.mem_2195_sv2v_reg  <= data_i[35];
    end 
    if(N5445) begin
      \nz.mem_2194_sv2v_reg  <= data_i[34];
    end 
    if(N5444) begin
      \nz.mem_2193_sv2v_reg  <= data_i[33];
    end 
    if(N5443) begin
      \nz.mem_2192_sv2v_reg  <= data_i[32];
    end 
    if(N5442) begin
      \nz.mem_2191_sv2v_reg  <= data_i[31];
    end 
    if(N5441) begin
      \nz.mem_2190_sv2v_reg  <= data_i[30];
    end 
    if(N5440) begin
      \nz.mem_2189_sv2v_reg  <= data_i[29];
    end 
    if(N5439) begin
      \nz.mem_2188_sv2v_reg  <= data_i[28];
    end 
    if(N5438) begin
      \nz.mem_2187_sv2v_reg  <= data_i[27];
    end 
    if(N5437) begin
      \nz.mem_2186_sv2v_reg  <= data_i[26];
    end 
    if(N5436) begin
      \nz.mem_2185_sv2v_reg  <= data_i[25];
    end 
    if(N5435) begin
      \nz.mem_2184_sv2v_reg  <= data_i[24];
    end 
    if(N5434) begin
      \nz.mem_2183_sv2v_reg  <= data_i[23];
    end 
    if(N5433) begin
      \nz.mem_2182_sv2v_reg  <= data_i[22];
    end 
    if(N5432) begin
      \nz.mem_2181_sv2v_reg  <= data_i[21];
    end 
    if(N5431) begin
      \nz.mem_2180_sv2v_reg  <= data_i[20];
    end 
    if(N5430) begin
      \nz.mem_2179_sv2v_reg  <= data_i[19];
    end 
    if(N5429) begin
      \nz.mem_2178_sv2v_reg  <= data_i[18];
    end 
    if(N5428) begin
      \nz.mem_2177_sv2v_reg  <= data_i[17];
    end 
    if(N5427) begin
      \nz.mem_2176_sv2v_reg  <= data_i[16];
    end 
    if(N5426) begin
      \nz.mem_2175_sv2v_reg  <= data_i[15];
    end 
    if(N5425) begin
      \nz.mem_2174_sv2v_reg  <= data_i[14];
    end 
    if(N5424) begin
      \nz.mem_2173_sv2v_reg  <= data_i[13];
    end 
    if(N5423) begin
      \nz.mem_2172_sv2v_reg  <= data_i[12];
    end 
    if(N5422) begin
      \nz.mem_2171_sv2v_reg  <= data_i[11];
    end 
    if(N5421) begin
      \nz.mem_2170_sv2v_reg  <= data_i[10];
    end 
    if(N5420) begin
      \nz.mem_2169_sv2v_reg  <= data_i[9];
    end 
    if(N5419) begin
      \nz.mem_2168_sv2v_reg  <= data_i[8];
    end 
    if(N5418) begin
      \nz.mem_2167_sv2v_reg  <= data_i[7];
    end 
    if(N5417) begin
      \nz.mem_2166_sv2v_reg  <= data_i[6];
    end 
    if(N5416) begin
      \nz.mem_2165_sv2v_reg  <= data_i[5];
    end 
    if(N5415) begin
      \nz.mem_2164_sv2v_reg  <= data_i[4];
    end 
    if(N5414) begin
      \nz.mem_2163_sv2v_reg  <= data_i[3];
    end 
    if(N5413) begin
      \nz.mem_2162_sv2v_reg  <= data_i[2];
    end 
    if(N5412) begin
      \nz.mem_2161_sv2v_reg  <= data_i[1];
    end 
    if(N5411) begin
      \nz.mem_2160_sv2v_reg  <= data_i[0];
    end 
    if(N5410) begin
      \nz.mem_2159_sv2v_reg  <= data_i[39];
    end 
    if(N5409) begin
      \nz.mem_2158_sv2v_reg  <= data_i[38];
    end 
    if(N5408) begin
      \nz.mem_2157_sv2v_reg  <= data_i[37];
    end 
    if(N5407) begin
      \nz.mem_2156_sv2v_reg  <= data_i[36];
    end 
    if(N5406) begin
      \nz.mem_2155_sv2v_reg  <= data_i[35];
    end 
    if(N5405) begin
      \nz.mem_2154_sv2v_reg  <= data_i[34];
    end 
    if(N5404) begin
      \nz.mem_2153_sv2v_reg  <= data_i[33];
    end 
    if(N5403) begin
      \nz.mem_2152_sv2v_reg  <= data_i[32];
    end 
    if(N5402) begin
      \nz.mem_2151_sv2v_reg  <= data_i[31];
    end 
    if(N5401) begin
      \nz.mem_2150_sv2v_reg  <= data_i[30];
    end 
    if(N5400) begin
      \nz.mem_2149_sv2v_reg  <= data_i[29];
    end 
    if(N5399) begin
      \nz.mem_2148_sv2v_reg  <= data_i[28];
    end 
    if(N5398) begin
      \nz.mem_2147_sv2v_reg  <= data_i[27];
    end 
    if(N5397) begin
      \nz.mem_2146_sv2v_reg  <= data_i[26];
    end 
    if(N5396) begin
      \nz.mem_2145_sv2v_reg  <= data_i[25];
    end 
    if(N5395) begin
      \nz.mem_2144_sv2v_reg  <= data_i[24];
    end 
    if(N5394) begin
      \nz.mem_2143_sv2v_reg  <= data_i[23];
    end 
    if(N5393) begin
      \nz.mem_2142_sv2v_reg  <= data_i[22];
    end 
    if(N5392) begin
      \nz.mem_2141_sv2v_reg  <= data_i[21];
    end 
    if(N5391) begin
      \nz.mem_2140_sv2v_reg  <= data_i[20];
    end 
    if(N5390) begin
      \nz.mem_2139_sv2v_reg  <= data_i[19];
    end 
    if(N5389) begin
      \nz.mem_2138_sv2v_reg  <= data_i[18];
    end 
    if(N5388) begin
      \nz.mem_2137_sv2v_reg  <= data_i[17];
    end 
    if(N5387) begin
      \nz.mem_2136_sv2v_reg  <= data_i[16];
    end 
    if(N5386) begin
      \nz.mem_2135_sv2v_reg  <= data_i[15];
    end 
    if(N5385) begin
      \nz.mem_2134_sv2v_reg  <= data_i[14];
    end 
    if(N5384) begin
      \nz.mem_2133_sv2v_reg  <= data_i[13];
    end 
    if(N5383) begin
      \nz.mem_2132_sv2v_reg  <= data_i[12];
    end 
    if(N5382) begin
      \nz.mem_2131_sv2v_reg  <= data_i[11];
    end 
    if(N5381) begin
      \nz.mem_2130_sv2v_reg  <= data_i[10];
    end 
    if(N5380) begin
      \nz.mem_2129_sv2v_reg  <= data_i[9];
    end 
    if(N5379) begin
      \nz.mem_2128_sv2v_reg  <= data_i[8];
    end 
    if(N5378) begin
      \nz.mem_2127_sv2v_reg  <= data_i[7];
    end 
    if(N5377) begin
      \nz.mem_2126_sv2v_reg  <= data_i[6];
    end 
    if(N5376) begin
      \nz.mem_2125_sv2v_reg  <= data_i[5];
    end 
    if(N5375) begin
      \nz.mem_2124_sv2v_reg  <= data_i[4];
    end 
    if(N5374) begin
      \nz.mem_2123_sv2v_reg  <= data_i[3];
    end 
    if(N5373) begin
      \nz.mem_2122_sv2v_reg  <= data_i[2];
    end 
    if(N5372) begin
      \nz.mem_2121_sv2v_reg  <= data_i[1];
    end 
    if(N5371) begin
      \nz.mem_2120_sv2v_reg  <= data_i[0];
    end 
    if(N5370) begin
      \nz.mem_2119_sv2v_reg  <= data_i[39];
    end 
    if(N5369) begin
      \nz.mem_2118_sv2v_reg  <= data_i[38];
    end 
    if(N5368) begin
      \nz.mem_2117_sv2v_reg  <= data_i[37];
    end 
    if(N5367) begin
      \nz.mem_2116_sv2v_reg  <= data_i[36];
    end 
    if(N5366) begin
      \nz.mem_2115_sv2v_reg  <= data_i[35];
    end 
    if(N5365) begin
      \nz.mem_2114_sv2v_reg  <= data_i[34];
    end 
    if(N5364) begin
      \nz.mem_2113_sv2v_reg  <= data_i[33];
    end 
    if(N5363) begin
      \nz.mem_2112_sv2v_reg  <= data_i[32];
    end 
    if(N5362) begin
      \nz.mem_2111_sv2v_reg  <= data_i[31];
    end 
    if(N5361) begin
      \nz.mem_2110_sv2v_reg  <= data_i[30];
    end 
    if(N5360) begin
      \nz.mem_2109_sv2v_reg  <= data_i[29];
    end 
    if(N5359) begin
      \nz.mem_2108_sv2v_reg  <= data_i[28];
    end 
    if(N5358) begin
      \nz.mem_2107_sv2v_reg  <= data_i[27];
    end 
    if(N5357) begin
      \nz.mem_2106_sv2v_reg  <= data_i[26];
    end 
    if(N5356) begin
      \nz.mem_2105_sv2v_reg  <= data_i[25];
    end 
    if(N5355) begin
      \nz.mem_2104_sv2v_reg  <= data_i[24];
    end 
    if(N5354) begin
      \nz.mem_2103_sv2v_reg  <= data_i[23];
    end 
    if(N5353) begin
      \nz.mem_2102_sv2v_reg  <= data_i[22];
    end 
    if(N5352) begin
      \nz.mem_2101_sv2v_reg  <= data_i[21];
    end 
    if(N5351) begin
      \nz.mem_2100_sv2v_reg  <= data_i[20];
    end 
    if(N5350) begin
      \nz.mem_2099_sv2v_reg  <= data_i[19];
    end 
    if(N5349) begin
      \nz.mem_2098_sv2v_reg  <= data_i[18];
    end 
    if(N5348) begin
      \nz.mem_2097_sv2v_reg  <= data_i[17];
    end 
    if(N5347) begin
      \nz.mem_2096_sv2v_reg  <= data_i[16];
    end 
    if(N5346) begin
      \nz.mem_2095_sv2v_reg  <= data_i[15];
    end 
    if(N5345) begin
      \nz.mem_2094_sv2v_reg  <= data_i[14];
    end 
    if(N5344) begin
      \nz.mem_2093_sv2v_reg  <= data_i[13];
    end 
    if(N5343) begin
      \nz.mem_2092_sv2v_reg  <= data_i[12];
    end 
    if(N5342) begin
      \nz.mem_2091_sv2v_reg  <= data_i[11];
    end 
    if(N5341) begin
      \nz.mem_2090_sv2v_reg  <= data_i[10];
    end 
    if(N5340) begin
      \nz.mem_2089_sv2v_reg  <= data_i[9];
    end 
    if(N5339) begin
      \nz.mem_2088_sv2v_reg  <= data_i[8];
    end 
    if(N5338) begin
      \nz.mem_2087_sv2v_reg  <= data_i[7];
    end 
    if(N5337) begin
      \nz.mem_2086_sv2v_reg  <= data_i[6];
    end 
    if(N5336) begin
      \nz.mem_2085_sv2v_reg  <= data_i[5];
    end 
    if(N5335) begin
      \nz.mem_2084_sv2v_reg  <= data_i[4];
    end 
    if(N5334) begin
      \nz.mem_2083_sv2v_reg  <= data_i[3];
    end 
    if(N5333) begin
      \nz.mem_2082_sv2v_reg  <= data_i[2];
    end 
    if(N5332) begin
      \nz.mem_2081_sv2v_reg  <= data_i[1];
    end 
    if(N5331) begin
      \nz.mem_2080_sv2v_reg  <= data_i[0];
    end 
    if(N5330) begin
      \nz.mem_2079_sv2v_reg  <= data_i[39];
    end 
    if(N5329) begin
      \nz.mem_2078_sv2v_reg  <= data_i[38];
    end 
    if(N5328) begin
      \nz.mem_2077_sv2v_reg  <= data_i[37];
    end 
    if(N5327) begin
      \nz.mem_2076_sv2v_reg  <= data_i[36];
    end 
    if(N5326) begin
      \nz.mem_2075_sv2v_reg  <= data_i[35];
    end 
    if(N5325) begin
      \nz.mem_2074_sv2v_reg  <= data_i[34];
    end 
    if(N5324) begin
      \nz.mem_2073_sv2v_reg  <= data_i[33];
    end 
    if(N5323) begin
      \nz.mem_2072_sv2v_reg  <= data_i[32];
    end 
    if(N5322) begin
      \nz.mem_2071_sv2v_reg  <= data_i[31];
    end 
    if(N5321) begin
      \nz.mem_2070_sv2v_reg  <= data_i[30];
    end 
    if(N5320) begin
      \nz.mem_2069_sv2v_reg  <= data_i[29];
    end 
    if(N5319) begin
      \nz.mem_2068_sv2v_reg  <= data_i[28];
    end 
    if(N5318) begin
      \nz.mem_2067_sv2v_reg  <= data_i[27];
    end 
    if(N5317) begin
      \nz.mem_2066_sv2v_reg  <= data_i[26];
    end 
    if(N5316) begin
      \nz.mem_2065_sv2v_reg  <= data_i[25];
    end 
    if(N5315) begin
      \nz.mem_2064_sv2v_reg  <= data_i[24];
    end 
    if(N5314) begin
      \nz.mem_2063_sv2v_reg  <= data_i[23];
    end 
    if(N5313) begin
      \nz.mem_2062_sv2v_reg  <= data_i[22];
    end 
    if(N5312) begin
      \nz.mem_2061_sv2v_reg  <= data_i[21];
    end 
    if(N5311) begin
      \nz.mem_2060_sv2v_reg  <= data_i[20];
    end 
    if(N5310) begin
      \nz.mem_2059_sv2v_reg  <= data_i[19];
    end 
    if(N5309) begin
      \nz.mem_2058_sv2v_reg  <= data_i[18];
    end 
    if(N5308) begin
      \nz.mem_2057_sv2v_reg  <= data_i[17];
    end 
    if(N5307) begin
      \nz.mem_2056_sv2v_reg  <= data_i[16];
    end 
    if(N5306) begin
      \nz.mem_2055_sv2v_reg  <= data_i[15];
    end 
    if(N5305) begin
      \nz.mem_2054_sv2v_reg  <= data_i[14];
    end 
    if(N5304) begin
      \nz.mem_2053_sv2v_reg  <= data_i[13];
    end 
    if(N5303) begin
      \nz.mem_2052_sv2v_reg  <= data_i[12];
    end 
    if(N5302) begin
      \nz.mem_2051_sv2v_reg  <= data_i[11];
    end 
    if(N5301) begin
      \nz.mem_2050_sv2v_reg  <= data_i[10];
    end 
    if(N5300) begin
      \nz.mem_2049_sv2v_reg  <= data_i[9];
    end 
    if(N5299) begin
      \nz.mem_2048_sv2v_reg  <= data_i[8];
    end 
    if(N5298) begin
      \nz.mem_2047_sv2v_reg  <= data_i[7];
    end 
    if(N5297) begin
      \nz.mem_2046_sv2v_reg  <= data_i[6];
    end 
    if(N5296) begin
      \nz.mem_2045_sv2v_reg  <= data_i[5];
    end 
    if(N5295) begin
      \nz.mem_2044_sv2v_reg  <= data_i[4];
    end 
    if(N5294) begin
      \nz.mem_2043_sv2v_reg  <= data_i[3];
    end 
    if(N5293) begin
      \nz.mem_2042_sv2v_reg  <= data_i[2];
    end 
    if(N5292) begin
      \nz.mem_2041_sv2v_reg  <= data_i[1];
    end 
    if(N5291) begin
      \nz.mem_2040_sv2v_reg  <= data_i[0];
    end 
    if(N5290) begin
      \nz.mem_2039_sv2v_reg  <= data_i[39];
    end 
    if(N5289) begin
      \nz.mem_2038_sv2v_reg  <= data_i[38];
    end 
    if(N5288) begin
      \nz.mem_2037_sv2v_reg  <= data_i[37];
    end 
    if(N5287) begin
      \nz.mem_2036_sv2v_reg  <= data_i[36];
    end 
    if(N5286) begin
      \nz.mem_2035_sv2v_reg  <= data_i[35];
    end 
    if(N5285) begin
      \nz.mem_2034_sv2v_reg  <= data_i[34];
    end 
    if(N5284) begin
      \nz.mem_2033_sv2v_reg  <= data_i[33];
    end 
    if(N5283) begin
      \nz.mem_2032_sv2v_reg  <= data_i[32];
    end 
    if(N5282) begin
      \nz.mem_2031_sv2v_reg  <= data_i[31];
    end 
    if(N5281) begin
      \nz.mem_2030_sv2v_reg  <= data_i[30];
    end 
    if(N5280) begin
      \nz.mem_2029_sv2v_reg  <= data_i[29];
    end 
    if(N5279) begin
      \nz.mem_2028_sv2v_reg  <= data_i[28];
    end 
    if(N5278) begin
      \nz.mem_2027_sv2v_reg  <= data_i[27];
    end 
    if(N5277) begin
      \nz.mem_2026_sv2v_reg  <= data_i[26];
    end 
    if(N5276) begin
      \nz.mem_2025_sv2v_reg  <= data_i[25];
    end 
    if(N5275) begin
      \nz.mem_2024_sv2v_reg  <= data_i[24];
    end 
    if(N5274) begin
      \nz.mem_2023_sv2v_reg  <= data_i[23];
    end 
    if(N5273) begin
      \nz.mem_2022_sv2v_reg  <= data_i[22];
    end 
    if(N5272) begin
      \nz.mem_2021_sv2v_reg  <= data_i[21];
    end 
    if(N5271) begin
      \nz.mem_2020_sv2v_reg  <= data_i[20];
    end 
    if(N5270) begin
      \nz.mem_2019_sv2v_reg  <= data_i[19];
    end 
    if(N5269) begin
      \nz.mem_2018_sv2v_reg  <= data_i[18];
    end 
    if(N5268) begin
      \nz.mem_2017_sv2v_reg  <= data_i[17];
    end 
    if(N5267) begin
      \nz.mem_2016_sv2v_reg  <= data_i[16];
    end 
    if(N5266) begin
      \nz.mem_2015_sv2v_reg  <= data_i[15];
    end 
    if(N5265) begin
      \nz.mem_2014_sv2v_reg  <= data_i[14];
    end 
    if(N5264) begin
      \nz.mem_2013_sv2v_reg  <= data_i[13];
    end 
    if(N5263) begin
      \nz.mem_2012_sv2v_reg  <= data_i[12];
    end 
    if(N5262) begin
      \nz.mem_2011_sv2v_reg  <= data_i[11];
    end 
    if(N5261) begin
      \nz.mem_2010_sv2v_reg  <= data_i[10];
    end 
    if(N5260) begin
      \nz.mem_2009_sv2v_reg  <= data_i[9];
    end 
    if(N5259) begin
      \nz.mem_2008_sv2v_reg  <= data_i[8];
    end 
    if(N5258) begin
      \nz.mem_2007_sv2v_reg  <= data_i[7];
    end 
    if(N5257) begin
      \nz.mem_2006_sv2v_reg  <= data_i[6];
    end 
    if(N5256) begin
      \nz.mem_2005_sv2v_reg  <= data_i[5];
    end 
    if(N5255) begin
      \nz.mem_2004_sv2v_reg  <= data_i[4];
    end 
    if(N5254) begin
      \nz.mem_2003_sv2v_reg  <= data_i[3];
    end 
    if(N5253) begin
      \nz.mem_2002_sv2v_reg  <= data_i[2];
    end 
    if(N5252) begin
      \nz.mem_2001_sv2v_reg  <= data_i[1];
    end 
    if(N5251) begin
      \nz.mem_2000_sv2v_reg  <= data_i[0];
    end 
    if(N5250) begin
      \nz.mem_1999_sv2v_reg  <= data_i[39];
    end 
    if(N5249) begin
      \nz.mem_1998_sv2v_reg  <= data_i[38];
    end 
    if(N5248) begin
      \nz.mem_1997_sv2v_reg  <= data_i[37];
    end 
    if(N5247) begin
      \nz.mem_1996_sv2v_reg  <= data_i[36];
    end 
    if(N5246) begin
      \nz.mem_1995_sv2v_reg  <= data_i[35];
    end 
    if(N5245) begin
      \nz.mem_1994_sv2v_reg  <= data_i[34];
    end 
    if(N5244) begin
      \nz.mem_1993_sv2v_reg  <= data_i[33];
    end 
    if(N5243) begin
      \nz.mem_1992_sv2v_reg  <= data_i[32];
    end 
    if(N5242) begin
      \nz.mem_1991_sv2v_reg  <= data_i[31];
    end 
    if(N5241) begin
      \nz.mem_1990_sv2v_reg  <= data_i[30];
    end 
    if(N5240) begin
      \nz.mem_1989_sv2v_reg  <= data_i[29];
    end 
    if(N5239) begin
      \nz.mem_1988_sv2v_reg  <= data_i[28];
    end 
    if(N5238) begin
      \nz.mem_1987_sv2v_reg  <= data_i[27];
    end 
    if(N5237) begin
      \nz.mem_1986_sv2v_reg  <= data_i[26];
    end 
    if(N5236) begin
      \nz.mem_1985_sv2v_reg  <= data_i[25];
    end 
    if(N5235) begin
      \nz.mem_1984_sv2v_reg  <= data_i[24];
    end 
    if(N5234) begin
      \nz.mem_1983_sv2v_reg  <= data_i[23];
    end 
    if(N5233) begin
      \nz.mem_1982_sv2v_reg  <= data_i[22];
    end 
    if(N5232) begin
      \nz.mem_1981_sv2v_reg  <= data_i[21];
    end 
    if(N5231) begin
      \nz.mem_1980_sv2v_reg  <= data_i[20];
    end 
    if(N5230) begin
      \nz.mem_1979_sv2v_reg  <= data_i[19];
    end 
    if(N5229) begin
      \nz.mem_1978_sv2v_reg  <= data_i[18];
    end 
    if(N5228) begin
      \nz.mem_1977_sv2v_reg  <= data_i[17];
    end 
    if(N5227) begin
      \nz.mem_1976_sv2v_reg  <= data_i[16];
    end 
    if(N5226) begin
      \nz.mem_1975_sv2v_reg  <= data_i[15];
    end 
    if(N5225) begin
      \nz.mem_1974_sv2v_reg  <= data_i[14];
    end 
    if(N5224) begin
      \nz.mem_1973_sv2v_reg  <= data_i[13];
    end 
    if(N5223) begin
      \nz.mem_1972_sv2v_reg  <= data_i[12];
    end 
    if(N5222) begin
      \nz.mem_1971_sv2v_reg  <= data_i[11];
    end 
    if(N5221) begin
      \nz.mem_1970_sv2v_reg  <= data_i[10];
    end 
    if(N5220) begin
      \nz.mem_1969_sv2v_reg  <= data_i[9];
    end 
    if(N5219) begin
      \nz.mem_1968_sv2v_reg  <= data_i[8];
    end 
    if(N5218) begin
      \nz.mem_1967_sv2v_reg  <= data_i[7];
    end 
    if(N5217) begin
      \nz.mem_1966_sv2v_reg  <= data_i[6];
    end 
    if(N5216) begin
      \nz.mem_1965_sv2v_reg  <= data_i[5];
    end 
    if(N5215) begin
      \nz.mem_1964_sv2v_reg  <= data_i[4];
    end 
    if(N5214) begin
      \nz.mem_1963_sv2v_reg  <= data_i[3];
    end 
    if(N5213) begin
      \nz.mem_1962_sv2v_reg  <= data_i[2];
    end 
    if(N5212) begin
      \nz.mem_1961_sv2v_reg  <= data_i[1];
    end 
    if(N5211) begin
      \nz.mem_1960_sv2v_reg  <= data_i[0];
    end 
    if(N5210) begin
      \nz.mem_1959_sv2v_reg  <= data_i[39];
    end 
    if(N5209) begin
      \nz.mem_1958_sv2v_reg  <= data_i[38];
    end 
    if(N5208) begin
      \nz.mem_1957_sv2v_reg  <= data_i[37];
    end 
    if(N5207) begin
      \nz.mem_1956_sv2v_reg  <= data_i[36];
    end 
    if(N5206) begin
      \nz.mem_1955_sv2v_reg  <= data_i[35];
    end 
    if(N5205) begin
      \nz.mem_1954_sv2v_reg  <= data_i[34];
    end 
    if(N5204) begin
      \nz.mem_1953_sv2v_reg  <= data_i[33];
    end 
    if(N5203) begin
      \nz.mem_1952_sv2v_reg  <= data_i[32];
    end 
    if(N5202) begin
      \nz.mem_1951_sv2v_reg  <= data_i[31];
    end 
    if(N5201) begin
      \nz.mem_1950_sv2v_reg  <= data_i[30];
    end 
    if(N5200) begin
      \nz.mem_1949_sv2v_reg  <= data_i[29];
    end 
    if(N5199) begin
      \nz.mem_1948_sv2v_reg  <= data_i[28];
    end 
    if(N5198) begin
      \nz.mem_1947_sv2v_reg  <= data_i[27];
    end 
    if(N5197) begin
      \nz.mem_1946_sv2v_reg  <= data_i[26];
    end 
    if(N5196) begin
      \nz.mem_1945_sv2v_reg  <= data_i[25];
    end 
    if(N5195) begin
      \nz.mem_1944_sv2v_reg  <= data_i[24];
    end 
    if(N5194) begin
      \nz.mem_1943_sv2v_reg  <= data_i[23];
    end 
    if(N5193) begin
      \nz.mem_1942_sv2v_reg  <= data_i[22];
    end 
    if(N5192) begin
      \nz.mem_1941_sv2v_reg  <= data_i[21];
    end 
    if(N5191) begin
      \nz.mem_1940_sv2v_reg  <= data_i[20];
    end 
    if(N5190) begin
      \nz.mem_1939_sv2v_reg  <= data_i[19];
    end 
    if(N5189) begin
      \nz.mem_1938_sv2v_reg  <= data_i[18];
    end 
    if(N5188) begin
      \nz.mem_1937_sv2v_reg  <= data_i[17];
    end 
    if(N5187) begin
      \nz.mem_1936_sv2v_reg  <= data_i[16];
    end 
    if(N5186) begin
      \nz.mem_1935_sv2v_reg  <= data_i[15];
    end 
    if(N5185) begin
      \nz.mem_1934_sv2v_reg  <= data_i[14];
    end 
    if(N5184) begin
      \nz.mem_1933_sv2v_reg  <= data_i[13];
    end 
    if(N5183) begin
      \nz.mem_1932_sv2v_reg  <= data_i[12];
    end 
    if(N5182) begin
      \nz.mem_1931_sv2v_reg  <= data_i[11];
    end 
    if(N5181) begin
      \nz.mem_1930_sv2v_reg  <= data_i[10];
    end 
    if(N5180) begin
      \nz.mem_1929_sv2v_reg  <= data_i[9];
    end 
    if(N5179) begin
      \nz.mem_1928_sv2v_reg  <= data_i[8];
    end 
    if(N5178) begin
      \nz.mem_1927_sv2v_reg  <= data_i[7];
    end 
    if(N5177) begin
      \nz.mem_1926_sv2v_reg  <= data_i[6];
    end 
    if(N5176) begin
      \nz.mem_1925_sv2v_reg  <= data_i[5];
    end 
    if(N5175) begin
      \nz.mem_1924_sv2v_reg  <= data_i[4];
    end 
    if(N5174) begin
      \nz.mem_1923_sv2v_reg  <= data_i[3];
    end 
    if(N5173) begin
      \nz.mem_1922_sv2v_reg  <= data_i[2];
    end 
    if(N5172) begin
      \nz.mem_1921_sv2v_reg  <= data_i[1];
    end 
    if(N5171) begin
      \nz.mem_1920_sv2v_reg  <= data_i[0];
    end 
    if(N5170) begin
      \nz.mem_1919_sv2v_reg  <= data_i[39];
    end 
    if(N5169) begin
      \nz.mem_1918_sv2v_reg  <= data_i[38];
    end 
    if(N5168) begin
      \nz.mem_1917_sv2v_reg  <= data_i[37];
    end 
    if(N5167) begin
      \nz.mem_1916_sv2v_reg  <= data_i[36];
    end 
    if(N5166) begin
      \nz.mem_1915_sv2v_reg  <= data_i[35];
    end 
    if(N5165) begin
      \nz.mem_1914_sv2v_reg  <= data_i[34];
    end 
    if(N5164) begin
      \nz.mem_1913_sv2v_reg  <= data_i[33];
    end 
    if(N5163) begin
      \nz.mem_1912_sv2v_reg  <= data_i[32];
    end 
    if(N5162) begin
      \nz.mem_1911_sv2v_reg  <= data_i[31];
    end 
    if(N5161) begin
      \nz.mem_1910_sv2v_reg  <= data_i[30];
    end 
    if(N5160) begin
      \nz.mem_1909_sv2v_reg  <= data_i[29];
    end 
    if(N5159) begin
      \nz.mem_1908_sv2v_reg  <= data_i[28];
    end 
    if(N5158) begin
      \nz.mem_1907_sv2v_reg  <= data_i[27];
    end 
    if(N5157) begin
      \nz.mem_1906_sv2v_reg  <= data_i[26];
    end 
    if(N5156) begin
      \nz.mem_1905_sv2v_reg  <= data_i[25];
    end 
    if(N5155) begin
      \nz.mem_1904_sv2v_reg  <= data_i[24];
    end 
    if(N5154) begin
      \nz.mem_1903_sv2v_reg  <= data_i[23];
    end 
    if(N5153) begin
      \nz.mem_1902_sv2v_reg  <= data_i[22];
    end 
    if(N5152) begin
      \nz.mem_1901_sv2v_reg  <= data_i[21];
    end 
    if(N5151) begin
      \nz.mem_1900_sv2v_reg  <= data_i[20];
    end 
    if(N5150) begin
      \nz.mem_1899_sv2v_reg  <= data_i[19];
    end 
    if(N5149) begin
      \nz.mem_1898_sv2v_reg  <= data_i[18];
    end 
    if(N5148) begin
      \nz.mem_1897_sv2v_reg  <= data_i[17];
    end 
    if(N5147) begin
      \nz.mem_1896_sv2v_reg  <= data_i[16];
    end 
    if(N5146) begin
      \nz.mem_1895_sv2v_reg  <= data_i[15];
    end 
    if(N5145) begin
      \nz.mem_1894_sv2v_reg  <= data_i[14];
    end 
    if(N5144) begin
      \nz.mem_1893_sv2v_reg  <= data_i[13];
    end 
    if(N5143) begin
      \nz.mem_1892_sv2v_reg  <= data_i[12];
    end 
    if(N5142) begin
      \nz.mem_1891_sv2v_reg  <= data_i[11];
    end 
    if(N5141) begin
      \nz.mem_1890_sv2v_reg  <= data_i[10];
    end 
    if(N5140) begin
      \nz.mem_1889_sv2v_reg  <= data_i[9];
    end 
    if(N5139) begin
      \nz.mem_1888_sv2v_reg  <= data_i[8];
    end 
    if(N5138) begin
      \nz.mem_1887_sv2v_reg  <= data_i[7];
    end 
    if(N5137) begin
      \nz.mem_1886_sv2v_reg  <= data_i[6];
    end 
    if(N5136) begin
      \nz.mem_1885_sv2v_reg  <= data_i[5];
    end 
    if(N5135) begin
      \nz.mem_1884_sv2v_reg  <= data_i[4];
    end 
    if(N5134) begin
      \nz.mem_1883_sv2v_reg  <= data_i[3];
    end 
    if(N5133) begin
      \nz.mem_1882_sv2v_reg  <= data_i[2];
    end 
    if(N5132) begin
      \nz.mem_1881_sv2v_reg  <= data_i[1];
    end 
    if(N5131) begin
      \nz.mem_1880_sv2v_reg  <= data_i[0];
    end 
    if(N5130) begin
      \nz.mem_1879_sv2v_reg  <= data_i[39];
    end 
    if(N5129) begin
      \nz.mem_1878_sv2v_reg  <= data_i[38];
    end 
    if(N5128) begin
      \nz.mem_1877_sv2v_reg  <= data_i[37];
    end 
    if(N5127) begin
      \nz.mem_1876_sv2v_reg  <= data_i[36];
    end 
    if(N5126) begin
      \nz.mem_1875_sv2v_reg  <= data_i[35];
    end 
    if(N5125) begin
      \nz.mem_1874_sv2v_reg  <= data_i[34];
    end 
    if(N5124) begin
      \nz.mem_1873_sv2v_reg  <= data_i[33];
    end 
    if(N5123) begin
      \nz.mem_1872_sv2v_reg  <= data_i[32];
    end 
    if(N5122) begin
      \nz.mem_1871_sv2v_reg  <= data_i[31];
    end 
    if(N5121) begin
      \nz.mem_1870_sv2v_reg  <= data_i[30];
    end 
    if(N5120) begin
      \nz.mem_1869_sv2v_reg  <= data_i[29];
    end 
    if(N5119) begin
      \nz.mem_1868_sv2v_reg  <= data_i[28];
    end 
    if(N5118) begin
      \nz.mem_1867_sv2v_reg  <= data_i[27];
    end 
    if(N5117) begin
      \nz.mem_1866_sv2v_reg  <= data_i[26];
    end 
    if(N5116) begin
      \nz.mem_1865_sv2v_reg  <= data_i[25];
    end 
    if(N5115) begin
      \nz.mem_1864_sv2v_reg  <= data_i[24];
    end 
    if(N5114) begin
      \nz.mem_1863_sv2v_reg  <= data_i[23];
    end 
    if(N5113) begin
      \nz.mem_1862_sv2v_reg  <= data_i[22];
    end 
    if(N5112) begin
      \nz.mem_1861_sv2v_reg  <= data_i[21];
    end 
    if(N5111) begin
      \nz.mem_1860_sv2v_reg  <= data_i[20];
    end 
    if(N5110) begin
      \nz.mem_1859_sv2v_reg  <= data_i[19];
    end 
    if(N5109) begin
      \nz.mem_1858_sv2v_reg  <= data_i[18];
    end 
    if(N5108) begin
      \nz.mem_1857_sv2v_reg  <= data_i[17];
    end 
    if(N5107) begin
      \nz.mem_1856_sv2v_reg  <= data_i[16];
    end 
    if(N5106) begin
      \nz.mem_1855_sv2v_reg  <= data_i[15];
    end 
    if(N5105) begin
      \nz.mem_1854_sv2v_reg  <= data_i[14];
    end 
    if(N5104) begin
      \nz.mem_1853_sv2v_reg  <= data_i[13];
    end 
    if(N5103) begin
      \nz.mem_1852_sv2v_reg  <= data_i[12];
    end 
    if(N5102) begin
      \nz.mem_1851_sv2v_reg  <= data_i[11];
    end 
    if(N5101) begin
      \nz.mem_1850_sv2v_reg  <= data_i[10];
    end 
    if(N5100) begin
      \nz.mem_1849_sv2v_reg  <= data_i[9];
    end 
    if(N5099) begin
      \nz.mem_1848_sv2v_reg  <= data_i[8];
    end 
    if(N5098) begin
      \nz.mem_1847_sv2v_reg  <= data_i[7];
    end 
    if(N5097) begin
      \nz.mem_1846_sv2v_reg  <= data_i[6];
    end 
    if(N5096) begin
      \nz.mem_1845_sv2v_reg  <= data_i[5];
    end 
    if(N5095) begin
      \nz.mem_1844_sv2v_reg  <= data_i[4];
    end 
    if(N5094) begin
      \nz.mem_1843_sv2v_reg  <= data_i[3];
    end 
    if(N5093) begin
      \nz.mem_1842_sv2v_reg  <= data_i[2];
    end 
    if(N5092) begin
      \nz.mem_1841_sv2v_reg  <= data_i[1];
    end 
    if(N5091) begin
      \nz.mem_1840_sv2v_reg  <= data_i[0];
    end 
    if(N5090) begin
      \nz.mem_1839_sv2v_reg  <= data_i[39];
    end 
    if(N5089) begin
      \nz.mem_1838_sv2v_reg  <= data_i[38];
    end 
    if(N5088) begin
      \nz.mem_1837_sv2v_reg  <= data_i[37];
    end 
    if(N5087) begin
      \nz.mem_1836_sv2v_reg  <= data_i[36];
    end 
    if(N5086) begin
      \nz.mem_1835_sv2v_reg  <= data_i[35];
    end 
    if(N5085) begin
      \nz.mem_1834_sv2v_reg  <= data_i[34];
    end 
    if(N5084) begin
      \nz.mem_1833_sv2v_reg  <= data_i[33];
    end 
    if(N5083) begin
      \nz.mem_1832_sv2v_reg  <= data_i[32];
    end 
    if(N5082) begin
      \nz.mem_1831_sv2v_reg  <= data_i[31];
    end 
    if(N5081) begin
      \nz.mem_1830_sv2v_reg  <= data_i[30];
    end 
    if(N5080) begin
      \nz.mem_1829_sv2v_reg  <= data_i[29];
    end 
    if(N5079) begin
      \nz.mem_1828_sv2v_reg  <= data_i[28];
    end 
    if(N5078) begin
      \nz.mem_1827_sv2v_reg  <= data_i[27];
    end 
    if(N5077) begin
      \nz.mem_1826_sv2v_reg  <= data_i[26];
    end 
    if(N5076) begin
      \nz.mem_1825_sv2v_reg  <= data_i[25];
    end 
    if(N5075) begin
      \nz.mem_1824_sv2v_reg  <= data_i[24];
    end 
    if(N5074) begin
      \nz.mem_1823_sv2v_reg  <= data_i[23];
    end 
    if(N5073) begin
      \nz.mem_1822_sv2v_reg  <= data_i[22];
    end 
    if(N5072) begin
      \nz.mem_1821_sv2v_reg  <= data_i[21];
    end 
    if(N5071) begin
      \nz.mem_1820_sv2v_reg  <= data_i[20];
    end 
    if(N5070) begin
      \nz.mem_1819_sv2v_reg  <= data_i[19];
    end 
    if(N5069) begin
      \nz.mem_1818_sv2v_reg  <= data_i[18];
    end 
    if(N5068) begin
      \nz.mem_1817_sv2v_reg  <= data_i[17];
    end 
    if(N5067) begin
      \nz.mem_1816_sv2v_reg  <= data_i[16];
    end 
    if(N5066) begin
      \nz.mem_1815_sv2v_reg  <= data_i[15];
    end 
    if(N5065) begin
      \nz.mem_1814_sv2v_reg  <= data_i[14];
    end 
    if(N5064) begin
      \nz.mem_1813_sv2v_reg  <= data_i[13];
    end 
    if(N5063) begin
      \nz.mem_1812_sv2v_reg  <= data_i[12];
    end 
    if(N5062) begin
      \nz.mem_1811_sv2v_reg  <= data_i[11];
    end 
    if(N5061) begin
      \nz.mem_1810_sv2v_reg  <= data_i[10];
    end 
    if(N5060) begin
      \nz.mem_1809_sv2v_reg  <= data_i[9];
    end 
    if(N5059) begin
      \nz.mem_1808_sv2v_reg  <= data_i[8];
    end 
    if(N5058) begin
      \nz.mem_1807_sv2v_reg  <= data_i[7];
    end 
    if(N5057) begin
      \nz.mem_1806_sv2v_reg  <= data_i[6];
    end 
    if(N5056) begin
      \nz.mem_1805_sv2v_reg  <= data_i[5];
    end 
    if(N5055) begin
      \nz.mem_1804_sv2v_reg  <= data_i[4];
    end 
    if(N5054) begin
      \nz.mem_1803_sv2v_reg  <= data_i[3];
    end 
    if(N5053) begin
      \nz.mem_1802_sv2v_reg  <= data_i[2];
    end 
    if(N5052) begin
      \nz.mem_1801_sv2v_reg  <= data_i[1];
    end 
    if(N5051) begin
      \nz.mem_1800_sv2v_reg  <= data_i[0];
    end 
    if(N5050) begin
      \nz.mem_1799_sv2v_reg  <= data_i[39];
    end 
    if(N5049) begin
      \nz.mem_1798_sv2v_reg  <= data_i[38];
    end 
    if(N5048) begin
      \nz.mem_1797_sv2v_reg  <= data_i[37];
    end 
    if(N5047) begin
      \nz.mem_1796_sv2v_reg  <= data_i[36];
    end 
    if(N5046) begin
      \nz.mem_1795_sv2v_reg  <= data_i[35];
    end 
    if(N5045) begin
      \nz.mem_1794_sv2v_reg  <= data_i[34];
    end 
    if(N5044) begin
      \nz.mem_1793_sv2v_reg  <= data_i[33];
    end 
    if(N5043) begin
      \nz.mem_1792_sv2v_reg  <= data_i[32];
    end 
    if(N5042) begin
      \nz.mem_1791_sv2v_reg  <= data_i[31];
    end 
    if(N5041) begin
      \nz.mem_1790_sv2v_reg  <= data_i[30];
    end 
    if(N5040) begin
      \nz.mem_1789_sv2v_reg  <= data_i[29];
    end 
    if(N5039) begin
      \nz.mem_1788_sv2v_reg  <= data_i[28];
    end 
    if(N5038) begin
      \nz.mem_1787_sv2v_reg  <= data_i[27];
    end 
    if(N5037) begin
      \nz.mem_1786_sv2v_reg  <= data_i[26];
    end 
    if(N5036) begin
      \nz.mem_1785_sv2v_reg  <= data_i[25];
    end 
    if(N5035) begin
      \nz.mem_1784_sv2v_reg  <= data_i[24];
    end 
    if(N5034) begin
      \nz.mem_1783_sv2v_reg  <= data_i[23];
    end 
    if(N5033) begin
      \nz.mem_1782_sv2v_reg  <= data_i[22];
    end 
    if(N5032) begin
      \nz.mem_1781_sv2v_reg  <= data_i[21];
    end 
    if(N5031) begin
      \nz.mem_1780_sv2v_reg  <= data_i[20];
    end 
    if(N5030) begin
      \nz.mem_1779_sv2v_reg  <= data_i[19];
    end 
    if(N5029) begin
      \nz.mem_1778_sv2v_reg  <= data_i[18];
    end 
    if(N5028) begin
      \nz.mem_1777_sv2v_reg  <= data_i[17];
    end 
    if(N5027) begin
      \nz.mem_1776_sv2v_reg  <= data_i[16];
    end 
    if(N5026) begin
      \nz.mem_1775_sv2v_reg  <= data_i[15];
    end 
    if(N5025) begin
      \nz.mem_1774_sv2v_reg  <= data_i[14];
    end 
    if(N5024) begin
      \nz.mem_1773_sv2v_reg  <= data_i[13];
    end 
    if(N5023) begin
      \nz.mem_1772_sv2v_reg  <= data_i[12];
    end 
    if(N5022) begin
      \nz.mem_1771_sv2v_reg  <= data_i[11];
    end 
    if(N5021) begin
      \nz.mem_1770_sv2v_reg  <= data_i[10];
    end 
    if(N5020) begin
      \nz.mem_1769_sv2v_reg  <= data_i[9];
    end 
    if(N5019) begin
      \nz.mem_1768_sv2v_reg  <= data_i[8];
    end 
    if(N5018) begin
      \nz.mem_1767_sv2v_reg  <= data_i[7];
    end 
    if(N5017) begin
      \nz.mem_1766_sv2v_reg  <= data_i[6];
    end 
    if(N5016) begin
      \nz.mem_1765_sv2v_reg  <= data_i[5];
    end 
    if(N5015) begin
      \nz.mem_1764_sv2v_reg  <= data_i[4];
    end 
    if(N5014) begin
      \nz.mem_1763_sv2v_reg  <= data_i[3];
    end 
    if(N5013) begin
      \nz.mem_1762_sv2v_reg  <= data_i[2];
    end 
    if(N5012) begin
      \nz.mem_1761_sv2v_reg  <= data_i[1];
    end 
    if(N5011) begin
      \nz.mem_1760_sv2v_reg  <= data_i[0];
    end 
    if(N5010) begin
      \nz.mem_1759_sv2v_reg  <= data_i[39];
    end 
    if(N5009) begin
      \nz.mem_1758_sv2v_reg  <= data_i[38];
    end 
    if(N5008) begin
      \nz.mem_1757_sv2v_reg  <= data_i[37];
    end 
    if(N5007) begin
      \nz.mem_1756_sv2v_reg  <= data_i[36];
    end 
    if(N5006) begin
      \nz.mem_1755_sv2v_reg  <= data_i[35];
    end 
    if(N5005) begin
      \nz.mem_1754_sv2v_reg  <= data_i[34];
    end 
    if(N5004) begin
      \nz.mem_1753_sv2v_reg  <= data_i[33];
    end 
    if(N5003) begin
      \nz.mem_1752_sv2v_reg  <= data_i[32];
    end 
    if(N5002) begin
      \nz.mem_1751_sv2v_reg  <= data_i[31];
    end 
    if(N5001) begin
      \nz.mem_1750_sv2v_reg  <= data_i[30];
    end 
    if(N5000) begin
      \nz.mem_1749_sv2v_reg  <= data_i[29];
    end 
    if(N4999) begin
      \nz.mem_1748_sv2v_reg  <= data_i[28];
    end 
    if(N4998) begin
      \nz.mem_1747_sv2v_reg  <= data_i[27];
    end 
    if(N4997) begin
      \nz.mem_1746_sv2v_reg  <= data_i[26];
    end 
    if(N4996) begin
      \nz.mem_1745_sv2v_reg  <= data_i[25];
    end 
    if(N4995) begin
      \nz.mem_1744_sv2v_reg  <= data_i[24];
    end 
    if(N4994) begin
      \nz.mem_1743_sv2v_reg  <= data_i[23];
    end 
    if(N4993) begin
      \nz.mem_1742_sv2v_reg  <= data_i[22];
    end 
    if(N4992) begin
      \nz.mem_1741_sv2v_reg  <= data_i[21];
    end 
    if(N4991) begin
      \nz.mem_1740_sv2v_reg  <= data_i[20];
    end 
    if(N4990) begin
      \nz.mem_1739_sv2v_reg  <= data_i[19];
    end 
    if(N4989) begin
      \nz.mem_1738_sv2v_reg  <= data_i[18];
    end 
    if(N4988) begin
      \nz.mem_1737_sv2v_reg  <= data_i[17];
    end 
    if(N4987) begin
      \nz.mem_1736_sv2v_reg  <= data_i[16];
    end 
    if(N4986) begin
      \nz.mem_1735_sv2v_reg  <= data_i[15];
    end 
    if(N4985) begin
      \nz.mem_1734_sv2v_reg  <= data_i[14];
    end 
    if(N4984) begin
      \nz.mem_1733_sv2v_reg  <= data_i[13];
    end 
    if(N4983) begin
      \nz.mem_1732_sv2v_reg  <= data_i[12];
    end 
    if(N4982) begin
      \nz.mem_1731_sv2v_reg  <= data_i[11];
    end 
    if(N4981) begin
      \nz.mem_1730_sv2v_reg  <= data_i[10];
    end 
    if(N4980) begin
      \nz.mem_1729_sv2v_reg  <= data_i[9];
    end 
    if(N4979) begin
      \nz.mem_1728_sv2v_reg  <= data_i[8];
    end 
    if(N4978) begin
      \nz.mem_1727_sv2v_reg  <= data_i[7];
    end 
    if(N4977) begin
      \nz.mem_1726_sv2v_reg  <= data_i[6];
    end 
    if(N4976) begin
      \nz.mem_1725_sv2v_reg  <= data_i[5];
    end 
    if(N4975) begin
      \nz.mem_1724_sv2v_reg  <= data_i[4];
    end 
    if(N4974) begin
      \nz.mem_1723_sv2v_reg  <= data_i[3];
    end 
    if(N4973) begin
      \nz.mem_1722_sv2v_reg  <= data_i[2];
    end 
    if(N4972) begin
      \nz.mem_1721_sv2v_reg  <= data_i[1];
    end 
    if(N4971) begin
      \nz.mem_1720_sv2v_reg  <= data_i[0];
    end 
    if(N4970) begin
      \nz.mem_1719_sv2v_reg  <= data_i[39];
    end 
    if(N4969) begin
      \nz.mem_1718_sv2v_reg  <= data_i[38];
    end 
    if(N4968) begin
      \nz.mem_1717_sv2v_reg  <= data_i[37];
    end 
    if(N4967) begin
      \nz.mem_1716_sv2v_reg  <= data_i[36];
    end 
    if(N4966) begin
      \nz.mem_1715_sv2v_reg  <= data_i[35];
    end 
    if(N4965) begin
      \nz.mem_1714_sv2v_reg  <= data_i[34];
    end 
    if(N4964) begin
      \nz.mem_1713_sv2v_reg  <= data_i[33];
    end 
    if(N4963) begin
      \nz.mem_1712_sv2v_reg  <= data_i[32];
    end 
    if(N4962) begin
      \nz.mem_1711_sv2v_reg  <= data_i[31];
    end 
    if(N4961) begin
      \nz.mem_1710_sv2v_reg  <= data_i[30];
    end 
    if(N4960) begin
      \nz.mem_1709_sv2v_reg  <= data_i[29];
    end 
    if(N4959) begin
      \nz.mem_1708_sv2v_reg  <= data_i[28];
    end 
    if(N4958) begin
      \nz.mem_1707_sv2v_reg  <= data_i[27];
    end 
    if(N4957) begin
      \nz.mem_1706_sv2v_reg  <= data_i[26];
    end 
    if(N4956) begin
      \nz.mem_1705_sv2v_reg  <= data_i[25];
    end 
    if(N4955) begin
      \nz.mem_1704_sv2v_reg  <= data_i[24];
    end 
    if(N4954) begin
      \nz.mem_1703_sv2v_reg  <= data_i[23];
    end 
    if(N4953) begin
      \nz.mem_1702_sv2v_reg  <= data_i[22];
    end 
    if(N4952) begin
      \nz.mem_1701_sv2v_reg  <= data_i[21];
    end 
    if(N4951) begin
      \nz.mem_1700_sv2v_reg  <= data_i[20];
    end 
    if(N4950) begin
      \nz.mem_1699_sv2v_reg  <= data_i[19];
    end 
    if(N4949) begin
      \nz.mem_1698_sv2v_reg  <= data_i[18];
    end 
    if(N4948) begin
      \nz.mem_1697_sv2v_reg  <= data_i[17];
    end 
    if(N4947) begin
      \nz.mem_1696_sv2v_reg  <= data_i[16];
    end 
    if(N4946) begin
      \nz.mem_1695_sv2v_reg  <= data_i[15];
    end 
    if(N4945) begin
      \nz.mem_1694_sv2v_reg  <= data_i[14];
    end 
    if(N4944) begin
      \nz.mem_1693_sv2v_reg  <= data_i[13];
    end 
    if(N4943) begin
      \nz.mem_1692_sv2v_reg  <= data_i[12];
    end 
    if(N4942) begin
      \nz.mem_1691_sv2v_reg  <= data_i[11];
    end 
    if(N4941) begin
      \nz.mem_1690_sv2v_reg  <= data_i[10];
    end 
    if(N4940) begin
      \nz.mem_1689_sv2v_reg  <= data_i[9];
    end 
    if(N4939) begin
      \nz.mem_1688_sv2v_reg  <= data_i[8];
    end 
    if(N4938) begin
      \nz.mem_1687_sv2v_reg  <= data_i[7];
    end 
    if(N4937) begin
      \nz.mem_1686_sv2v_reg  <= data_i[6];
    end 
    if(N4936) begin
      \nz.mem_1685_sv2v_reg  <= data_i[5];
    end 
    if(N4935) begin
      \nz.mem_1684_sv2v_reg  <= data_i[4];
    end 
    if(N4934) begin
      \nz.mem_1683_sv2v_reg  <= data_i[3];
    end 
    if(N4933) begin
      \nz.mem_1682_sv2v_reg  <= data_i[2];
    end 
    if(N4932) begin
      \nz.mem_1681_sv2v_reg  <= data_i[1];
    end 
    if(N4931) begin
      \nz.mem_1680_sv2v_reg  <= data_i[0];
    end 
    if(N4930) begin
      \nz.mem_1679_sv2v_reg  <= data_i[39];
    end 
    if(N4929) begin
      \nz.mem_1678_sv2v_reg  <= data_i[38];
    end 
    if(N4928) begin
      \nz.mem_1677_sv2v_reg  <= data_i[37];
    end 
    if(N4927) begin
      \nz.mem_1676_sv2v_reg  <= data_i[36];
    end 
    if(N4926) begin
      \nz.mem_1675_sv2v_reg  <= data_i[35];
    end 
    if(N4925) begin
      \nz.mem_1674_sv2v_reg  <= data_i[34];
    end 
    if(N4924) begin
      \nz.mem_1673_sv2v_reg  <= data_i[33];
    end 
    if(N4923) begin
      \nz.mem_1672_sv2v_reg  <= data_i[32];
    end 
    if(N4922) begin
      \nz.mem_1671_sv2v_reg  <= data_i[31];
    end 
    if(N4921) begin
      \nz.mem_1670_sv2v_reg  <= data_i[30];
    end 
    if(N4920) begin
      \nz.mem_1669_sv2v_reg  <= data_i[29];
    end 
    if(N4919) begin
      \nz.mem_1668_sv2v_reg  <= data_i[28];
    end 
    if(N4918) begin
      \nz.mem_1667_sv2v_reg  <= data_i[27];
    end 
    if(N4917) begin
      \nz.mem_1666_sv2v_reg  <= data_i[26];
    end 
    if(N4916) begin
      \nz.mem_1665_sv2v_reg  <= data_i[25];
    end 
    if(N4915) begin
      \nz.mem_1664_sv2v_reg  <= data_i[24];
    end 
    if(N4914) begin
      \nz.mem_1663_sv2v_reg  <= data_i[23];
    end 
    if(N4913) begin
      \nz.mem_1662_sv2v_reg  <= data_i[22];
    end 
    if(N4912) begin
      \nz.mem_1661_sv2v_reg  <= data_i[21];
    end 
    if(N4911) begin
      \nz.mem_1660_sv2v_reg  <= data_i[20];
    end 
    if(N4910) begin
      \nz.mem_1659_sv2v_reg  <= data_i[19];
    end 
    if(N4909) begin
      \nz.mem_1658_sv2v_reg  <= data_i[18];
    end 
    if(N4908) begin
      \nz.mem_1657_sv2v_reg  <= data_i[17];
    end 
    if(N4907) begin
      \nz.mem_1656_sv2v_reg  <= data_i[16];
    end 
    if(N4906) begin
      \nz.mem_1655_sv2v_reg  <= data_i[15];
    end 
    if(N4905) begin
      \nz.mem_1654_sv2v_reg  <= data_i[14];
    end 
    if(N4904) begin
      \nz.mem_1653_sv2v_reg  <= data_i[13];
    end 
    if(N4903) begin
      \nz.mem_1652_sv2v_reg  <= data_i[12];
    end 
    if(N4902) begin
      \nz.mem_1651_sv2v_reg  <= data_i[11];
    end 
    if(N4901) begin
      \nz.mem_1650_sv2v_reg  <= data_i[10];
    end 
    if(N4900) begin
      \nz.mem_1649_sv2v_reg  <= data_i[9];
    end 
    if(N4899) begin
      \nz.mem_1648_sv2v_reg  <= data_i[8];
    end 
    if(N4898) begin
      \nz.mem_1647_sv2v_reg  <= data_i[7];
    end 
    if(N4897) begin
      \nz.mem_1646_sv2v_reg  <= data_i[6];
    end 
    if(N4896) begin
      \nz.mem_1645_sv2v_reg  <= data_i[5];
    end 
    if(N4895) begin
      \nz.mem_1644_sv2v_reg  <= data_i[4];
    end 
    if(N4894) begin
      \nz.mem_1643_sv2v_reg  <= data_i[3];
    end 
    if(N4893) begin
      \nz.mem_1642_sv2v_reg  <= data_i[2];
    end 
    if(N4892) begin
      \nz.mem_1641_sv2v_reg  <= data_i[1];
    end 
    if(N4891) begin
      \nz.mem_1640_sv2v_reg  <= data_i[0];
    end 
    if(N4890) begin
      \nz.mem_1639_sv2v_reg  <= data_i[39];
    end 
    if(N4889) begin
      \nz.mem_1638_sv2v_reg  <= data_i[38];
    end 
    if(N4888) begin
      \nz.mem_1637_sv2v_reg  <= data_i[37];
    end 
    if(N4887) begin
      \nz.mem_1636_sv2v_reg  <= data_i[36];
    end 
    if(N4886) begin
      \nz.mem_1635_sv2v_reg  <= data_i[35];
    end 
    if(N4885) begin
      \nz.mem_1634_sv2v_reg  <= data_i[34];
    end 
    if(N4884) begin
      \nz.mem_1633_sv2v_reg  <= data_i[33];
    end 
    if(N4883) begin
      \nz.mem_1632_sv2v_reg  <= data_i[32];
    end 
    if(N4882) begin
      \nz.mem_1631_sv2v_reg  <= data_i[31];
    end 
    if(N4881) begin
      \nz.mem_1630_sv2v_reg  <= data_i[30];
    end 
    if(N4880) begin
      \nz.mem_1629_sv2v_reg  <= data_i[29];
    end 
    if(N4879) begin
      \nz.mem_1628_sv2v_reg  <= data_i[28];
    end 
    if(N4878) begin
      \nz.mem_1627_sv2v_reg  <= data_i[27];
    end 
    if(N4877) begin
      \nz.mem_1626_sv2v_reg  <= data_i[26];
    end 
    if(N4876) begin
      \nz.mem_1625_sv2v_reg  <= data_i[25];
    end 
    if(N4875) begin
      \nz.mem_1624_sv2v_reg  <= data_i[24];
    end 
    if(N4874) begin
      \nz.mem_1623_sv2v_reg  <= data_i[23];
    end 
    if(N4873) begin
      \nz.mem_1622_sv2v_reg  <= data_i[22];
    end 
    if(N4872) begin
      \nz.mem_1621_sv2v_reg  <= data_i[21];
    end 
    if(N4871) begin
      \nz.mem_1620_sv2v_reg  <= data_i[20];
    end 
    if(N4870) begin
      \nz.mem_1619_sv2v_reg  <= data_i[19];
    end 
    if(N4869) begin
      \nz.mem_1618_sv2v_reg  <= data_i[18];
    end 
    if(N4868) begin
      \nz.mem_1617_sv2v_reg  <= data_i[17];
    end 
    if(N4867) begin
      \nz.mem_1616_sv2v_reg  <= data_i[16];
    end 
    if(N4866) begin
      \nz.mem_1615_sv2v_reg  <= data_i[15];
    end 
    if(N4865) begin
      \nz.mem_1614_sv2v_reg  <= data_i[14];
    end 
    if(N4864) begin
      \nz.mem_1613_sv2v_reg  <= data_i[13];
    end 
    if(N4863) begin
      \nz.mem_1612_sv2v_reg  <= data_i[12];
    end 
    if(N4862) begin
      \nz.mem_1611_sv2v_reg  <= data_i[11];
    end 
    if(N4861) begin
      \nz.mem_1610_sv2v_reg  <= data_i[10];
    end 
    if(N4860) begin
      \nz.mem_1609_sv2v_reg  <= data_i[9];
    end 
    if(N4859) begin
      \nz.mem_1608_sv2v_reg  <= data_i[8];
    end 
    if(N4858) begin
      \nz.mem_1607_sv2v_reg  <= data_i[7];
    end 
    if(N4857) begin
      \nz.mem_1606_sv2v_reg  <= data_i[6];
    end 
    if(N4856) begin
      \nz.mem_1605_sv2v_reg  <= data_i[5];
    end 
    if(N4855) begin
      \nz.mem_1604_sv2v_reg  <= data_i[4];
    end 
    if(N4854) begin
      \nz.mem_1603_sv2v_reg  <= data_i[3];
    end 
    if(N4853) begin
      \nz.mem_1602_sv2v_reg  <= data_i[2];
    end 
    if(N4852) begin
      \nz.mem_1601_sv2v_reg  <= data_i[1];
    end 
    if(N4851) begin
      \nz.mem_1600_sv2v_reg  <= data_i[0];
    end 
    if(N4850) begin
      \nz.mem_1599_sv2v_reg  <= data_i[39];
    end 
    if(N4849) begin
      \nz.mem_1598_sv2v_reg  <= data_i[38];
    end 
    if(N4848) begin
      \nz.mem_1597_sv2v_reg  <= data_i[37];
    end 
    if(N4847) begin
      \nz.mem_1596_sv2v_reg  <= data_i[36];
    end 
    if(N4846) begin
      \nz.mem_1595_sv2v_reg  <= data_i[35];
    end 
    if(N4845) begin
      \nz.mem_1594_sv2v_reg  <= data_i[34];
    end 
    if(N4844) begin
      \nz.mem_1593_sv2v_reg  <= data_i[33];
    end 
    if(N4843) begin
      \nz.mem_1592_sv2v_reg  <= data_i[32];
    end 
    if(N4842) begin
      \nz.mem_1591_sv2v_reg  <= data_i[31];
    end 
    if(N4841) begin
      \nz.mem_1590_sv2v_reg  <= data_i[30];
    end 
    if(N4840) begin
      \nz.mem_1589_sv2v_reg  <= data_i[29];
    end 
    if(N4839) begin
      \nz.mem_1588_sv2v_reg  <= data_i[28];
    end 
    if(N4838) begin
      \nz.mem_1587_sv2v_reg  <= data_i[27];
    end 
    if(N4837) begin
      \nz.mem_1586_sv2v_reg  <= data_i[26];
    end 
    if(N4836) begin
      \nz.mem_1585_sv2v_reg  <= data_i[25];
    end 
    if(N4835) begin
      \nz.mem_1584_sv2v_reg  <= data_i[24];
    end 
    if(N4834) begin
      \nz.mem_1583_sv2v_reg  <= data_i[23];
    end 
    if(N4833) begin
      \nz.mem_1582_sv2v_reg  <= data_i[22];
    end 
    if(N4832) begin
      \nz.mem_1581_sv2v_reg  <= data_i[21];
    end 
    if(N4831) begin
      \nz.mem_1580_sv2v_reg  <= data_i[20];
    end 
    if(N4830) begin
      \nz.mem_1579_sv2v_reg  <= data_i[19];
    end 
    if(N4829) begin
      \nz.mem_1578_sv2v_reg  <= data_i[18];
    end 
    if(N4828) begin
      \nz.mem_1577_sv2v_reg  <= data_i[17];
    end 
    if(N4827) begin
      \nz.mem_1576_sv2v_reg  <= data_i[16];
    end 
    if(N4826) begin
      \nz.mem_1575_sv2v_reg  <= data_i[15];
    end 
    if(N4825) begin
      \nz.mem_1574_sv2v_reg  <= data_i[14];
    end 
    if(N4824) begin
      \nz.mem_1573_sv2v_reg  <= data_i[13];
    end 
    if(N4823) begin
      \nz.mem_1572_sv2v_reg  <= data_i[12];
    end 
    if(N4822) begin
      \nz.mem_1571_sv2v_reg  <= data_i[11];
    end 
    if(N4821) begin
      \nz.mem_1570_sv2v_reg  <= data_i[10];
    end 
    if(N4820) begin
      \nz.mem_1569_sv2v_reg  <= data_i[9];
    end 
    if(N4819) begin
      \nz.mem_1568_sv2v_reg  <= data_i[8];
    end 
    if(N4818) begin
      \nz.mem_1567_sv2v_reg  <= data_i[7];
    end 
    if(N4817) begin
      \nz.mem_1566_sv2v_reg  <= data_i[6];
    end 
    if(N4816) begin
      \nz.mem_1565_sv2v_reg  <= data_i[5];
    end 
    if(N4815) begin
      \nz.mem_1564_sv2v_reg  <= data_i[4];
    end 
    if(N4814) begin
      \nz.mem_1563_sv2v_reg  <= data_i[3];
    end 
    if(N4813) begin
      \nz.mem_1562_sv2v_reg  <= data_i[2];
    end 
    if(N4812) begin
      \nz.mem_1561_sv2v_reg  <= data_i[1];
    end 
    if(N4811) begin
      \nz.mem_1560_sv2v_reg  <= data_i[0];
    end 
    if(N4810) begin
      \nz.mem_1559_sv2v_reg  <= data_i[39];
    end 
    if(N4809) begin
      \nz.mem_1558_sv2v_reg  <= data_i[38];
    end 
    if(N4808) begin
      \nz.mem_1557_sv2v_reg  <= data_i[37];
    end 
    if(N4807) begin
      \nz.mem_1556_sv2v_reg  <= data_i[36];
    end 
    if(N4806) begin
      \nz.mem_1555_sv2v_reg  <= data_i[35];
    end 
    if(N4805) begin
      \nz.mem_1554_sv2v_reg  <= data_i[34];
    end 
    if(N4804) begin
      \nz.mem_1553_sv2v_reg  <= data_i[33];
    end 
    if(N4803) begin
      \nz.mem_1552_sv2v_reg  <= data_i[32];
    end 
    if(N4802) begin
      \nz.mem_1551_sv2v_reg  <= data_i[31];
    end 
    if(N4801) begin
      \nz.mem_1550_sv2v_reg  <= data_i[30];
    end 
    if(N4800) begin
      \nz.mem_1549_sv2v_reg  <= data_i[29];
    end 
    if(N4799) begin
      \nz.mem_1548_sv2v_reg  <= data_i[28];
    end 
    if(N4798) begin
      \nz.mem_1547_sv2v_reg  <= data_i[27];
    end 
    if(N4797) begin
      \nz.mem_1546_sv2v_reg  <= data_i[26];
    end 
    if(N4796) begin
      \nz.mem_1545_sv2v_reg  <= data_i[25];
    end 
    if(N4795) begin
      \nz.mem_1544_sv2v_reg  <= data_i[24];
    end 
    if(N4794) begin
      \nz.mem_1543_sv2v_reg  <= data_i[23];
    end 
    if(N4793) begin
      \nz.mem_1542_sv2v_reg  <= data_i[22];
    end 
    if(N4792) begin
      \nz.mem_1541_sv2v_reg  <= data_i[21];
    end 
    if(N4791) begin
      \nz.mem_1540_sv2v_reg  <= data_i[20];
    end 
    if(N4790) begin
      \nz.mem_1539_sv2v_reg  <= data_i[19];
    end 
    if(N4789) begin
      \nz.mem_1538_sv2v_reg  <= data_i[18];
    end 
    if(N4788) begin
      \nz.mem_1537_sv2v_reg  <= data_i[17];
    end 
    if(N4787) begin
      \nz.mem_1536_sv2v_reg  <= data_i[16];
    end 
    if(N4786) begin
      \nz.mem_1535_sv2v_reg  <= data_i[15];
    end 
    if(N4785) begin
      \nz.mem_1534_sv2v_reg  <= data_i[14];
    end 
    if(N4784) begin
      \nz.mem_1533_sv2v_reg  <= data_i[13];
    end 
    if(N4783) begin
      \nz.mem_1532_sv2v_reg  <= data_i[12];
    end 
    if(N4782) begin
      \nz.mem_1531_sv2v_reg  <= data_i[11];
    end 
    if(N4781) begin
      \nz.mem_1530_sv2v_reg  <= data_i[10];
    end 
    if(N4780) begin
      \nz.mem_1529_sv2v_reg  <= data_i[9];
    end 
    if(N4779) begin
      \nz.mem_1528_sv2v_reg  <= data_i[8];
    end 
    if(N4778) begin
      \nz.mem_1527_sv2v_reg  <= data_i[7];
    end 
    if(N4777) begin
      \nz.mem_1526_sv2v_reg  <= data_i[6];
    end 
    if(N4776) begin
      \nz.mem_1525_sv2v_reg  <= data_i[5];
    end 
    if(N4775) begin
      \nz.mem_1524_sv2v_reg  <= data_i[4];
    end 
    if(N4774) begin
      \nz.mem_1523_sv2v_reg  <= data_i[3];
    end 
    if(N4773) begin
      \nz.mem_1522_sv2v_reg  <= data_i[2];
    end 
    if(N4772) begin
      \nz.mem_1521_sv2v_reg  <= data_i[1];
    end 
    if(N4771) begin
      \nz.mem_1520_sv2v_reg  <= data_i[0];
    end 
    if(N4770) begin
      \nz.mem_1519_sv2v_reg  <= data_i[39];
    end 
    if(N4769) begin
      \nz.mem_1518_sv2v_reg  <= data_i[38];
    end 
    if(N4768) begin
      \nz.mem_1517_sv2v_reg  <= data_i[37];
    end 
    if(N4767) begin
      \nz.mem_1516_sv2v_reg  <= data_i[36];
    end 
    if(N4766) begin
      \nz.mem_1515_sv2v_reg  <= data_i[35];
    end 
    if(N4765) begin
      \nz.mem_1514_sv2v_reg  <= data_i[34];
    end 
    if(N4764) begin
      \nz.mem_1513_sv2v_reg  <= data_i[33];
    end 
    if(N4763) begin
      \nz.mem_1512_sv2v_reg  <= data_i[32];
    end 
    if(N4762) begin
      \nz.mem_1511_sv2v_reg  <= data_i[31];
    end 
    if(N4761) begin
      \nz.mem_1510_sv2v_reg  <= data_i[30];
    end 
    if(N4760) begin
      \nz.mem_1509_sv2v_reg  <= data_i[29];
    end 
    if(N4759) begin
      \nz.mem_1508_sv2v_reg  <= data_i[28];
    end 
    if(N4758) begin
      \nz.mem_1507_sv2v_reg  <= data_i[27];
    end 
    if(N4757) begin
      \nz.mem_1506_sv2v_reg  <= data_i[26];
    end 
    if(N4756) begin
      \nz.mem_1505_sv2v_reg  <= data_i[25];
    end 
    if(N4755) begin
      \nz.mem_1504_sv2v_reg  <= data_i[24];
    end 
    if(N4754) begin
      \nz.mem_1503_sv2v_reg  <= data_i[23];
    end 
    if(N4753) begin
      \nz.mem_1502_sv2v_reg  <= data_i[22];
    end 
    if(N4752) begin
      \nz.mem_1501_sv2v_reg  <= data_i[21];
    end 
    if(N4751) begin
      \nz.mem_1500_sv2v_reg  <= data_i[20];
    end 
    if(N4750) begin
      \nz.mem_1499_sv2v_reg  <= data_i[19];
    end 
    if(N4749) begin
      \nz.mem_1498_sv2v_reg  <= data_i[18];
    end 
    if(N4748) begin
      \nz.mem_1497_sv2v_reg  <= data_i[17];
    end 
    if(N4747) begin
      \nz.mem_1496_sv2v_reg  <= data_i[16];
    end 
    if(N4746) begin
      \nz.mem_1495_sv2v_reg  <= data_i[15];
    end 
    if(N4745) begin
      \nz.mem_1494_sv2v_reg  <= data_i[14];
    end 
    if(N4744) begin
      \nz.mem_1493_sv2v_reg  <= data_i[13];
    end 
    if(N4743) begin
      \nz.mem_1492_sv2v_reg  <= data_i[12];
    end 
    if(N4742) begin
      \nz.mem_1491_sv2v_reg  <= data_i[11];
    end 
    if(N4741) begin
      \nz.mem_1490_sv2v_reg  <= data_i[10];
    end 
    if(N4740) begin
      \nz.mem_1489_sv2v_reg  <= data_i[9];
    end 
    if(N4739) begin
      \nz.mem_1488_sv2v_reg  <= data_i[8];
    end 
    if(N4738) begin
      \nz.mem_1487_sv2v_reg  <= data_i[7];
    end 
    if(N4737) begin
      \nz.mem_1486_sv2v_reg  <= data_i[6];
    end 
    if(N4736) begin
      \nz.mem_1485_sv2v_reg  <= data_i[5];
    end 
    if(N4735) begin
      \nz.mem_1484_sv2v_reg  <= data_i[4];
    end 
    if(N4734) begin
      \nz.mem_1483_sv2v_reg  <= data_i[3];
    end 
    if(N4733) begin
      \nz.mem_1482_sv2v_reg  <= data_i[2];
    end 
    if(N4732) begin
      \nz.mem_1481_sv2v_reg  <= data_i[1];
    end 
    if(N4731) begin
      \nz.mem_1480_sv2v_reg  <= data_i[0];
    end 
    if(N4730) begin
      \nz.mem_1479_sv2v_reg  <= data_i[39];
    end 
    if(N4729) begin
      \nz.mem_1478_sv2v_reg  <= data_i[38];
    end 
    if(N4728) begin
      \nz.mem_1477_sv2v_reg  <= data_i[37];
    end 
    if(N4727) begin
      \nz.mem_1476_sv2v_reg  <= data_i[36];
    end 
    if(N4726) begin
      \nz.mem_1475_sv2v_reg  <= data_i[35];
    end 
    if(N4725) begin
      \nz.mem_1474_sv2v_reg  <= data_i[34];
    end 
    if(N4724) begin
      \nz.mem_1473_sv2v_reg  <= data_i[33];
    end 
    if(N4723) begin
      \nz.mem_1472_sv2v_reg  <= data_i[32];
    end 
    if(N4722) begin
      \nz.mem_1471_sv2v_reg  <= data_i[31];
    end 
    if(N4721) begin
      \nz.mem_1470_sv2v_reg  <= data_i[30];
    end 
    if(N4720) begin
      \nz.mem_1469_sv2v_reg  <= data_i[29];
    end 
    if(N4719) begin
      \nz.mem_1468_sv2v_reg  <= data_i[28];
    end 
    if(N4718) begin
      \nz.mem_1467_sv2v_reg  <= data_i[27];
    end 
    if(N4717) begin
      \nz.mem_1466_sv2v_reg  <= data_i[26];
    end 
    if(N4716) begin
      \nz.mem_1465_sv2v_reg  <= data_i[25];
    end 
    if(N4715) begin
      \nz.mem_1464_sv2v_reg  <= data_i[24];
    end 
    if(N4714) begin
      \nz.mem_1463_sv2v_reg  <= data_i[23];
    end 
    if(N4713) begin
      \nz.mem_1462_sv2v_reg  <= data_i[22];
    end 
    if(N4712) begin
      \nz.mem_1461_sv2v_reg  <= data_i[21];
    end 
    if(N4711) begin
      \nz.mem_1460_sv2v_reg  <= data_i[20];
    end 
    if(N4710) begin
      \nz.mem_1459_sv2v_reg  <= data_i[19];
    end 
    if(N4709) begin
      \nz.mem_1458_sv2v_reg  <= data_i[18];
    end 
    if(N4708) begin
      \nz.mem_1457_sv2v_reg  <= data_i[17];
    end 
    if(N4707) begin
      \nz.mem_1456_sv2v_reg  <= data_i[16];
    end 
    if(N4706) begin
      \nz.mem_1455_sv2v_reg  <= data_i[15];
    end 
    if(N4705) begin
      \nz.mem_1454_sv2v_reg  <= data_i[14];
    end 
    if(N4704) begin
      \nz.mem_1453_sv2v_reg  <= data_i[13];
    end 
    if(N4703) begin
      \nz.mem_1452_sv2v_reg  <= data_i[12];
    end 
    if(N4702) begin
      \nz.mem_1451_sv2v_reg  <= data_i[11];
    end 
    if(N4701) begin
      \nz.mem_1450_sv2v_reg  <= data_i[10];
    end 
    if(N4700) begin
      \nz.mem_1449_sv2v_reg  <= data_i[9];
    end 
    if(N4699) begin
      \nz.mem_1448_sv2v_reg  <= data_i[8];
    end 
    if(N4698) begin
      \nz.mem_1447_sv2v_reg  <= data_i[7];
    end 
    if(N4697) begin
      \nz.mem_1446_sv2v_reg  <= data_i[6];
    end 
    if(N4696) begin
      \nz.mem_1445_sv2v_reg  <= data_i[5];
    end 
    if(N4695) begin
      \nz.mem_1444_sv2v_reg  <= data_i[4];
    end 
    if(N4694) begin
      \nz.mem_1443_sv2v_reg  <= data_i[3];
    end 
    if(N4693) begin
      \nz.mem_1442_sv2v_reg  <= data_i[2];
    end 
    if(N4692) begin
      \nz.mem_1441_sv2v_reg  <= data_i[1];
    end 
    if(N4691) begin
      \nz.mem_1440_sv2v_reg  <= data_i[0];
    end 
    if(N4690) begin
      \nz.mem_1439_sv2v_reg  <= data_i[39];
    end 
    if(N4689) begin
      \nz.mem_1438_sv2v_reg  <= data_i[38];
    end 
    if(N4688) begin
      \nz.mem_1437_sv2v_reg  <= data_i[37];
    end 
    if(N4687) begin
      \nz.mem_1436_sv2v_reg  <= data_i[36];
    end 
    if(N4686) begin
      \nz.mem_1435_sv2v_reg  <= data_i[35];
    end 
    if(N4685) begin
      \nz.mem_1434_sv2v_reg  <= data_i[34];
    end 
    if(N4684) begin
      \nz.mem_1433_sv2v_reg  <= data_i[33];
    end 
    if(N4683) begin
      \nz.mem_1432_sv2v_reg  <= data_i[32];
    end 
    if(N4682) begin
      \nz.mem_1431_sv2v_reg  <= data_i[31];
    end 
    if(N4681) begin
      \nz.mem_1430_sv2v_reg  <= data_i[30];
    end 
    if(N4680) begin
      \nz.mem_1429_sv2v_reg  <= data_i[29];
    end 
    if(N4679) begin
      \nz.mem_1428_sv2v_reg  <= data_i[28];
    end 
    if(N4678) begin
      \nz.mem_1427_sv2v_reg  <= data_i[27];
    end 
    if(N4677) begin
      \nz.mem_1426_sv2v_reg  <= data_i[26];
    end 
    if(N4676) begin
      \nz.mem_1425_sv2v_reg  <= data_i[25];
    end 
    if(N4675) begin
      \nz.mem_1424_sv2v_reg  <= data_i[24];
    end 
    if(N4674) begin
      \nz.mem_1423_sv2v_reg  <= data_i[23];
    end 
    if(N4673) begin
      \nz.mem_1422_sv2v_reg  <= data_i[22];
    end 
    if(N4672) begin
      \nz.mem_1421_sv2v_reg  <= data_i[21];
    end 
    if(N4671) begin
      \nz.mem_1420_sv2v_reg  <= data_i[20];
    end 
    if(N4670) begin
      \nz.mem_1419_sv2v_reg  <= data_i[19];
    end 
    if(N4669) begin
      \nz.mem_1418_sv2v_reg  <= data_i[18];
    end 
    if(N4668) begin
      \nz.mem_1417_sv2v_reg  <= data_i[17];
    end 
    if(N4667) begin
      \nz.mem_1416_sv2v_reg  <= data_i[16];
    end 
    if(N4666) begin
      \nz.mem_1415_sv2v_reg  <= data_i[15];
    end 
    if(N4665) begin
      \nz.mem_1414_sv2v_reg  <= data_i[14];
    end 
    if(N4664) begin
      \nz.mem_1413_sv2v_reg  <= data_i[13];
    end 
    if(N4663) begin
      \nz.mem_1412_sv2v_reg  <= data_i[12];
    end 
    if(N4662) begin
      \nz.mem_1411_sv2v_reg  <= data_i[11];
    end 
    if(N4661) begin
      \nz.mem_1410_sv2v_reg  <= data_i[10];
    end 
    if(N4660) begin
      \nz.mem_1409_sv2v_reg  <= data_i[9];
    end 
    if(N4659) begin
      \nz.mem_1408_sv2v_reg  <= data_i[8];
    end 
    if(N4658) begin
      \nz.mem_1407_sv2v_reg  <= data_i[7];
    end 
    if(N4657) begin
      \nz.mem_1406_sv2v_reg  <= data_i[6];
    end 
    if(N4656) begin
      \nz.mem_1405_sv2v_reg  <= data_i[5];
    end 
    if(N4655) begin
      \nz.mem_1404_sv2v_reg  <= data_i[4];
    end 
    if(N4654) begin
      \nz.mem_1403_sv2v_reg  <= data_i[3];
    end 
    if(N4653) begin
      \nz.mem_1402_sv2v_reg  <= data_i[2];
    end 
    if(N4652) begin
      \nz.mem_1401_sv2v_reg  <= data_i[1];
    end 
    if(N4651) begin
      \nz.mem_1400_sv2v_reg  <= data_i[0];
    end 
    if(N4650) begin
      \nz.mem_1399_sv2v_reg  <= data_i[39];
    end 
    if(N4649) begin
      \nz.mem_1398_sv2v_reg  <= data_i[38];
    end 
    if(N4648) begin
      \nz.mem_1397_sv2v_reg  <= data_i[37];
    end 
    if(N4647) begin
      \nz.mem_1396_sv2v_reg  <= data_i[36];
    end 
    if(N4646) begin
      \nz.mem_1395_sv2v_reg  <= data_i[35];
    end 
    if(N4645) begin
      \nz.mem_1394_sv2v_reg  <= data_i[34];
    end 
    if(N4644) begin
      \nz.mem_1393_sv2v_reg  <= data_i[33];
    end 
    if(N4643) begin
      \nz.mem_1392_sv2v_reg  <= data_i[32];
    end 
    if(N4642) begin
      \nz.mem_1391_sv2v_reg  <= data_i[31];
    end 
    if(N4641) begin
      \nz.mem_1390_sv2v_reg  <= data_i[30];
    end 
    if(N4640) begin
      \nz.mem_1389_sv2v_reg  <= data_i[29];
    end 
    if(N4639) begin
      \nz.mem_1388_sv2v_reg  <= data_i[28];
    end 
    if(N4638) begin
      \nz.mem_1387_sv2v_reg  <= data_i[27];
    end 
    if(N4637) begin
      \nz.mem_1386_sv2v_reg  <= data_i[26];
    end 
    if(N4636) begin
      \nz.mem_1385_sv2v_reg  <= data_i[25];
    end 
    if(N4635) begin
      \nz.mem_1384_sv2v_reg  <= data_i[24];
    end 
    if(N4634) begin
      \nz.mem_1383_sv2v_reg  <= data_i[23];
    end 
    if(N4633) begin
      \nz.mem_1382_sv2v_reg  <= data_i[22];
    end 
    if(N4632) begin
      \nz.mem_1381_sv2v_reg  <= data_i[21];
    end 
    if(N4631) begin
      \nz.mem_1380_sv2v_reg  <= data_i[20];
    end 
    if(N4630) begin
      \nz.mem_1379_sv2v_reg  <= data_i[19];
    end 
    if(N4629) begin
      \nz.mem_1378_sv2v_reg  <= data_i[18];
    end 
    if(N4628) begin
      \nz.mem_1377_sv2v_reg  <= data_i[17];
    end 
    if(N4627) begin
      \nz.mem_1376_sv2v_reg  <= data_i[16];
    end 
    if(N4626) begin
      \nz.mem_1375_sv2v_reg  <= data_i[15];
    end 
    if(N4625) begin
      \nz.mem_1374_sv2v_reg  <= data_i[14];
    end 
    if(N4624) begin
      \nz.mem_1373_sv2v_reg  <= data_i[13];
    end 
    if(N4623) begin
      \nz.mem_1372_sv2v_reg  <= data_i[12];
    end 
    if(N4622) begin
      \nz.mem_1371_sv2v_reg  <= data_i[11];
    end 
    if(N4621) begin
      \nz.mem_1370_sv2v_reg  <= data_i[10];
    end 
    if(N4620) begin
      \nz.mem_1369_sv2v_reg  <= data_i[9];
    end 
    if(N4619) begin
      \nz.mem_1368_sv2v_reg  <= data_i[8];
    end 
    if(N4618) begin
      \nz.mem_1367_sv2v_reg  <= data_i[7];
    end 
    if(N4617) begin
      \nz.mem_1366_sv2v_reg  <= data_i[6];
    end 
    if(N4616) begin
      \nz.mem_1365_sv2v_reg  <= data_i[5];
    end 
    if(N4615) begin
      \nz.mem_1364_sv2v_reg  <= data_i[4];
    end 
    if(N4614) begin
      \nz.mem_1363_sv2v_reg  <= data_i[3];
    end 
    if(N4613) begin
      \nz.mem_1362_sv2v_reg  <= data_i[2];
    end 
    if(N4612) begin
      \nz.mem_1361_sv2v_reg  <= data_i[1];
    end 
    if(N4611) begin
      \nz.mem_1360_sv2v_reg  <= data_i[0];
    end 
    if(N4610) begin
      \nz.mem_1359_sv2v_reg  <= data_i[39];
    end 
    if(N4609) begin
      \nz.mem_1358_sv2v_reg  <= data_i[38];
    end 
    if(N4608) begin
      \nz.mem_1357_sv2v_reg  <= data_i[37];
    end 
    if(N4607) begin
      \nz.mem_1356_sv2v_reg  <= data_i[36];
    end 
    if(N4606) begin
      \nz.mem_1355_sv2v_reg  <= data_i[35];
    end 
    if(N4605) begin
      \nz.mem_1354_sv2v_reg  <= data_i[34];
    end 
    if(N4604) begin
      \nz.mem_1353_sv2v_reg  <= data_i[33];
    end 
    if(N4603) begin
      \nz.mem_1352_sv2v_reg  <= data_i[32];
    end 
    if(N4602) begin
      \nz.mem_1351_sv2v_reg  <= data_i[31];
    end 
    if(N4601) begin
      \nz.mem_1350_sv2v_reg  <= data_i[30];
    end 
    if(N4600) begin
      \nz.mem_1349_sv2v_reg  <= data_i[29];
    end 
    if(N4599) begin
      \nz.mem_1348_sv2v_reg  <= data_i[28];
    end 
    if(N4598) begin
      \nz.mem_1347_sv2v_reg  <= data_i[27];
    end 
    if(N4597) begin
      \nz.mem_1346_sv2v_reg  <= data_i[26];
    end 
    if(N4596) begin
      \nz.mem_1345_sv2v_reg  <= data_i[25];
    end 
    if(N4595) begin
      \nz.mem_1344_sv2v_reg  <= data_i[24];
    end 
    if(N4594) begin
      \nz.mem_1343_sv2v_reg  <= data_i[23];
    end 
    if(N4593) begin
      \nz.mem_1342_sv2v_reg  <= data_i[22];
    end 
    if(N4592) begin
      \nz.mem_1341_sv2v_reg  <= data_i[21];
    end 
    if(N4591) begin
      \nz.mem_1340_sv2v_reg  <= data_i[20];
    end 
    if(N4590) begin
      \nz.mem_1339_sv2v_reg  <= data_i[19];
    end 
    if(N4589) begin
      \nz.mem_1338_sv2v_reg  <= data_i[18];
    end 
    if(N4588) begin
      \nz.mem_1337_sv2v_reg  <= data_i[17];
    end 
    if(N4587) begin
      \nz.mem_1336_sv2v_reg  <= data_i[16];
    end 
    if(N4586) begin
      \nz.mem_1335_sv2v_reg  <= data_i[15];
    end 
    if(N4585) begin
      \nz.mem_1334_sv2v_reg  <= data_i[14];
    end 
    if(N4584) begin
      \nz.mem_1333_sv2v_reg  <= data_i[13];
    end 
    if(N4583) begin
      \nz.mem_1332_sv2v_reg  <= data_i[12];
    end 
    if(N4582) begin
      \nz.mem_1331_sv2v_reg  <= data_i[11];
    end 
    if(N4581) begin
      \nz.mem_1330_sv2v_reg  <= data_i[10];
    end 
    if(N4580) begin
      \nz.mem_1329_sv2v_reg  <= data_i[9];
    end 
    if(N4579) begin
      \nz.mem_1328_sv2v_reg  <= data_i[8];
    end 
    if(N4578) begin
      \nz.mem_1327_sv2v_reg  <= data_i[7];
    end 
    if(N4577) begin
      \nz.mem_1326_sv2v_reg  <= data_i[6];
    end 
    if(N4576) begin
      \nz.mem_1325_sv2v_reg  <= data_i[5];
    end 
    if(N4575) begin
      \nz.mem_1324_sv2v_reg  <= data_i[4];
    end 
    if(N4574) begin
      \nz.mem_1323_sv2v_reg  <= data_i[3];
    end 
    if(N4573) begin
      \nz.mem_1322_sv2v_reg  <= data_i[2];
    end 
    if(N4572) begin
      \nz.mem_1321_sv2v_reg  <= data_i[1];
    end 
    if(N4571) begin
      \nz.mem_1320_sv2v_reg  <= data_i[0];
    end 
    if(N4570) begin
      \nz.mem_1319_sv2v_reg  <= data_i[39];
    end 
    if(N4569) begin
      \nz.mem_1318_sv2v_reg  <= data_i[38];
    end 
    if(N4568) begin
      \nz.mem_1317_sv2v_reg  <= data_i[37];
    end 
    if(N4567) begin
      \nz.mem_1316_sv2v_reg  <= data_i[36];
    end 
    if(N4566) begin
      \nz.mem_1315_sv2v_reg  <= data_i[35];
    end 
    if(N4565) begin
      \nz.mem_1314_sv2v_reg  <= data_i[34];
    end 
    if(N4564) begin
      \nz.mem_1313_sv2v_reg  <= data_i[33];
    end 
    if(N4563) begin
      \nz.mem_1312_sv2v_reg  <= data_i[32];
    end 
    if(N4562) begin
      \nz.mem_1311_sv2v_reg  <= data_i[31];
    end 
    if(N4561) begin
      \nz.mem_1310_sv2v_reg  <= data_i[30];
    end 
    if(N4560) begin
      \nz.mem_1309_sv2v_reg  <= data_i[29];
    end 
    if(N4559) begin
      \nz.mem_1308_sv2v_reg  <= data_i[28];
    end 
    if(N4558) begin
      \nz.mem_1307_sv2v_reg  <= data_i[27];
    end 
    if(N4557) begin
      \nz.mem_1306_sv2v_reg  <= data_i[26];
    end 
    if(N4556) begin
      \nz.mem_1305_sv2v_reg  <= data_i[25];
    end 
    if(N4555) begin
      \nz.mem_1304_sv2v_reg  <= data_i[24];
    end 
    if(N4554) begin
      \nz.mem_1303_sv2v_reg  <= data_i[23];
    end 
    if(N4553) begin
      \nz.mem_1302_sv2v_reg  <= data_i[22];
    end 
    if(N4552) begin
      \nz.mem_1301_sv2v_reg  <= data_i[21];
    end 
    if(N4551) begin
      \nz.mem_1300_sv2v_reg  <= data_i[20];
    end 
    if(N4550) begin
      \nz.mem_1299_sv2v_reg  <= data_i[19];
    end 
    if(N4549) begin
      \nz.mem_1298_sv2v_reg  <= data_i[18];
    end 
    if(N4548) begin
      \nz.mem_1297_sv2v_reg  <= data_i[17];
    end 
    if(N4547) begin
      \nz.mem_1296_sv2v_reg  <= data_i[16];
    end 
    if(N4546) begin
      \nz.mem_1295_sv2v_reg  <= data_i[15];
    end 
    if(N4545) begin
      \nz.mem_1294_sv2v_reg  <= data_i[14];
    end 
    if(N4544) begin
      \nz.mem_1293_sv2v_reg  <= data_i[13];
    end 
    if(N4543) begin
      \nz.mem_1292_sv2v_reg  <= data_i[12];
    end 
    if(N4542) begin
      \nz.mem_1291_sv2v_reg  <= data_i[11];
    end 
    if(N4541) begin
      \nz.mem_1290_sv2v_reg  <= data_i[10];
    end 
    if(N4540) begin
      \nz.mem_1289_sv2v_reg  <= data_i[9];
    end 
    if(N4539) begin
      \nz.mem_1288_sv2v_reg  <= data_i[8];
    end 
    if(N4538) begin
      \nz.mem_1287_sv2v_reg  <= data_i[7];
    end 
    if(N4537) begin
      \nz.mem_1286_sv2v_reg  <= data_i[6];
    end 
    if(N4536) begin
      \nz.mem_1285_sv2v_reg  <= data_i[5];
    end 
    if(N4535) begin
      \nz.mem_1284_sv2v_reg  <= data_i[4];
    end 
    if(N4534) begin
      \nz.mem_1283_sv2v_reg  <= data_i[3];
    end 
    if(N4533) begin
      \nz.mem_1282_sv2v_reg  <= data_i[2];
    end 
    if(N4532) begin
      \nz.mem_1281_sv2v_reg  <= data_i[1];
    end 
    if(N4531) begin
      \nz.mem_1280_sv2v_reg  <= data_i[0];
    end 
    if(N4530) begin
      \nz.mem_1279_sv2v_reg  <= data_i[39];
    end 
    if(N4529) begin
      \nz.mem_1278_sv2v_reg  <= data_i[38];
    end 
    if(N4528) begin
      \nz.mem_1277_sv2v_reg  <= data_i[37];
    end 
    if(N4527) begin
      \nz.mem_1276_sv2v_reg  <= data_i[36];
    end 
    if(N4526) begin
      \nz.mem_1275_sv2v_reg  <= data_i[35];
    end 
    if(N4525) begin
      \nz.mem_1274_sv2v_reg  <= data_i[34];
    end 
    if(N4524) begin
      \nz.mem_1273_sv2v_reg  <= data_i[33];
    end 
    if(N4523) begin
      \nz.mem_1272_sv2v_reg  <= data_i[32];
    end 
    if(N4522) begin
      \nz.mem_1271_sv2v_reg  <= data_i[31];
    end 
    if(N4521) begin
      \nz.mem_1270_sv2v_reg  <= data_i[30];
    end 
    if(N4520) begin
      \nz.mem_1269_sv2v_reg  <= data_i[29];
    end 
    if(N4519) begin
      \nz.mem_1268_sv2v_reg  <= data_i[28];
    end 
    if(N4518) begin
      \nz.mem_1267_sv2v_reg  <= data_i[27];
    end 
    if(N4517) begin
      \nz.mem_1266_sv2v_reg  <= data_i[26];
    end 
    if(N4516) begin
      \nz.mem_1265_sv2v_reg  <= data_i[25];
    end 
    if(N4515) begin
      \nz.mem_1264_sv2v_reg  <= data_i[24];
    end 
    if(N4514) begin
      \nz.mem_1263_sv2v_reg  <= data_i[23];
    end 
    if(N4513) begin
      \nz.mem_1262_sv2v_reg  <= data_i[22];
    end 
    if(N4512) begin
      \nz.mem_1261_sv2v_reg  <= data_i[21];
    end 
    if(N4511) begin
      \nz.mem_1260_sv2v_reg  <= data_i[20];
    end 
    if(N4510) begin
      \nz.mem_1259_sv2v_reg  <= data_i[19];
    end 
    if(N4509) begin
      \nz.mem_1258_sv2v_reg  <= data_i[18];
    end 
    if(N4508) begin
      \nz.mem_1257_sv2v_reg  <= data_i[17];
    end 
    if(N4507) begin
      \nz.mem_1256_sv2v_reg  <= data_i[16];
    end 
    if(N4506) begin
      \nz.mem_1255_sv2v_reg  <= data_i[15];
    end 
    if(N4505) begin
      \nz.mem_1254_sv2v_reg  <= data_i[14];
    end 
    if(N4504) begin
      \nz.mem_1253_sv2v_reg  <= data_i[13];
    end 
    if(N4503) begin
      \nz.mem_1252_sv2v_reg  <= data_i[12];
    end 
    if(N4502) begin
      \nz.mem_1251_sv2v_reg  <= data_i[11];
    end 
    if(N4501) begin
      \nz.mem_1250_sv2v_reg  <= data_i[10];
    end 
    if(N4500) begin
      \nz.mem_1249_sv2v_reg  <= data_i[9];
    end 
    if(N4499) begin
      \nz.mem_1248_sv2v_reg  <= data_i[8];
    end 
    if(N4498) begin
      \nz.mem_1247_sv2v_reg  <= data_i[7];
    end 
    if(N4497) begin
      \nz.mem_1246_sv2v_reg  <= data_i[6];
    end 
    if(N4496) begin
      \nz.mem_1245_sv2v_reg  <= data_i[5];
    end 
    if(N4495) begin
      \nz.mem_1244_sv2v_reg  <= data_i[4];
    end 
    if(N4494) begin
      \nz.mem_1243_sv2v_reg  <= data_i[3];
    end 
    if(N4493) begin
      \nz.mem_1242_sv2v_reg  <= data_i[2];
    end 
    if(N4492) begin
      \nz.mem_1241_sv2v_reg  <= data_i[1];
    end 
    if(N4491) begin
      \nz.mem_1240_sv2v_reg  <= data_i[0];
    end 
    if(N4490) begin
      \nz.mem_1239_sv2v_reg  <= data_i[39];
    end 
    if(N4489) begin
      \nz.mem_1238_sv2v_reg  <= data_i[38];
    end 
    if(N4488) begin
      \nz.mem_1237_sv2v_reg  <= data_i[37];
    end 
    if(N4487) begin
      \nz.mem_1236_sv2v_reg  <= data_i[36];
    end 
    if(N4486) begin
      \nz.mem_1235_sv2v_reg  <= data_i[35];
    end 
    if(N4485) begin
      \nz.mem_1234_sv2v_reg  <= data_i[34];
    end 
    if(N4484) begin
      \nz.mem_1233_sv2v_reg  <= data_i[33];
    end 
    if(N4483) begin
      \nz.mem_1232_sv2v_reg  <= data_i[32];
    end 
    if(N4482) begin
      \nz.mem_1231_sv2v_reg  <= data_i[31];
    end 
    if(N4481) begin
      \nz.mem_1230_sv2v_reg  <= data_i[30];
    end 
    if(N4480) begin
      \nz.mem_1229_sv2v_reg  <= data_i[29];
    end 
    if(N4479) begin
      \nz.mem_1228_sv2v_reg  <= data_i[28];
    end 
    if(N4478) begin
      \nz.mem_1227_sv2v_reg  <= data_i[27];
    end 
    if(N4477) begin
      \nz.mem_1226_sv2v_reg  <= data_i[26];
    end 
    if(N4476) begin
      \nz.mem_1225_sv2v_reg  <= data_i[25];
    end 
    if(N4475) begin
      \nz.mem_1224_sv2v_reg  <= data_i[24];
    end 
    if(N4474) begin
      \nz.mem_1223_sv2v_reg  <= data_i[23];
    end 
    if(N4473) begin
      \nz.mem_1222_sv2v_reg  <= data_i[22];
    end 
    if(N4472) begin
      \nz.mem_1221_sv2v_reg  <= data_i[21];
    end 
    if(N4471) begin
      \nz.mem_1220_sv2v_reg  <= data_i[20];
    end 
    if(N4470) begin
      \nz.mem_1219_sv2v_reg  <= data_i[19];
    end 
    if(N4469) begin
      \nz.mem_1218_sv2v_reg  <= data_i[18];
    end 
    if(N4468) begin
      \nz.mem_1217_sv2v_reg  <= data_i[17];
    end 
    if(N4467) begin
      \nz.mem_1216_sv2v_reg  <= data_i[16];
    end 
    if(N4466) begin
      \nz.mem_1215_sv2v_reg  <= data_i[15];
    end 
    if(N4465) begin
      \nz.mem_1214_sv2v_reg  <= data_i[14];
    end 
    if(N4464) begin
      \nz.mem_1213_sv2v_reg  <= data_i[13];
    end 
    if(N4463) begin
      \nz.mem_1212_sv2v_reg  <= data_i[12];
    end 
    if(N4462) begin
      \nz.mem_1211_sv2v_reg  <= data_i[11];
    end 
    if(N4461) begin
      \nz.mem_1210_sv2v_reg  <= data_i[10];
    end 
    if(N4460) begin
      \nz.mem_1209_sv2v_reg  <= data_i[9];
    end 
    if(N4459) begin
      \nz.mem_1208_sv2v_reg  <= data_i[8];
    end 
    if(N4458) begin
      \nz.mem_1207_sv2v_reg  <= data_i[7];
    end 
    if(N4457) begin
      \nz.mem_1206_sv2v_reg  <= data_i[6];
    end 
    if(N4456) begin
      \nz.mem_1205_sv2v_reg  <= data_i[5];
    end 
    if(N4455) begin
      \nz.mem_1204_sv2v_reg  <= data_i[4];
    end 
    if(N4454) begin
      \nz.mem_1203_sv2v_reg  <= data_i[3];
    end 
    if(N4453) begin
      \nz.mem_1202_sv2v_reg  <= data_i[2];
    end 
    if(N4452) begin
      \nz.mem_1201_sv2v_reg  <= data_i[1];
    end 
    if(N4451) begin
      \nz.mem_1200_sv2v_reg  <= data_i[0];
    end 
    if(N4450) begin
      \nz.mem_1199_sv2v_reg  <= data_i[39];
    end 
    if(N4449) begin
      \nz.mem_1198_sv2v_reg  <= data_i[38];
    end 
    if(N4448) begin
      \nz.mem_1197_sv2v_reg  <= data_i[37];
    end 
    if(N4447) begin
      \nz.mem_1196_sv2v_reg  <= data_i[36];
    end 
    if(N4446) begin
      \nz.mem_1195_sv2v_reg  <= data_i[35];
    end 
    if(N4445) begin
      \nz.mem_1194_sv2v_reg  <= data_i[34];
    end 
    if(N4444) begin
      \nz.mem_1193_sv2v_reg  <= data_i[33];
    end 
    if(N4443) begin
      \nz.mem_1192_sv2v_reg  <= data_i[32];
    end 
    if(N4442) begin
      \nz.mem_1191_sv2v_reg  <= data_i[31];
    end 
    if(N4441) begin
      \nz.mem_1190_sv2v_reg  <= data_i[30];
    end 
    if(N4440) begin
      \nz.mem_1189_sv2v_reg  <= data_i[29];
    end 
    if(N4439) begin
      \nz.mem_1188_sv2v_reg  <= data_i[28];
    end 
    if(N4438) begin
      \nz.mem_1187_sv2v_reg  <= data_i[27];
    end 
    if(N4437) begin
      \nz.mem_1186_sv2v_reg  <= data_i[26];
    end 
    if(N4436) begin
      \nz.mem_1185_sv2v_reg  <= data_i[25];
    end 
    if(N4435) begin
      \nz.mem_1184_sv2v_reg  <= data_i[24];
    end 
    if(N4434) begin
      \nz.mem_1183_sv2v_reg  <= data_i[23];
    end 
    if(N4433) begin
      \nz.mem_1182_sv2v_reg  <= data_i[22];
    end 
    if(N4432) begin
      \nz.mem_1181_sv2v_reg  <= data_i[21];
    end 
    if(N4431) begin
      \nz.mem_1180_sv2v_reg  <= data_i[20];
    end 
    if(N4430) begin
      \nz.mem_1179_sv2v_reg  <= data_i[19];
    end 
    if(N4429) begin
      \nz.mem_1178_sv2v_reg  <= data_i[18];
    end 
    if(N4428) begin
      \nz.mem_1177_sv2v_reg  <= data_i[17];
    end 
    if(N4427) begin
      \nz.mem_1176_sv2v_reg  <= data_i[16];
    end 
    if(N4426) begin
      \nz.mem_1175_sv2v_reg  <= data_i[15];
    end 
    if(N4425) begin
      \nz.mem_1174_sv2v_reg  <= data_i[14];
    end 
    if(N4424) begin
      \nz.mem_1173_sv2v_reg  <= data_i[13];
    end 
    if(N4423) begin
      \nz.mem_1172_sv2v_reg  <= data_i[12];
    end 
    if(N4422) begin
      \nz.mem_1171_sv2v_reg  <= data_i[11];
    end 
    if(N4421) begin
      \nz.mem_1170_sv2v_reg  <= data_i[10];
    end 
    if(N4420) begin
      \nz.mem_1169_sv2v_reg  <= data_i[9];
    end 
    if(N4419) begin
      \nz.mem_1168_sv2v_reg  <= data_i[8];
    end 
    if(N4418) begin
      \nz.mem_1167_sv2v_reg  <= data_i[7];
    end 
    if(N4417) begin
      \nz.mem_1166_sv2v_reg  <= data_i[6];
    end 
    if(N4416) begin
      \nz.mem_1165_sv2v_reg  <= data_i[5];
    end 
    if(N4415) begin
      \nz.mem_1164_sv2v_reg  <= data_i[4];
    end 
    if(N4414) begin
      \nz.mem_1163_sv2v_reg  <= data_i[3];
    end 
    if(N4413) begin
      \nz.mem_1162_sv2v_reg  <= data_i[2];
    end 
    if(N4412) begin
      \nz.mem_1161_sv2v_reg  <= data_i[1];
    end 
    if(N4411) begin
      \nz.mem_1160_sv2v_reg  <= data_i[0];
    end 
    if(N4410) begin
      \nz.mem_1159_sv2v_reg  <= data_i[39];
    end 
    if(N4409) begin
      \nz.mem_1158_sv2v_reg  <= data_i[38];
    end 
    if(N4408) begin
      \nz.mem_1157_sv2v_reg  <= data_i[37];
    end 
    if(N4407) begin
      \nz.mem_1156_sv2v_reg  <= data_i[36];
    end 
    if(N4406) begin
      \nz.mem_1155_sv2v_reg  <= data_i[35];
    end 
    if(N4405) begin
      \nz.mem_1154_sv2v_reg  <= data_i[34];
    end 
    if(N4404) begin
      \nz.mem_1153_sv2v_reg  <= data_i[33];
    end 
    if(N4403) begin
      \nz.mem_1152_sv2v_reg  <= data_i[32];
    end 
    if(N4402) begin
      \nz.mem_1151_sv2v_reg  <= data_i[31];
    end 
    if(N4401) begin
      \nz.mem_1150_sv2v_reg  <= data_i[30];
    end 
    if(N4400) begin
      \nz.mem_1149_sv2v_reg  <= data_i[29];
    end 
    if(N4399) begin
      \nz.mem_1148_sv2v_reg  <= data_i[28];
    end 
    if(N4398) begin
      \nz.mem_1147_sv2v_reg  <= data_i[27];
    end 
    if(N4397) begin
      \nz.mem_1146_sv2v_reg  <= data_i[26];
    end 
    if(N4396) begin
      \nz.mem_1145_sv2v_reg  <= data_i[25];
    end 
    if(N4395) begin
      \nz.mem_1144_sv2v_reg  <= data_i[24];
    end 
    if(N4394) begin
      \nz.mem_1143_sv2v_reg  <= data_i[23];
    end 
    if(N4393) begin
      \nz.mem_1142_sv2v_reg  <= data_i[22];
    end 
    if(N4392) begin
      \nz.mem_1141_sv2v_reg  <= data_i[21];
    end 
    if(N4391) begin
      \nz.mem_1140_sv2v_reg  <= data_i[20];
    end 
    if(N4390) begin
      \nz.mem_1139_sv2v_reg  <= data_i[19];
    end 
    if(N4389) begin
      \nz.mem_1138_sv2v_reg  <= data_i[18];
    end 
    if(N4388) begin
      \nz.mem_1137_sv2v_reg  <= data_i[17];
    end 
    if(N4387) begin
      \nz.mem_1136_sv2v_reg  <= data_i[16];
    end 
    if(N4386) begin
      \nz.mem_1135_sv2v_reg  <= data_i[15];
    end 
    if(N4385) begin
      \nz.mem_1134_sv2v_reg  <= data_i[14];
    end 
    if(N4384) begin
      \nz.mem_1133_sv2v_reg  <= data_i[13];
    end 
    if(N4383) begin
      \nz.mem_1132_sv2v_reg  <= data_i[12];
    end 
    if(N4382) begin
      \nz.mem_1131_sv2v_reg  <= data_i[11];
    end 
    if(N4381) begin
      \nz.mem_1130_sv2v_reg  <= data_i[10];
    end 
    if(N4380) begin
      \nz.mem_1129_sv2v_reg  <= data_i[9];
    end 
    if(N4379) begin
      \nz.mem_1128_sv2v_reg  <= data_i[8];
    end 
    if(N4378) begin
      \nz.mem_1127_sv2v_reg  <= data_i[7];
    end 
    if(N4377) begin
      \nz.mem_1126_sv2v_reg  <= data_i[6];
    end 
    if(N4376) begin
      \nz.mem_1125_sv2v_reg  <= data_i[5];
    end 
    if(N4375) begin
      \nz.mem_1124_sv2v_reg  <= data_i[4];
    end 
    if(N4374) begin
      \nz.mem_1123_sv2v_reg  <= data_i[3];
    end 
    if(N4373) begin
      \nz.mem_1122_sv2v_reg  <= data_i[2];
    end 
    if(N4372) begin
      \nz.mem_1121_sv2v_reg  <= data_i[1];
    end 
    if(N4371) begin
      \nz.mem_1120_sv2v_reg  <= data_i[0];
    end 
    if(N4370) begin
      \nz.mem_1119_sv2v_reg  <= data_i[39];
    end 
    if(N4369) begin
      \nz.mem_1118_sv2v_reg  <= data_i[38];
    end 
    if(N4368) begin
      \nz.mem_1117_sv2v_reg  <= data_i[37];
    end 
    if(N4367) begin
      \nz.mem_1116_sv2v_reg  <= data_i[36];
    end 
    if(N4366) begin
      \nz.mem_1115_sv2v_reg  <= data_i[35];
    end 
    if(N4365) begin
      \nz.mem_1114_sv2v_reg  <= data_i[34];
    end 
    if(N4364) begin
      \nz.mem_1113_sv2v_reg  <= data_i[33];
    end 
    if(N4363) begin
      \nz.mem_1112_sv2v_reg  <= data_i[32];
    end 
    if(N4362) begin
      \nz.mem_1111_sv2v_reg  <= data_i[31];
    end 
    if(N4361) begin
      \nz.mem_1110_sv2v_reg  <= data_i[30];
    end 
    if(N4360) begin
      \nz.mem_1109_sv2v_reg  <= data_i[29];
    end 
    if(N4359) begin
      \nz.mem_1108_sv2v_reg  <= data_i[28];
    end 
    if(N4358) begin
      \nz.mem_1107_sv2v_reg  <= data_i[27];
    end 
    if(N4357) begin
      \nz.mem_1106_sv2v_reg  <= data_i[26];
    end 
    if(N4356) begin
      \nz.mem_1105_sv2v_reg  <= data_i[25];
    end 
    if(N4355) begin
      \nz.mem_1104_sv2v_reg  <= data_i[24];
    end 
    if(N4354) begin
      \nz.mem_1103_sv2v_reg  <= data_i[23];
    end 
    if(N4353) begin
      \nz.mem_1102_sv2v_reg  <= data_i[22];
    end 
    if(N4352) begin
      \nz.mem_1101_sv2v_reg  <= data_i[21];
    end 
    if(N4351) begin
      \nz.mem_1100_sv2v_reg  <= data_i[20];
    end 
    if(N4350) begin
      \nz.mem_1099_sv2v_reg  <= data_i[19];
    end 
    if(N4349) begin
      \nz.mem_1098_sv2v_reg  <= data_i[18];
    end 
    if(N4348) begin
      \nz.mem_1097_sv2v_reg  <= data_i[17];
    end 
    if(N4347) begin
      \nz.mem_1096_sv2v_reg  <= data_i[16];
    end 
    if(N4346) begin
      \nz.mem_1095_sv2v_reg  <= data_i[15];
    end 
    if(N4345) begin
      \nz.mem_1094_sv2v_reg  <= data_i[14];
    end 
    if(N4344) begin
      \nz.mem_1093_sv2v_reg  <= data_i[13];
    end 
    if(N4343) begin
      \nz.mem_1092_sv2v_reg  <= data_i[12];
    end 
    if(N4342) begin
      \nz.mem_1091_sv2v_reg  <= data_i[11];
    end 
    if(N4341) begin
      \nz.mem_1090_sv2v_reg  <= data_i[10];
    end 
    if(N4340) begin
      \nz.mem_1089_sv2v_reg  <= data_i[9];
    end 
    if(N4339) begin
      \nz.mem_1088_sv2v_reg  <= data_i[8];
    end 
    if(N4338) begin
      \nz.mem_1087_sv2v_reg  <= data_i[7];
    end 
    if(N4337) begin
      \nz.mem_1086_sv2v_reg  <= data_i[6];
    end 
    if(N4336) begin
      \nz.mem_1085_sv2v_reg  <= data_i[5];
    end 
    if(N4335) begin
      \nz.mem_1084_sv2v_reg  <= data_i[4];
    end 
    if(N4334) begin
      \nz.mem_1083_sv2v_reg  <= data_i[3];
    end 
    if(N4333) begin
      \nz.mem_1082_sv2v_reg  <= data_i[2];
    end 
    if(N4332) begin
      \nz.mem_1081_sv2v_reg  <= data_i[1];
    end 
    if(N4331) begin
      \nz.mem_1080_sv2v_reg  <= data_i[0];
    end 
    if(N4330) begin
      \nz.mem_1079_sv2v_reg  <= data_i[39];
    end 
    if(N4329) begin
      \nz.mem_1078_sv2v_reg  <= data_i[38];
    end 
    if(N4328) begin
      \nz.mem_1077_sv2v_reg  <= data_i[37];
    end 
    if(N4327) begin
      \nz.mem_1076_sv2v_reg  <= data_i[36];
    end 
    if(N4326) begin
      \nz.mem_1075_sv2v_reg  <= data_i[35];
    end 
    if(N4325) begin
      \nz.mem_1074_sv2v_reg  <= data_i[34];
    end 
    if(N4324) begin
      \nz.mem_1073_sv2v_reg  <= data_i[33];
    end 
    if(N4323) begin
      \nz.mem_1072_sv2v_reg  <= data_i[32];
    end 
    if(N4322) begin
      \nz.mem_1071_sv2v_reg  <= data_i[31];
    end 
    if(N4321) begin
      \nz.mem_1070_sv2v_reg  <= data_i[30];
    end 
    if(N4320) begin
      \nz.mem_1069_sv2v_reg  <= data_i[29];
    end 
    if(N4319) begin
      \nz.mem_1068_sv2v_reg  <= data_i[28];
    end 
    if(N4318) begin
      \nz.mem_1067_sv2v_reg  <= data_i[27];
    end 
    if(N4317) begin
      \nz.mem_1066_sv2v_reg  <= data_i[26];
    end 
    if(N4316) begin
      \nz.mem_1065_sv2v_reg  <= data_i[25];
    end 
    if(N4315) begin
      \nz.mem_1064_sv2v_reg  <= data_i[24];
    end 
    if(N4314) begin
      \nz.mem_1063_sv2v_reg  <= data_i[23];
    end 
    if(N4313) begin
      \nz.mem_1062_sv2v_reg  <= data_i[22];
    end 
    if(N4312) begin
      \nz.mem_1061_sv2v_reg  <= data_i[21];
    end 
    if(N4311) begin
      \nz.mem_1060_sv2v_reg  <= data_i[20];
    end 
    if(N4310) begin
      \nz.mem_1059_sv2v_reg  <= data_i[19];
    end 
    if(N4309) begin
      \nz.mem_1058_sv2v_reg  <= data_i[18];
    end 
    if(N4308) begin
      \nz.mem_1057_sv2v_reg  <= data_i[17];
    end 
    if(N4307) begin
      \nz.mem_1056_sv2v_reg  <= data_i[16];
    end 
    if(N4306) begin
      \nz.mem_1055_sv2v_reg  <= data_i[15];
    end 
    if(N4305) begin
      \nz.mem_1054_sv2v_reg  <= data_i[14];
    end 
    if(N4304) begin
      \nz.mem_1053_sv2v_reg  <= data_i[13];
    end 
    if(N4303) begin
      \nz.mem_1052_sv2v_reg  <= data_i[12];
    end 
    if(N4302) begin
      \nz.mem_1051_sv2v_reg  <= data_i[11];
    end 
    if(N4301) begin
      \nz.mem_1050_sv2v_reg  <= data_i[10];
    end 
    if(N4300) begin
      \nz.mem_1049_sv2v_reg  <= data_i[9];
    end 
    if(N4299) begin
      \nz.mem_1048_sv2v_reg  <= data_i[8];
    end 
    if(N4298) begin
      \nz.mem_1047_sv2v_reg  <= data_i[7];
    end 
    if(N4297) begin
      \nz.mem_1046_sv2v_reg  <= data_i[6];
    end 
    if(N4296) begin
      \nz.mem_1045_sv2v_reg  <= data_i[5];
    end 
    if(N4295) begin
      \nz.mem_1044_sv2v_reg  <= data_i[4];
    end 
    if(N4294) begin
      \nz.mem_1043_sv2v_reg  <= data_i[3];
    end 
    if(N4293) begin
      \nz.mem_1042_sv2v_reg  <= data_i[2];
    end 
    if(N4292) begin
      \nz.mem_1041_sv2v_reg  <= data_i[1];
    end 
    if(N4291) begin
      \nz.mem_1040_sv2v_reg  <= data_i[0];
    end 
    if(N4290) begin
      \nz.mem_1039_sv2v_reg  <= data_i[39];
    end 
    if(N4289) begin
      \nz.mem_1038_sv2v_reg  <= data_i[38];
    end 
    if(N4288) begin
      \nz.mem_1037_sv2v_reg  <= data_i[37];
    end 
    if(N4287) begin
      \nz.mem_1036_sv2v_reg  <= data_i[36];
    end 
    if(N4286) begin
      \nz.mem_1035_sv2v_reg  <= data_i[35];
    end 
    if(N4285) begin
      \nz.mem_1034_sv2v_reg  <= data_i[34];
    end 
    if(N4284) begin
      \nz.mem_1033_sv2v_reg  <= data_i[33];
    end 
    if(N4283) begin
      \nz.mem_1032_sv2v_reg  <= data_i[32];
    end 
    if(N4282) begin
      \nz.mem_1031_sv2v_reg  <= data_i[31];
    end 
    if(N4281) begin
      \nz.mem_1030_sv2v_reg  <= data_i[30];
    end 
    if(N4280) begin
      \nz.mem_1029_sv2v_reg  <= data_i[29];
    end 
    if(N4279) begin
      \nz.mem_1028_sv2v_reg  <= data_i[28];
    end 
    if(N4278) begin
      \nz.mem_1027_sv2v_reg  <= data_i[27];
    end 
    if(N4277) begin
      \nz.mem_1026_sv2v_reg  <= data_i[26];
    end 
    if(N4276) begin
      \nz.mem_1025_sv2v_reg  <= data_i[25];
    end 
    if(N4275) begin
      \nz.mem_1024_sv2v_reg  <= data_i[24];
    end 
    if(N4274) begin
      \nz.mem_1023_sv2v_reg  <= data_i[23];
    end 
    if(N4273) begin
      \nz.mem_1022_sv2v_reg  <= data_i[22];
    end 
    if(N4272) begin
      \nz.mem_1021_sv2v_reg  <= data_i[21];
    end 
    if(N4271) begin
      \nz.mem_1020_sv2v_reg  <= data_i[20];
    end 
    if(N4270) begin
      \nz.mem_1019_sv2v_reg  <= data_i[19];
    end 
    if(N4269) begin
      \nz.mem_1018_sv2v_reg  <= data_i[18];
    end 
    if(N4268) begin
      \nz.mem_1017_sv2v_reg  <= data_i[17];
    end 
    if(N4267) begin
      \nz.mem_1016_sv2v_reg  <= data_i[16];
    end 
    if(N4266) begin
      \nz.mem_1015_sv2v_reg  <= data_i[15];
    end 
    if(N4265) begin
      \nz.mem_1014_sv2v_reg  <= data_i[14];
    end 
    if(N4264) begin
      \nz.mem_1013_sv2v_reg  <= data_i[13];
    end 
    if(N4263) begin
      \nz.mem_1012_sv2v_reg  <= data_i[12];
    end 
    if(N4262) begin
      \nz.mem_1011_sv2v_reg  <= data_i[11];
    end 
    if(N4261) begin
      \nz.mem_1010_sv2v_reg  <= data_i[10];
    end 
    if(N4260) begin
      \nz.mem_1009_sv2v_reg  <= data_i[9];
    end 
    if(N4259) begin
      \nz.mem_1008_sv2v_reg  <= data_i[8];
    end 
    if(N4258) begin
      \nz.mem_1007_sv2v_reg  <= data_i[7];
    end 
    if(N4257) begin
      \nz.mem_1006_sv2v_reg  <= data_i[6];
    end 
    if(N4256) begin
      \nz.mem_1005_sv2v_reg  <= data_i[5];
    end 
    if(N4255) begin
      \nz.mem_1004_sv2v_reg  <= data_i[4];
    end 
    if(N4254) begin
      \nz.mem_1003_sv2v_reg  <= data_i[3];
    end 
    if(N4253) begin
      \nz.mem_1002_sv2v_reg  <= data_i[2];
    end 
    if(N4252) begin
      \nz.mem_1001_sv2v_reg  <= data_i[1];
    end 
    if(N4251) begin
      \nz.mem_1000_sv2v_reg  <= data_i[0];
    end 
    if(N4250) begin
      \nz.mem_999_sv2v_reg  <= data_i[39];
    end 
    if(N4249) begin
      \nz.mem_998_sv2v_reg  <= data_i[38];
    end 
    if(N4248) begin
      \nz.mem_997_sv2v_reg  <= data_i[37];
    end 
    if(N4247) begin
      \nz.mem_996_sv2v_reg  <= data_i[36];
    end 
    if(N4246) begin
      \nz.mem_995_sv2v_reg  <= data_i[35];
    end 
    if(N4245) begin
      \nz.mem_994_sv2v_reg  <= data_i[34];
    end 
    if(N4244) begin
      \nz.mem_993_sv2v_reg  <= data_i[33];
    end 
    if(N4243) begin
      \nz.mem_992_sv2v_reg  <= data_i[32];
    end 
    if(N4242) begin
      \nz.mem_991_sv2v_reg  <= data_i[31];
    end 
    if(N4241) begin
      \nz.mem_990_sv2v_reg  <= data_i[30];
    end 
    if(N4240) begin
      \nz.mem_989_sv2v_reg  <= data_i[29];
    end 
    if(N4239) begin
      \nz.mem_988_sv2v_reg  <= data_i[28];
    end 
    if(N4238) begin
      \nz.mem_987_sv2v_reg  <= data_i[27];
    end 
    if(N4237) begin
      \nz.mem_986_sv2v_reg  <= data_i[26];
    end 
    if(N4236) begin
      \nz.mem_985_sv2v_reg  <= data_i[25];
    end 
    if(N4235) begin
      \nz.mem_984_sv2v_reg  <= data_i[24];
    end 
    if(N4234) begin
      \nz.mem_983_sv2v_reg  <= data_i[23];
    end 
    if(N4233) begin
      \nz.mem_982_sv2v_reg  <= data_i[22];
    end 
    if(N4232) begin
      \nz.mem_981_sv2v_reg  <= data_i[21];
    end 
    if(N4231) begin
      \nz.mem_980_sv2v_reg  <= data_i[20];
    end 
    if(N4230) begin
      \nz.mem_979_sv2v_reg  <= data_i[19];
    end 
    if(N4229) begin
      \nz.mem_978_sv2v_reg  <= data_i[18];
    end 
    if(N4228) begin
      \nz.mem_977_sv2v_reg  <= data_i[17];
    end 
    if(N4227) begin
      \nz.mem_976_sv2v_reg  <= data_i[16];
    end 
    if(N4226) begin
      \nz.mem_975_sv2v_reg  <= data_i[15];
    end 
    if(N4225) begin
      \nz.mem_974_sv2v_reg  <= data_i[14];
    end 
    if(N4224) begin
      \nz.mem_973_sv2v_reg  <= data_i[13];
    end 
    if(N4223) begin
      \nz.mem_972_sv2v_reg  <= data_i[12];
    end 
    if(N4222) begin
      \nz.mem_971_sv2v_reg  <= data_i[11];
    end 
    if(N4221) begin
      \nz.mem_970_sv2v_reg  <= data_i[10];
    end 
    if(N4220) begin
      \nz.mem_969_sv2v_reg  <= data_i[9];
    end 
    if(N4219) begin
      \nz.mem_968_sv2v_reg  <= data_i[8];
    end 
    if(N4218) begin
      \nz.mem_967_sv2v_reg  <= data_i[7];
    end 
    if(N4217) begin
      \nz.mem_966_sv2v_reg  <= data_i[6];
    end 
    if(N4216) begin
      \nz.mem_965_sv2v_reg  <= data_i[5];
    end 
    if(N4215) begin
      \nz.mem_964_sv2v_reg  <= data_i[4];
    end 
    if(N4214) begin
      \nz.mem_963_sv2v_reg  <= data_i[3];
    end 
    if(N4213) begin
      \nz.mem_962_sv2v_reg  <= data_i[2];
    end 
    if(N4212) begin
      \nz.mem_961_sv2v_reg  <= data_i[1];
    end 
    if(N4211) begin
      \nz.mem_960_sv2v_reg  <= data_i[0];
    end 
    if(N4210) begin
      \nz.mem_959_sv2v_reg  <= data_i[39];
    end 
    if(N4209) begin
      \nz.mem_958_sv2v_reg  <= data_i[38];
    end 
    if(N4208) begin
      \nz.mem_957_sv2v_reg  <= data_i[37];
    end 
    if(N4207) begin
      \nz.mem_956_sv2v_reg  <= data_i[36];
    end 
    if(N4206) begin
      \nz.mem_955_sv2v_reg  <= data_i[35];
    end 
    if(N4205) begin
      \nz.mem_954_sv2v_reg  <= data_i[34];
    end 
    if(N4204) begin
      \nz.mem_953_sv2v_reg  <= data_i[33];
    end 
    if(N4203) begin
      \nz.mem_952_sv2v_reg  <= data_i[32];
    end 
    if(N4202) begin
      \nz.mem_951_sv2v_reg  <= data_i[31];
    end 
    if(N4201) begin
      \nz.mem_950_sv2v_reg  <= data_i[30];
    end 
    if(N4200) begin
      \nz.mem_949_sv2v_reg  <= data_i[29];
    end 
    if(N4199) begin
      \nz.mem_948_sv2v_reg  <= data_i[28];
    end 
    if(N4198) begin
      \nz.mem_947_sv2v_reg  <= data_i[27];
    end 
    if(N4197) begin
      \nz.mem_946_sv2v_reg  <= data_i[26];
    end 
    if(N4196) begin
      \nz.mem_945_sv2v_reg  <= data_i[25];
    end 
    if(N4195) begin
      \nz.mem_944_sv2v_reg  <= data_i[24];
    end 
    if(N4194) begin
      \nz.mem_943_sv2v_reg  <= data_i[23];
    end 
    if(N4193) begin
      \nz.mem_942_sv2v_reg  <= data_i[22];
    end 
    if(N4192) begin
      \nz.mem_941_sv2v_reg  <= data_i[21];
    end 
    if(N4191) begin
      \nz.mem_940_sv2v_reg  <= data_i[20];
    end 
    if(N4190) begin
      \nz.mem_939_sv2v_reg  <= data_i[19];
    end 
    if(N4189) begin
      \nz.mem_938_sv2v_reg  <= data_i[18];
    end 
    if(N4188) begin
      \nz.mem_937_sv2v_reg  <= data_i[17];
    end 
    if(N4187) begin
      \nz.mem_936_sv2v_reg  <= data_i[16];
    end 
    if(N4186) begin
      \nz.mem_935_sv2v_reg  <= data_i[15];
    end 
    if(N4185) begin
      \nz.mem_934_sv2v_reg  <= data_i[14];
    end 
    if(N4184) begin
      \nz.mem_933_sv2v_reg  <= data_i[13];
    end 
    if(N4183) begin
      \nz.mem_932_sv2v_reg  <= data_i[12];
    end 
    if(N4182) begin
      \nz.mem_931_sv2v_reg  <= data_i[11];
    end 
    if(N4181) begin
      \nz.mem_930_sv2v_reg  <= data_i[10];
    end 
    if(N4180) begin
      \nz.mem_929_sv2v_reg  <= data_i[9];
    end 
    if(N4179) begin
      \nz.mem_928_sv2v_reg  <= data_i[8];
    end 
    if(N4178) begin
      \nz.mem_927_sv2v_reg  <= data_i[7];
    end 
    if(N4177) begin
      \nz.mem_926_sv2v_reg  <= data_i[6];
    end 
    if(N4176) begin
      \nz.mem_925_sv2v_reg  <= data_i[5];
    end 
    if(N4175) begin
      \nz.mem_924_sv2v_reg  <= data_i[4];
    end 
    if(N4174) begin
      \nz.mem_923_sv2v_reg  <= data_i[3];
    end 
    if(N4173) begin
      \nz.mem_922_sv2v_reg  <= data_i[2];
    end 
    if(N4172) begin
      \nz.mem_921_sv2v_reg  <= data_i[1];
    end 
    if(N4171) begin
      \nz.mem_920_sv2v_reg  <= data_i[0];
    end 
    if(N4170) begin
      \nz.mem_919_sv2v_reg  <= data_i[39];
    end 
    if(N4169) begin
      \nz.mem_918_sv2v_reg  <= data_i[38];
    end 
    if(N4168) begin
      \nz.mem_917_sv2v_reg  <= data_i[37];
    end 
    if(N4167) begin
      \nz.mem_916_sv2v_reg  <= data_i[36];
    end 
    if(N4166) begin
      \nz.mem_915_sv2v_reg  <= data_i[35];
    end 
    if(N4165) begin
      \nz.mem_914_sv2v_reg  <= data_i[34];
    end 
    if(N4164) begin
      \nz.mem_913_sv2v_reg  <= data_i[33];
    end 
    if(N4163) begin
      \nz.mem_912_sv2v_reg  <= data_i[32];
    end 
    if(N4162) begin
      \nz.mem_911_sv2v_reg  <= data_i[31];
    end 
    if(N4161) begin
      \nz.mem_910_sv2v_reg  <= data_i[30];
    end 
    if(N4160) begin
      \nz.mem_909_sv2v_reg  <= data_i[29];
    end 
    if(N4159) begin
      \nz.mem_908_sv2v_reg  <= data_i[28];
    end 
    if(N4158) begin
      \nz.mem_907_sv2v_reg  <= data_i[27];
    end 
    if(N4157) begin
      \nz.mem_906_sv2v_reg  <= data_i[26];
    end 
    if(N4156) begin
      \nz.mem_905_sv2v_reg  <= data_i[25];
    end 
    if(N4155) begin
      \nz.mem_904_sv2v_reg  <= data_i[24];
    end 
    if(N4154) begin
      \nz.mem_903_sv2v_reg  <= data_i[23];
    end 
    if(N4153) begin
      \nz.mem_902_sv2v_reg  <= data_i[22];
    end 
    if(N4152) begin
      \nz.mem_901_sv2v_reg  <= data_i[21];
    end 
    if(N4151) begin
      \nz.mem_900_sv2v_reg  <= data_i[20];
    end 
    if(N4150) begin
      \nz.mem_899_sv2v_reg  <= data_i[19];
    end 
    if(N4149) begin
      \nz.mem_898_sv2v_reg  <= data_i[18];
    end 
    if(N4148) begin
      \nz.mem_897_sv2v_reg  <= data_i[17];
    end 
    if(N4147) begin
      \nz.mem_896_sv2v_reg  <= data_i[16];
    end 
    if(N4146) begin
      \nz.mem_895_sv2v_reg  <= data_i[15];
    end 
    if(N4145) begin
      \nz.mem_894_sv2v_reg  <= data_i[14];
    end 
    if(N4144) begin
      \nz.mem_893_sv2v_reg  <= data_i[13];
    end 
    if(N4143) begin
      \nz.mem_892_sv2v_reg  <= data_i[12];
    end 
    if(N4142) begin
      \nz.mem_891_sv2v_reg  <= data_i[11];
    end 
    if(N4141) begin
      \nz.mem_890_sv2v_reg  <= data_i[10];
    end 
    if(N4140) begin
      \nz.mem_889_sv2v_reg  <= data_i[9];
    end 
    if(N4139) begin
      \nz.mem_888_sv2v_reg  <= data_i[8];
    end 
    if(N4138) begin
      \nz.mem_887_sv2v_reg  <= data_i[7];
    end 
    if(N4137) begin
      \nz.mem_886_sv2v_reg  <= data_i[6];
    end 
    if(N4136) begin
      \nz.mem_885_sv2v_reg  <= data_i[5];
    end 
    if(N4135) begin
      \nz.mem_884_sv2v_reg  <= data_i[4];
    end 
    if(N4134) begin
      \nz.mem_883_sv2v_reg  <= data_i[3];
    end 
    if(N4133) begin
      \nz.mem_882_sv2v_reg  <= data_i[2];
    end 
    if(N4132) begin
      \nz.mem_881_sv2v_reg  <= data_i[1];
    end 
    if(N4131) begin
      \nz.mem_880_sv2v_reg  <= data_i[0];
    end 
    if(N4130) begin
      \nz.mem_879_sv2v_reg  <= data_i[39];
    end 
    if(N4129) begin
      \nz.mem_878_sv2v_reg  <= data_i[38];
    end 
    if(N4128) begin
      \nz.mem_877_sv2v_reg  <= data_i[37];
    end 
    if(N4127) begin
      \nz.mem_876_sv2v_reg  <= data_i[36];
    end 
    if(N4126) begin
      \nz.mem_875_sv2v_reg  <= data_i[35];
    end 
    if(N4125) begin
      \nz.mem_874_sv2v_reg  <= data_i[34];
    end 
    if(N4124) begin
      \nz.mem_873_sv2v_reg  <= data_i[33];
    end 
    if(N4123) begin
      \nz.mem_872_sv2v_reg  <= data_i[32];
    end 
    if(N4122) begin
      \nz.mem_871_sv2v_reg  <= data_i[31];
    end 
    if(N4121) begin
      \nz.mem_870_sv2v_reg  <= data_i[30];
    end 
    if(N4120) begin
      \nz.mem_869_sv2v_reg  <= data_i[29];
    end 
    if(N4119) begin
      \nz.mem_868_sv2v_reg  <= data_i[28];
    end 
    if(N4118) begin
      \nz.mem_867_sv2v_reg  <= data_i[27];
    end 
    if(N4117) begin
      \nz.mem_866_sv2v_reg  <= data_i[26];
    end 
    if(N4116) begin
      \nz.mem_865_sv2v_reg  <= data_i[25];
    end 
    if(N4115) begin
      \nz.mem_864_sv2v_reg  <= data_i[24];
    end 
    if(N4114) begin
      \nz.mem_863_sv2v_reg  <= data_i[23];
    end 
    if(N4113) begin
      \nz.mem_862_sv2v_reg  <= data_i[22];
    end 
    if(N4112) begin
      \nz.mem_861_sv2v_reg  <= data_i[21];
    end 
    if(N4111) begin
      \nz.mem_860_sv2v_reg  <= data_i[20];
    end 
    if(N4110) begin
      \nz.mem_859_sv2v_reg  <= data_i[19];
    end 
    if(N4109) begin
      \nz.mem_858_sv2v_reg  <= data_i[18];
    end 
    if(N4108) begin
      \nz.mem_857_sv2v_reg  <= data_i[17];
    end 
    if(N4107) begin
      \nz.mem_856_sv2v_reg  <= data_i[16];
    end 
    if(N4106) begin
      \nz.mem_855_sv2v_reg  <= data_i[15];
    end 
    if(N4105) begin
      \nz.mem_854_sv2v_reg  <= data_i[14];
    end 
    if(N4104) begin
      \nz.mem_853_sv2v_reg  <= data_i[13];
    end 
    if(N4103) begin
      \nz.mem_852_sv2v_reg  <= data_i[12];
    end 
    if(N4102) begin
      \nz.mem_851_sv2v_reg  <= data_i[11];
    end 
    if(N4101) begin
      \nz.mem_850_sv2v_reg  <= data_i[10];
    end 
    if(N4100) begin
      \nz.mem_849_sv2v_reg  <= data_i[9];
    end 
    if(N4099) begin
      \nz.mem_848_sv2v_reg  <= data_i[8];
    end 
    if(N4098) begin
      \nz.mem_847_sv2v_reg  <= data_i[7];
    end 
    if(N4097) begin
      \nz.mem_846_sv2v_reg  <= data_i[6];
    end 
    if(N4096) begin
      \nz.mem_845_sv2v_reg  <= data_i[5];
    end 
    if(N4095) begin
      \nz.mem_844_sv2v_reg  <= data_i[4];
    end 
    if(N4094) begin
      \nz.mem_843_sv2v_reg  <= data_i[3];
    end 
    if(N4093) begin
      \nz.mem_842_sv2v_reg  <= data_i[2];
    end 
    if(N4092) begin
      \nz.mem_841_sv2v_reg  <= data_i[1];
    end 
    if(N4091) begin
      \nz.mem_840_sv2v_reg  <= data_i[0];
    end 
    if(N4090) begin
      \nz.mem_839_sv2v_reg  <= data_i[39];
    end 
    if(N4089) begin
      \nz.mem_838_sv2v_reg  <= data_i[38];
    end 
    if(N4088) begin
      \nz.mem_837_sv2v_reg  <= data_i[37];
    end 
    if(N4087) begin
      \nz.mem_836_sv2v_reg  <= data_i[36];
    end 
    if(N4086) begin
      \nz.mem_835_sv2v_reg  <= data_i[35];
    end 
    if(N4085) begin
      \nz.mem_834_sv2v_reg  <= data_i[34];
    end 
    if(N4084) begin
      \nz.mem_833_sv2v_reg  <= data_i[33];
    end 
    if(N4083) begin
      \nz.mem_832_sv2v_reg  <= data_i[32];
    end 
    if(N4082) begin
      \nz.mem_831_sv2v_reg  <= data_i[31];
    end 
    if(N4081) begin
      \nz.mem_830_sv2v_reg  <= data_i[30];
    end 
    if(N4080) begin
      \nz.mem_829_sv2v_reg  <= data_i[29];
    end 
    if(N4079) begin
      \nz.mem_828_sv2v_reg  <= data_i[28];
    end 
    if(N4078) begin
      \nz.mem_827_sv2v_reg  <= data_i[27];
    end 
    if(N4077) begin
      \nz.mem_826_sv2v_reg  <= data_i[26];
    end 
    if(N4076) begin
      \nz.mem_825_sv2v_reg  <= data_i[25];
    end 
    if(N4075) begin
      \nz.mem_824_sv2v_reg  <= data_i[24];
    end 
    if(N4074) begin
      \nz.mem_823_sv2v_reg  <= data_i[23];
    end 
    if(N4073) begin
      \nz.mem_822_sv2v_reg  <= data_i[22];
    end 
    if(N4072) begin
      \nz.mem_821_sv2v_reg  <= data_i[21];
    end 
    if(N4071) begin
      \nz.mem_820_sv2v_reg  <= data_i[20];
    end 
    if(N4070) begin
      \nz.mem_819_sv2v_reg  <= data_i[19];
    end 
    if(N4069) begin
      \nz.mem_818_sv2v_reg  <= data_i[18];
    end 
    if(N4068) begin
      \nz.mem_817_sv2v_reg  <= data_i[17];
    end 
    if(N4067) begin
      \nz.mem_816_sv2v_reg  <= data_i[16];
    end 
    if(N4066) begin
      \nz.mem_815_sv2v_reg  <= data_i[15];
    end 
    if(N4065) begin
      \nz.mem_814_sv2v_reg  <= data_i[14];
    end 
    if(N4064) begin
      \nz.mem_813_sv2v_reg  <= data_i[13];
    end 
    if(N4063) begin
      \nz.mem_812_sv2v_reg  <= data_i[12];
    end 
    if(N4062) begin
      \nz.mem_811_sv2v_reg  <= data_i[11];
    end 
    if(N4061) begin
      \nz.mem_810_sv2v_reg  <= data_i[10];
    end 
    if(N4060) begin
      \nz.mem_809_sv2v_reg  <= data_i[9];
    end 
    if(N4059) begin
      \nz.mem_808_sv2v_reg  <= data_i[8];
    end 
    if(N4058) begin
      \nz.mem_807_sv2v_reg  <= data_i[7];
    end 
    if(N4057) begin
      \nz.mem_806_sv2v_reg  <= data_i[6];
    end 
    if(N4056) begin
      \nz.mem_805_sv2v_reg  <= data_i[5];
    end 
    if(N4055) begin
      \nz.mem_804_sv2v_reg  <= data_i[4];
    end 
    if(N4054) begin
      \nz.mem_803_sv2v_reg  <= data_i[3];
    end 
    if(N4053) begin
      \nz.mem_802_sv2v_reg  <= data_i[2];
    end 
    if(N4052) begin
      \nz.mem_801_sv2v_reg  <= data_i[1];
    end 
    if(N4051) begin
      \nz.mem_800_sv2v_reg  <= data_i[0];
    end 
    if(N4050) begin
      \nz.mem_799_sv2v_reg  <= data_i[39];
    end 
    if(N4049) begin
      \nz.mem_798_sv2v_reg  <= data_i[38];
    end 
    if(N4048) begin
      \nz.mem_797_sv2v_reg  <= data_i[37];
    end 
    if(N4047) begin
      \nz.mem_796_sv2v_reg  <= data_i[36];
    end 
    if(N4046) begin
      \nz.mem_795_sv2v_reg  <= data_i[35];
    end 
    if(N4045) begin
      \nz.mem_794_sv2v_reg  <= data_i[34];
    end 
    if(N4044) begin
      \nz.mem_793_sv2v_reg  <= data_i[33];
    end 
    if(N4043) begin
      \nz.mem_792_sv2v_reg  <= data_i[32];
    end 
    if(N4042) begin
      \nz.mem_791_sv2v_reg  <= data_i[31];
    end 
    if(N4041) begin
      \nz.mem_790_sv2v_reg  <= data_i[30];
    end 
    if(N4040) begin
      \nz.mem_789_sv2v_reg  <= data_i[29];
    end 
    if(N4039) begin
      \nz.mem_788_sv2v_reg  <= data_i[28];
    end 
    if(N4038) begin
      \nz.mem_787_sv2v_reg  <= data_i[27];
    end 
    if(N4037) begin
      \nz.mem_786_sv2v_reg  <= data_i[26];
    end 
    if(N4036) begin
      \nz.mem_785_sv2v_reg  <= data_i[25];
    end 
    if(N4035) begin
      \nz.mem_784_sv2v_reg  <= data_i[24];
    end 
    if(N4034) begin
      \nz.mem_783_sv2v_reg  <= data_i[23];
    end 
    if(N4033) begin
      \nz.mem_782_sv2v_reg  <= data_i[22];
    end 
    if(N4032) begin
      \nz.mem_781_sv2v_reg  <= data_i[21];
    end 
    if(N4031) begin
      \nz.mem_780_sv2v_reg  <= data_i[20];
    end 
    if(N4030) begin
      \nz.mem_779_sv2v_reg  <= data_i[19];
    end 
    if(N4029) begin
      \nz.mem_778_sv2v_reg  <= data_i[18];
    end 
    if(N4028) begin
      \nz.mem_777_sv2v_reg  <= data_i[17];
    end 
    if(N4027) begin
      \nz.mem_776_sv2v_reg  <= data_i[16];
    end 
    if(N4026) begin
      \nz.mem_775_sv2v_reg  <= data_i[15];
    end 
    if(N4025) begin
      \nz.mem_774_sv2v_reg  <= data_i[14];
    end 
    if(N4024) begin
      \nz.mem_773_sv2v_reg  <= data_i[13];
    end 
    if(N4023) begin
      \nz.mem_772_sv2v_reg  <= data_i[12];
    end 
    if(N4022) begin
      \nz.mem_771_sv2v_reg  <= data_i[11];
    end 
    if(N4021) begin
      \nz.mem_770_sv2v_reg  <= data_i[10];
    end 
    if(N4020) begin
      \nz.mem_769_sv2v_reg  <= data_i[9];
    end 
    if(N4019) begin
      \nz.mem_768_sv2v_reg  <= data_i[8];
    end 
    if(N4018) begin
      \nz.mem_767_sv2v_reg  <= data_i[7];
    end 
    if(N4017) begin
      \nz.mem_766_sv2v_reg  <= data_i[6];
    end 
    if(N4016) begin
      \nz.mem_765_sv2v_reg  <= data_i[5];
    end 
    if(N4015) begin
      \nz.mem_764_sv2v_reg  <= data_i[4];
    end 
    if(N4014) begin
      \nz.mem_763_sv2v_reg  <= data_i[3];
    end 
    if(N4013) begin
      \nz.mem_762_sv2v_reg  <= data_i[2];
    end 
    if(N4012) begin
      \nz.mem_761_sv2v_reg  <= data_i[1];
    end 
    if(N4011) begin
      \nz.mem_760_sv2v_reg  <= data_i[0];
    end 
    if(N4010) begin
      \nz.mem_759_sv2v_reg  <= data_i[39];
    end 
    if(N4009) begin
      \nz.mem_758_sv2v_reg  <= data_i[38];
    end 
    if(N4008) begin
      \nz.mem_757_sv2v_reg  <= data_i[37];
    end 
    if(N4007) begin
      \nz.mem_756_sv2v_reg  <= data_i[36];
    end 
    if(N4006) begin
      \nz.mem_755_sv2v_reg  <= data_i[35];
    end 
    if(N4005) begin
      \nz.mem_754_sv2v_reg  <= data_i[34];
    end 
    if(N4004) begin
      \nz.mem_753_sv2v_reg  <= data_i[33];
    end 
    if(N4003) begin
      \nz.mem_752_sv2v_reg  <= data_i[32];
    end 
    if(N4002) begin
      \nz.mem_751_sv2v_reg  <= data_i[31];
    end 
    if(N4001) begin
      \nz.mem_750_sv2v_reg  <= data_i[30];
    end 
    if(N4000) begin
      \nz.mem_749_sv2v_reg  <= data_i[29];
    end 
    if(N3999) begin
      \nz.mem_748_sv2v_reg  <= data_i[28];
    end 
    if(N3998) begin
      \nz.mem_747_sv2v_reg  <= data_i[27];
    end 
    if(N3997) begin
      \nz.mem_746_sv2v_reg  <= data_i[26];
    end 
    if(N3996) begin
      \nz.mem_745_sv2v_reg  <= data_i[25];
    end 
    if(N3995) begin
      \nz.mem_744_sv2v_reg  <= data_i[24];
    end 
    if(N3994) begin
      \nz.mem_743_sv2v_reg  <= data_i[23];
    end 
    if(N3993) begin
      \nz.mem_742_sv2v_reg  <= data_i[22];
    end 
    if(N3992) begin
      \nz.mem_741_sv2v_reg  <= data_i[21];
    end 
    if(N3991) begin
      \nz.mem_740_sv2v_reg  <= data_i[20];
    end 
    if(N3990) begin
      \nz.mem_739_sv2v_reg  <= data_i[19];
    end 
    if(N3989) begin
      \nz.mem_738_sv2v_reg  <= data_i[18];
    end 
    if(N3988) begin
      \nz.mem_737_sv2v_reg  <= data_i[17];
    end 
    if(N3987) begin
      \nz.mem_736_sv2v_reg  <= data_i[16];
    end 
    if(N3986) begin
      \nz.mem_735_sv2v_reg  <= data_i[15];
    end 
    if(N3985) begin
      \nz.mem_734_sv2v_reg  <= data_i[14];
    end 
    if(N3984) begin
      \nz.mem_733_sv2v_reg  <= data_i[13];
    end 
    if(N3983) begin
      \nz.mem_732_sv2v_reg  <= data_i[12];
    end 
    if(N3982) begin
      \nz.mem_731_sv2v_reg  <= data_i[11];
    end 
    if(N3981) begin
      \nz.mem_730_sv2v_reg  <= data_i[10];
    end 
    if(N3980) begin
      \nz.mem_729_sv2v_reg  <= data_i[9];
    end 
    if(N3979) begin
      \nz.mem_728_sv2v_reg  <= data_i[8];
    end 
    if(N3978) begin
      \nz.mem_727_sv2v_reg  <= data_i[7];
    end 
    if(N3977) begin
      \nz.mem_726_sv2v_reg  <= data_i[6];
    end 
    if(N3976) begin
      \nz.mem_725_sv2v_reg  <= data_i[5];
    end 
    if(N3975) begin
      \nz.mem_724_sv2v_reg  <= data_i[4];
    end 
    if(N3974) begin
      \nz.mem_723_sv2v_reg  <= data_i[3];
    end 
    if(N3973) begin
      \nz.mem_722_sv2v_reg  <= data_i[2];
    end 
    if(N3972) begin
      \nz.mem_721_sv2v_reg  <= data_i[1];
    end 
    if(N3971) begin
      \nz.mem_720_sv2v_reg  <= data_i[0];
    end 
    if(N3970) begin
      \nz.mem_719_sv2v_reg  <= data_i[39];
    end 
    if(N3969) begin
      \nz.mem_718_sv2v_reg  <= data_i[38];
    end 
    if(N3968) begin
      \nz.mem_717_sv2v_reg  <= data_i[37];
    end 
    if(N3967) begin
      \nz.mem_716_sv2v_reg  <= data_i[36];
    end 
    if(N3966) begin
      \nz.mem_715_sv2v_reg  <= data_i[35];
    end 
    if(N3965) begin
      \nz.mem_714_sv2v_reg  <= data_i[34];
    end 
    if(N3964) begin
      \nz.mem_713_sv2v_reg  <= data_i[33];
    end 
    if(N3963) begin
      \nz.mem_712_sv2v_reg  <= data_i[32];
    end 
    if(N3962) begin
      \nz.mem_711_sv2v_reg  <= data_i[31];
    end 
    if(N3961) begin
      \nz.mem_710_sv2v_reg  <= data_i[30];
    end 
    if(N3960) begin
      \nz.mem_709_sv2v_reg  <= data_i[29];
    end 
    if(N3959) begin
      \nz.mem_708_sv2v_reg  <= data_i[28];
    end 
    if(N3958) begin
      \nz.mem_707_sv2v_reg  <= data_i[27];
    end 
    if(N3957) begin
      \nz.mem_706_sv2v_reg  <= data_i[26];
    end 
    if(N3956) begin
      \nz.mem_705_sv2v_reg  <= data_i[25];
    end 
    if(N3955) begin
      \nz.mem_704_sv2v_reg  <= data_i[24];
    end 
    if(N3954) begin
      \nz.mem_703_sv2v_reg  <= data_i[23];
    end 
    if(N3953) begin
      \nz.mem_702_sv2v_reg  <= data_i[22];
    end 
    if(N3952) begin
      \nz.mem_701_sv2v_reg  <= data_i[21];
    end 
    if(N3951) begin
      \nz.mem_700_sv2v_reg  <= data_i[20];
    end 
    if(N3950) begin
      \nz.mem_699_sv2v_reg  <= data_i[19];
    end 
    if(N3949) begin
      \nz.mem_698_sv2v_reg  <= data_i[18];
    end 
    if(N3948) begin
      \nz.mem_697_sv2v_reg  <= data_i[17];
    end 
    if(N3947) begin
      \nz.mem_696_sv2v_reg  <= data_i[16];
    end 
    if(N3946) begin
      \nz.mem_695_sv2v_reg  <= data_i[15];
    end 
    if(N3945) begin
      \nz.mem_694_sv2v_reg  <= data_i[14];
    end 
    if(N3944) begin
      \nz.mem_693_sv2v_reg  <= data_i[13];
    end 
    if(N3943) begin
      \nz.mem_692_sv2v_reg  <= data_i[12];
    end 
    if(N3942) begin
      \nz.mem_691_sv2v_reg  <= data_i[11];
    end 
    if(N3941) begin
      \nz.mem_690_sv2v_reg  <= data_i[10];
    end 
    if(N3940) begin
      \nz.mem_689_sv2v_reg  <= data_i[9];
    end 
    if(N3939) begin
      \nz.mem_688_sv2v_reg  <= data_i[8];
    end 
    if(N3938) begin
      \nz.mem_687_sv2v_reg  <= data_i[7];
    end 
    if(N3937) begin
      \nz.mem_686_sv2v_reg  <= data_i[6];
    end 
    if(N3936) begin
      \nz.mem_685_sv2v_reg  <= data_i[5];
    end 
    if(N3935) begin
      \nz.mem_684_sv2v_reg  <= data_i[4];
    end 
    if(N3934) begin
      \nz.mem_683_sv2v_reg  <= data_i[3];
    end 
    if(N3933) begin
      \nz.mem_682_sv2v_reg  <= data_i[2];
    end 
    if(N3932) begin
      \nz.mem_681_sv2v_reg  <= data_i[1];
    end 
    if(N3931) begin
      \nz.mem_680_sv2v_reg  <= data_i[0];
    end 
    if(N3930) begin
      \nz.mem_679_sv2v_reg  <= data_i[39];
    end 
    if(N3929) begin
      \nz.mem_678_sv2v_reg  <= data_i[38];
    end 
    if(N3928) begin
      \nz.mem_677_sv2v_reg  <= data_i[37];
    end 
    if(N3927) begin
      \nz.mem_676_sv2v_reg  <= data_i[36];
    end 
    if(N3926) begin
      \nz.mem_675_sv2v_reg  <= data_i[35];
    end 
    if(N3925) begin
      \nz.mem_674_sv2v_reg  <= data_i[34];
    end 
    if(N3924) begin
      \nz.mem_673_sv2v_reg  <= data_i[33];
    end 
    if(N3923) begin
      \nz.mem_672_sv2v_reg  <= data_i[32];
    end 
    if(N3922) begin
      \nz.mem_671_sv2v_reg  <= data_i[31];
    end 
    if(N3921) begin
      \nz.mem_670_sv2v_reg  <= data_i[30];
    end 
    if(N3920) begin
      \nz.mem_669_sv2v_reg  <= data_i[29];
    end 
    if(N3919) begin
      \nz.mem_668_sv2v_reg  <= data_i[28];
    end 
    if(N3918) begin
      \nz.mem_667_sv2v_reg  <= data_i[27];
    end 
    if(N3917) begin
      \nz.mem_666_sv2v_reg  <= data_i[26];
    end 
    if(N3916) begin
      \nz.mem_665_sv2v_reg  <= data_i[25];
    end 
    if(N3915) begin
      \nz.mem_664_sv2v_reg  <= data_i[24];
    end 
    if(N3914) begin
      \nz.mem_663_sv2v_reg  <= data_i[23];
    end 
    if(N3913) begin
      \nz.mem_662_sv2v_reg  <= data_i[22];
    end 
    if(N3912) begin
      \nz.mem_661_sv2v_reg  <= data_i[21];
    end 
    if(N3911) begin
      \nz.mem_660_sv2v_reg  <= data_i[20];
    end 
    if(N3910) begin
      \nz.mem_659_sv2v_reg  <= data_i[19];
    end 
    if(N3909) begin
      \nz.mem_658_sv2v_reg  <= data_i[18];
    end 
    if(N3908) begin
      \nz.mem_657_sv2v_reg  <= data_i[17];
    end 
    if(N3907) begin
      \nz.mem_656_sv2v_reg  <= data_i[16];
    end 
    if(N3906) begin
      \nz.mem_655_sv2v_reg  <= data_i[15];
    end 
    if(N3905) begin
      \nz.mem_654_sv2v_reg  <= data_i[14];
    end 
    if(N3904) begin
      \nz.mem_653_sv2v_reg  <= data_i[13];
    end 
    if(N3903) begin
      \nz.mem_652_sv2v_reg  <= data_i[12];
    end 
    if(N3902) begin
      \nz.mem_651_sv2v_reg  <= data_i[11];
    end 
    if(N3901) begin
      \nz.mem_650_sv2v_reg  <= data_i[10];
    end 
    if(N3900) begin
      \nz.mem_649_sv2v_reg  <= data_i[9];
    end 
    if(N3899) begin
      \nz.mem_648_sv2v_reg  <= data_i[8];
    end 
    if(N3898) begin
      \nz.mem_647_sv2v_reg  <= data_i[7];
    end 
    if(N3897) begin
      \nz.mem_646_sv2v_reg  <= data_i[6];
    end 
    if(N3896) begin
      \nz.mem_645_sv2v_reg  <= data_i[5];
    end 
    if(N3895) begin
      \nz.mem_644_sv2v_reg  <= data_i[4];
    end 
    if(N3894) begin
      \nz.mem_643_sv2v_reg  <= data_i[3];
    end 
    if(N3893) begin
      \nz.mem_642_sv2v_reg  <= data_i[2];
    end 
    if(N3892) begin
      \nz.mem_641_sv2v_reg  <= data_i[1];
    end 
    if(N3891) begin
      \nz.mem_640_sv2v_reg  <= data_i[0];
    end 
    if(N3890) begin
      \nz.mem_639_sv2v_reg  <= data_i[39];
    end 
    if(N3889) begin
      \nz.mem_638_sv2v_reg  <= data_i[38];
    end 
    if(N3888) begin
      \nz.mem_637_sv2v_reg  <= data_i[37];
    end 
    if(N3887) begin
      \nz.mem_636_sv2v_reg  <= data_i[36];
    end 
    if(N3886) begin
      \nz.mem_635_sv2v_reg  <= data_i[35];
    end 
    if(N3885) begin
      \nz.mem_634_sv2v_reg  <= data_i[34];
    end 
    if(N3884) begin
      \nz.mem_633_sv2v_reg  <= data_i[33];
    end 
    if(N3883) begin
      \nz.mem_632_sv2v_reg  <= data_i[32];
    end 
    if(N3882) begin
      \nz.mem_631_sv2v_reg  <= data_i[31];
    end 
    if(N3881) begin
      \nz.mem_630_sv2v_reg  <= data_i[30];
    end 
    if(N3880) begin
      \nz.mem_629_sv2v_reg  <= data_i[29];
    end 
    if(N3879) begin
      \nz.mem_628_sv2v_reg  <= data_i[28];
    end 
    if(N3878) begin
      \nz.mem_627_sv2v_reg  <= data_i[27];
    end 
    if(N3877) begin
      \nz.mem_626_sv2v_reg  <= data_i[26];
    end 
    if(N3876) begin
      \nz.mem_625_sv2v_reg  <= data_i[25];
    end 
    if(N3875) begin
      \nz.mem_624_sv2v_reg  <= data_i[24];
    end 
    if(N3874) begin
      \nz.mem_623_sv2v_reg  <= data_i[23];
    end 
    if(N3873) begin
      \nz.mem_622_sv2v_reg  <= data_i[22];
    end 
    if(N3872) begin
      \nz.mem_621_sv2v_reg  <= data_i[21];
    end 
    if(N3871) begin
      \nz.mem_620_sv2v_reg  <= data_i[20];
    end 
    if(N3870) begin
      \nz.mem_619_sv2v_reg  <= data_i[19];
    end 
    if(N3869) begin
      \nz.mem_618_sv2v_reg  <= data_i[18];
    end 
    if(N3868) begin
      \nz.mem_617_sv2v_reg  <= data_i[17];
    end 
    if(N3867) begin
      \nz.mem_616_sv2v_reg  <= data_i[16];
    end 
    if(N3866) begin
      \nz.mem_615_sv2v_reg  <= data_i[15];
    end 
    if(N3865) begin
      \nz.mem_614_sv2v_reg  <= data_i[14];
    end 
    if(N3864) begin
      \nz.mem_613_sv2v_reg  <= data_i[13];
    end 
    if(N3863) begin
      \nz.mem_612_sv2v_reg  <= data_i[12];
    end 
    if(N3862) begin
      \nz.mem_611_sv2v_reg  <= data_i[11];
    end 
    if(N3861) begin
      \nz.mem_610_sv2v_reg  <= data_i[10];
    end 
    if(N3860) begin
      \nz.mem_609_sv2v_reg  <= data_i[9];
    end 
    if(N3859) begin
      \nz.mem_608_sv2v_reg  <= data_i[8];
    end 
    if(N3858) begin
      \nz.mem_607_sv2v_reg  <= data_i[7];
    end 
    if(N3857) begin
      \nz.mem_606_sv2v_reg  <= data_i[6];
    end 
    if(N3856) begin
      \nz.mem_605_sv2v_reg  <= data_i[5];
    end 
    if(N3855) begin
      \nz.mem_604_sv2v_reg  <= data_i[4];
    end 
    if(N3854) begin
      \nz.mem_603_sv2v_reg  <= data_i[3];
    end 
    if(N3853) begin
      \nz.mem_602_sv2v_reg  <= data_i[2];
    end 
    if(N3852) begin
      \nz.mem_601_sv2v_reg  <= data_i[1];
    end 
    if(N3851) begin
      \nz.mem_600_sv2v_reg  <= data_i[0];
    end 
    if(N3850) begin
      \nz.mem_599_sv2v_reg  <= data_i[39];
    end 
    if(N3849) begin
      \nz.mem_598_sv2v_reg  <= data_i[38];
    end 
    if(N3848) begin
      \nz.mem_597_sv2v_reg  <= data_i[37];
    end 
    if(N3847) begin
      \nz.mem_596_sv2v_reg  <= data_i[36];
    end 
    if(N3846) begin
      \nz.mem_595_sv2v_reg  <= data_i[35];
    end 
    if(N3845) begin
      \nz.mem_594_sv2v_reg  <= data_i[34];
    end 
    if(N3844) begin
      \nz.mem_593_sv2v_reg  <= data_i[33];
    end 
    if(N3843) begin
      \nz.mem_592_sv2v_reg  <= data_i[32];
    end 
    if(N3842) begin
      \nz.mem_591_sv2v_reg  <= data_i[31];
    end 
    if(N3841) begin
      \nz.mem_590_sv2v_reg  <= data_i[30];
    end 
    if(N3840) begin
      \nz.mem_589_sv2v_reg  <= data_i[29];
    end 
    if(N3839) begin
      \nz.mem_588_sv2v_reg  <= data_i[28];
    end 
    if(N3838) begin
      \nz.mem_587_sv2v_reg  <= data_i[27];
    end 
    if(N3837) begin
      \nz.mem_586_sv2v_reg  <= data_i[26];
    end 
    if(N3836) begin
      \nz.mem_585_sv2v_reg  <= data_i[25];
    end 
    if(N3835) begin
      \nz.mem_584_sv2v_reg  <= data_i[24];
    end 
    if(N3834) begin
      \nz.mem_583_sv2v_reg  <= data_i[23];
    end 
    if(N3833) begin
      \nz.mem_582_sv2v_reg  <= data_i[22];
    end 
    if(N3832) begin
      \nz.mem_581_sv2v_reg  <= data_i[21];
    end 
    if(N3831) begin
      \nz.mem_580_sv2v_reg  <= data_i[20];
    end 
    if(N3830) begin
      \nz.mem_579_sv2v_reg  <= data_i[19];
    end 
    if(N3829) begin
      \nz.mem_578_sv2v_reg  <= data_i[18];
    end 
    if(N3828) begin
      \nz.mem_577_sv2v_reg  <= data_i[17];
    end 
    if(N3827) begin
      \nz.mem_576_sv2v_reg  <= data_i[16];
    end 
    if(N3826) begin
      \nz.mem_575_sv2v_reg  <= data_i[15];
    end 
    if(N3825) begin
      \nz.mem_574_sv2v_reg  <= data_i[14];
    end 
    if(N3824) begin
      \nz.mem_573_sv2v_reg  <= data_i[13];
    end 
    if(N3823) begin
      \nz.mem_572_sv2v_reg  <= data_i[12];
    end 
    if(N3822) begin
      \nz.mem_571_sv2v_reg  <= data_i[11];
    end 
    if(N3821) begin
      \nz.mem_570_sv2v_reg  <= data_i[10];
    end 
    if(N3820) begin
      \nz.mem_569_sv2v_reg  <= data_i[9];
    end 
    if(N3819) begin
      \nz.mem_568_sv2v_reg  <= data_i[8];
    end 
    if(N3818) begin
      \nz.mem_567_sv2v_reg  <= data_i[7];
    end 
    if(N3817) begin
      \nz.mem_566_sv2v_reg  <= data_i[6];
    end 
    if(N3816) begin
      \nz.mem_565_sv2v_reg  <= data_i[5];
    end 
    if(N3815) begin
      \nz.mem_564_sv2v_reg  <= data_i[4];
    end 
    if(N3814) begin
      \nz.mem_563_sv2v_reg  <= data_i[3];
    end 
    if(N3813) begin
      \nz.mem_562_sv2v_reg  <= data_i[2];
    end 
    if(N3812) begin
      \nz.mem_561_sv2v_reg  <= data_i[1];
    end 
    if(N3811) begin
      \nz.mem_560_sv2v_reg  <= data_i[0];
    end 
    if(N3810) begin
      \nz.mem_559_sv2v_reg  <= data_i[39];
    end 
    if(N3809) begin
      \nz.mem_558_sv2v_reg  <= data_i[38];
    end 
    if(N3808) begin
      \nz.mem_557_sv2v_reg  <= data_i[37];
    end 
    if(N3807) begin
      \nz.mem_556_sv2v_reg  <= data_i[36];
    end 
    if(N3806) begin
      \nz.mem_555_sv2v_reg  <= data_i[35];
    end 
    if(N3805) begin
      \nz.mem_554_sv2v_reg  <= data_i[34];
    end 
    if(N3804) begin
      \nz.mem_553_sv2v_reg  <= data_i[33];
    end 
    if(N3803) begin
      \nz.mem_552_sv2v_reg  <= data_i[32];
    end 
    if(N3802) begin
      \nz.mem_551_sv2v_reg  <= data_i[31];
    end 
    if(N3801) begin
      \nz.mem_550_sv2v_reg  <= data_i[30];
    end 
    if(N3800) begin
      \nz.mem_549_sv2v_reg  <= data_i[29];
    end 
    if(N3799) begin
      \nz.mem_548_sv2v_reg  <= data_i[28];
    end 
    if(N3798) begin
      \nz.mem_547_sv2v_reg  <= data_i[27];
    end 
    if(N3797) begin
      \nz.mem_546_sv2v_reg  <= data_i[26];
    end 
    if(N3796) begin
      \nz.mem_545_sv2v_reg  <= data_i[25];
    end 
    if(N3795) begin
      \nz.mem_544_sv2v_reg  <= data_i[24];
    end 
    if(N3794) begin
      \nz.mem_543_sv2v_reg  <= data_i[23];
    end 
    if(N3793) begin
      \nz.mem_542_sv2v_reg  <= data_i[22];
    end 
    if(N3792) begin
      \nz.mem_541_sv2v_reg  <= data_i[21];
    end 
    if(N3791) begin
      \nz.mem_540_sv2v_reg  <= data_i[20];
    end 
    if(N3790) begin
      \nz.mem_539_sv2v_reg  <= data_i[19];
    end 
    if(N3789) begin
      \nz.mem_538_sv2v_reg  <= data_i[18];
    end 
    if(N3788) begin
      \nz.mem_537_sv2v_reg  <= data_i[17];
    end 
    if(N3787) begin
      \nz.mem_536_sv2v_reg  <= data_i[16];
    end 
    if(N3786) begin
      \nz.mem_535_sv2v_reg  <= data_i[15];
    end 
    if(N3785) begin
      \nz.mem_534_sv2v_reg  <= data_i[14];
    end 
    if(N3784) begin
      \nz.mem_533_sv2v_reg  <= data_i[13];
    end 
    if(N3783) begin
      \nz.mem_532_sv2v_reg  <= data_i[12];
    end 
    if(N3782) begin
      \nz.mem_531_sv2v_reg  <= data_i[11];
    end 
    if(N3781) begin
      \nz.mem_530_sv2v_reg  <= data_i[10];
    end 
    if(N3780) begin
      \nz.mem_529_sv2v_reg  <= data_i[9];
    end 
    if(N3779) begin
      \nz.mem_528_sv2v_reg  <= data_i[8];
    end 
    if(N3778) begin
      \nz.mem_527_sv2v_reg  <= data_i[7];
    end 
    if(N3777) begin
      \nz.mem_526_sv2v_reg  <= data_i[6];
    end 
    if(N3776) begin
      \nz.mem_525_sv2v_reg  <= data_i[5];
    end 
    if(N3775) begin
      \nz.mem_524_sv2v_reg  <= data_i[4];
    end 
    if(N3774) begin
      \nz.mem_523_sv2v_reg  <= data_i[3];
    end 
    if(N3773) begin
      \nz.mem_522_sv2v_reg  <= data_i[2];
    end 
    if(N3772) begin
      \nz.mem_521_sv2v_reg  <= data_i[1];
    end 
    if(N3771) begin
      \nz.mem_520_sv2v_reg  <= data_i[0];
    end 
    if(N3770) begin
      \nz.mem_519_sv2v_reg  <= data_i[39];
    end 
    if(N3769) begin
      \nz.mem_518_sv2v_reg  <= data_i[38];
    end 
    if(N3768) begin
      \nz.mem_517_sv2v_reg  <= data_i[37];
    end 
    if(N3767) begin
      \nz.mem_516_sv2v_reg  <= data_i[36];
    end 
    if(N3766) begin
      \nz.mem_515_sv2v_reg  <= data_i[35];
    end 
    if(N3765) begin
      \nz.mem_514_sv2v_reg  <= data_i[34];
    end 
    if(N3764) begin
      \nz.mem_513_sv2v_reg  <= data_i[33];
    end 
    if(N3763) begin
      \nz.mem_512_sv2v_reg  <= data_i[32];
    end 
    if(N3762) begin
      \nz.mem_511_sv2v_reg  <= data_i[31];
    end 
    if(N3761) begin
      \nz.mem_510_sv2v_reg  <= data_i[30];
    end 
    if(N3760) begin
      \nz.mem_509_sv2v_reg  <= data_i[29];
    end 
    if(N3759) begin
      \nz.mem_508_sv2v_reg  <= data_i[28];
    end 
    if(N3758) begin
      \nz.mem_507_sv2v_reg  <= data_i[27];
    end 
    if(N3757) begin
      \nz.mem_506_sv2v_reg  <= data_i[26];
    end 
    if(N3756) begin
      \nz.mem_505_sv2v_reg  <= data_i[25];
    end 
    if(N3755) begin
      \nz.mem_504_sv2v_reg  <= data_i[24];
    end 
    if(N3754) begin
      \nz.mem_503_sv2v_reg  <= data_i[23];
    end 
    if(N3753) begin
      \nz.mem_502_sv2v_reg  <= data_i[22];
    end 
    if(N3752) begin
      \nz.mem_501_sv2v_reg  <= data_i[21];
    end 
    if(N3751) begin
      \nz.mem_500_sv2v_reg  <= data_i[20];
    end 
    if(N3750) begin
      \nz.mem_499_sv2v_reg  <= data_i[19];
    end 
    if(N3749) begin
      \nz.mem_498_sv2v_reg  <= data_i[18];
    end 
    if(N3748) begin
      \nz.mem_497_sv2v_reg  <= data_i[17];
    end 
    if(N3747) begin
      \nz.mem_496_sv2v_reg  <= data_i[16];
    end 
    if(N3746) begin
      \nz.mem_495_sv2v_reg  <= data_i[15];
    end 
    if(N3745) begin
      \nz.mem_494_sv2v_reg  <= data_i[14];
    end 
    if(N3744) begin
      \nz.mem_493_sv2v_reg  <= data_i[13];
    end 
    if(N3743) begin
      \nz.mem_492_sv2v_reg  <= data_i[12];
    end 
    if(N3742) begin
      \nz.mem_491_sv2v_reg  <= data_i[11];
    end 
    if(N3741) begin
      \nz.mem_490_sv2v_reg  <= data_i[10];
    end 
    if(N3740) begin
      \nz.mem_489_sv2v_reg  <= data_i[9];
    end 
    if(N3739) begin
      \nz.mem_488_sv2v_reg  <= data_i[8];
    end 
    if(N3738) begin
      \nz.mem_487_sv2v_reg  <= data_i[7];
    end 
    if(N3737) begin
      \nz.mem_486_sv2v_reg  <= data_i[6];
    end 
    if(N3736) begin
      \nz.mem_485_sv2v_reg  <= data_i[5];
    end 
    if(N3735) begin
      \nz.mem_484_sv2v_reg  <= data_i[4];
    end 
    if(N3734) begin
      \nz.mem_483_sv2v_reg  <= data_i[3];
    end 
    if(N3733) begin
      \nz.mem_482_sv2v_reg  <= data_i[2];
    end 
    if(N3732) begin
      \nz.mem_481_sv2v_reg  <= data_i[1];
    end 
    if(N3731) begin
      \nz.mem_480_sv2v_reg  <= data_i[0];
    end 
    if(N3730) begin
      \nz.mem_479_sv2v_reg  <= data_i[39];
    end 
    if(N3729) begin
      \nz.mem_478_sv2v_reg  <= data_i[38];
    end 
    if(N3728) begin
      \nz.mem_477_sv2v_reg  <= data_i[37];
    end 
    if(N3727) begin
      \nz.mem_476_sv2v_reg  <= data_i[36];
    end 
    if(N3726) begin
      \nz.mem_475_sv2v_reg  <= data_i[35];
    end 
    if(N3725) begin
      \nz.mem_474_sv2v_reg  <= data_i[34];
    end 
    if(N3724) begin
      \nz.mem_473_sv2v_reg  <= data_i[33];
    end 
    if(N3723) begin
      \nz.mem_472_sv2v_reg  <= data_i[32];
    end 
    if(N3722) begin
      \nz.mem_471_sv2v_reg  <= data_i[31];
    end 
    if(N3721) begin
      \nz.mem_470_sv2v_reg  <= data_i[30];
    end 
    if(N3720) begin
      \nz.mem_469_sv2v_reg  <= data_i[29];
    end 
    if(N3719) begin
      \nz.mem_468_sv2v_reg  <= data_i[28];
    end 
    if(N3718) begin
      \nz.mem_467_sv2v_reg  <= data_i[27];
    end 
    if(N3717) begin
      \nz.mem_466_sv2v_reg  <= data_i[26];
    end 
    if(N3716) begin
      \nz.mem_465_sv2v_reg  <= data_i[25];
    end 
    if(N3715) begin
      \nz.mem_464_sv2v_reg  <= data_i[24];
    end 
    if(N3714) begin
      \nz.mem_463_sv2v_reg  <= data_i[23];
    end 
    if(N3713) begin
      \nz.mem_462_sv2v_reg  <= data_i[22];
    end 
    if(N3712) begin
      \nz.mem_461_sv2v_reg  <= data_i[21];
    end 
    if(N3711) begin
      \nz.mem_460_sv2v_reg  <= data_i[20];
    end 
    if(N3710) begin
      \nz.mem_459_sv2v_reg  <= data_i[19];
    end 
    if(N3709) begin
      \nz.mem_458_sv2v_reg  <= data_i[18];
    end 
    if(N3708) begin
      \nz.mem_457_sv2v_reg  <= data_i[17];
    end 
    if(N3707) begin
      \nz.mem_456_sv2v_reg  <= data_i[16];
    end 
    if(N3706) begin
      \nz.mem_455_sv2v_reg  <= data_i[15];
    end 
    if(N3705) begin
      \nz.mem_454_sv2v_reg  <= data_i[14];
    end 
    if(N3704) begin
      \nz.mem_453_sv2v_reg  <= data_i[13];
    end 
    if(N3703) begin
      \nz.mem_452_sv2v_reg  <= data_i[12];
    end 
    if(N3702) begin
      \nz.mem_451_sv2v_reg  <= data_i[11];
    end 
    if(N3701) begin
      \nz.mem_450_sv2v_reg  <= data_i[10];
    end 
    if(N3700) begin
      \nz.mem_449_sv2v_reg  <= data_i[9];
    end 
    if(N3699) begin
      \nz.mem_448_sv2v_reg  <= data_i[8];
    end 
    if(N3698) begin
      \nz.mem_447_sv2v_reg  <= data_i[7];
    end 
    if(N3697) begin
      \nz.mem_446_sv2v_reg  <= data_i[6];
    end 
    if(N3696) begin
      \nz.mem_445_sv2v_reg  <= data_i[5];
    end 
    if(N3695) begin
      \nz.mem_444_sv2v_reg  <= data_i[4];
    end 
    if(N3694) begin
      \nz.mem_443_sv2v_reg  <= data_i[3];
    end 
    if(N3693) begin
      \nz.mem_442_sv2v_reg  <= data_i[2];
    end 
    if(N3692) begin
      \nz.mem_441_sv2v_reg  <= data_i[1];
    end 
    if(N3691) begin
      \nz.mem_440_sv2v_reg  <= data_i[0];
    end 
    if(N3690) begin
      \nz.mem_439_sv2v_reg  <= data_i[39];
    end 
    if(N3689) begin
      \nz.mem_438_sv2v_reg  <= data_i[38];
    end 
    if(N3688) begin
      \nz.mem_437_sv2v_reg  <= data_i[37];
    end 
    if(N3687) begin
      \nz.mem_436_sv2v_reg  <= data_i[36];
    end 
    if(N3686) begin
      \nz.mem_435_sv2v_reg  <= data_i[35];
    end 
    if(N3685) begin
      \nz.mem_434_sv2v_reg  <= data_i[34];
    end 
    if(N3684) begin
      \nz.mem_433_sv2v_reg  <= data_i[33];
    end 
    if(N3683) begin
      \nz.mem_432_sv2v_reg  <= data_i[32];
    end 
    if(N3682) begin
      \nz.mem_431_sv2v_reg  <= data_i[31];
    end 
    if(N3681) begin
      \nz.mem_430_sv2v_reg  <= data_i[30];
    end 
    if(N3680) begin
      \nz.mem_429_sv2v_reg  <= data_i[29];
    end 
    if(N3679) begin
      \nz.mem_428_sv2v_reg  <= data_i[28];
    end 
    if(N3678) begin
      \nz.mem_427_sv2v_reg  <= data_i[27];
    end 
    if(N3677) begin
      \nz.mem_426_sv2v_reg  <= data_i[26];
    end 
    if(N3676) begin
      \nz.mem_425_sv2v_reg  <= data_i[25];
    end 
    if(N3675) begin
      \nz.mem_424_sv2v_reg  <= data_i[24];
    end 
    if(N3674) begin
      \nz.mem_423_sv2v_reg  <= data_i[23];
    end 
    if(N3673) begin
      \nz.mem_422_sv2v_reg  <= data_i[22];
    end 
    if(N3672) begin
      \nz.mem_421_sv2v_reg  <= data_i[21];
    end 
    if(N3671) begin
      \nz.mem_420_sv2v_reg  <= data_i[20];
    end 
    if(N3670) begin
      \nz.mem_419_sv2v_reg  <= data_i[19];
    end 
    if(N3669) begin
      \nz.mem_418_sv2v_reg  <= data_i[18];
    end 
    if(N3668) begin
      \nz.mem_417_sv2v_reg  <= data_i[17];
    end 
    if(N3667) begin
      \nz.mem_416_sv2v_reg  <= data_i[16];
    end 
    if(N3666) begin
      \nz.mem_415_sv2v_reg  <= data_i[15];
    end 
    if(N3665) begin
      \nz.mem_414_sv2v_reg  <= data_i[14];
    end 
    if(N3664) begin
      \nz.mem_413_sv2v_reg  <= data_i[13];
    end 
    if(N3663) begin
      \nz.mem_412_sv2v_reg  <= data_i[12];
    end 
    if(N3662) begin
      \nz.mem_411_sv2v_reg  <= data_i[11];
    end 
    if(N3661) begin
      \nz.mem_410_sv2v_reg  <= data_i[10];
    end 
    if(N3660) begin
      \nz.mem_409_sv2v_reg  <= data_i[9];
    end 
    if(N3659) begin
      \nz.mem_408_sv2v_reg  <= data_i[8];
    end 
    if(N3658) begin
      \nz.mem_407_sv2v_reg  <= data_i[7];
    end 
    if(N3657) begin
      \nz.mem_406_sv2v_reg  <= data_i[6];
    end 
    if(N3656) begin
      \nz.mem_405_sv2v_reg  <= data_i[5];
    end 
    if(N3655) begin
      \nz.mem_404_sv2v_reg  <= data_i[4];
    end 
    if(N3654) begin
      \nz.mem_403_sv2v_reg  <= data_i[3];
    end 
    if(N3653) begin
      \nz.mem_402_sv2v_reg  <= data_i[2];
    end 
    if(N3652) begin
      \nz.mem_401_sv2v_reg  <= data_i[1];
    end 
    if(N3651) begin
      \nz.mem_400_sv2v_reg  <= data_i[0];
    end 
    if(N3650) begin
      \nz.mem_399_sv2v_reg  <= data_i[39];
    end 
    if(N3649) begin
      \nz.mem_398_sv2v_reg  <= data_i[38];
    end 
    if(N3648) begin
      \nz.mem_397_sv2v_reg  <= data_i[37];
    end 
    if(N3647) begin
      \nz.mem_396_sv2v_reg  <= data_i[36];
    end 
    if(N3646) begin
      \nz.mem_395_sv2v_reg  <= data_i[35];
    end 
    if(N3645) begin
      \nz.mem_394_sv2v_reg  <= data_i[34];
    end 
    if(N3644) begin
      \nz.mem_393_sv2v_reg  <= data_i[33];
    end 
    if(N3643) begin
      \nz.mem_392_sv2v_reg  <= data_i[32];
    end 
    if(N3642) begin
      \nz.mem_391_sv2v_reg  <= data_i[31];
    end 
    if(N3641) begin
      \nz.mem_390_sv2v_reg  <= data_i[30];
    end 
    if(N3640) begin
      \nz.mem_389_sv2v_reg  <= data_i[29];
    end 
    if(N3639) begin
      \nz.mem_388_sv2v_reg  <= data_i[28];
    end 
    if(N3638) begin
      \nz.mem_387_sv2v_reg  <= data_i[27];
    end 
    if(N3637) begin
      \nz.mem_386_sv2v_reg  <= data_i[26];
    end 
    if(N3636) begin
      \nz.mem_385_sv2v_reg  <= data_i[25];
    end 
    if(N3635) begin
      \nz.mem_384_sv2v_reg  <= data_i[24];
    end 
    if(N3634) begin
      \nz.mem_383_sv2v_reg  <= data_i[23];
    end 
    if(N3633) begin
      \nz.mem_382_sv2v_reg  <= data_i[22];
    end 
    if(N3632) begin
      \nz.mem_381_sv2v_reg  <= data_i[21];
    end 
    if(N3631) begin
      \nz.mem_380_sv2v_reg  <= data_i[20];
    end 
    if(N3630) begin
      \nz.mem_379_sv2v_reg  <= data_i[19];
    end 
    if(N3629) begin
      \nz.mem_378_sv2v_reg  <= data_i[18];
    end 
    if(N3628) begin
      \nz.mem_377_sv2v_reg  <= data_i[17];
    end 
    if(N3627) begin
      \nz.mem_376_sv2v_reg  <= data_i[16];
    end 
    if(N3626) begin
      \nz.mem_375_sv2v_reg  <= data_i[15];
    end 
    if(N3625) begin
      \nz.mem_374_sv2v_reg  <= data_i[14];
    end 
    if(N3624) begin
      \nz.mem_373_sv2v_reg  <= data_i[13];
    end 
    if(N3623) begin
      \nz.mem_372_sv2v_reg  <= data_i[12];
    end 
    if(N3622) begin
      \nz.mem_371_sv2v_reg  <= data_i[11];
    end 
    if(N3621) begin
      \nz.mem_370_sv2v_reg  <= data_i[10];
    end 
    if(N3620) begin
      \nz.mem_369_sv2v_reg  <= data_i[9];
    end 
    if(N3619) begin
      \nz.mem_368_sv2v_reg  <= data_i[8];
    end 
    if(N3618) begin
      \nz.mem_367_sv2v_reg  <= data_i[7];
    end 
    if(N3617) begin
      \nz.mem_366_sv2v_reg  <= data_i[6];
    end 
    if(N3616) begin
      \nz.mem_365_sv2v_reg  <= data_i[5];
    end 
    if(N3615) begin
      \nz.mem_364_sv2v_reg  <= data_i[4];
    end 
    if(N3614) begin
      \nz.mem_363_sv2v_reg  <= data_i[3];
    end 
    if(N3613) begin
      \nz.mem_362_sv2v_reg  <= data_i[2];
    end 
    if(N3612) begin
      \nz.mem_361_sv2v_reg  <= data_i[1];
    end 
    if(N3611) begin
      \nz.mem_360_sv2v_reg  <= data_i[0];
    end 
    if(N3610) begin
      \nz.mem_359_sv2v_reg  <= data_i[39];
    end 
    if(N3609) begin
      \nz.mem_358_sv2v_reg  <= data_i[38];
    end 
    if(N3608) begin
      \nz.mem_357_sv2v_reg  <= data_i[37];
    end 
    if(N3607) begin
      \nz.mem_356_sv2v_reg  <= data_i[36];
    end 
    if(N3606) begin
      \nz.mem_355_sv2v_reg  <= data_i[35];
    end 
    if(N3605) begin
      \nz.mem_354_sv2v_reg  <= data_i[34];
    end 
    if(N3604) begin
      \nz.mem_353_sv2v_reg  <= data_i[33];
    end 
    if(N3603) begin
      \nz.mem_352_sv2v_reg  <= data_i[32];
    end 
    if(N3602) begin
      \nz.mem_351_sv2v_reg  <= data_i[31];
    end 
    if(N3601) begin
      \nz.mem_350_sv2v_reg  <= data_i[30];
    end 
    if(N3600) begin
      \nz.mem_349_sv2v_reg  <= data_i[29];
    end 
    if(N3599) begin
      \nz.mem_348_sv2v_reg  <= data_i[28];
    end 
    if(N3598) begin
      \nz.mem_347_sv2v_reg  <= data_i[27];
    end 
    if(N3597) begin
      \nz.mem_346_sv2v_reg  <= data_i[26];
    end 
    if(N3596) begin
      \nz.mem_345_sv2v_reg  <= data_i[25];
    end 
    if(N3595) begin
      \nz.mem_344_sv2v_reg  <= data_i[24];
    end 
    if(N3594) begin
      \nz.mem_343_sv2v_reg  <= data_i[23];
    end 
    if(N3593) begin
      \nz.mem_342_sv2v_reg  <= data_i[22];
    end 
    if(N3592) begin
      \nz.mem_341_sv2v_reg  <= data_i[21];
    end 
    if(N3591) begin
      \nz.mem_340_sv2v_reg  <= data_i[20];
    end 
    if(N3590) begin
      \nz.mem_339_sv2v_reg  <= data_i[19];
    end 
    if(N3589) begin
      \nz.mem_338_sv2v_reg  <= data_i[18];
    end 
    if(N3588) begin
      \nz.mem_337_sv2v_reg  <= data_i[17];
    end 
    if(N3587) begin
      \nz.mem_336_sv2v_reg  <= data_i[16];
    end 
    if(N3586) begin
      \nz.mem_335_sv2v_reg  <= data_i[15];
    end 
    if(N3585) begin
      \nz.mem_334_sv2v_reg  <= data_i[14];
    end 
    if(N3584) begin
      \nz.mem_333_sv2v_reg  <= data_i[13];
    end 
    if(N3583) begin
      \nz.mem_332_sv2v_reg  <= data_i[12];
    end 
    if(N3582) begin
      \nz.mem_331_sv2v_reg  <= data_i[11];
    end 
    if(N3581) begin
      \nz.mem_330_sv2v_reg  <= data_i[10];
    end 
    if(N3580) begin
      \nz.mem_329_sv2v_reg  <= data_i[9];
    end 
    if(N3579) begin
      \nz.mem_328_sv2v_reg  <= data_i[8];
    end 
    if(N3578) begin
      \nz.mem_327_sv2v_reg  <= data_i[7];
    end 
    if(N3577) begin
      \nz.mem_326_sv2v_reg  <= data_i[6];
    end 
    if(N3576) begin
      \nz.mem_325_sv2v_reg  <= data_i[5];
    end 
    if(N3575) begin
      \nz.mem_324_sv2v_reg  <= data_i[4];
    end 
    if(N3574) begin
      \nz.mem_323_sv2v_reg  <= data_i[3];
    end 
    if(N3573) begin
      \nz.mem_322_sv2v_reg  <= data_i[2];
    end 
    if(N3572) begin
      \nz.mem_321_sv2v_reg  <= data_i[1];
    end 
    if(N3571) begin
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N3570) begin
      \nz.mem_319_sv2v_reg  <= data_i[39];
    end 
    if(N3569) begin
      \nz.mem_318_sv2v_reg  <= data_i[38];
    end 
    if(N3568) begin
      \nz.mem_317_sv2v_reg  <= data_i[37];
    end 
    if(N3567) begin
      \nz.mem_316_sv2v_reg  <= data_i[36];
    end 
    if(N3566) begin
      \nz.mem_315_sv2v_reg  <= data_i[35];
    end 
    if(N3565) begin
      \nz.mem_314_sv2v_reg  <= data_i[34];
    end 
    if(N3564) begin
      \nz.mem_313_sv2v_reg  <= data_i[33];
    end 
    if(N3563) begin
      \nz.mem_312_sv2v_reg  <= data_i[32];
    end 
    if(N3562) begin
      \nz.mem_311_sv2v_reg  <= data_i[31];
    end 
    if(N3561) begin
      \nz.mem_310_sv2v_reg  <= data_i[30];
    end 
    if(N3560) begin
      \nz.mem_309_sv2v_reg  <= data_i[29];
    end 
    if(N3559) begin
      \nz.mem_308_sv2v_reg  <= data_i[28];
    end 
    if(N3558) begin
      \nz.mem_307_sv2v_reg  <= data_i[27];
    end 
    if(N3557) begin
      \nz.mem_306_sv2v_reg  <= data_i[26];
    end 
    if(N3556) begin
      \nz.mem_305_sv2v_reg  <= data_i[25];
    end 
    if(N3555) begin
      \nz.mem_304_sv2v_reg  <= data_i[24];
    end 
    if(N3554) begin
      \nz.mem_303_sv2v_reg  <= data_i[23];
    end 
    if(N3553) begin
      \nz.mem_302_sv2v_reg  <= data_i[22];
    end 
    if(N3552) begin
      \nz.mem_301_sv2v_reg  <= data_i[21];
    end 
    if(N3551) begin
      \nz.mem_300_sv2v_reg  <= data_i[20];
    end 
    if(N3550) begin
      \nz.mem_299_sv2v_reg  <= data_i[19];
    end 
    if(N3549) begin
      \nz.mem_298_sv2v_reg  <= data_i[18];
    end 
    if(N3548) begin
      \nz.mem_297_sv2v_reg  <= data_i[17];
    end 
    if(N3547) begin
      \nz.mem_296_sv2v_reg  <= data_i[16];
    end 
    if(N3546) begin
      \nz.mem_295_sv2v_reg  <= data_i[15];
    end 
    if(N3545) begin
      \nz.mem_294_sv2v_reg  <= data_i[14];
    end 
    if(N3544) begin
      \nz.mem_293_sv2v_reg  <= data_i[13];
    end 
    if(N3543) begin
      \nz.mem_292_sv2v_reg  <= data_i[12];
    end 
    if(N3542) begin
      \nz.mem_291_sv2v_reg  <= data_i[11];
    end 
    if(N3541) begin
      \nz.mem_290_sv2v_reg  <= data_i[10];
    end 
    if(N3540) begin
      \nz.mem_289_sv2v_reg  <= data_i[9];
    end 
    if(N3539) begin
      \nz.mem_288_sv2v_reg  <= data_i[8];
    end 
    if(N3538) begin
      \nz.mem_287_sv2v_reg  <= data_i[7];
    end 
    if(N3537) begin
      \nz.mem_286_sv2v_reg  <= data_i[6];
    end 
    if(N3536) begin
      \nz.mem_285_sv2v_reg  <= data_i[5];
    end 
    if(N3535) begin
      \nz.mem_284_sv2v_reg  <= data_i[4];
    end 
    if(N3534) begin
      \nz.mem_283_sv2v_reg  <= data_i[3];
    end 
    if(N3533) begin
      \nz.mem_282_sv2v_reg  <= data_i[2];
    end 
    if(N3532) begin
      \nz.mem_281_sv2v_reg  <= data_i[1];
    end 
    if(N3531) begin
      \nz.mem_280_sv2v_reg  <= data_i[0];
    end 
    if(N3530) begin
      \nz.mem_279_sv2v_reg  <= data_i[39];
    end 
    if(N3529) begin
      \nz.mem_278_sv2v_reg  <= data_i[38];
    end 
    if(N3528) begin
      \nz.mem_277_sv2v_reg  <= data_i[37];
    end 
    if(N3527) begin
      \nz.mem_276_sv2v_reg  <= data_i[36];
    end 
    if(N3526) begin
      \nz.mem_275_sv2v_reg  <= data_i[35];
    end 
    if(N3525) begin
      \nz.mem_274_sv2v_reg  <= data_i[34];
    end 
    if(N3524) begin
      \nz.mem_273_sv2v_reg  <= data_i[33];
    end 
    if(N3523) begin
      \nz.mem_272_sv2v_reg  <= data_i[32];
    end 
    if(N3522) begin
      \nz.mem_271_sv2v_reg  <= data_i[31];
    end 
    if(N3521) begin
      \nz.mem_270_sv2v_reg  <= data_i[30];
    end 
    if(N3520) begin
      \nz.mem_269_sv2v_reg  <= data_i[29];
    end 
    if(N3519) begin
      \nz.mem_268_sv2v_reg  <= data_i[28];
    end 
    if(N3518) begin
      \nz.mem_267_sv2v_reg  <= data_i[27];
    end 
    if(N3517) begin
      \nz.mem_266_sv2v_reg  <= data_i[26];
    end 
    if(N3516) begin
      \nz.mem_265_sv2v_reg  <= data_i[25];
    end 
    if(N3515) begin
      \nz.mem_264_sv2v_reg  <= data_i[24];
    end 
    if(N3514) begin
      \nz.mem_263_sv2v_reg  <= data_i[23];
    end 
    if(N3513) begin
      \nz.mem_262_sv2v_reg  <= data_i[22];
    end 
    if(N3512) begin
      \nz.mem_261_sv2v_reg  <= data_i[21];
    end 
    if(N3511) begin
      \nz.mem_260_sv2v_reg  <= data_i[20];
    end 
    if(N3510) begin
      \nz.mem_259_sv2v_reg  <= data_i[19];
    end 
    if(N3509) begin
      \nz.mem_258_sv2v_reg  <= data_i[18];
    end 
    if(N3508) begin
      \nz.mem_257_sv2v_reg  <= data_i[17];
    end 
    if(N3507) begin
      \nz.mem_256_sv2v_reg  <= data_i[16];
    end 
    if(N3506) begin
      \nz.mem_255_sv2v_reg  <= data_i[15];
    end 
    if(N3505) begin
      \nz.mem_254_sv2v_reg  <= data_i[14];
    end 
    if(N3504) begin
      \nz.mem_253_sv2v_reg  <= data_i[13];
    end 
    if(N3503) begin
      \nz.mem_252_sv2v_reg  <= data_i[12];
    end 
    if(N3502) begin
      \nz.mem_251_sv2v_reg  <= data_i[11];
    end 
    if(N3501) begin
      \nz.mem_250_sv2v_reg  <= data_i[10];
    end 
    if(N3500) begin
      \nz.mem_249_sv2v_reg  <= data_i[9];
    end 
    if(N3499) begin
      \nz.mem_248_sv2v_reg  <= data_i[8];
    end 
    if(N3498) begin
      \nz.mem_247_sv2v_reg  <= data_i[7];
    end 
    if(N3497) begin
      \nz.mem_246_sv2v_reg  <= data_i[6];
    end 
    if(N3496) begin
      \nz.mem_245_sv2v_reg  <= data_i[5];
    end 
    if(N3495) begin
      \nz.mem_244_sv2v_reg  <= data_i[4];
    end 
    if(N3494) begin
      \nz.mem_243_sv2v_reg  <= data_i[3];
    end 
    if(N3493) begin
      \nz.mem_242_sv2v_reg  <= data_i[2];
    end 
    if(N3492) begin
      \nz.mem_241_sv2v_reg  <= data_i[1];
    end 
    if(N3491) begin
      \nz.mem_240_sv2v_reg  <= data_i[0];
    end 
    if(N3490) begin
      \nz.mem_239_sv2v_reg  <= data_i[39];
    end 
    if(N3489) begin
      \nz.mem_238_sv2v_reg  <= data_i[38];
    end 
    if(N3488) begin
      \nz.mem_237_sv2v_reg  <= data_i[37];
    end 
    if(N3487) begin
      \nz.mem_236_sv2v_reg  <= data_i[36];
    end 
    if(N3486) begin
      \nz.mem_235_sv2v_reg  <= data_i[35];
    end 
    if(N3485) begin
      \nz.mem_234_sv2v_reg  <= data_i[34];
    end 
    if(N3484) begin
      \nz.mem_233_sv2v_reg  <= data_i[33];
    end 
    if(N3483) begin
      \nz.mem_232_sv2v_reg  <= data_i[32];
    end 
    if(N3482) begin
      \nz.mem_231_sv2v_reg  <= data_i[31];
    end 
    if(N3481) begin
      \nz.mem_230_sv2v_reg  <= data_i[30];
    end 
    if(N3480) begin
      \nz.mem_229_sv2v_reg  <= data_i[29];
    end 
    if(N3479) begin
      \nz.mem_228_sv2v_reg  <= data_i[28];
    end 
    if(N3478) begin
      \nz.mem_227_sv2v_reg  <= data_i[27];
    end 
    if(N3477) begin
      \nz.mem_226_sv2v_reg  <= data_i[26];
    end 
    if(N3476) begin
      \nz.mem_225_sv2v_reg  <= data_i[25];
    end 
    if(N3475) begin
      \nz.mem_224_sv2v_reg  <= data_i[24];
    end 
    if(N3474) begin
      \nz.mem_223_sv2v_reg  <= data_i[23];
    end 
    if(N3473) begin
      \nz.mem_222_sv2v_reg  <= data_i[22];
    end 
    if(N3472) begin
      \nz.mem_221_sv2v_reg  <= data_i[21];
    end 
    if(N3471) begin
      \nz.mem_220_sv2v_reg  <= data_i[20];
    end 
    if(N3470) begin
      \nz.mem_219_sv2v_reg  <= data_i[19];
    end 
    if(N3469) begin
      \nz.mem_218_sv2v_reg  <= data_i[18];
    end 
    if(N3468) begin
      \nz.mem_217_sv2v_reg  <= data_i[17];
    end 
    if(N3467) begin
      \nz.mem_216_sv2v_reg  <= data_i[16];
    end 
    if(N3466) begin
      \nz.mem_215_sv2v_reg  <= data_i[15];
    end 
    if(N3465) begin
      \nz.mem_214_sv2v_reg  <= data_i[14];
    end 
    if(N3464) begin
      \nz.mem_213_sv2v_reg  <= data_i[13];
    end 
    if(N3463) begin
      \nz.mem_212_sv2v_reg  <= data_i[12];
    end 
    if(N3462) begin
      \nz.mem_211_sv2v_reg  <= data_i[11];
    end 
    if(N3461) begin
      \nz.mem_210_sv2v_reg  <= data_i[10];
    end 
    if(N3460) begin
      \nz.mem_209_sv2v_reg  <= data_i[9];
    end 
    if(N3459) begin
      \nz.mem_208_sv2v_reg  <= data_i[8];
    end 
    if(N3458) begin
      \nz.mem_207_sv2v_reg  <= data_i[7];
    end 
    if(N3457) begin
      \nz.mem_206_sv2v_reg  <= data_i[6];
    end 
    if(N3456) begin
      \nz.mem_205_sv2v_reg  <= data_i[5];
    end 
    if(N3455) begin
      \nz.mem_204_sv2v_reg  <= data_i[4];
    end 
    if(N3454) begin
      \nz.mem_203_sv2v_reg  <= data_i[3];
    end 
    if(N3453) begin
      \nz.mem_202_sv2v_reg  <= data_i[2];
    end 
    if(N3452) begin
      \nz.mem_201_sv2v_reg  <= data_i[1];
    end 
    if(N3451) begin
      \nz.mem_200_sv2v_reg  <= data_i[0];
    end 
    if(N3450) begin
      \nz.mem_199_sv2v_reg  <= data_i[39];
    end 
    if(N3449) begin
      \nz.mem_198_sv2v_reg  <= data_i[38];
    end 
    if(N3448) begin
      \nz.mem_197_sv2v_reg  <= data_i[37];
    end 
    if(N3447) begin
      \nz.mem_196_sv2v_reg  <= data_i[36];
    end 
    if(N3446) begin
      \nz.mem_195_sv2v_reg  <= data_i[35];
    end 
    if(N3445) begin
      \nz.mem_194_sv2v_reg  <= data_i[34];
    end 
    if(N3444) begin
      \nz.mem_193_sv2v_reg  <= data_i[33];
    end 
    if(N3443) begin
      \nz.mem_192_sv2v_reg  <= data_i[32];
    end 
    if(N3442) begin
      \nz.mem_191_sv2v_reg  <= data_i[31];
    end 
    if(N3441) begin
      \nz.mem_190_sv2v_reg  <= data_i[30];
    end 
    if(N3440) begin
      \nz.mem_189_sv2v_reg  <= data_i[29];
    end 
    if(N3439) begin
      \nz.mem_188_sv2v_reg  <= data_i[28];
    end 
    if(N3438) begin
      \nz.mem_187_sv2v_reg  <= data_i[27];
    end 
    if(N3437) begin
      \nz.mem_186_sv2v_reg  <= data_i[26];
    end 
    if(N3436) begin
      \nz.mem_185_sv2v_reg  <= data_i[25];
    end 
    if(N3435) begin
      \nz.mem_184_sv2v_reg  <= data_i[24];
    end 
    if(N3434) begin
      \nz.mem_183_sv2v_reg  <= data_i[23];
    end 
    if(N3433) begin
      \nz.mem_182_sv2v_reg  <= data_i[22];
    end 
    if(N3432) begin
      \nz.mem_181_sv2v_reg  <= data_i[21];
    end 
    if(N3431) begin
      \nz.mem_180_sv2v_reg  <= data_i[20];
    end 
    if(N3430) begin
      \nz.mem_179_sv2v_reg  <= data_i[19];
    end 
    if(N3429) begin
      \nz.mem_178_sv2v_reg  <= data_i[18];
    end 
    if(N3428) begin
      \nz.mem_177_sv2v_reg  <= data_i[17];
    end 
    if(N3427) begin
      \nz.mem_176_sv2v_reg  <= data_i[16];
    end 
    if(N3426) begin
      \nz.mem_175_sv2v_reg  <= data_i[15];
    end 
    if(N3425) begin
      \nz.mem_174_sv2v_reg  <= data_i[14];
    end 
    if(N3424) begin
      \nz.mem_173_sv2v_reg  <= data_i[13];
    end 
    if(N3423) begin
      \nz.mem_172_sv2v_reg  <= data_i[12];
    end 
    if(N3422) begin
      \nz.mem_171_sv2v_reg  <= data_i[11];
    end 
    if(N3421) begin
      \nz.mem_170_sv2v_reg  <= data_i[10];
    end 
    if(N3420) begin
      \nz.mem_169_sv2v_reg  <= data_i[9];
    end 
    if(N3419) begin
      \nz.mem_168_sv2v_reg  <= data_i[8];
    end 
    if(N3418) begin
      \nz.mem_167_sv2v_reg  <= data_i[7];
    end 
    if(N3417) begin
      \nz.mem_166_sv2v_reg  <= data_i[6];
    end 
    if(N3416) begin
      \nz.mem_165_sv2v_reg  <= data_i[5];
    end 
    if(N3415) begin
      \nz.mem_164_sv2v_reg  <= data_i[4];
    end 
    if(N3414) begin
      \nz.mem_163_sv2v_reg  <= data_i[3];
    end 
    if(N3413) begin
      \nz.mem_162_sv2v_reg  <= data_i[2];
    end 
    if(N3412) begin
      \nz.mem_161_sv2v_reg  <= data_i[1];
    end 
    if(N3411) begin
      \nz.mem_160_sv2v_reg  <= data_i[0];
    end 
    if(N3410) begin
      \nz.mem_159_sv2v_reg  <= data_i[39];
    end 
    if(N3409) begin
      \nz.mem_158_sv2v_reg  <= data_i[38];
    end 
    if(N3408) begin
      \nz.mem_157_sv2v_reg  <= data_i[37];
    end 
    if(N3407) begin
      \nz.mem_156_sv2v_reg  <= data_i[36];
    end 
    if(N3406) begin
      \nz.mem_155_sv2v_reg  <= data_i[35];
    end 
    if(N3405) begin
      \nz.mem_154_sv2v_reg  <= data_i[34];
    end 
    if(N3404) begin
      \nz.mem_153_sv2v_reg  <= data_i[33];
    end 
    if(N3403) begin
      \nz.mem_152_sv2v_reg  <= data_i[32];
    end 
    if(N3402) begin
      \nz.mem_151_sv2v_reg  <= data_i[31];
    end 
    if(N3401) begin
      \nz.mem_150_sv2v_reg  <= data_i[30];
    end 
    if(N3400) begin
      \nz.mem_149_sv2v_reg  <= data_i[29];
    end 
    if(N3399) begin
      \nz.mem_148_sv2v_reg  <= data_i[28];
    end 
    if(N3398) begin
      \nz.mem_147_sv2v_reg  <= data_i[27];
    end 
    if(N3397) begin
      \nz.mem_146_sv2v_reg  <= data_i[26];
    end 
    if(N3396) begin
      \nz.mem_145_sv2v_reg  <= data_i[25];
    end 
    if(N3395) begin
      \nz.mem_144_sv2v_reg  <= data_i[24];
    end 
    if(N3394) begin
      \nz.mem_143_sv2v_reg  <= data_i[23];
    end 
    if(N3393) begin
      \nz.mem_142_sv2v_reg  <= data_i[22];
    end 
    if(N3392) begin
      \nz.mem_141_sv2v_reg  <= data_i[21];
    end 
    if(N3391) begin
      \nz.mem_140_sv2v_reg  <= data_i[20];
    end 
    if(N3390) begin
      \nz.mem_139_sv2v_reg  <= data_i[19];
    end 
    if(N3389) begin
      \nz.mem_138_sv2v_reg  <= data_i[18];
    end 
    if(N3388) begin
      \nz.mem_137_sv2v_reg  <= data_i[17];
    end 
    if(N3387) begin
      \nz.mem_136_sv2v_reg  <= data_i[16];
    end 
    if(N3386) begin
      \nz.mem_135_sv2v_reg  <= data_i[15];
    end 
    if(N3385) begin
      \nz.mem_134_sv2v_reg  <= data_i[14];
    end 
    if(N3384) begin
      \nz.mem_133_sv2v_reg  <= data_i[13];
    end 
    if(N3383) begin
      \nz.mem_132_sv2v_reg  <= data_i[12];
    end 
    if(N3382) begin
      \nz.mem_131_sv2v_reg  <= data_i[11];
    end 
    if(N3381) begin
      \nz.mem_130_sv2v_reg  <= data_i[10];
    end 
    if(N3380) begin
      \nz.mem_129_sv2v_reg  <= data_i[9];
    end 
    if(N3379) begin
      \nz.mem_128_sv2v_reg  <= data_i[8];
    end 
    if(N3378) begin
      \nz.mem_127_sv2v_reg  <= data_i[7];
    end 
    if(N3377) begin
      \nz.mem_126_sv2v_reg  <= data_i[6];
    end 
    if(N3376) begin
      \nz.mem_125_sv2v_reg  <= data_i[5];
    end 
    if(N3375) begin
      \nz.mem_124_sv2v_reg  <= data_i[4];
    end 
    if(N3374) begin
      \nz.mem_123_sv2v_reg  <= data_i[3];
    end 
    if(N3373) begin
      \nz.mem_122_sv2v_reg  <= data_i[2];
    end 
    if(N3372) begin
      \nz.mem_121_sv2v_reg  <= data_i[1];
    end 
    if(N3371) begin
      \nz.mem_120_sv2v_reg  <= data_i[0];
    end 
    if(N3370) begin
      \nz.mem_119_sv2v_reg  <= data_i[39];
    end 
    if(N3369) begin
      \nz.mem_118_sv2v_reg  <= data_i[38];
    end 
    if(N3368) begin
      \nz.mem_117_sv2v_reg  <= data_i[37];
    end 
    if(N3367) begin
      \nz.mem_116_sv2v_reg  <= data_i[36];
    end 
    if(N3366) begin
      \nz.mem_115_sv2v_reg  <= data_i[35];
    end 
    if(N3365) begin
      \nz.mem_114_sv2v_reg  <= data_i[34];
    end 
    if(N3364) begin
      \nz.mem_113_sv2v_reg  <= data_i[33];
    end 
    if(N3363) begin
      \nz.mem_112_sv2v_reg  <= data_i[32];
    end 
    if(N3362) begin
      \nz.mem_111_sv2v_reg  <= data_i[31];
    end 
    if(N3361) begin
      \nz.mem_110_sv2v_reg  <= data_i[30];
    end 
    if(N3360) begin
      \nz.mem_109_sv2v_reg  <= data_i[29];
    end 
    if(N3359) begin
      \nz.mem_108_sv2v_reg  <= data_i[28];
    end 
    if(N3358) begin
      \nz.mem_107_sv2v_reg  <= data_i[27];
    end 
    if(N3357) begin
      \nz.mem_106_sv2v_reg  <= data_i[26];
    end 
    if(N3356) begin
      \nz.mem_105_sv2v_reg  <= data_i[25];
    end 
    if(N3355) begin
      \nz.mem_104_sv2v_reg  <= data_i[24];
    end 
    if(N3354) begin
      \nz.mem_103_sv2v_reg  <= data_i[23];
    end 
    if(N3353) begin
      \nz.mem_102_sv2v_reg  <= data_i[22];
    end 
    if(N3352) begin
      \nz.mem_101_sv2v_reg  <= data_i[21];
    end 
    if(N3351) begin
      \nz.mem_100_sv2v_reg  <= data_i[20];
    end 
    if(N3350) begin
      \nz.mem_99_sv2v_reg  <= data_i[19];
    end 
    if(N3349) begin
      \nz.mem_98_sv2v_reg  <= data_i[18];
    end 
    if(N3348) begin
      \nz.mem_97_sv2v_reg  <= data_i[17];
    end 
    if(N3347) begin
      \nz.mem_96_sv2v_reg  <= data_i[16];
    end 
    if(N3346) begin
      \nz.mem_95_sv2v_reg  <= data_i[15];
    end 
    if(N3345) begin
      \nz.mem_94_sv2v_reg  <= data_i[14];
    end 
    if(N3344) begin
      \nz.mem_93_sv2v_reg  <= data_i[13];
    end 
    if(N3343) begin
      \nz.mem_92_sv2v_reg  <= data_i[12];
    end 
    if(N3342) begin
      \nz.mem_91_sv2v_reg  <= data_i[11];
    end 
    if(N3341) begin
      \nz.mem_90_sv2v_reg  <= data_i[10];
    end 
    if(N3340) begin
      \nz.mem_89_sv2v_reg  <= data_i[9];
    end 
    if(N3339) begin
      \nz.mem_88_sv2v_reg  <= data_i[8];
    end 
    if(N3338) begin
      \nz.mem_87_sv2v_reg  <= data_i[7];
    end 
    if(N3337) begin
      \nz.mem_86_sv2v_reg  <= data_i[6];
    end 
    if(N3336) begin
      \nz.mem_85_sv2v_reg  <= data_i[5];
    end 
    if(N3335) begin
      \nz.mem_84_sv2v_reg  <= data_i[4];
    end 
    if(N3334) begin
      \nz.mem_83_sv2v_reg  <= data_i[3];
    end 
    if(N3333) begin
      \nz.mem_82_sv2v_reg  <= data_i[2];
    end 
    if(N3332) begin
      \nz.mem_81_sv2v_reg  <= data_i[1];
    end 
    if(N3331) begin
      \nz.mem_80_sv2v_reg  <= data_i[0];
    end 
    if(N3330) begin
      \nz.mem_79_sv2v_reg  <= data_i[39];
    end 
    if(N3329) begin
      \nz.mem_78_sv2v_reg  <= data_i[38];
    end 
    if(N3328) begin
      \nz.mem_77_sv2v_reg  <= data_i[37];
    end 
    if(N3327) begin
      \nz.mem_76_sv2v_reg  <= data_i[36];
    end 
    if(N3326) begin
      \nz.mem_75_sv2v_reg  <= data_i[35];
    end 
    if(N3325) begin
      \nz.mem_74_sv2v_reg  <= data_i[34];
    end 
    if(N3324) begin
      \nz.mem_73_sv2v_reg  <= data_i[33];
    end 
    if(N3323) begin
      \nz.mem_72_sv2v_reg  <= data_i[32];
    end 
    if(N3322) begin
      \nz.mem_71_sv2v_reg  <= data_i[31];
    end 
    if(N3321) begin
      \nz.mem_70_sv2v_reg  <= data_i[30];
    end 
    if(N3320) begin
      \nz.mem_69_sv2v_reg  <= data_i[29];
    end 
    if(N3319) begin
      \nz.mem_68_sv2v_reg  <= data_i[28];
    end 
    if(N3318) begin
      \nz.mem_67_sv2v_reg  <= data_i[27];
    end 
    if(N3317) begin
      \nz.mem_66_sv2v_reg  <= data_i[26];
    end 
    if(N3316) begin
      \nz.mem_65_sv2v_reg  <= data_i[25];
    end 
    if(N3315) begin
      \nz.mem_64_sv2v_reg  <= data_i[24];
    end 
    if(N3314) begin
      \nz.mem_63_sv2v_reg  <= data_i[23];
    end 
    if(N3313) begin
      \nz.mem_62_sv2v_reg  <= data_i[22];
    end 
    if(N3312) begin
      \nz.mem_61_sv2v_reg  <= data_i[21];
    end 
    if(N3311) begin
      \nz.mem_60_sv2v_reg  <= data_i[20];
    end 
    if(N3310) begin
      \nz.mem_59_sv2v_reg  <= data_i[19];
    end 
    if(N3309) begin
      \nz.mem_58_sv2v_reg  <= data_i[18];
    end 
    if(N3308) begin
      \nz.mem_57_sv2v_reg  <= data_i[17];
    end 
    if(N3307) begin
      \nz.mem_56_sv2v_reg  <= data_i[16];
    end 
    if(N3306) begin
      \nz.mem_55_sv2v_reg  <= data_i[15];
    end 
    if(N3305) begin
      \nz.mem_54_sv2v_reg  <= data_i[14];
    end 
    if(N3304) begin
      \nz.mem_53_sv2v_reg  <= data_i[13];
    end 
    if(N3303) begin
      \nz.mem_52_sv2v_reg  <= data_i[12];
    end 
    if(N3302) begin
      \nz.mem_51_sv2v_reg  <= data_i[11];
    end 
    if(N3301) begin
      \nz.mem_50_sv2v_reg  <= data_i[10];
    end 
    if(N3300) begin
      \nz.mem_49_sv2v_reg  <= data_i[9];
    end 
    if(N3299) begin
      \nz.mem_48_sv2v_reg  <= data_i[8];
    end 
    if(N3298) begin
      \nz.mem_47_sv2v_reg  <= data_i[7];
    end 
    if(N3297) begin
      \nz.mem_46_sv2v_reg  <= data_i[6];
    end 
    if(N3296) begin
      \nz.mem_45_sv2v_reg  <= data_i[5];
    end 
    if(N3295) begin
      \nz.mem_44_sv2v_reg  <= data_i[4];
    end 
    if(N3294) begin
      \nz.mem_43_sv2v_reg  <= data_i[3];
    end 
    if(N3293) begin
      \nz.mem_42_sv2v_reg  <= data_i[2];
    end 
    if(N3292) begin
      \nz.mem_41_sv2v_reg  <= data_i[1];
    end 
    if(N3291) begin
      \nz.mem_40_sv2v_reg  <= data_i[0];
    end 
    if(N3290) begin
      \nz.mem_39_sv2v_reg  <= data_i[39];
    end 
    if(N3289) begin
      \nz.mem_38_sv2v_reg  <= data_i[38];
    end 
    if(N3288) begin
      \nz.mem_37_sv2v_reg  <= data_i[37];
    end 
    if(N3287) begin
      \nz.mem_36_sv2v_reg  <= data_i[36];
    end 
    if(N3286) begin
      \nz.mem_35_sv2v_reg  <= data_i[35];
    end 
    if(N3285) begin
      \nz.mem_34_sv2v_reg  <= data_i[34];
    end 
    if(N3284) begin
      \nz.mem_33_sv2v_reg  <= data_i[33];
    end 
    if(N3283) begin
      \nz.mem_32_sv2v_reg  <= data_i[32];
    end 
    if(N3282) begin
      \nz.mem_31_sv2v_reg  <= data_i[31];
    end 
    if(N3281) begin
      \nz.mem_30_sv2v_reg  <= data_i[30];
    end 
    if(N3280) begin
      \nz.mem_29_sv2v_reg  <= data_i[29];
    end 
    if(N3279) begin
      \nz.mem_28_sv2v_reg  <= data_i[28];
    end 
    if(N3278) begin
      \nz.mem_27_sv2v_reg  <= data_i[27];
    end 
    if(N3277) begin
      \nz.mem_26_sv2v_reg  <= data_i[26];
    end 
    if(N3276) begin
      \nz.mem_25_sv2v_reg  <= data_i[25];
    end 
    if(N3275) begin
      \nz.mem_24_sv2v_reg  <= data_i[24];
    end 
    if(N3274) begin
      \nz.mem_23_sv2v_reg  <= data_i[23];
    end 
    if(N3273) begin
      \nz.mem_22_sv2v_reg  <= data_i[22];
    end 
    if(N3272) begin
      \nz.mem_21_sv2v_reg  <= data_i[21];
    end 
    if(N3271) begin
      \nz.mem_20_sv2v_reg  <= data_i[20];
    end 
    if(N3270) begin
      \nz.mem_19_sv2v_reg  <= data_i[19];
    end 
    if(N3269) begin
      \nz.mem_18_sv2v_reg  <= data_i[18];
    end 
    if(N3268) begin
      \nz.mem_17_sv2v_reg  <= data_i[17];
    end 
    if(N3267) begin
      \nz.mem_16_sv2v_reg  <= data_i[16];
    end 
    if(N3266) begin
      \nz.mem_15_sv2v_reg  <= data_i[15];
    end 
    if(N3265) begin
      \nz.mem_14_sv2v_reg  <= data_i[14];
    end 
    if(N3264) begin
      \nz.mem_13_sv2v_reg  <= data_i[13];
    end 
    if(N3263) begin
      \nz.mem_12_sv2v_reg  <= data_i[12];
    end 
    if(N3262) begin
      \nz.mem_11_sv2v_reg  <= data_i[11];
    end 
    if(N3261) begin
      \nz.mem_10_sv2v_reg  <= data_i[10];
    end 
    if(N3260) begin
      \nz.mem_9_sv2v_reg  <= data_i[9];
    end 
    if(N3259) begin
      \nz.mem_8_sv2v_reg  <= data_i[8];
    end 
    if(N3258) begin
      \nz.mem_7_sv2v_reg  <= data_i[7];
    end 
    if(N3257) begin
      \nz.mem_6_sv2v_reg  <= data_i[6];
    end 
    if(N3256) begin
      \nz.mem_5_sv2v_reg  <= data_i[5];
    end 
    if(N3255) begin
      \nz.mem_4_sv2v_reg  <= data_i[4];
    end 
    if(N3254) begin
      \nz.mem_3_sv2v_reg  <= data_i[3];
    end 
    if(N3253) begin
      \nz.mem_2_sv2v_reg  <= data_i[2];
    end 
    if(N3252) begin
      \nz.mem_1_sv2v_reg  <= data_i[1];
    end 
    if(N3251) begin
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p40_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [39:0] data_i;
  input [5:0] addr_i;
  input [39:0] w_mask_i;
  output [39:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [39:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p40_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_dff_en_width_p8_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  wire [7:0] data_o;
  reg data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_7_sv2v_reg <= data_i[7];
      data_o_6_sv2v_reg <= data_i[6];
      data_o_5_sv2v_reg <= data_i[5];
      data_o_4_sv2v_reg <= data_i[4];
      data_o_3_sv2v_reg <= data_i[3];
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p8
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input en_i;
  wire [7:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p8_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1_verbose_p0
(
  clk_i,
  v_i,
  reset_i,
  data_i,
  addr_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input v_i;
  input reset_i;
  input w_i;
  wire [7:0] data_o,\nz.addr_r ,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,\nz.read_en ,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,
  N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,
  N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,
  N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,
  N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,
  N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,
  N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,
  N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,
  N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,
  N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,
  N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,
  N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
  N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,
  N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,
  N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,
  N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,
  N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,
  N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,
  N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,
  N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,
  N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,
  N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,
  N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,
  N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,
  N531,N532,\nz.llr.read_en_r ,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095;
  wire [2047:0] \nz.mem ;
  reg \nz.addr_r_7_sv2v_reg ,\nz.addr_r_6_sv2v_reg ,\nz.addr_r_5_sv2v_reg ,
  \nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,\nz.addr_r_2_sv2v_reg ,
  \nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,\nz.mem_2047_sv2v_reg ,\nz.mem_2046_sv2v_reg ,
  \nz.mem_2045_sv2v_reg ,\nz.mem_2044_sv2v_reg ,\nz.mem_2043_sv2v_reg ,
  \nz.mem_2042_sv2v_reg ,\nz.mem_2041_sv2v_reg ,\nz.mem_2040_sv2v_reg ,\nz.mem_2039_sv2v_reg ,
  \nz.mem_2038_sv2v_reg ,\nz.mem_2037_sv2v_reg ,\nz.mem_2036_sv2v_reg ,
  \nz.mem_2035_sv2v_reg ,\nz.mem_2034_sv2v_reg ,\nz.mem_2033_sv2v_reg ,\nz.mem_2032_sv2v_reg ,
  \nz.mem_2031_sv2v_reg ,\nz.mem_2030_sv2v_reg ,\nz.mem_2029_sv2v_reg ,
  \nz.mem_2028_sv2v_reg ,\nz.mem_2027_sv2v_reg ,\nz.mem_2026_sv2v_reg ,\nz.mem_2025_sv2v_reg ,
  \nz.mem_2024_sv2v_reg ,\nz.mem_2023_sv2v_reg ,\nz.mem_2022_sv2v_reg ,
  \nz.mem_2021_sv2v_reg ,\nz.mem_2020_sv2v_reg ,\nz.mem_2019_sv2v_reg ,\nz.mem_2018_sv2v_reg ,
  \nz.mem_2017_sv2v_reg ,\nz.mem_2016_sv2v_reg ,\nz.mem_2015_sv2v_reg ,
  \nz.mem_2014_sv2v_reg ,\nz.mem_2013_sv2v_reg ,\nz.mem_2012_sv2v_reg ,\nz.mem_2011_sv2v_reg ,
  \nz.mem_2010_sv2v_reg ,\nz.mem_2009_sv2v_reg ,\nz.mem_2008_sv2v_reg ,
  \nz.mem_2007_sv2v_reg ,\nz.mem_2006_sv2v_reg ,\nz.mem_2005_sv2v_reg ,\nz.mem_2004_sv2v_reg ,
  \nz.mem_2003_sv2v_reg ,\nz.mem_2002_sv2v_reg ,\nz.mem_2001_sv2v_reg ,
  \nz.mem_2000_sv2v_reg ,\nz.mem_1999_sv2v_reg ,\nz.mem_1998_sv2v_reg ,\nz.mem_1997_sv2v_reg ,
  \nz.mem_1996_sv2v_reg ,\nz.mem_1995_sv2v_reg ,\nz.mem_1994_sv2v_reg ,
  \nz.mem_1993_sv2v_reg ,\nz.mem_1992_sv2v_reg ,\nz.mem_1991_sv2v_reg ,\nz.mem_1990_sv2v_reg ,
  \nz.mem_1989_sv2v_reg ,\nz.mem_1988_sv2v_reg ,\nz.mem_1987_sv2v_reg ,
  \nz.mem_1986_sv2v_reg ,\nz.mem_1985_sv2v_reg ,\nz.mem_1984_sv2v_reg ,\nz.mem_1983_sv2v_reg ,
  \nz.mem_1982_sv2v_reg ,\nz.mem_1981_sv2v_reg ,\nz.mem_1980_sv2v_reg ,
  \nz.mem_1979_sv2v_reg ,\nz.mem_1978_sv2v_reg ,\nz.mem_1977_sv2v_reg ,\nz.mem_1976_sv2v_reg ,
  \nz.mem_1975_sv2v_reg ,\nz.mem_1974_sv2v_reg ,\nz.mem_1973_sv2v_reg ,
  \nz.mem_1972_sv2v_reg ,\nz.mem_1971_sv2v_reg ,\nz.mem_1970_sv2v_reg ,
  \nz.mem_1969_sv2v_reg ,\nz.mem_1968_sv2v_reg ,\nz.mem_1967_sv2v_reg ,\nz.mem_1966_sv2v_reg ,
  \nz.mem_1965_sv2v_reg ,\nz.mem_1964_sv2v_reg ,\nz.mem_1963_sv2v_reg ,
  \nz.mem_1962_sv2v_reg ,\nz.mem_1961_sv2v_reg ,\nz.mem_1960_sv2v_reg ,\nz.mem_1959_sv2v_reg ,
  \nz.mem_1958_sv2v_reg ,\nz.mem_1957_sv2v_reg ,\nz.mem_1956_sv2v_reg ,
  \nz.mem_1955_sv2v_reg ,\nz.mem_1954_sv2v_reg ,\nz.mem_1953_sv2v_reg ,\nz.mem_1952_sv2v_reg ,
  \nz.mem_1951_sv2v_reg ,\nz.mem_1950_sv2v_reg ,\nz.mem_1949_sv2v_reg ,
  \nz.mem_1948_sv2v_reg ,\nz.mem_1947_sv2v_reg ,\nz.mem_1946_sv2v_reg ,\nz.mem_1945_sv2v_reg ,
  \nz.mem_1944_sv2v_reg ,\nz.mem_1943_sv2v_reg ,\nz.mem_1942_sv2v_reg ,
  \nz.mem_1941_sv2v_reg ,\nz.mem_1940_sv2v_reg ,\nz.mem_1939_sv2v_reg ,\nz.mem_1938_sv2v_reg ,
  \nz.mem_1937_sv2v_reg ,\nz.mem_1936_sv2v_reg ,\nz.mem_1935_sv2v_reg ,
  \nz.mem_1934_sv2v_reg ,\nz.mem_1933_sv2v_reg ,\nz.mem_1932_sv2v_reg ,\nz.mem_1931_sv2v_reg ,
  \nz.mem_1930_sv2v_reg ,\nz.mem_1929_sv2v_reg ,\nz.mem_1928_sv2v_reg ,
  \nz.mem_1927_sv2v_reg ,\nz.mem_1926_sv2v_reg ,\nz.mem_1925_sv2v_reg ,\nz.mem_1924_sv2v_reg ,
  \nz.mem_1923_sv2v_reg ,\nz.mem_1922_sv2v_reg ,\nz.mem_1921_sv2v_reg ,
  \nz.mem_1920_sv2v_reg ,\nz.mem_1919_sv2v_reg ,\nz.mem_1918_sv2v_reg ,\nz.mem_1917_sv2v_reg ,
  \nz.mem_1916_sv2v_reg ,\nz.mem_1915_sv2v_reg ,\nz.mem_1914_sv2v_reg ,
  \nz.mem_1913_sv2v_reg ,\nz.mem_1912_sv2v_reg ,\nz.mem_1911_sv2v_reg ,\nz.mem_1910_sv2v_reg ,
  \nz.mem_1909_sv2v_reg ,\nz.mem_1908_sv2v_reg ,\nz.mem_1907_sv2v_reg ,
  \nz.mem_1906_sv2v_reg ,\nz.mem_1905_sv2v_reg ,\nz.mem_1904_sv2v_reg ,\nz.mem_1903_sv2v_reg ,
  \nz.mem_1902_sv2v_reg ,\nz.mem_1901_sv2v_reg ,\nz.mem_1900_sv2v_reg ,
  \nz.mem_1899_sv2v_reg ,\nz.mem_1898_sv2v_reg ,\nz.mem_1897_sv2v_reg ,\nz.mem_1896_sv2v_reg ,
  \nz.mem_1895_sv2v_reg ,\nz.mem_1894_sv2v_reg ,\nz.mem_1893_sv2v_reg ,
  \nz.mem_1892_sv2v_reg ,\nz.mem_1891_sv2v_reg ,\nz.mem_1890_sv2v_reg ,
  \nz.mem_1889_sv2v_reg ,\nz.mem_1888_sv2v_reg ,\nz.mem_1887_sv2v_reg ,\nz.mem_1886_sv2v_reg ,
  \nz.mem_1885_sv2v_reg ,\nz.mem_1884_sv2v_reg ,\nz.mem_1883_sv2v_reg ,
  \nz.mem_1882_sv2v_reg ,\nz.mem_1881_sv2v_reg ,\nz.mem_1880_sv2v_reg ,\nz.mem_1879_sv2v_reg ,
  \nz.mem_1878_sv2v_reg ,\nz.mem_1877_sv2v_reg ,\nz.mem_1876_sv2v_reg ,
  \nz.mem_1875_sv2v_reg ,\nz.mem_1874_sv2v_reg ,\nz.mem_1873_sv2v_reg ,\nz.mem_1872_sv2v_reg ,
  \nz.mem_1871_sv2v_reg ,\nz.mem_1870_sv2v_reg ,\nz.mem_1869_sv2v_reg ,
  \nz.mem_1868_sv2v_reg ,\nz.mem_1867_sv2v_reg ,\nz.mem_1866_sv2v_reg ,\nz.mem_1865_sv2v_reg ,
  \nz.mem_1864_sv2v_reg ,\nz.mem_1863_sv2v_reg ,\nz.mem_1862_sv2v_reg ,
  \nz.mem_1861_sv2v_reg ,\nz.mem_1860_sv2v_reg ,\nz.mem_1859_sv2v_reg ,\nz.mem_1858_sv2v_reg ,
  \nz.mem_1857_sv2v_reg ,\nz.mem_1856_sv2v_reg ,\nz.mem_1855_sv2v_reg ,
  \nz.mem_1854_sv2v_reg ,\nz.mem_1853_sv2v_reg ,\nz.mem_1852_sv2v_reg ,\nz.mem_1851_sv2v_reg ,
  \nz.mem_1850_sv2v_reg ,\nz.mem_1849_sv2v_reg ,\nz.mem_1848_sv2v_reg ,
  \nz.mem_1847_sv2v_reg ,\nz.mem_1846_sv2v_reg ,\nz.mem_1845_sv2v_reg ,\nz.mem_1844_sv2v_reg ,
  \nz.mem_1843_sv2v_reg ,\nz.mem_1842_sv2v_reg ,\nz.mem_1841_sv2v_reg ,
  \nz.mem_1840_sv2v_reg ,\nz.mem_1839_sv2v_reg ,\nz.mem_1838_sv2v_reg ,\nz.mem_1837_sv2v_reg ,
  \nz.mem_1836_sv2v_reg ,\nz.mem_1835_sv2v_reg ,\nz.mem_1834_sv2v_reg ,
  \nz.mem_1833_sv2v_reg ,\nz.mem_1832_sv2v_reg ,\nz.mem_1831_sv2v_reg ,\nz.mem_1830_sv2v_reg ,
  \nz.mem_1829_sv2v_reg ,\nz.mem_1828_sv2v_reg ,\nz.mem_1827_sv2v_reg ,
  \nz.mem_1826_sv2v_reg ,\nz.mem_1825_sv2v_reg ,\nz.mem_1824_sv2v_reg ,\nz.mem_1823_sv2v_reg ,
  \nz.mem_1822_sv2v_reg ,\nz.mem_1821_sv2v_reg ,\nz.mem_1820_sv2v_reg ,
  \nz.mem_1819_sv2v_reg ,\nz.mem_1818_sv2v_reg ,\nz.mem_1817_sv2v_reg ,\nz.mem_1816_sv2v_reg ,
  \nz.mem_1815_sv2v_reg ,\nz.mem_1814_sv2v_reg ,\nz.mem_1813_sv2v_reg ,
  \nz.mem_1812_sv2v_reg ,\nz.mem_1811_sv2v_reg ,\nz.mem_1810_sv2v_reg ,
  \nz.mem_1809_sv2v_reg ,\nz.mem_1808_sv2v_reg ,\nz.mem_1807_sv2v_reg ,\nz.mem_1806_sv2v_reg ,
  \nz.mem_1805_sv2v_reg ,\nz.mem_1804_sv2v_reg ,\nz.mem_1803_sv2v_reg ,
  \nz.mem_1802_sv2v_reg ,\nz.mem_1801_sv2v_reg ,\nz.mem_1800_sv2v_reg ,\nz.mem_1799_sv2v_reg ,
  \nz.mem_1798_sv2v_reg ,\nz.mem_1797_sv2v_reg ,\nz.mem_1796_sv2v_reg ,
  \nz.mem_1795_sv2v_reg ,\nz.mem_1794_sv2v_reg ,\nz.mem_1793_sv2v_reg ,\nz.mem_1792_sv2v_reg ,
  \nz.mem_1791_sv2v_reg ,\nz.mem_1790_sv2v_reg ,\nz.mem_1789_sv2v_reg ,
  \nz.mem_1788_sv2v_reg ,\nz.mem_1787_sv2v_reg ,\nz.mem_1786_sv2v_reg ,\nz.mem_1785_sv2v_reg ,
  \nz.mem_1784_sv2v_reg ,\nz.mem_1783_sv2v_reg ,\nz.mem_1782_sv2v_reg ,
  \nz.mem_1781_sv2v_reg ,\nz.mem_1780_sv2v_reg ,\nz.mem_1779_sv2v_reg ,\nz.mem_1778_sv2v_reg ,
  \nz.mem_1777_sv2v_reg ,\nz.mem_1776_sv2v_reg ,\nz.mem_1775_sv2v_reg ,
  \nz.mem_1774_sv2v_reg ,\nz.mem_1773_sv2v_reg ,\nz.mem_1772_sv2v_reg ,\nz.mem_1771_sv2v_reg ,
  \nz.mem_1770_sv2v_reg ,\nz.mem_1769_sv2v_reg ,\nz.mem_1768_sv2v_reg ,
  \nz.mem_1767_sv2v_reg ,\nz.mem_1766_sv2v_reg ,\nz.mem_1765_sv2v_reg ,\nz.mem_1764_sv2v_reg ,
  \nz.mem_1763_sv2v_reg ,\nz.mem_1762_sv2v_reg ,\nz.mem_1761_sv2v_reg ,
  \nz.mem_1760_sv2v_reg ,\nz.mem_1759_sv2v_reg ,\nz.mem_1758_sv2v_reg ,\nz.mem_1757_sv2v_reg ,
  \nz.mem_1756_sv2v_reg ,\nz.mem_1755_sv2v_reg ,\nz.mem_1754_sv2v_reg ,
  \nz.mem_1753_sv2v_reg ,\nz.mem_1752_sv2v_reg ,\nz.mem_1751_sv2v_reg ,\nz.mem_1750_sv2v_reg ,
  \nz.mem_1749_sv2v_reg ,\nz.mem_1748_sv2v_reg ,\nz.mem_1747_sv2v_reg ,
  \nz.mem_1746_sv2v_reg ,\nz.mem_1745_sv2v_reg ,\nz.mem_1744_sv2v_reg ,\nz.mem_1743_sv2v_reg ,
  \nz.mem_1742_sv2v_reg ,\nz.mem_1741_sv2v_reg ,\nz.mem_1740_sv2v_reg ,
  \nz.mem_1739_sv2v_reg ,\nz.mem_1738_sv2v_reg ,\nz.mem_1737_sv2v_reg ,\nz.mem_1736_sv2v_reg ,
  \nz.mem_1735_sv2v_reg ,\nz.mem_1734_sv2v_reg ,\nz.mem_1733_sv2v_reg ,
  \nz.mem_1732_sv2v_reg ,\nz.mem_1731_sv2v_reg ,\nz.mem_1730_sv2v_reg ,
  \nz.mem_1729_sv2v_reg ,\nz.mem_1728_sv2v_reg ,\nz.mem_1727_sv2v_reg ,\nz.mem_1726_sv2v_reg ,
  \nz.mem_1725_sv2v_reg ,\nz.mem_1724_sv2v_reg ,\nz.mem_1723_sv2v_reg ,
  \nz.mem_1722_sv2v_reg ,\nz.mem_1721_sv2v_reg ,\nz.mem_1720_sv2v_reg ,\nz.mem_1719_sv2v_reg ,
  \nz.mem_1718_sv2v_reg ,\nz.mem_1717_sv2v_reg ,\nz.mem_1716_sv2v_reg ,
  \nz.mem_1715_sv2v_reg ,\nz.mem_1714_sv2v_reg ,\nz.mem_1713_sv2v_reg ,\nz.mem_1712_sv2v_reg ,
  \nz.mem_1711_sv2v_reg ,\nz.mem_1710_sv2v_reg ,\nz.mem_1709_sv2v_reg ,
  \nz.mem_1708_sv2v_reg ,\nz.mem_1707_sv2v_reg ,\nz.mem_1706_sv2v_reg ,\nz.mem_1705_sv2v_reg ,
  \nz.mem_1704_sv2v_reg ,\nz.mem_1703_sv2v_reg ,\nz.mem_1702_sv2v_reg ,
  \nz.mem_1701_sv2v_reg ,\nz.mem_1700_sv2v_reg ,\nz.mem_1699_sv2v_reg ,\nz.mem_1698_sv2v_reg ,
  \nz.mem_1697_sv2v_reg ,\nz.mem_1696_sv2v_reg ,\nz.mem_1695_sv2v_reg ,
  \nz.mem_1694_sv2v_reg ,\nz.mem_1693_sv2v_reg ,\nz.mem_1692_sv2v_reg ,\nz.mem_1691_sv2v_reg ,
  \nz.mem_1690_sv2v_reg ,\nz.mem_1689_sv2v_reg ,\nz.mem_1688_sv2v_reg ,
  \nz.mem_1687_sv2v_reg ,\nz.mem_1686_sv2v_reg ,\nz.mem_1685_sv2v_reg ,\nz.mem_1684_sv2v_reg ,
  \nz.mem_1683_sv2v_reg ,\nz.mem_1682_sv2v_reg ,\nz.mem_1681_sv2v_reg ,
  \nz.mem_1680_sv2v_reg ,\nz.mem_1679_sv2v_reg ,\nz.mem_1678_sv2v_reg ,\nz.mem_1677_sv2v_reg ,
  \nz.mem_1676_sv2v_reg ,\nz.mem_1675_sv2v_reg ,\nz.mem_1674_sv2v_reg ,
  \nz.mem_1673_sv2v_reg ,\nz.mem_1672_sv2v_reg ,\nz.mem_1671_sv2v_reg ,\nz.mem_1670_sv2v_reg ,
  \nz.mem_1669_sv2v_reg ,\nz.mem_1668_sv2v_reg ,\nz.mem_1667_sv2v_reg ,
  \nz.mem_1666_sv2v_reg ,\nz.mem_1665_sv2v_reg ,\nz.mem_1664_sv2v_reg ,\nz.mem_1663_sv2v_reg ,
  \nz.mem_1662_sv2v_reg ,\nz.mem_1661_sv2v_reg ,\nz.mem_1660_sv2v_reg ,
  \nz.mem_1659_sv2v_reg ,\nz.mem_1658_sv2v_reg ,\nz.mem_1657_sv2v_reg ,\nz.mem_1656_sv2v_reg ,
  \nz.mem_1655_sv2v_reg ,\nz.mem_1654_sv2v_reg ,\nz.mem_1653_sv2v_reg ,
  \nz.mem_1652_sv2v_reg ,\nz.mem_1651_sv2v_reg ,\nz.mem_1650_sv2v_reg ,
  \nz.mem_1649_sv2v_reg ,\nz.mem_1648_sv2v_reg ,\nz.mem_1647_sv2v_reg ,\nz.mem_1646_sv2v_reg ,
  \nz.mem_1645_sv2v_reg ,\nz.mem_1644_sv2v_reg ,\nz.mem_1643_sv2v_reg ,
  \nz.mem_1642_sv2v_reg ,\nz.mem_1641_sv2v_reg ,\nz.mem_1640_sv2v_reg ,\nz.mem_1639_sv2v_reg ,
  \nz.mem_1638_sv2v_reg ,\nz.mem_1637_sv2v_reg ,\nz.mem_1636_sv2v_reg ,
  \nz.mem_1635_sv2v_reg ,\nz.mem_1634_sv2v_reg ,\nz.mem_1633_sv2v_reg ,\nz.mem_1632_sv2v_reg ,
  \nz.mem_1631_sv2v_reg ,\nz.mem_1630_sv2v_reg ,\nz.mem_1629_sv2v_reg ,
  \nz.mem_1628_sv2v_reg ,\nz.mem_1627_sv2v_reg ,\nz.mem_1626_sv2v_reg ,\nz.mem_1625_sv2v_reg ,
  \nz.mem_1624_sv2v_reg ,\nz.mem_1623_sv2v_reg ,\nz.mem_1622_sv2v_reg ,
  \nz.mem_1621_sv2v_reg ,\nz.mem_1620_sv2v_reg ,\nz.mem_1619_sv2v_reg ,\nz.mem_1618_sv2v_reg ,
  \nz.mem_1617_sv2v_reg ,\nz.mem_1616_sv2v_reg ,\nz.mem_1615_sv2v_reg ,
  \nz.mem_1614_sv2v_reg ,\nz.mem_1613_sv2v_reg ,\nz.mem_1612_sv2v_reg ,\nz.mem_1611_sv2v_reg ,
  \nz.mem_1610_sv2v_reg ,\nz.mem_1609_sv2v_reg ,\nz.mem_1608_sv2v_reg ,
  \nz.mem_1607_sv2v_reg ,\nz.mem_1606_sv2v_reg ,\nz.mem_1605_sv2v_reg ,\nz.mem_1604_sv2v_reg ,
  \nz.mem_1603_sv2v_reg ,\nz.mem_1602_sv2v_reg ,\nz.mem_1601_sv2v_reg ,
  \nz.mem_1600_sv2v_reg ,\nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,
  \nz.mem_1596_sv2v_reg ,\nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,
  \nz.mem_1593_sv2v_reg ,\nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,
  \nz.mem_1589_sv2v_reg ,\nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,
  \nz.mem_1586_sv2v_reg ,\nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,
  \nz.mem_1582_sv2v_reg ,\nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,
  \nz.mem_1579_sv2v_reg ,\nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,
  \nz.mem_1575_sv2v_reg ,\nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,
  \nz.mem_1572_sv2v_reg ,\nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,
  \nz.mem_1569_sv2v_reg ,\nz.mem_1568_sv2v_reg ,\nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,
  \nz.mem_1565_sv2v_reg ,\nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,
  \nz.mem_1562_sv2v_reg ,\nz.mem_1561_sv2v_reg ,\nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,
  \nz.mem_1558_sv2v_reg ,\nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,
  \nz.mem_1555_sv2v_reg ,\nz.mem_1554_sv2v_reg ,\nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,
  \nz.mem_1551_sv2v_reg ,\nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,
  \nz.mem_1548_sv2v_reg ,\nz.mem_1547_sv2v_reg ,\nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,
  \nz.mem_1544_sv2v_reg ,\nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,
  \nz.mem_1541_sv2v_reg ,\nz.mem_1540_sv2v_reg ,\nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,
  \nz.mem_1537_sv2v_reg ,\nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,
  \nz.mem_1534_sv2v_reg ,\nz.mem_1533_sv2v_reg ,\nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,
  \nz.mem_1530_sv2v_reg ,\nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,
  \nz.mem_1527_sv2v_reg ,\nz.mem_1526_sv2v_reg ,\nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,
  \nz.mem_1523_sv2v_reg ,\nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,
  \nz.mem_1520_sv2v_reg ,\nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,
  \nz.mem_1516_sv2v_reg ,\nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,
  \nz.mem_1513_sv2v_reg ,\nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,
  \nz.mem_1509_sv2v_reg ,\nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,
  \nz.mem_1506_sv2v_reg ,\nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,
  \nz.mem_1502_sv2v_reg ,\nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,
  \nz.mem_1499_sv2v_reg ,\nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,
  \nz.mem_1495_sv2v_reg ,\nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,
  \nz.mem_1492_sv2v_reg ,\nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,
  \nz.mem_1489_sv2v_reg ,\nz.mem_1488_sv2v_reg ,\nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,
  \nz.mem_1485_sv2v_reg ,\nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,
  \nz.mem_1482_sv2v_reg ,\nz.mem_1481_sv2v_reg ,\nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,
  \nz.mem_1478_sv2v_reg ,\nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,
  \nz.mem_1475_sv2v_reg ,\nz.mem_1474_sv2v_reg ,\nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,
  \nz.mem_1471_sv2v_reg ,\nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,
  \nz.mem_1468_sv2v_reg ,\nz.mem_1467_sv2v_reg ,\nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,
  \nz.mem_1464_sv2v_reg ,\nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,
  \nz.mem_1461_sv2v_reg ,\nz.mem_1460_sv2v_reg ,\nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,
  \nz.mem_1457_sv2v_reg ,\nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,
  \nz.mem_1454_sv2v_reg ,\nz.mem_1453_sv2v_reg ,\nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,
  \nz.mem_1450_sv2v_reg ,\nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,
  \nz.mem_1447_sv2v_reg ,\nz.mem_1446_sv2v_reg ,\nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,
  \nz.mem_1443_sv2v_reg ,\nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,
  \nz.mem_1440_sv2v_reg ,\nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,
  \nz.mem_1436_sv2v_reg ,\nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,
  \nz.mem_1433_sv2v_reg ,\nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,
  \nz.mem_1429_sv2v_reg ,\nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,
  \nz.mem_1426_sv2v_reg ,\nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,
  \nz.mem_1422_sv2v_reg ,\nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,
  \nz.mem_1419_sv2v_reg ,\nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,
  \nz.mem_1415_sv2v_reg ,\nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,
  \nz.mem_1412_sv2v_reg ,\nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,
  \nz.mem_1409_sv2v_reg ,\nz.mem_1408_sv2v_reg ,\nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,
  \nz.mem_1405_sv2v_reg ,\nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,
  \nz.mem_1402_sv2v_reg ,\nz.mem_1401_sv2v_reg ,\nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,
  \nz.mem_1398_sv2v_reg ,\nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,
  \nz.mem_1395_sv2v_reg ,\nz.mem_1394_sv2v_reg ,\nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,
  \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,
  \nz.mem_1388_sv2v_reg ,\nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,
  \nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,
  \nz.mem_1381_sv2v_reg ,\nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,
  \nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,
  \nz.mem_1374_sv2v_reg ,\nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,
  \nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,
  \nz.mem_1367_sv2v_reg ,\nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,
  \nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,
  \nz.mem_1360_sv2v_reg ,\nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,
  \nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,
  \nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,
  \nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,
  \nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,
  \nz.mem_1329_sv2v_reg ,\nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,
  \nz.mem_1322_sv2v_reg ,\nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,
  \nz.mem_1315_sv2v_reg ,\nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,
  \nz.mem_1308_sv2v_reg ,\nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,
  \nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,
  \nz.mem_1301_sv2v_reg ,\nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,
  \nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,
  \nz.mem_1294_sv2v_reg ,\nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,
  \nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,
  \nz.mem_1287_sv2v_reg ,\nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,
  \nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,
  \nz.mem_1280_sv2v_reg ,\nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,
  \nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,
  \nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,
  \nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,
  \nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,
  \nz.mem_1249_sv2v_reg ,\nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,
  \nz.mem_1242_sv2v_reg ,\nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,
  \nz.mem_1235_sv2v_reg ,\nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,
  \nz.mem_1228_sv2v_reg ,\nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,
  \nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,
  \nz.mem_1221_sv2v_reg ,\nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,
  \nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,
  \nz.mem_1214_sv2v_reg ,\nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,
  \nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,
  \nz.mem_1207_sv2v_reg ,\nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,
  \nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,
  \nz.mem_1200_sv2v_reg ,\nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,
  \nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,
  \nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,
  \nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,
  \nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,
  \nz.mem_1169_sv2v_reg ,\nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,
  \nz.mem_1162_sv2v_reg ,\nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,
  \nz.mem_1155_sv2v_reg ,\nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,
  \nz.mem_1148_sv2v_reg ,\nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,
  \nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,
  \nz.mem_1141_sv2v_reg ,\nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,
  \nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,
  \nz.mem_1134_sv2v_reg ,\nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,
  \nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,
  \nz.mem_1127_sv2v_reg ,\nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,
  \nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,
  \nz.mem_1120_sv2v_reg ,\nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,
  \nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,
  \nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,
  \nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,
  \nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,
  \nz.mem_1089_sv2v_reg ,\nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,
  \nz.mem_1082_sv2v_reg ,\nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,
  \nz.mem_1075_sv2v_reg ,\nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,
  \nz.mem_1068_sv2v_reg ,\nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,
  \nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,
  \nz.mem_1061_sv2v_reg ,\nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,
  \nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,
  \nz.mem_1054_sv2v_reg ,\nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,
  \nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,
  \nz.mem_1047_sv2v_reg ,\nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,
  \nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,
  \nz.mem_1040_sv2v_reg ,\nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,
  \nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,
  \nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,
  \nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,
  \nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,
  \nz.mem_1009_sv2v_reg ,\nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,
  \nz.mem_1002_sv2v_reg ,\nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,
  \nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,
  \nz.mem_991_sv2v_reg ,\nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,
  \nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,
  \nz.mem_980_sv2v_reg ,\nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,
  \nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,
  \nz.mem_973_sv2v_reg ,\nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,
  \nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,
  \nz.mem_962_sv2v_reg ,\nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,
  \nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,
  \nz.mem_951_sv2v_reg ,\nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,
  \nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,
  \nz.mem_940_sv2v_reg ,\nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,
  \nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,
  \nz.mem_933_sv2v_reg ,\nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,
  \nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,
  \nz.mem_922_sv2v_reg ,\nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,
  \nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,
  \nz.mem_911_sv2v_reg ,\nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,
  \nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,
  \nz.mem_900_sv2v_reg ,\nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,
  \nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,
  \nz.mem_893_sv2v_reg ,\nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,
  \nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,
  \nz.mem_882_sv2v_reg ,\nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,
  \nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,
  \nz.mem_871_sv2v_reg ,\nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,
  \nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,
  \nz.mem_860_sv2v_reg ,\nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,
  \nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,
  \nz.mem_853_sv2v_reg ,\nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,
  \nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,
  \nz.mem_842_sv2v_reg ,\nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,
  \nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,
  \nz.mem_831_sv2v_reg ,\nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,
  \nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,
  \nz.mem_820_sv2v_reg ,\nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,
  \nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,
  \nz.mem_813_sv2v_reg ,\nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,
  \nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,
  \nz.mem_802_sv2v_reg ,\nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,
  \nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,
  \nz.mem_791_sv2v_reg ,\nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,
  \nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,
  \nz.mem_780_sv2v_reg ,\nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,
  \nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,
  \nz.mem_773_sv2v_reg ,\nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,
  \nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,
  \nz.mem_762_sv2v_reg ,\nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,
  \nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,
  \nz.mem_751_sv2v_reg ,\nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,
  \nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,
  \nz.mem_740_sv2v_reg ,\nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,
  \nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,
  \nz.mem_733_sv2v_reg ,\nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,
  \nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,
  \nz.mem_722_sv2v_reg ,\nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,
  \nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,
  \nz.mem_711_sv2v_reg ,\nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,
  \nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,
  \nz.mem_700_sv2v_reg ,\nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,
  \nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,
  \nz.mem_693_sv2v_reg ,\nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,
  \nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,
  \nz.mem_682_sv2v_reg ,\nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,
  \nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,
  \nz.mem_671_sv2v_reg ,\nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,
  \nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,
  \nz.mem_660_sv2v_reg ,\nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,
  \nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,
  \nz.mem_653_sv2v_reg ,\nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,
  \nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,
  \nz.mem_642_sv2v_reg ,\nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,
  \nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,
  \nz.mem_631_sv2v_reg ,\nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,
  \nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,
  \nz.mem_620_sv2v_reg ,\nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,
  \nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,
  \nz.mem_613_sv2v_reg ,\nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,
  \nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,
  \nz.mem_602_sv2v_reg ,\nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,
  \nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,
  \nz.mem_591_sv2v_reg ,\nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,
  \nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,
  \nz.mem_580_sv2v_reg ,\nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,
  \nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,
  \nz.mem_573_sv2v_reg ,\nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,
  \nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,
  \nz.mem_562_sv2v_reg ,\nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,
  \nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,
  \nz.mem_551_sv2v_reg ,\nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,
  \nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,
  \nz.mem_540_sv2v_reg ,\nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,
  \nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,
  \nz.mem_533_sv2v_reg ,\nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,
  \nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,
  \nz.mem_522_sv2v_reg ,\nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,
  \nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,
  \nz.mem_511_sv2v_reg ,\nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,
  \nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,
  \nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,
  \nz.mem_493_sv2v_reg ,\nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,
  \nz.mem_482_sv2v_reg ,\nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,
  \nz.mem_471_sv2v_reg ,\nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,
  \nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,
  \nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,
  \nz.mem_453_sv2v_reg ,\nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,
  \nz.mem_442_sv2v_reg ,\nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,
  \nz.mem_431_sv2v_reg ,\nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,
  \nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,
  \nz.mem_413_sv2v_reg ,\nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,
  \nz.mem_402_sv2v_reg ,\nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,
  \nz.mem_391_sv2v_reg ,\nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,
  \nz.mem_373_sv2v_reg ,\nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,
  \nz.mem_362_sv2v_reg ,\nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,
  \nz.mem_351_sv2v_reg ,\nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,
  \nz.mem_333_sv2v_reg ,\nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,
  \nz.mem_322_sv2v_reg ,\nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,
  \nz.mem_311_sv2v_reg ,\nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,
  \nz.mem_293_sv2v_reg ,\nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,
  \nz.mem_282_sv2v_reg ,\nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,
  \nz.mem_271_sv2v_reg ,\nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,
  \nz.mem_253_sv2v_reg ,\nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,
  \nz.mem_242_sv2v_reg ,\nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,
  \nz.mem_231_sv2v_reg ,\nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,
  \nz.mem_213_sv2v_reg ,\nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,
  \nz.mem_202_sv2v_reg ,\nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,
  \nz.mem_191_sv2v_reg ,\nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,
  \nz.mem_173_sv2v_reg ,\nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,
  \nz.mem_162_sv2v_reg ,\nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,
  \nz.mem_151_sv2v_reg ,\nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,
  \nz.mem_133_sv2v_reg ,\nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,
  \nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,
  \nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,
  \nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,
  \nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,
  \nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,
  \nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,
  \nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,
  \nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [7] = \nz.addr_r_7_sv2v_reg ;
  assign \nz.addr_r [6] = \nz.addr_r_6_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [2047] = \nz.mem_2047_sv2v_reg ;
  assign \nz.mem [2046] = \nz.mem_2046_sv2v_reg ;
  assign \nz.mem [2045] = \nz.mem_2045_sv2v_reg ;
  assign \nz.mem [2044] = \nz.mem_2044_sv2v_reg ;
  assign \nz.mem [2043] = \nz.mem_2043_sv2v_reg ;
  assign \nz.mem [2042] = \nz.mem_2042_sv2v_reg ;
  assign \nz.mem [2041] = \nz.mem_2041_sv2v_reg ;
  assign \nz.mem [2040] = \nz.mem_2040_sv2v_reg ;
  assign \nz.mem [2039] = \nz.mem_2039_sv2v_reg ;
  assign \nz.mem [2038] = \nz.mem_2038_sv2v_reg ;
  assign \nz.mem [2037] = \nz.mem_2037_sv2v_reg ;
  assign \nz.mem [2036] = \nz.mem_2036_sv2v_reg ;
  assign \nz.mem [2035] = \nz.mem_2035_sv2v_reg ;
  assign \nz.mem [2034] = \nz.mem_2034_sv2v_reg ;
  assign \nz.mem [2033] = \nz.mem_2033_sv2v_reg ;
  assign \nz.mem [2032] = \nz.mem_2032_sv2v_reg ;
  assign \nz.mem [2031] = \nz.mem_2031_sv2v_reg ;
  assign \nz.mem [2030] = \nz.mem_2030_sv2v_reg ;
  assign \nz.mem [2029] = \nz.mem_2029_sv2v_reg ;
  assign \nz.mem [2028] = \nz.mem_2028_sv2v_reg ;
  assign \nz.mem [2027] = \nz.mem_2027_sv2v_reg ;
  assign \nz.mem [2026] = \nz.mem_2026_sv2v_reg ;
  assign \nz.mem [2025] = \nz.mem_2025_sv2v_reg ;
  assign \nz.mem [2024] = \nz.mem_2024_sv2v_reg ;
  assign \nz.mem [2023] = \nz.mem_2023_sv2v_reg ;
  assign \nz.mem [2022] = \nz.mem_2022_sv2v_reg ;
  assign \nz.mem [2021] = \nz.mem_2021_sv2v_reg ;
  assign \nz.mem [2020] = \nz.mem_2020_sv2v_reg ;
  assign \nz.mem [2019] = \nz.mem_2019_sv2v_reg ;
  assign \nz.mem [2018] = \nz.mem_2018_sv2v_reg ;
  assign \nz.mem [2017] = \nz.mem_2017_sv2v_reg ;
  assign \nz.mem [2016] = \nz.mem_2016_sv2v_reg ;
  assign \nz.mem [2015] = \nz.mem_2015_sv2v_reg ;
  assign \nz.mem [2014] = \nz.mem_2014_sv2v_reg ;
  assign \nz.mem [2013] = \nz.mem_2013_sv2v_reg ;
  assign \nz.mem [2012] = \nz.mem_2012_sv2v_reg ;
  assign \nz.mem [2011] = \nz.mem_2011_sv2v_reg ;
  assign \nz.mem [2010] = \nz.mem_2010_sv2v_reg ;
  assign \nz.mem [2009] = \nz.mem_2009_sv2v_reg ;
  assign \nz.mem [2008] = \nz.mem_2008_sv2v_reg ;
  assign \nz.mem [2007] = \nz.mem_2007_sv2v_reg ;
  assign \nz.mem [2006] = \nz.mem_2006_sv2v_reg ;
  assign \nz.mem [2005] = \nz.mem_2005_sv2v_reg ;
  assign \nz.mem [2004] = \nz.mem_2004_sv2v_reg ;
  assign \nz.mem [2003] = \nz.mem_2003_sv2v_reg ;
  assign \nz.mem [2002] = \nz.mem_2002_sv2v_reg ;
  assign \nz.mem [2001] = \nz.mem_2001_sv2v_reg ;
  assign \nz.mem [2000] = \nz.mem_2000_sv2v_reg ;
  assign \nz.mem [1999] = \nz.mem_1999_sv2v_reg ;
  assign \nz.mem [1998] = \nz.mem_1998_sv2v_reg ;
  assign \nz.mem [1997] = \nz.mem_1997_sv2v_reg ;
  assign \nz.mem [1996] = \nz.mem_1996_sv2v_reg ;
  assign \nz.mem [1995] = \nz.mem_1995_sv2v_reg ;
  assign \nz.mem [1994] = \nz.mem_1994_sv2v_reg ;
  assign \nz.mem [1993] = \nz.mem_1993_sv2v_reg ;
  assign \nz.mem [1992] = \nz.mem_1992_sv2v_reg ;
  assign \nz.mem [1991] = \nz.mem_1991_sv2v_reg ;
  assign \nz.mem [1990] = \nz.mem_1990_sv2v_reg ;
  assign \nz.mem [1989] = \nz.mem_1989_sv2v_reg ;
  assign \nz.mem [1988] = \nz.mem_1988_sv2v_reg ;
  assign \nz.mem [1987] = \nz.mem_1987_sv2v_reg ;
  assign \nz.mem [1986] = \nz.mem_1986_sv2v_reg ;
  assign \nz.mem [1985] = \nz.mem_1985_sv2v_reg ;
  assign \nz.mem [1984] = \nz.mem_1984_sv2v_reg ;
  assign \nz.mem [1983] = \nz.mem_1983_sv2v_reg ;
  assign \nz.mem [1982] = \nz.mem_1982_sv2v_reg ;
  assign \nz.mem [1981] = \nz.mem_1981_sv2v_reg ;
  assign \nz.mem [1980] = \nz.mem_1980_sv2v_reg ;
  assign \nz.mem [1979] = \nz.mem_1979_sv2v_reg ;
  assign \nz.mem [1978] = \nz.mem_1978_sv2v_reg ;
  assign \nz.mem [1977] = \nz.mem_1977_sv2v_reg ;
  assign \nz.mem [1976] = \nz.mem_1976_sv2v_reg ;
  assign \nz.mem [1975] = \nz.mem_1975_sv2v_reg ;
  assign \nz.mem [1974] = \nz.mem_1974_sv2v_reg ;
  assign \nz.mem [1973] = \nz.mem_1973_sv2v_reg ;
  assign \nz.mem [1972] = \nz.mem_1972_sv2v_reg ;
  assign \nz.mem [1971] = \nz.mem_1971_sv2v_reg ;
  assign \nz.mem [1970] = \nz.mem_1970_sv2v_reg ;
  assign \nz.mem [1969] = \nz.mem_1969_sv2v_reg ;
  assign \nz.mem [1968] = \nz.mem_1968_sv2v_reg ;
  assign \nz.mem [1967] = \nz.mem_1967_sv2v_reg ;
  assign \nz.mem [1966] = \nz.mem_1966_sv2v_reg ;
  assign \nz.mem [1965] = \nz.mem_1965_sv2v_reg ;
  assign \nz.mem [1964] = \nz.mem_1964_sv2v_reg ;
  assign \nz.mem [1963] = \nz.mem_1963_sv2v_reg ;
  assign \nz.mem [1962] = \nz.mem_1962_sv2v_reg ;
  assign \nz.mem [1961] = \nz.mem_1961_sv2v_reg ;
  assign \nz.mem [1960] = \nz.mem_1960_sv2v_reg ;
  assign \nz.mem [1959] = \nz.mem_1959_sv2v_reg ;
  assign \nz.mem [1958] = \nz.mem_1958_sv2v_reg ;
  assign \nz.mem [1957] = \nz.mem_1957_sv2v_reg ;
  assign \nz.mem [1956] = \nz.mem_1956_sv2v_reg ;
  assign \nz.mem [1955] = \nz.mem_1955_sv2v_reg ;
  assign \nz.mem [1954] = \nz.mem_1954_sv2v_reg ;
  assign \nz.mem [1953] = \nz.mem_1953_sv2v_reg ;
  assign \nz.mem [1952] = \nz.mem_1952_sv2v_reg ;
  assign \nz.mem [1951] = \nz.mem_1951_sv2v_reg ;
  assign \nz.mem [1950] = \nz.mem_1950_sv2v_reg ;
  assign \nz.mem [1949] = \nz.mem_1949_sv2v_reg ;
  assign \nz.mem [1948] = \nz.mem_1948_sv2v_reg ;
  assign \nz.mem [1947] = \nz.mem_1947_sv2v_reg ;
  assign \nz.mem [1946] = \nz.mem_1946_sv2v_reg ;
  assign \nz.mem [1945] = \nz.mem_1945_sv2v_reg ;
  assign \nz.mem [1944] = \nz.mem_1944_sv2v_reg ;
  assign \nz.mem [1943] = \nz.mem_1943_sv2v_reg ;
  assign \nz.mem [1942] = \nz.mem_1942_sv2v_reg ;
  assign \nz.mem [1941] = \nz.mem_1941_sv2v_reg ;
  assign \nz.mem [1940] = \nz.mem_1940_sv2v_reg ;
  assign \nz.mem [1939] = \nz.mem_1939_sv2v_reg ;
  assign \nz.mem [1938] = \nz.mem_1938_sv2v_reg ;
  assign \nz.mem [1937] = \nz.mem_1937_sv2v_reg ;
  assign \nz.mem [1936] = \nz.mem_1936_sv2v_reg ;
  assign \nz.mem [1935] = \nz.mem_1935_sv2v_reg ;
  assign \nz.mem [1934] = \nz.mem_1934_sv2v_reg ;
  assign \nz.mem [1933] = \nz.mem_1933_sv2v_reg ;
  assign \nz.mem [1932] = \nz.mem_1932_sv2v_reg ;
  assign \nz.mem [1931] = \nz.mem_1931_sv2v_reg ;
  assign \nz.mem [1930] = \nz.mem_1930_sv2v_reg ;
  assign \nz.mem [1929] = \nz.mem_1929_sv2v_reg ;
  assign \nz.mem [1928] = \nz.mem_1928_sv2v_reg ;
  assign \nz.mem [1927] = \nz.mem_1927_sv2v_reg ;
  assign \nz.mem [1926] = \nz.mem_1926_sv2v_reg ;
  assign \nz.mem [1925] = \nz.mem_1925_sv2v_reg ;
  assign \nz.mem [1924] = \nz.mem_1924_sv2v_reg ;
  assign \nz.mem [1923] = \nz.mem_1923_sv2v_reg ;
  assign \nz.mem [1922] = \nz.mem_1922_sv2v_reg ;
  assign \nz.mem [1921] = \nz.mem_1921_sv2v_reg ;
  assign \nz.mem [1920] = \nz.mem_1920_sv2v_reg ;
  assign \nz.mem [1919] = \nz.mem_1919_sv2v_reg ;
  assign \nz.mem [1918] = \nz.mem_1918_sv2v_reg ;
  assign \nz.mem [1917] = \nz.mem_1917_sv2v_reg ;
  assign \nz.mem [1916] = \nz.mem_1916_sv2v_reg ;
  assign \nz.mem [1915] = \nz.mem_1915_sv2v_reg ;
  assign \nz.mem [1914] = \nz.mem_1914_sv2v_reg ;
  assign \nz.mem [1913] = \nz.mem_1913_sv2v_reg ;
  assign \nz.mem [1912] = \nz.mem_1912_sv2v_reg ;
  assign \nz.mem [1911] = \nz.mem_1911_sv2v_reg ;
  assign \nz.mem [1910] = \nz.mem_1910_sv2v_reg ;
  assign \nz.mem [1909] = \nz.mem_1909_sv2v_reg ;
  assign \nz.mem [1908] = \nz.mem_1908_sv2v_reg ;
  assign \nz.mem [1907] = \nz.mem_1907_sv2v_reg ;
  assign \nz.mem [1906] = \nz.mem_1906_sv2v_reg ;
  assign \nz.mem [1905] = \nz.mem_1905_sv2v_reg ;
  assign \nz.mem [1904] = \nz.mem_1904_sv2v_reg ;
  assign \nz.mem [1903] = \nz.mem_1903_sv2v_reg ;
  assign \nz.mem [1902] = \nz.mem_1902_sv2v_reg ;
  assign \nz.mem [1901] = \nz.mem_1901_sv2v_reg ;
  assign \nz.mem [1900] = \nz.mem_1900_sv2v_reg ;
  assign \nz.mem [1899] = \nz.mem_1899_sv2v_reg ;
  assign \nz.mem [1898] = \nz.mem_1898_sv2v_reg ;
  assign \nz.mem [1897] = \nz.mem_1897_sv2v_reg ;
  assign \nz.mem [1896] = \nz.mem_1896_sv2v_reg ;
  assign \nz.mem [1895] = \nz.mem_1895_sv2v_reg ;
  assign \nz.mem [1894] = \nz.mem_1894_sv2v_reg ;
  assign \nz.mem [1893] = \nz.mem_1893_sv2v_reg ;
  assign \nz.mem [1892] = \nz.mem_1892_sv2v_reg ;
  assign \nz.mem [1891] = \nz.mem_1891_sv2v_reg ;
  assign \nz.mem [1890] = \nz.mem_1890_sv2v_reg ;
  assign \nz.mem [1889] = \nz.mem_1889_sv2v_reg ;
  assign \nz.mem [1888] = \nz.mem_1888_sv2v_reg ;
  assign \nz.mem [1887] = \nz.mem_1887_sv2v_reg ;
  assign \nz.mem [1886] = \nz.mem_1886_sv2v_reg ;
  assign \nz.mem [1885] = \nz.mem_1885_sv2v_reg ;
  assign \nz.mem [1884] = \nz.mem_1884_sv2v_reg ;
  assign \nz.mem [1883] = \nz.mem_1883_sv2v_reg ;
  assign \nz.mem [1882] = \nz.mem_1882_sv2v_reg ;
  assign \nz.mem [1881] = \nz.mem_1881_sv2v_reg ;
  assign \nz.mem [1880] = \nz.mem_1880_sv2v_reg ;
  assign \nz.mem [1879] = \nz.mem_1879_sv2v_reg ;
  assign \nz.mem [1878] = \nz.mem_1878_sv2v_reg ;
  assign \nz.mem [1877] = \nz.mem_1877_sv2v_reg ;
  assign \nz.mem [1876] = \nz.mem_1876_sv2v_reg ;
  assign \nz.mem [1875] = \nz.mem_1875_sv2v_reg ;
  assign \nz.mem [1874] = \nz.mem_1874_sv2v_reg ;
  assign \nz.mem [1873] = \nz.mem_1873_sv2v_reg ;
  assign \nz.mem [1872] = \nz.mem_1872_sv2v_reg ;
  assign \nz.mem [1871] = \nz.mem_1871_sv2v_reg ;
  assign \nz.mem [1870] = \nz.mem_1870_sv2v_reg ;
  assign \nz.mem [1869] = \nz.mem_1869_sv2v_reg ;
  assign \nz.mem [1868] = \nz.mem_1868_sv2v_reg ;
  assign \nz.mem [1867] = \nz.mem_1867_sv2v_reg ;
  assign \nz.mem [1866] = \nz.mem_1866_sv2v_reg ;
  assign \nz.mem [1865] = \nz.mem_1865_sv2v_reg ;
  assign \nz.mem [1864] = \nz.mem_1864_sv2v_reg ;
  assign \nz.mem [1863] = \nz.mem_1863_sv2v_reg ;
  assign \nz.mem [1862] = \nz.mem_1862_sv2v_reg ;
  assign \nz.mem [1861] = \nz.mem_1861_sv2v_reg ;
  assign \nz.mem [1860] = \nz.mem_1860_sv2v_reg ;
  assign \nz.mem [1859] = \nz.mem_1859_sv2v_reg ;
  assign \nz.mem [1858] = \nz.mem_1858_sv2v_reg ;
  assign \nz.mem [1857] = \nz.mem_1857_sv2v_reg ;
  assign \nz.mem [1856] = \nz.mem_1856_sv2v_reg ;
  assign \nz.mem [1855] = \nz.mem_1855_sv2v_reg ;
  assign \nz.mem [1854] = \nz.mem_1854_sv2v_reg ;
  assign \nz.mem [1853] = \nz.mem_1853_sv2v_reg ;
  assign \nz.mem [1852] = \nz.mem_1852_sv2v_reg ;
  assign \nz.mem [1851] = \nz.mem_1851_sv2v_reg ;
  assign \nz.mem [1850] = \nz.mem_1850_sv2v_reg ;
  assign \nz.mem [1849] = \nz.mem_1849_sv2v_reg ;
  assign \nz.mem [1848] = \nz.mem_1848_sv2v_reg ;
  assign \nz.mem [1847] = \nz.mem_1847_sv2v_reg ;
  assign \nz.mem [1846] = \nz.mem_1846_sv2v_reg ;
  assign \nz.mem [1845] = \nz.mem_1845_sv2v_reg ;
  assign \nz.mem [1844] = \nz.mem_1844_sv2v_reg ;
  assign \nz.mem [1843] = \nz.mem_1843_sv2v_reg ;
  assign \nz.mem [1842] = \nz.mem_1842_sv2v_reg ;
  assign \nz.mem [1841] = \nz.mem_1841_sv2v_reg ;
  assign \nz.mem [1840] = \nz.mem_1840_sv2v_reg ;
  assign \nz.mem [1839] = \nz.mem_1839_sv2v_reg ;
  assign \nz.mem [1838] = \nz.mem_1838_sv2v_reg ;
  assign \nz.mem [1837] = \nz.mem_1837_sv2v_reg ;
  assign \nz.mem [1836] = \nz.mem_1836_sv2v_reg ;
  assign \nz.mem [1835] = \nz.mem_1835_sv2v_reg ;
  assign \nz.mem [1834] = \nz.mem_1834_sv2v_reg ;
  assign \nz.mem [1833] = \nz.mem_1833_sv2v_reg ;
  assign \nz.mem [1832] = \nz.mem_1832_sv2v_reg ;
  assign \nz.mem [1831] = \nz.mem_1831_sv2v_reg ;
  assign \nz.mem [1830] = \nz.mem_1830_sv2v_reg ;
  assign \nz.mem [1829] = \nz.mem_1829_sv2v_reg ;
  assign \nz.mem [1828] = \nz.mem_1828_sv2v_reg ;
  assign \nz.mem [1827] = \nz.mem_1827_sv2v_reg ;
  assign \nz.mem [1826] = \nz.mem_1826_sv2v_reg ;
  assign \nz.mem [1825] = \nz.mem_1825_sv2v_reg ;
  assign \nz.mem [1824] = \nz.mem_1824_sv2v_reg ;
  assign \nz.mem [1823] = \nz.mem_1823_sv2v_reg ;
  assign \nz.mem [1822] = \nz.mem_1822_sv2v_reg ;
  assign \nz.mem [1821] = \nz.mem_1821_sv2v_reg ;
  assign \nz.mem [1820] = \nz.mem_1820_sv2v_reg ;
  assign \nz.mem [1819] = \nz.mem_1819_sv2v_reg ;
  assign \nz.mem [1818] = \nz.mem_1818_sv2v_reg ;
  assign \nz.mem [1817] = \nz.mem_1817_sv2v_reg ;
  assign \nz.mem [1816] = \nz.mem_1816_sv2v_reg ;
  assign \nz.mem [1815] = \nz.mem_1815_sv2v_reg ;
  assign \nz.mem [1814] = \nz.mem_1814_sv2v_reg ;
  assign \nz.mem [1813] = \nz.mem_1813_sv2v_reg ;
  assign \nz.mem [1812] = \nz.mem_1812_sv2v_reg ;
  assign \nz.mem [1811] = \nz.mem_1811_sv2v_reg ;
  assign \nz.mem [1810] = \nz.mem_1810_sv2v_reg ;
  assign \nz.mem [1809] = \nz.mem_1809_sv2v_reg ;
  assign \nz.mem [1808] = \nz.mem_1808_sv2v_reg ;
  assign \nz.mem [1807] = \nz.mem_1807_sv2v_reg ;
  assign \nz.mem [1806] = \nz.mem_1806_sv2v_reg ;
  assign \nz.mem [1805] = \nz.mem_1805_sv2v_reg ;
  assign \nz.mem [1804] = \nz.mem_1804_sv2v_reg ;
  assign \nz.mem [1803] = \nz.mem_1803_sv2v_reg ;
  assign \nz.mem [1802] = \nz.mem_1802_sv2v_reg ;
  assign \nz.mem [1801] = \nz.mem_1801_sv2v_reg ;
  assign \nz.mem [1800] = \nz.mem_1800_sv2v_reg ;
  assign \nz.mem [1799] = \nz.mem_1799_sv2v_reg ;
  assign \nz.mem [1798] = \nz.mem_1798_sv2v_reg ;
  assign \nz.mem [1797] = \nz.mem_1797_sv2v_reg ;
  assign \nz.mem [1796] = \nz.mem_1796_sv2v_reg ;
  assign \nz.mem [1795] = \nz.mem_1795_sv2v_reg ;
  assign \nz.mem [1794] = \nz.mem_1794_sv2v_reg ;
  assign \nz.mem [1793] = \nz.mem_1793_sv2v_reg ;
  assign \nz.mem [1792] = \nz.mem_1792_sv2v_reg ;
  assign \nz.mem [1791] = \nz.mem_1791_sv2v_reg ;
  assign \nz.mem [1790] = \nz.mem_1790_sv2v_reg ;
  assign \nz.mem [1789] = \nz.mem_1789_sv2v_reg ;
  assign \nz.mem [1788] = \nz.mem_1788_sv2v_reg ;
  assign \nz.mem [1787] = \nz.mem_1787_sv2v_reg ;
  assign \nz.mem [1786] = \nz.mem_1786_sv2v_reg ;
  assign \nz.mem [1785] = \nz.mem_1785_sv2v_reg ;
  assign \nz.mem [1784] = \nz.mem_1784_sv2v_reg ;
  assign \nz.mem [1783] = \nz.mem_1783_sv2v_reg ;
  assign \nz.mem [1782] = \nz.mem_1782_sv2v_reg ;
  assign \nz.mem [1781] = \nz.mem_1781_sv2v_reg ;
  assign \nz.mem [1780] = \nz.mem_1780_sv2v_reg ;
  assign \nz.mem [1779] = \nz.mem_1779_sv2v_reg ;
  assign \nz.mem [1778] = \nz.mem_1778_sv2v_reg ;
  assign \nz.mem [1777] = \nz.mem_1777_sv2v_reg ;
  assign \nz.mem [1776] = \nz.mem_1776_sv2v_reg ;
  assign \nz.mem [1775] = \nz.mem_1775_sv2v_reg ;
  assign \nz.mem [1774] = \nz.mem_1774_sv2v_reg ;
  assign \nz.mem [1773] = \nz.mem_1773_sv2v_reg ;
  assign \nz.mem [1772] = \nz.mem_1772_sv2v_reg ;
  assign \nz.mem [1771] = \nz.mem_1771_sv2v_reg ;
  assign \nz.mem [1770] = \nz.mem_1770_sv2v_reg ;
  assign \nz.mem [1769] = \nz.mem_1769_sv2v_reg ;
  assign \nz.mem [1768] = \nz.mem_1768_sv2v_reg ;
  assign \nz.mem [1767] = \nz.mem_1767_sv2v_reg ;
  assign \nz.mem [1766] = \nz.mem_1766_sv2v_reg ;
  assign \nz.mem [1765] = \nz.mem_1765_sv2v_reg ;
  assign \nz.mem [1764] = \nz.mem_1764_sv2v_reg ;
  assign \nz.mem [1763] = \nz.mem_1763_sv2v_reg ;
  assign \nz.mem [1762] = \nz.mem_1762_sv2v_reg ;
  assign \nz.mem [1761] = \nz.mem_1761_sv2v_reg ;
  assign \nz.mem [1760] = \nz.mem_1760_sv2v_reg ;
  assign \nz.mem [1759] = \nz.mem_1759_sv2v_reg ;
  assign \nz.mem [1758] = \nz.mem_1758_sv2v_reg ;
  assign \nz.mem [1757] = \nz.mem_1757_sv2v_reg ;
  assign \nz.mem [1756] = \nz.mem_1756_sv2v_reg ;
  assign \nz.mem [1755] = \nz.mem_1755_sv2v_reg ;
  assign \nz.mem [1754] = \nz.mem_1754_sv2v_reg ;
  assign \nz.mem [1753] = \nz.mem_1753_sv2v_reg ;
  assign \nz.mem [1752] = \nz.mem_1752_sv2v_reg ;
  assign \nz.mem [1751] = \nz.mem_1751_sv2v_reg ;
  assign \nz.mem [1750] = \nz.mem_1750_sv2v_reg ;
  assign \nz.mem [1749] = \nz.mem_1749_sv2v_reg ;
  assign \nz.mem [1748] = \nz.mem_1748_sv2v_reg ;
  assign \nz.mem [1747] = \nz.mem_1747_sv2v_reg ;
  assign \nz.mem [1746] = \nz.mem_1746_sv2v_reg ;
  assign \nz.mem [1745] = \nz.mem_1745_sv2v_reg ;
  assign \nz.mem [1744] = \nz.mem_1744_sv2v_reg ;
  assign \nz.mem [1743] = \nz.mem_1743_sv2v_reg ;
  assign \nz.mem [1742] = \nz.mem_1742_sv2v_reg ;
  assign \nz.mem [1741] = \nz.mem_1741_sv2v_reg ;
  assign \nz.mem [1740] = \nz.mem_1740_sv2v_reg ;
  assign \nz.mem [1739] = \nz.mem_1739_sv2v_reg ;
  assign \nz.mem [1738] = \nz.mem_1738_sv2v_reg ;
  assign \nz.mem [1737] = \nz.mem_1737_sv2v_reg ;
  assign \nz.mem [1736] = \nz.mem_1736_sv2v_reg ;
  assign \nz.mem [1735] = \nz.mem_1735_sv2v_reg ;
  assign \nz.mem [1734] = \nz.mem_1734_sv2v_reg ;
  assign \nz.mem [1733] = \nz.mem_1733_sv2v_reg ;
  assign \nz.mem [1732] = \nz.mem_1732_sv2v_reg ;
  assign \nz.mem [1731] = \nz.mem_1731_sv2v_reg ;
  assign \nz.mem [1730] = \nz.mem_1730_sv2v_reg ;
  assign \nz.mem [1729] = \nz.mem_1729_sv2v_reg ;
  assign \nz.mem [1728] = \nz.mem_1728_sv2v_reg ;
  assign \nz.mem [1727] = \nz.mem_1727_sv2v_reg ;
  assign \nz.mem [1726] = \nz.mem_1726_sv2v_reg ;
  assign \nz.mem [1725] = \nz.mem_1725_sv2v_reg ;
  assign \nz.mem [1724] = \nz.mem_1724_sv2v_reg ;
  assign \nz.mem [1723] = \nz.mem_1723_sv2v_reg ;
  assign \nz.mem [1722] = \nz.mem_1722_sv2v_reg ;
  assign \nz.mem [1721] = \nz.mem_1721_sv2v_reg ;
  assign \nz.mem [1720] = \nz.mem_1720_sv2v_reg ;
  assign \nz.mem [1719] = \nz.mem_1719_sv2v_reg ;
  assign \nz.mem [1718] = \nz.mem_1718_sv2v_reg ;
  assign \nz.mem [1717] = \nz.mem_1717_sv2v_reg ;
  assign \nz.mem [1716] = \nz.mem_1716_sv2v_reg ;
  assign \nz.mem [1715] = \nz.mem_1715_sv2v_reg ;
  assign \nz.mem [1714] = \nz.mem_1714_sv2v_reg ;
  assign \nz.mem [1713] = \nz.mem_1713_sv2v_reg ;
  assign \nz.mem [1712] = \nz.mem_1712_sv2v_reg ;
  assign \nz.mem [1711] = \nz.mem_1711_sv2v_reg ;
  assign \nz.mem [1710] = \nz.mem_1710_sv2v_reg ;
  assign \nz.mem [1709] = \nz.mem_1709_sv2v_reg ;
  assign \nz.mem [1708] = \nz.mem_1708_sv2v_reg ;
  assign \nz.mem [1707] = \nz.mem_1707_sv2v_reg ;
  assign \nz.mem [1706] = \nz.mem_1706_sv2v_reg ;
  assign \nz.mem [1705] = \nz.mem_1705_sv2v_reg ;
  assign \nz.mem [1704] = \nz.mem_1704_sv2v_reg ;
  assign \nz.mem [1703] = \nz.mem_1703_sv2v_reg ;
  assign \nz.mem [1702] = \nz.mem_1702_sv2v_reg ;
  assign \nz.mem [1701] = \nz.mem_1701_sv2v_reg ;
  assign \nz.mem [1700] = \nz.mem_1700_sv2v_reg ;
  assign \nz.mem [1699] = \nz.mem_1699_sv2v_reg ;
  assign \nz.mem [1698] = \nz.mem_1698_sv2v_reg ;
  assign \nz.mem [1697] = \nz.mem_1697_sv2v_reg ;
  assign \nz.mem [1696] = \nz.mem_1696_sv2v_reg ;
  assign \nz.mem [1695] = \nz.mem_1695_sv2v_reg ;
  assign \nz.mem [1694] = \nz.mem_1694_sv2v_reg ;
  assign \nz.mem [1693] = \nz.mem_1693_sv2v_reg ;
  assign \nz.mem [1692] = \nz.mem_1692_sv2v_reg ;
  assign \nz.mem [1691] = \nz.mem_1691_sv2v_reg ;
  assign \nz.mem [1690] = \nz.mem_1690_sv2v_reg ;
  assign \nz.mem [1689] = \nz.mem_1689_sv2v_reg ;
  assign \nz.mem [1688] = \nz.mem_1688_sv2v_reg ;
  assign \nz.mem [1687] = \nz.mem_1687_sv2v_reg ;
  assign \nz.mem [1686] = \nz.mem_1686_sv2v_reg ;
  assign \nz.mem [1685] = \nz.mem_1685_sv2v_reg ;
  assign \nz.mem [1684] = \nz.mem_1684_sv2v_reg ;
  assign \nz.mem [1683] = \nz.mem_1683_sv2v_reg ;
  assign \nz.mem [1682] = \nz.mem_1682_sv2v_reg ;
  assign \nz.mem [1681] = \nz.mem_1681_sv2v_reg ;
  assign \nz.mem [1680] = \nz.mem_1680_sv2v_reg ;
  assign \nz.mem [1679] = \nz.mem_1679_sv2v_reg ;
  assign \nz.mem [1678] = \nz.mem_1678_sv2v_reg ;
  assign \nz.mem [1677] = \nz.mem_1677_sv2v_reg ;
  assign \nz.mem [1676] = \nz.mem_1676_sv2v_reg ;
  assign \nz.mem [1675] = \nz.mem_1675_sv2v_reg ;
  assign \nz.mem [1674] = \nz.mem_1674_sv2v_reg ;
  assign \nz.mem [1673] = \nz.mem_1673_sv2v_reg ;
  assign \nz.mem [1672] = \nz.mem_1672_sv2v_reg ;
  assign \nz.mem [1671] = \nz.mem_1671_sv2v_reg ;
  assign \nz.mem [1670] = \nz.mem_1670_sv2v_reg ;
  assign \nz.mem [1669] = \nz.mem_1669_sv2v_reg ;
  assign \nz.mem [1668] = \nz.mem_1668_sv2v_reg ;
  assign \nz.mem [1667] = \nz.mem_1667_sv2v_reg ;
  assign \nz.mem [1666] = \nz.mem_1666_sv2v_reg ;
  assign \nz.mem [1665] = \nz.mem_1665_sv2v_reg ;
  assign \nz.mem [1664] = \nz.mem_1664_sv2v_reg ;
  assign \nz.mem [1663] = \nz.mem_1663_sv2v_reg ;
  assign \nz.mem [1662] = \nz.mem_1662_sv2v_reg ;
  assign \nz.mem [1661] = \nz.mem_1661_sv2v_reg ;
  assign \nz.mem [1660] = \nz.mem_1660_sv2v_reg ;
  assign \nz.mem [1659] = \nz.mem_1659_sv2v_reg ;
  assign \nz.mem [1658] = \nz.mem_1658_sv2v_reg ;
  assign \nz.mem [1657] = \nz.mem_1657_sv2v_reg ;
  assign \nz.mem [1656] = \nz.mem_1656_sv2v_reg ;
  assign \nz.mem [1655] = \nz.mem_1655_sv2v_reg ;
  assign \nz.mem [1654] = \nz.mem_1654_sv2v_reg ;
  assign \nz.mem [1653] = \nz.mem_1653_sv2v_reg ;
  assign \nz.mem [1652] = \nz.mem_1652_sv2v_reg ;
  assign \nz.mem [1651] = \nz.mem_1651_sv2v_reg ;
  assign \nz.mem [1650] = \nz.mem_1650_sv2v_reg ;
  assign \nz.mem [1649] = \nz.mem_1649_sv2v_reg ;
  assign \nz.mem [1648] = \nz.mem_1648_sv2v_reg ;
  assign \nz.mem [1647] = \nz.mem_1647_sv2v_reg ;
  assign \nz.mem [1646] = \nz.mem_1646_sv2v_reg ;
  assign \nz.mem [1645] = \nz.mem_1645_sv2v_reg ;
  assign \nz.mem [1644] = \nz.mem_1644_sv2v_reg ;
  assign \nz.mem [1643] = \nz.mem_1643_sv2v_reg ;
  assign \nz.mem [1642] = \nz.mem_1642_sv2v_reg ;
  assign \nz.mem [1641] = \nz.mem_1641_sv2v_reg ;
  assign \nz.mem [1640] = \nz.mem_1640_sv2v_reg ;
  assign \nz.mem [1639] = \nz.mem_1639_sv2v_reg ;
  assign \nz.mem [1638] = \nz.mem_1638_sv2v_reg ;
  assign \nz.mem [1637] = \nz.mem_1637_sv2v_reg ;
  assign \nz.mem [1636] = \nz.mem_1636_sv2v_reg ;
  assign \nz.mem [1635] = \nz.mem_1635_sv2v_reg ;
  assign \nz.mem [1634] = \nz.mem_1634_sv2v_reg ;
  assign \nz.mem [1633] = \nz.mem_1633_sv2v_reg ;
  assign \nz.mem [1632] = \nz.mem_1632_sv2v_reg ;
  assign \nz.mem [1631] = \nz.mem_1631_sv2v_reg ;
  assign \nz.mem [1630] = \nz.mem_1630_sv2v_reg ;
  assign \nz.mem [1629] = \nz.mem_1629_sv2v_reg ;
  assign \nz.mem [1628] = \nz.mem_1628_sv2v_reg ;
  assign \nz.mem [1627] = \nz.mem_1627_sv2v_reg ;
  assign \nz.mem [1626] = \nz.mem_1626_sv2v_reg ;
  assign \nz.mem [1625] = \nz.mem_1625_sv2v_reg ;
  assign \nz.mem [1624] = \nz.mem_1624_sv2v_reg ;
  assign \nz.mem [1623] = \nz.mem_1623_sv2v_reg ;
  assign \nz.mem [1622] = \nz.mem_1622_sv2v_reg ;
  assign \nz.mem [1621] = \nz.mem_1621_sv2v_reg ;
  assign \nz.mem [1620] = \nz.mem_1620_sv2v_reg ;
  assign \nz.mem [1619] = \nz.mem_1619_sv2v_reg ;
  assign \nz.mem [1618] = \nz.mem_1618_sv2v_reg ;
  assign \nz.mem [1617] = \nz.mem_1617_sv2v_reg ;
  assign \nz.mem [1616] = \nz.mem_1616_sv2v_reg ;
  assign \nz.mem [1615] = \nz.mem_1615_sv2v_reg ;
  assign \nz.mem [1614] = \nz.mem_1614_sv2v_reg ;
  assign \nz.mem [1613] = \nz.mem_1613_sv2v_reg ;
  assign \nz.mem [1612] = \nz.mem_1612_sv2v_reg ;
  assign \nz.mem [1611] = \nz.mem_1611_sv2v_reg ;
  assign \nz.mem [1610] = \nz.mem_1610_sv2v_reg ;
  assign \nz.mem [1609] = \nz.mem_1609_sv2v_reg ;
  assign \nz.mem [1608] = \nz.mem_1608_sv2v_reg ;
  assign \nz.mem [1607] = \nz.mem_1607_sv2v_reg ;
  assign \nz.mem [1606] = \nz.mem_1606_sv2v_reg ;
  assign \nz.mem [1605] = \nz.mem_1605_sv2v_reg ;
  assign \nz.mem [1604] = \nz.mem_1604_sv2v_reg ;
  assign \nz.mem [1603] = \nz.mem_1603_sv2v_reg ;
  assign \nz.mem [1602] = \nz.mem_1602_sv2v_reg ;
  assign \nz.mem [1601] = \nz.mem_1601_sv2v_reg ;
  assign \nz.mem [1600] = \nz.mem_1600_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [7] = (N277)? \nz.mem [7] : 
                            (N279)? \nz.mem [15] : 
                            (N281)? \nz.mem [23] : 
                            (N283)? \nz.mem [31] : 
                            (N285)? \nz.mem [39] : 
                            (N287)? \nz.mem [47] : 
                            (N289)? \nz.mem [55] : 
                            (N291)? \nz.mem [63] : 
                            (N293)? \nz.mem [71] : 
                            (N295)? \nz.mem [79] : 
                            (N297)? \nz.mem [87] : 
                            (N299)? \nz.mem [95] : 
                            (N301)? \nz.mem [103] : 
                            (N303)? \nz.mem [111] : 
                            (N305)? \nz.mem [119] : 
                            (N307)? \nz.mem [127] : 
                            (N309)? \nz.mem [135] : 
                            (N311)? \nz.mem [143] : 
                            (N313)? \nz.mem [151] : 
                            (N315)? \nz.mem [159] : 
                            (N317)? \nz.mem [167] : 
                            (N319)? \nz.mem [175] : 
                            (N321)? \nz.mem [183] : 
                            (N323)? \nz.mem [191] : 
                            (N325)? \nz.mem [199] : 
                            (N327)? \nz.mem [207] : 
                            (N329)? \nz.mem [215] : 
                            (N331)? \nz.mem [223] : 
                            (N333)? \nz.mem [231] : 
                            (N335)? \nz.mem [239] : 
                            (N337)? \nz.mem [247] : 
                            (N339)? \nz.mem [255] : 
                            (N341)? \nz.mem [263] : 
                            (N343)? \nz.mem [271] : 
                            (N345)? \nz.mem [279] : 
                            (N347)? \nz.mem [287] : 
                            (N349)? \nz.mem [295] : 
                            (N351)? \nz.mem [303] : 
                            (N353)? \nz.mem [311] : 
                            (N355)? \nz.mem [319] : 
                            (N357)? \nz.mem [327] : 
                            (N359)? \nz.mem [335] : 
                            (N361)? \nz.mem [343] : 
                            (N363)? \nz.mem [351] : 
                            (N365)? \nz.mem [359] : 
                            (N367)? \nz.mem [367] : 
                            (N369)? \nz.mem [375] : 
                            (N371)? \nz.mem [383] : 
                            (N373)? \nz.mem [391] : 
                            (N375)? \nz.mem [399] : 
                            (N377)? \nz.mem [407] : 
                            (N379)? \nz.mem [415] : 
                            (N381)? \nz.mem [423] : 
                            (N383)? \nz.mem [431] : 
                            (N385)? \nz.mem [439] : 
                            (N387)? \nz.mem [447] : 
                            (N389)? \nz.mem [455] : 
                            (N391)? \nz.mem [463] : 
                            (N393)? \nz.mem [471] : 
                            (N395)? \nz.mem [479] : 
                            (N397)? \nz.mem [487] : 
                            (N399)? \nz.mem [495] : 
                            (N401)? \nz.mem [503] : 
                            (N403)? \nz.mem [511] : 
                            (N405)? \nz.mem [519] : 
                            (N407)? \nz.mem [527] : 
                            (N409)? \nz.mem [535] : 
                            (N411)? \nz.mem [543] : 
                            (N413)? \nz.mem [551] : 
                            (N415)? \nz.mem [559] : 
                            (N417)? \nz.mem [567] : 
                            (N419)? \nz.mem [575] : 
                            (N421)? \nz.mem [583] : 
                            (N423)? \nz.mem [591] : 
                            (N425)? \nz.mem [599] : 
                            (N427)? \nz.mem [607] : 
                            (N429)? \nz.mem [615] : 
                            (N431)? \nz.mem [623] : 
                            (N433)? \nz.mem [631] : 
                            (N435)? \nz.mem [639] : 
                            (N437)? \nz.mem [647] : 
                            (N439)? \nz.mem [655] : 
                            (N441)? \nz.mem [663] : 
                            (N443)? \nz.mem [671] : 
                            (N445)? \nz.mem [679] : 
                            (N447)? \nz.mem [687] : 
                            (N449)? \nz.mem [695] : 
                            (N451)? \nz.mem [703] : 
                            (N453)? \nz.mem [711] : 
                            (N455)? \nz.mem [719] : 
                            (N457)? \nz.mem [727] : 
                            (N459)? \nz.mem [735] : 
                            (N461)? \nz.mem [743] : 
                            (N463)? \nz.mem [751] : 
                            (N465)? \nz.mem [759] : 
                            (N467)? \nz.mem [767] : 
                            (N469)? \nz.mem [775] : 
                            (N471)? \nz.mem [783] : 
                            (N473)? \nz.mem [791] : 
                            (N475)? \nz.mem [799] : 
                            (N477)? \nz.mem [807] : 
                            (N479)? \nz.mem [815] : 
                            (N481)? \nz.mem [823] : 
                            (N483)? \nz.mem [831] : 
                            (N485)? \nz.mem [839] : 
                            (N487)? \nz.mem [847] : 
                            (N489)? \nz.mem [855] : 
                            (N491)? \nz.mem [863] : 
                            (N493)? \nz.mem [871] : 
                            (N495)? \nz.mem [879] : 
                            (N497)? \nz.mem [887] : 
                            (N499)? \nz.mem [895] : 
                            (N501)? \nz.mem [903] : 
                            (N503)? \nz.mem [911] : 
                            (N505)? \nz.mem [919] : 
                            (N507)? \nz.mem [927] : 
                            (N509)? \nz.mem [935] : 
                            (N511)? \nz.mem [943] : 
                            (N513)? \nz.mem [951] : 
                            (N515)? \nz.mem [959] : 
                            (N517)? \nz.mem [967] : 
                            (N519)? \nz.mem [975] : 
                            (N521)? \nz.mem [983] : 
                            (N523)? \nz.mem [991] : 
                            (N525)? \nz.mem [999] : 
                            (N527)? \nz.mem [1007] : 
                            (N529)? \nz.mem [1015] : 
                            (N531)? \nz.mem [1023] : 
                            (N278)? \nz.mem [1031] : 
                            (N280)? \nz.mem [1039] : 
                            (N282)? \nz.mem [1047] : 
                            (N284)? \nz.mem [1055] : 
                            (N286)? \nz.mem [1063] : 
                            (N288)? \nz.mem [1071] : 
                            (N290)? \nz.mem [1079] : 
                            (N292)? \nz.mem [1087] : 
                            (N294)? \nz.mem [1095] : 
                            (N296)? \nz.mem [1103] : 
                            (N298)? \nz.mem [1111] : 
                            (N300)? \nz.mem [1119] : 
                            (N302)? \nz.mem [1127] : 
                            (N304)? \nz.mem [1135] : 
                            (N306)? \nz.mem [1143] : 
                            (N308)? \nz.mem [1151] : 
                            (N310)? \nz.mem [1159] : 
                            (N312)? \nz.mem [1167] : 
                            (N314)? \nz.mem [1175] : 
                            (N316)? \nz.mem [1183] : 
                            (N318)? \nz.mem [1191] : 
                            (N320)? \nz.mem [1199] : 
                            (N322)? \nz.mem [1207] : 
                            (N324)? \nz.mem [1215] : 
                            (N326)? \nz.mem [1223] : 
                            (N328)? \nz.mem [1231] : 
                            (N330)? \nz.mem [1239] : 
                            (N332)? \nz.mem [1247] : 
                            (N334)? \nz.mem [1255] : 
                            (N336)? \nz.mem [1263] : 
                            (N338)? \nz.mem [1271] : 
                            (N340)? \nz.mem [1279] : 
                            (N342)? \nz.mem [1287] : 
                            (N344)? \nz.mem [1295] : 
                            (N346)? \nz.mem [1303] : 
                            (N348)? \nz.mem [1311] : 
                            (N350)? \nz.mem [1319] : 
                            (N352)? \nz.mem [1327] : 
                            (N354)? \nz.mem [1335] : 
                            (N356)? \nz.mem [1343] : 
                            (N358)? \nz.mem [1351] : 
                            (N360)? \nz.mem [1359] : 
                            (N362)? \nz.mem [1367] : 
                            (N364)? \nz.mem [1375] : 
                            (N366)? \nz.mem [1383] : 
                            (N368)? \nz.mem [1391] : 
                            (N370)? \nz.mem [1399] : 
                            (N372)? \nz.mem [1407] : 
                            (N374)? \nz.mem [1415] : 
                            (N376)? \nz.mem [1423] : 
                            (N378)? \nz.mem [1431] : 
                            (N380)? \nz.mem [1439] : 
                            (N382)? \nz.mem [1447] : 
                            (N384)? \nz.mem [1455] : 
                            (N386)? \nz.mem [1463] : 
                            (N388)? \nz.mem [1471] : 
                            (N390)? \nz.mem [1479] : 
                            (N392)? \nz.mem [1487] : 
                            (N394)? \nz.mem [1495] : 
                            (N396)? \nz.mem [1503] : 
                            (N398)? \nz.mem [1511] : 
                            (N400)? \nz.mem [1519] : 
                            (N402)? \nz.mem [1527] : 
                            (N404)? \nz.mem [1535] : 
                            (N406)? \nz.mem [1543] : 
                            (N408)? \nz.mem [1551] : 
                            (N410)? \nz.mem [1559] : 
                            (N412)? \nz.mem [1567] : 
                            (N414)? \nz.mem [1575] : 
                            (N416)? \nz.mem [1583] : 
                            (N418)? \nz.mem [1591] : 
                            (N420)? \nz.mem [1599] : 
                            (N422)? \nz.mem [1607] : 
                            (N424)? \nz.mem [1615] : 
                            (N426)? \nz.mem [1623] : 
                            (N428)? \nz.mem [1631] : 
                            (N430)? \nz.mem [1639] : 
                            (N432)? \nz.mem [1647] : 
                            (N434)? \nz.mem [1655] : 
                            (N436)? \nz.mem [1663] : 
                            (N438)? \nz.mem [1671] : 
                            (N440)? \nz.mem [1679] : 
                            (N442)? \nz.mem [1687] : 
                            (N444)? \nz.mem [1695] : 
                            (N446)? \nz.mem [1703] : 
                            (N448)? \nz.mem [1711] : 
                            (N450)? \nz.mem [1719] : 
                            (N452)? \nz.mem [1727] : 
                            (N454)? \nz.mem [1735] : 
                            (N456)? \nz.mem [1743] : 
                            (N458)? \nz.mem [1751] : 
                            (N460)? \nz.mem [1759] : 
                            (N462)? \nz.mem [1767] : 
                            (N464)? \nz.mem [1775] : 
                            (N466)? \nz.mem [1783] : 
                            (N468)? \nz.mem [1791] : 
                            (N470)? \nz.mem [1799] : 
                            (N472)? \nz.mem [1807] : 
                            (N474)? \nz.mem [1815] : 
                            (N476)? \nz.mem [1823] : 
                            (N478)? \nz.mem [1831] : 
                            (N480)? \nz.mem [1839] : 
                            (N482)? \nz.mem [1847] : 
                            (N484)? \nz.mem [1855] : 
                            (N486)? \nz.mem [1863] : 
                            (N488)? \nz.mem [1871] : 
                            (N490)? \nz.mem [1879] : 
                            (N492)? \nz.mem [1887] : 
                            (N494)? \nz.mem [1895] : 
                            (N496)? \nz.mem [1903] : 
                            (N498)? \nz.mem [1911] : 
                            (N500)? \nz.mem [1919] : 
                            (N502)? \nz.mem [1927] : 
                            (N504)? \nz.mem [1935] : 
                            (N506)? \nz.mem [1943] : 
                            (N508)? \nz.mem [1951] : 
                            (N510)? \nz.mem [1959] : 
                            (N512)? \nz.mem [1967] : 
                            (N514)? \nz.mem [1975] : 
                            (N516)? \nz.mem [1983] : 
                            (N518)? \nz.mem [1991] : 
                            (N520)? \nz.mem [1999] : 
                            (N522)? \nz.mem [2007] : 
                            (N524)? \nz.mem [2015] : 
                            (N526)? \nz.mem [2023] : 
                            (N528)? \nz.mem [2031] : 
                            (N530)? \nz.mem [2039] : 
                            (N532)? \nz.mem [2047] : 1'b0;
  assign \nz.data_out [6] = (N277)? \nz.mem [6] : 
                            (N279)? \nz.mem [14] : 
                            (N281)? \nz.mem [22] : 
                            (N283)? \nz.mem [30] : 
                            (N285)? \nz.mem [38] : 
                            (N287)? \nz.mem [46] : 
                            (N289)? \nz.mem [54] : 
                            (N291)? \nz.mem [62] : 
                            (N293)? \nz.mem [70] : 
                            (N295)? \nz.mem [78] : 
                            (N297)? \nz.mem [86] : 
                            (N299)? \nz.mem [94] : 
                            (N301)? \nz.mem [102] : 
                            (N303)? \nz.mem [110] : 
                            (N305)? \nz.mem [118] : 
                            (N307)? \nz.mem [126] : 
                            (N309)? \nz.mem [134] : 
                            (N311)? \nz.mem [142] : 
                            (N313)? \nz.mem [150] : 
                            (N315)? \nz.mem [158] : 
                            (N317)? \nz.mem [166] : 
                            (N319)? \nz.mem [174] : 
                            (N321)? \nz.mem [182] : 
                            (N323)? \nz.mem [190] : 
                            (N325)? \nz.mem [198] : 
                            (N327)? \nz.mem [206] : 
                            (N329)? \nz.mem [214] : 
                            (N331)? \nz.mem [222] : 
                            (N333)? \nz.mem [230] : 
                            (N335)? \nz.mem [238] : 
                            (N337)? \nz.mem [246] : 
                            (N339)? \nz.mem [254] : 
                            (N341)? \nz.mem [262] : 
                            (N343)? \nz.mem [270] : 
                            (N345)? \nz.mem [278] : 
                            (N347)? \nz.mem [286] : 
                            (N349)? \nz.mem [294] : 
                            (N351)? \nz.mem [302] : 
                            (N353)? \nz.mem [310] : 
                            (N355)? \nz.mem [318] : 
                            (N357)? \nz.mem [326] : 
                            (N359)? \nz.mem [334] : 
                            (N361)? \nz.mem [342] : 
                            (N363)? \nz.mem [350] : 
                            (N365)? \nz.mem [358] : 
                            (N367)? \nz.mem [366] : 
                            (N369)? \nz.mem [374] : 
                            (N371)? \nz.mem [382] : 
                            (N373)? \nz.mem [390] : 
                            (N375)? \nz.mem [398] : 
                            (N377)? \nz.mem [406] : 
                            (N379)? \nz.mem [414] : 
                            (N381)? \nz.mem [422] : 
                            (N383)? \nz.mem [430] : 
                            (N385)? \nz.mem [438] : 
                            (N387)? \nz.mem [446] : 
                            (N389)? \nz.mem [454] : 
                            (N391)? \nz.mem [462] : 
                            (N393)? \nz.mem [470] : 
                            (N395)? \nz.mem [478] : 
                            (N397)? \nz.mem [486] : 
                            (N399)? \nz.mem [494] : 
                            (N401)? \nz.mem [502] : 
                            (N403)? \nz.mem [510] : 
                            (N405)? \nz.mem [518] : 
                            (N407)? \nz.mem [526] : 
                            (N409)? \nz.mem [534] : 
                            (N411)? \nz.mem [542] : 
                            (N413)? \nz.mem [550] : 
                            (N415)? \nz.mem [558] : 
                            (N417)? \nz.mem [566] : 
                            (N419)? \nz.mem [574] : 
                            (N421)? \nz.mem [582] : 
                            (N423)? \nz.mem [590] : 
                            (N425)? \nz.mem [598] : 
                            (N427)? \nz.mem [606] : 
                            (N429)? \nz.mem [614] : 
                            (N431)? \nz.mem [622] : 
                            (N433)? \nz.mem [630] : 
                            (N435)? \nz.mem [638] : 
                            (N437)? \nz.mem [646] : 
                            (N439)? \nz.mem [654] : 
                            (N441)? \nz.mem [662] : 
                            (N443)? \nz.mem [670] : 
                            (N445)? \nz.mem [678] : 
                            (N447)? \nz.mem [686] : 
                            (N449)? \nz.mem [694] : 
                            (N451)? \nz.mem [702] : 
                            (N453)? \nz.mem [710] : 
                            (N455)? \nz.mem [718] : 
                            (N457)? \nz.mem [726] : 
                            (N459)? \nz.mem [734] : 
                            (N461)? \nz.mem [742] : 
                            (N463)? \nz.mem [750] : 
                            (N465)? \nz.mem [758] : 
                            (N467)? \nz.mem [766] : 
                            (N469)? \nz.mem [774] : 
                            (N471)? \nz.mem [782] : 
                            (N473)? \nz.mem [790] : 
                            (N475)? \nz.mem [798] : 
                            (N477)? \nz.mem [806] : 
                            (N479)? \nz.mem [814] : 
                            (N481)? \nz.mem [822] : 
                            (N483)? \nz.mem [830] : 
                            (N485)? \nz.mem [838] : 
                            (N487)? \nz.mem [846] : 
                            (N489)? \nz.mem [854] : 
                            (N491)? \nz.mem [862] : 
                            (N493)? \nz.mem [870] : 
                            (N495)? \nz.mem [878] : 
                            (N497)? \nz.mem [886] : 
                            (N499)? \nz.mem [894] : 
                            (N501)? \nz.mem [902] : 
                            (N503)? \nz.mem [910] : 
                            (N505)? \nz.mem [918] : 
                            (N507)? \nz.mem [926] : 
                            (N509)? \nz.mem [934] : 
                            (N511)? \nz.mem [942] : 
                            (N513)? \nz.mem [950] : 
                            (N515)? \nz.mem [958] : 
                            (N517)? \nz.mem [966] : 
                            (N519)? \nz.mem [974] : 
                            (N521)? \nz.mem [982] : 
                            (N523)? \nz.mem [990] : 
                            (N525)? \nz.mem [998] : 
                            (N527)? \nz.mem [1006] : 
                            (N529)? \nz.mem [1014] : 
                            (N531)? \nz.mem [1022] : 
                            (N278)? \nz.mem [1030] : 
                            (N280)? \nz.mem [1038] : 
                            (N282)? \nz.mem [1046] : 
                            (N284)? \nz.mem [1054] : 
                            (N286)? \nz.mem [1062] : 
                            (N288)? \nz.mem [1070] : 
                            (N290)? \nz.mem [1078] : 
                            (N292)? \nz.mem [1086] : 
                            (N294)? \nz.mem [1094] : 
                            (N296)? \nz.mem [1102] : 
                            (N298)? \nz.mem [1110] : 
                            (N300)? \nz.mem [1118] : 
                            (N302)? \nz.mem [1126] : 
                            (N304)? \nz.mem [1134] : 
                            (N306)? \nz.mem [1142] : 
                            (N308)? \nz.mem [1150] : 
                            (N310)? \nz.mem [1158] : 
                            (N312)? \nz.mem [1166] : 
                            (N314)? \nz.mem [1174] : 
                            (N316)? \nz.mem [1182] : 
                            (N318)? \nz.mem [1190] : 
                            (N320)? \nz.mem [1198] : 
                            (N322)? \nz.mem [1206] : 
                            (N324)? \nz.mem [1214] : 
                            (N326)? \nz.mem [1222] : 
                            (N328)? \nz.mem [1230] : 
                            (N330)? \nz.mem [1238] : 
                            (N332)? \nz.mem [1246] : 
                            (N334)? \nz.mem [1254] : 
                            (N336)? \nz.mem [1262] : 
                            (N338)? \nz.mem [1270] : 
                            (N340)? \nz.mem [1278] : 
                            (N342)? \nz.mem [1286] : 
                            (N344)? \nz.mem [1294] : 
                            (N346)? \nz.mem [1302] : 
                            (N348)? \nz.mem [1310] : 
                            (N350)? \nz.mem [1318] : 
                            (N352)? \nz.mem [1326] : 
                            (N354)? \nz.mem [1334] : 
                            (N356)? \nz.mem [1342] : 
                            (N358)? \nz.mem [1350] : 
                            (N360)? \nz.mem [1358] : 
                            (N362)? \nz.mem [1366] : 
                            (N364)? \nz.mem [1374] : 
                            (N366)? \nz.mem [1382] : 
                            (N368)? \nz.mem [1390] : 
                            (N370)? \nz.mem [1398] : 
                            (N372)? \nz.mem [1406] : 
                            (N374)? \nz.mem [1414] : 
                            (N376)? \nz.mem [1422] : 
                            (N378)? \nz.mem [1430] : 
                            (N380)? \nz.mem [1438] : 
                            (N382)? \nz.mem [1446] : 
                            (N384)? \nz.mem [1454] : 
                            (N386)? \nz.mem [1462] : 
                            (N388)? \nz.mem [1470] : 
                            (N390)? \nz.mem [1478] : 
                            (N392)? \nz.mem [1486] : 
                            (N394)? \nz.mem [1494] : 
                            (N396)? \nz.mem [1502] : 
                            (N398)? \nz.mem [1510] : 
                            (N400)? \nz.mem [1518] : 
                            (N402)? \nz.mem [1526] : 
                            (N404)? \nz.mem [1534] : 
                            (N406)? \nz.mem [1542] : 
                            (N408)? \nz.mem [1550] : 
                            (N410)? \nz.mem [1558] : 
                            (N412)? \nz.mem [1566] : 
                            (N414)? \nz.mem [1574] : 
                            (N416)? \nz.mem [1582] : 
                            (N418)? \nz.mem [1590] : 
                            (N420)? \nz.mem [1598] : 
                            (N422)? \nz.mem [1606] : 
                            (N424)? \nz.mem [1614] : 
                            (N426)? \nz.mem [1622] : 
                            (N428)? \nz.mem [1630] : 
                            (N430)? \nz.mem [1638] : 
                            (N432)? \nz.mem [1646] : 
                            (N434)? \nz.mem [1654] : 
                            (N436)? \nz.mem [1662] : 
                            (N438)? \nz.mem [1670] : 
                            (N440)? \nz.mem [1678] : 
                            (N442)? \nz.mem [1686] : 
                            (N444)? \nz.mem [1694] : 
                            (N446)? \nz.mem [1702] : 
                            (N448)? \nz.mem [1710] : 
                            (N450)? \nz.mem [1718] : 
                            (N452)? \nz.mem [1726] : 
                            (N454)? \nz.mem [1734] : 
                            (N456)? \nz.mem [1742] : 
                            (N458)? \nz.mem [1750] : 
                            (N460)? \nz.mem [1758] : 
                            (N462)? \nz.mem [1766] : 
                            (N464)? \nz.mem [1774] : 
                            (N466)? \nz.mem [1782] : 
                            (N468)? \nz.mem [1790] : 
                            (N470)? \nz.mem [1798] : 
                            (N472)? \nz.mem [1806] : 
                            (N474)? \nz.mem [1814] : 
                            (N476)? \nz.mem [1822] : 
                            (N478)? \nz.mem [1830] : 
                            (N480)? \nz.mem [1838] : 
                            (N482)? \nz.mem [1846] : 
                            (N484)? \nz.mem [1854] : 
                            (N486)? \nz.mem [1862] : 
                            (N488)? \nz.mem [1870] : 
                            (N490)? \nz.mem [1878] : 
                            (N492)? \nz.mem [1886] : 
                            (N494)? \nz.mem [1894] : 
                            (N496)? \nz.mem [1902] : 
                            (N498)? \nz.mem [1910] : 
                            (N500)? \nz.mem [1918] : 
                            (N502)? \nz.mem [1926] : 
                            (N504)? \nz.mem [1934] : 
                            (N506)? \nz.mem [1942] : 
                            (N508)? \nz.mem [1950] : 
                            (N510)? \nz.mem [1958] : 
                            (N512)? \nz.mem [1966] : 
                            (N514)? \nz.mem [1974] : 
                            (N516)? \nz.mem [1982] : 
                            (N518)? \nz.mem [1990] : 
                            (N520)? \nz.mem [1998] : 
                            (N522)? \nz.mem [2006] : 
                            (N524)? \nz.mem [2014] : 
                            (N526)? \nz.mem [2022] : 
                            (N528)? \nz.mem [2030] : 
                            (N530)? \nz.mem [2038] : 
                            (N532)? \nz.mem [2046] : 1'b0;
  assign \nz.data_out [5] = (N277)? \nz.mem [5] : 
                            (N279)? \nz.mem [13] : 
                            (N281)? \nz.mem [21] : 
                            (N283)? \nz.mem [29] : 
                            (N285)? \nz.mem [37] : 
                            (N287)? \nz.mem [45] : 
                            (N289)? \nz.mem [53] : 
                            (N291)? \nz.mem [61] : 
                            (N293)? \nz.mem [69] : 
                            (N295)? \nz.mem [77] : 
                            (N297)? \nz.mem [85] : 
                            (N299)? \nz.mem [93] : 
                            (N301)? \nz.mem [101] : 
                            (N303)? \nz.mem [109] : 
                            (N305)? \nz.mem [117] : 
                            (N307)? \nz.mem [125] : 
                            (N309)? \nz.mem [133] : 
                            (N311)? \nz.mem [141] : 
                            (N313)? \nz.mem [149] : 
                            (N315)? \nz.mem [157] : 
                            (N317)? \nz.mem [165] : 
                            (N319)? \nz.mem [173] : 
                            (N321)? \nz.mem [181] : 
                            (N323)? \nz.mem [189] : 
                            (N325)? \nz.mem [197] : 
                            (N327)? \nz.mem [205] : 
                            (N329)? \nz.mem [213] : 
                            (N331)? \nz.mem [221] : 
                            (N333)? \nz.mem [229] : 
                            (N335)? \nz.mem [237] : 
                            (N337)? \nz.mem [245] : 
                            (N339)? \nz.mem [253] : 
                            (N341)? \nz.mem [261] : 
                            (N343)? \nz.mem [269] : 
                            (N345)? \nz.mem [277] : 
                            (N347)? \nz.mem [285] : 
                            (N349)? \nz.mem [293] : 
                            (N351)? \nz.mem [301] : 
                            (N353)? \nz.mem [309] : 
                            (N355)? \nz.mem [317] : 
                            (N357)? \nz.mem [325] : 
                            (N359)? \nz.mem [333] : 
                            (N361)? \nz.mem [341] : 
                            (N363)? \nz.mem [349] : 
                            (N365)? \nz.mem [357] : 
                            (N367)? \nz.mem [365] : 
                            (N369)? \nz.mem [373] : 
                            (N371)? \nz.mem [381] : 
                            (N373)? \nz.mem [389] : 
                            (N375)? \nz.mem [397] : 
                            (N377)? \nz.mem [405] : 
                            (N379)? \nz.mem [413] : 
                            (N381)? \nz.mem [421] : 
                            (N383)? \nz.mem [429] : 
                            (N385)? \nz.mem [437] : 
                            (N387)? \nz.mem [445] : 
                            (N389)? \nz.mem [453] : 
                            (N391)? \nz.mem [461] : 
                            (N393)? \nz.mem [469] : 
                            (N395)? \nz.mem [477] : 
                            (N397)? \nz.mem [485] : 
                            (N399)? \nz.mem [493] : 
                            (N401)? \nz.mem [501] : 
                            (N403)? \nz.mem [509] : 
                            (N405)? \nz.mem [517] : 
                            (N407)? \nz.mem [525] : 
                            (N409)? \nz.mem [533] : 
                            (N411)? \nz.mem [541] : 
                            (N413)? \nz.mem [549] : 
                            (N415)? \nz.mem [557] : 
                            (N417)? \nz.mem [565] : 
                            (N419)? \nz.mem [573] : 
                            (N421)? \nz.mem [581] : 
                            (N423)? \nz.mem [589] : 
                            (N425)? \nz.mem [597] : 
                            (N427)? \nz.mem [605] : 
                            (N429)? \nz.mem [613] : 
                            (N431)? \nz.mem [621] : 
                            (N433)? \nz.mem [629] : 
                            (N435)? \nz.mem [637] : 
                            (N437)? \nz.mem [645] : 
                            (N439)? \nz.mem [653] : 
                            (N441)? \nz.mem [661] : 
                            (N443)? \nz.mem [669] : 
                            (N445)? \nz.mem [677] : 
                            (N447)? \nz.mem [685] : 
                            (N449)? \nz.mem [693] : 
                            (N451)? \nz.mem [701] : 
                            (N453)? \nz.mem [709] : 
                            (N455)? \nz.mem [717] : 
                            (N457)? \nz.mem [725] : 
                            (N459)? \nz.mem [733] : 
                            (N461)? \nz.mem [741] : 
                            (N463)? \nz.mem [749] : 
                            (N465)? \nz.mem [757] : 
                            (N467)? \nz.mem [765] : 
                            (N469)? \nz.mem [773] : 
                            (N471)? \nz.mem [781] : 
                            (N473)? \nz.mem [789] : 
                            (N475)? \nz.mem [797] : 
                            (N477)? \nz.mem [805] : 
                            (N479)? \nz.mem [813] : 
                            (N481)? \nz.mem [821] : 
                            (N483)? \nz.mem [829] : 
                            (N485)? \nz.mem [837] : 
                            (N487)? \nz.mem [845] : 
                            (N489)? \nz.mem [853] : 
                            (N491)? \nz.mem [861] : 
                            (N493)? \nz.mem [869] : 
                            (N495)? \nz.mem [877] : 
                            (N497)? \nz.mem [885] : 
                            (N499)? \nz.mem [893] : 
                            (N501)? \nz.mem [901] : 
                            (N503)? \nz.mem [909] : 
                            (N505)? \nz.mem [917] : 
                            (N507)? \nz.mem [925] : 
                            (N509)? \nz.mem [933] : 
                            (N511)? \nz.mem [941] : 
                            (N513)? \nz.mem [949] : 
                            (N515)? \nz.mem [957] : 
                            (N517)? \nz.mem [965] : 
                            (N519)? \nz.mem [973] : 
                            (N521)? \nz.mem [981] : 
                            (N523)? \nz.mem [989] : 
                            (N525)? \nz.mem [997] : 
                            (N527)? \nz.mem [1005] : 
                            (N529)? \nz.mem [1013] : 
                            (N531)? \nz.mem [1021] : 
                            (N278)? \nz.mem [1029] : 
                            (N280)? \nz.mem [1037] : 
                            (N282)? \nz.mem [1045] : 
                            (N284)? \nz.mem [1053] : 
                            (N286)? \nz.mem [1061] : 
                            (N288)? \nz.mem [1069] : 
                            (N290)? \nz.mem [1077] : 
                            (N292)? \nz.mem [1085] : 
                            (N294)? \nz.mem [1093] : 
                            (N296)? \nz.mem [1101] : 
                            (N298)? \nz.mem [1109] : 
                            (N300)? \nz.mem [1117] : 
                            (N302)? \nz.mem [1125] : 
                            (N304)? \nz.mem [1133] : 
                            (N306)? \nz.mem [1141] : 
                            (N308)? \nz.mem [1149] : 
                            (N310)? \nz.mem [1157] : 
                            (N312)? \nz.mem [1165] : 
                            (N314)? \nz.mem [1173] : 
                            (N316)? \nz.mem [1181] : 
                            (N318)? \nz.mem [1189] : 
                            (N320)? \nz.mem [1197] : 
                            (N322)? \nz.mem [1205] : 
                            (N324)? \nz.mem [1213] : 
                            (N326)? \nz.mem [1221] : 
                            (N328)? \nz.mem [1229] : 
                            (N330)? \nz.mem [1237] : 
                            (N332)? \nz.mem [1245] : 
                            (N334)? \nz.mem [1253] : 
                            (N336)? \nz.mem [1261] : 
                            (N338)? \nz.mem [1269] : 
                            (N340)? \nz.mem [1277] : 
                            (N342)? \nz.mem [1285] : 
                            (N344)? \nz.mem [1293] : 
                            (N346)? \nz.mem [1301] : 
                            (N348)? \nz.mem [1309] : 
                            (N350)? \nz.mem [1317] : 
                            (N352)? \nz.mem [1325] : 
                            (N354)? \nz.mem [1333] : 
                            (N356)? \nz.mem [1341] : 
                            (N358)? \nz.mem [1349] : 
                            (N360)? \nz.mem [1357] : 
                            (N362)? \nz.mem [1365] : 
                            (N364)? \nz.mem [1373] : 
                            (N366)? \nz.mem [1381] : 
                            (N368)? \nz.mem [1389] : 
                            (N370)? \nz.mem [1397] : 
                            (N372)? \nz.mem [1405] : 
                            (N374)? \nz.mem [1413] : 
                            (N376)? \nz.mem [1421] : 
                            (N378)? \nz.mem [1429] : 
                            (N380)? \nz.mem [1437] : 
                            (N382)? \nz.mem [1445] : 
                            (N384)? \nz.mem [1453] : 
                            (N386)? \nz.mem [1461] : 
                            (N388)? \nz.mem [1469] : 
                            (N390)? \nz.mem [1477] : 
                            (N392)? \nz.mem [1485] : 
                            (N394)? \nz.mem [1493] : 
                            (N396)? \nz.mem [1501] : 
                            (N398)? \nz.mem [1509] : 
                            (N400)? \nz.mem [1517] : 
                            (N402)? \nz.mem [1525] : 
                            (N404)? \nz.mem [1533] : 
                            (N406)? \nz.mem [1541] : 
                            (N408)? \nz.mem [1549] : 
                            (N410)? \nz.mem [1557] : 
                            (N412)? \nz.mem [1565] : 
                            (N414)? \nz.mem [1573] : 
                            (N416)? \nz.mem [1581] : 
                            (N418)? \nz.mem [1589] : 
                            (N420)? \nz.mem [1597] : 
                            (N422)? \nz.mem [1605] : 
                            (N424)? \nz.mem [1613] : 
                            (N426)? \nz.mem [1621] : 
                            (N428)? \nz.mem [1629] : 
                            (N430)? \nz.mem [1637] : 
                            (N432)? \nz.mem [1645] : 
                            (N434)? \nz.mem [1653] : 
                            (N436)? \nz.mem [1661] : 
                            (N438)? \nz.mem [1669] : 
                            (N440)? \nz.mem [1677] : 
                            (N442)? \nz.mem [1685] : 
                            (N444)? \nz.mem [1693] : 
                            (N446)? \nz.mem [1701] : 
                            (N448)? \nz.mem [1709] : 
                            (N450)? \nz.mem [1717] : 
                            (N452)? \nz.mem [1725] : 
                            (N454)? \nz.mem [1733] : 
                            (N456)? \nz.mem [1741] : 
                            (N458)? \nz.mem [1749] : 
                            (N460)? \nz.mem [1757] : 
                            (N462)? \nz.mem [1765] : 
                            (N464)? \nz.mem [1773] : 
                            (N466)? \nz.mem [1781] : 
                            (N468)? \nz.mem [1789] : 
                            (N470)? \nz.mem [1797] : 
                            (N472)? \nz.mem [1805] : 
                            (N474)? \nz.mem [1813] : 
                            (N476)? \nz.mem [1821] : 
                            (N478)? \nz.mem [1829] : 
                            (N480)? \nz.mem [1837] : 
                            (N482)? \nz.mem [1845] : 
                            (N484)? \nz.mem [1853] : 
                            (N486)? \nz.mem [1861] : 
                            (N488)? \nz.mem [1869] : 
                            (N490)? \nz.mem [1877] : 
                            (N492)? \nz.mem [1885] : 
                            (N494)? \nz.mem [1893] : 
                            (N496)? \nz.mem [1901] : 
                            (N498)? \nz.mem [1909] : 
                            (N500)? \nz.mem [1917] : 
                            (N502)? \nz.mem [1925] : 
                            (N504)? \nz.mem [1933] : 
                            (N506)? \nz.mem [1941] : 
                            (N508)? \nz.mem [1949] : 
                            (N510)? \nz.mem [1957] : 
                            (N512)? \nz.mem [1965] : 
                            (N514)? \nz.mem [1973] : 
                            (N516)? \nz.mem [1981] : 
                            (N518)? \nz.mem [1989] : 
                            (N520)? \nz.mem [1997] : 
                            (N522)? \nz.mem [2005] : 
                            (N524)? \nz.mem [2013] : 
                            (N526)? \nz.mem [2021] : 
                            (N528)? \nz.mem [2029] : 
                            (N530)? \nz.mem [2037] : 
                            (N532)? \nz.mem [2045] : 1'b0;
  assign \nz.data_out [4] = (N277)? \nz.mem [4] : 
                            (N279)? \nz.mem [12] : 
                            (N281)? \nz.mem [20] : 
                            (N283)? \nz.mem [28] : 
                            (N285)? \nz.mem [36] : 
                            (N287)? \nz.mem [44] : 
                            (N289)? \nz.mem [52] : 
                            (N291)? \nz.mem [60] : 
                            (N293)? \nz.mem [68] : 
                            (N295)? \nz.mem [76] : 
                            (N297)? \nz.mem [84] : 
                            (N299)? \nz.mem [92] : 
                            (N301)? \nz.mem [100] : 
                            (N303)? \nz.mem [108] : 
                            (N305)? \nz.mem [116] : 
                            (N307)? \nz.mem [124] : 
                            (N309)? \nz.mem [132] : 
                            (N311)? \nz.mem [140] : 
                            (N313)? \nz.mem [148] : 
                            (N315)? \nz.mem [156] : 
                            (N317)? \nz.mem [164] : 
                            (N319)? \nz.mem [172] : 
                            (N321)? \nz.mem [180] : 
                            (N323)? \nz.mem [188] : 
                            (N325)? \nz.mem [196] : 
                            (N327)? \nz.mem [204] : 
                            (N329)? \nz.mem [212] : 
                            (N331)? \nz.mem [220] : 
                            (N333)? \nz.mem [228] : 
                            (N335)? \nz.mem [236] : 
                            (N337)? \nz.mem [244] : 
                            (N339)? \nz.mem [252] : 
                            (N341)? \nz.mem [260] : 
                            (N343)? \nz.mem [268] : 
                            (N345)? \nz.mem [276] : 
                            (N347)? \nz.mem [284] : 
                            (N349)? \nz.mem [292] : 
                            (N351)? \nz.mem [300] : 
                            (N353)? \nz.mem [308] : 
                            (N355)? \nz.mem [316] : 
                            (N357)? \nz.mem [324] : 
                            (N359)? \nz.mem [332] : 
                            (N361)? \nz.mem [340] : 
                            (N363)? \nz.mem [348] : 
                            (N365)? \nz.mem [356] : 
                            (N367)? \nz.mem [364] : 
                            (N369)? \nz.mem [372] : 
                            (N371)? \nz.mem [380] : 
                            (N373)? \nz.mem [388] : 
                            (N375)? \nz.mem [396] : 
                            (N377)? \nz.mem [404] : 
                            (N379)? \nz.mem [412] : 
                            (N381)? \nz.mem [420] : 
                            (N383)? \nz.mem [428] : 
                            (N385)? \nz.mem [436] : 
                            (N387)? \nz.mem [444] : 
                            (N389)? \nz.mem [452] : 
                            (N391)? \nz.mem [460] : 
                            (N393)? \nz.mem [468] : 
                            (N395)? \nz.mem [476] : 
                            (N397)? \nz.mem [484] : 
                            (N399)? \nz.mem [492] : 
                            (N401)? \nz.mem [500] : 
                            (N403)? \nz.mem [508] : 
                            (N405)? \nz.mem [516] : 
                            (N407)? \nz.mem [524] : 
                            (N409)? \nz.mem [532] : 
                            (N411)? \nz.mem [540] : 
                            (N413)? \nz.mem [548] : 
                            (N415)? \nz.mem [556] : 
                            (N417)? \nz.mem [564] : 
                            (N419)? \nz.mem [572] : 
                            (N421)? \nz.mem [580] : 
                            (N423)? \nz.mem [588] : 
                            (N425)? \nz.mem [596] : 
                            (N427)? \nz.mem [604] : 
                            (N429)? \nz.mem [612] : 
                            (N431)? \nz.mem [620] : 
                            (N433)? \nz.mem [628] : 
                            (N435)? \nz.mem [636] : 
                            (N437)? \nz.mem [644] : 
                            (N439)? \nz.mem [652] : 
                            (N441)? \nz.mem [660] : 
                            (N443)? \nz.mem [668] : 
                            (N445)? \nz.mem [676] : 
                            (N447)? \nz.mem [684] : 
                            (N449)? \nz.mem [692] : 
                            (N451)? \nz.mem [700] : 
                            (N453)? \nz.mem [708] : 
                            (N455)? \nz.mem [716] : 
                            (N457)? \nz.mem [724] : 
                            (N459)? \nz.mem [732] : 
                            (N461)? \nz.mem [740] : 
                            (N463)? \nz.mem [748] : 
                            (N465)? \nz.mem [756] : 
                            (N467)? \nz.mem [764] : 
                            (N469)? \nz.mem [772] : 
                            (N471)? \nz.mem [780] : 
                            (N473)? \nz.mem [788] : 
                            (N475)? \nz.mem [796] : 
                            (N477)? \nz.mem [804] : 
                            (N479)? \nz.mem [812] : 
                            (N481)? \nz.mem [820] : 
                            (N483)? \nz.mem [828] : 
                            (N485)? \nz.mem [836] : 
                            (N487)? \nz.mem [844] : 
                            (N489)? \nz.mem [852] : 
                            (N491)? \nz.mem [860] : 
                            (N493)? \nz.mem [868] : 
                            (N495)? \nz.mem [876] : 
                            (N497)? \nz.mem [884] : 
                            (N499)? \nz.mem [892] : 
                            (N501)? \nz.mem [900] : 
                            (N503)? \nz.mem [908] : 
                            (N505)? \nz.mem [916] : 
                            (N507)? \nz.mem [924] : 
                            (N509)? \nz.mem [932] : 
                            (N511)? \nz.mem [940] : 
                            (N513)? \nz.mem [948] : 
                            (N515)? \nz.mem [956] : 
                            (N517)? \nz.mem [964] : 
                            (N519)? \nz.mem [972] : 
                            (N521)? \nz.mem [980] : 
                            (N523)? \nz.mem [988] : 
                            (N525)? \nz.mem [996] : 
                            (N527)? \nz.mem [1004] : 
                            (N529)? \nz.mem [1012] : 
                            (N531)? \nz.mem [1020] : 
                            (N278)? \nz.mem [1028] : 
                            (N280)? \nz.mem [1036] : 
                            (N282)? \nz.mem [1044] : 
                            (N284)? \nz.mem [1052] : 
                            (N286)? \nz.mem [1060] : 
                            (N288)? \nz.mem [1068] : 
                            (N290)? \nz.mem [1076] : 
                            (N292)? \nz.mem [1084] : 
                            (N294)? \nz.mem [1092] : 
                            (N296)? \nz.mem [1100] : 
                            (N298)? \nz.mem [1108] : 
                            (N300)? \nz.mem [1116] : 
                            (N302)? \nz.mem [1124] : 
                            (N304)? \nz.mem [1132] : 
                            (N306)? \nz.mem [1140] : 
                            (N308)? \nz.mem [1148] : 
                            (N310)? \nz.mem [1156] : 
                            (N312)? \nz.mem [1164] : 
                            (N314)? \nz.mem [1172] : 
                            (N316)? \nz.mem [1180] : 
                            (N318)? \nz.mem [1188] : 
                            (N320)? \nz.mem [1196] : 
                            (N322)? \nz.mem [1204] : 
                            (N324)? \nz.mem [1212] : 
                            (N326)? \nz.mem [1220] : 
                            (N328)? \nz.mem [1228] : 
                            (N330)? \nz.mem [1236] : 
                            (N332)? \nz.mem [1244] : 
                            (N334)? \nz.mem [1252] : 
                            (N336)? \nz.mem [1260] : 
                            (N338)? \nz.mem [1268] : 
                            (N340)? \nz.mem [1276] : 
                            (N342)? \nz.mem [1284] : 
                            (N344)? \nz.mem [1292] : 
                            (N346)? \nz.mem [1300] : 
                            (N348)? \nz.mem [1308] : 
                            (N350)? \nz.mem [1316] : 
                            (N352)? \nz.mem [1324] : 
                            (N354)? \nz.mem [1332] : 
                            (N356)? \nz.mem [1340] : 
                            (N358)? \nz.mem [1348] : 
                            (N360)? \nz.mem [1356] : 
                            (N362)? \nz.mem [1364] : 
                            (N364)? \nz.mem [1372] : 
                            (N366)? \nz.mem [1380] : 
                            (N368)? \nz.mem [1388] : 
                            (N370)? \nz.mem [1396] : 
                            (N372)? \nz.mem [1404] : 
                            (N374)? \nz.mem [1412] : 
                            (N376)? \nz.mem [1420] : 
                            (N378)? \nz.mem [1428] : 
                            (N380)? \nz.mem [1436] : 
                            (N382)? \nz.mem [1444] : 
                            (N384)? \nz.mem [1452] : 
                            (N386)? \nz.mem [1460] : 
                            (N388)? \nz.mem [1468] : 
                            (N390)? \nz.mem [1476] : 
                            (N392)? \nz.mem [1484] : 
                            (N394)? \nz.mem [1492] : 
                            (N396)? \nz.mem [1500] : 
                            (N398)? \nz.mem [1508] : 
                            (N400)? \nz.mem [1516] : 
                            (N402)? \nz.mem [1524] : 
                            (N404)? \nz.mem [1532] : 
                            (N406)? \nz.mem [1540] : 
                            (N408)? \nz.mem [1548] : 
                            (N410)? \nz.mem [1556] : 
                            (N412)? \nz.mem [1564] : 
                            (N414)? \nz.mem [1572] : 
                            (N416)? \nz.mem [1580] : 
                            (N418)? \nz.mem [1588] : 
                            (N420)? \nz.mem [1596] : 
                            (N422)? \nz.mem [1604] : 
                            (N424)? \nz.mem [1612] : 
                            (N426)? \nz.mem [1620] : 
                            (N428)? \nz.mem [1628] : 
                            (N430)? \nz.mem [1636] : 
                            (N432)? \nz.mem [1644] : 
                            (N434)? \nz.mem [1652] : 
                            (N436)? \nz.mem [1660] : 
                            (N438)? \nz.mem [1668] : 
                            (N440)? \nz.mem [1676] : 
                            (N442)? \nz.mem [1684] : 
                            (N444)? \nz.mem [1692] : 
                            (N446)? \nz.mem [1700] : 
                            (N448)? \nz.mem [1708] : 
                            (N450)? \nz.mem [1716] : 
                            (N452)? \nz.mem [1724] : 
                            (N454)? \nz.mem [1732] : 
                            (N456)? \nz.mem [1740] : 
                            (N458)? \nz.mem [1748] : 
                            (N460)? \nz.mem [1756] : 
                            (N462)? \nz.mem [1764] : 
                            (N464)? \nz.mem [1772] : 
                            (N466)? \nz.mem [1780] : 
                            (N468)? \nz.mem [1788] : 
                            (N470)? \nz.mem [1796] : 
                            (N472)? \nz.mem [1804] : 
                            (N474)? \nz.mem [1812] : 
                            (N476)? \nz.mem [1820] : 
                            (N478)? \nz.mem [1828] : 
                            (N480)? \nz.mem [1836] : 
                            (N482)? \nz.mem [1844] : 
                            (N484)? \nz.mem [1852] : 
                            (N486)? \nz.mem [1860] : 
                            (N488)? \nz.mem [1868] : 
                            (N490)? \nz.mem [1876] : 
                            (N492)? \nz.mem [1884] : 
                            (N494)? \nz.mem [1892] : 
                            (N496)? \nz.mem [1900] : 
                            (N498)? \nz.mem [1908] : 
                            (N500)? \nz.mem [1916] : 
                            (N502)? \nz.mem [1924] : 
                            (N504)? \nz.mem [1932] : 
                            (N506)? \nz.mem [1940] : 
                            (N508)? \nz.mem [1948] : 
                            (N510)? \nz.mem [1956] : 
                            (N512)? \nz.mem [1964] : 
                            (N514)? \nz.mem [1972] : 
                            (N516)? \nz.mem [1980] : 
                            (N518)? \nz.mem [1988] : 
                            (N520)? \nz.mem [1996] : 
                            (N522)? \nz.mem [2004] : 
                            (N524)? \nz.mem [2012] : 
                            (N526)? \nz.mem [2020] : 
                            (N528)? \nz.mem [2028] : 
                            (N530)? \nz.mem [2036] : 
                            (N532)? \nz.mem [2044] : 1'b0;
  assign \nz.data_out [3] = (N277)? \nz.mem [3] : 
                            (N279)? \nz.mem [11] : 
                            (N281)? \nz.mem [19] : 
                            (N283)? \nz.mem [27] : 
                            (N285)? \nz.mem [35] : 
                            (N287)? \nz.mem [43] : 
                            (N289)? \nz.mem [51] : 
                            (N291)? \nz.mem [59] : 
                            (N293)? \nz.mem [67] : 
                            (N295)? \nz.mem [75] : 
                            (N297)? \nz.mem [83] : 
                            (N299)? \nz.mem [91] : 
                            (N301)? \nz.mem [99] : 
                            (N303)? \nz.mem [107] : 
                            (N305)? \nz.mem [115] : 
                            (N307)? \nz.mem [123] : 
                            (N309)? \nz.mem [131] : 
                            (N311)? \nz.mem [139] : 
                            (N313)? \nz.mem [147] : 
                            (N315)? \nz.mem [155] : 
                            (N317)? \nz.mem [163] : 
                            (N319)? \nz.mem [171] : 
                            (N321)? \nz.mem [179] : 
                            (N323)? \nz.mem [187] : 
                            (N325)? \nz.mem [195] : 
                            (N327)? \nz.mem [203] : 
                            (N329)? \nz.mem [211] : 
                            (N331)? \nz.mem [219] : 
                            (N333)? \nz.mem [227] : 
                            (N335)? \nz.mem [235] : 
                            (N337)? \nz.mem [243] : 
                            (N339)? \nz.mem [251] : 
                            (N341)? \nz.mem [259] : 
                            (N343)? \nz.mem [267] : 
                            (N345)? \nz.mem [275] : 
                            (N347)? \nz.mem [283] : 
                            (N349)? \nz.mem [291] : 
                            (N351)? \nz.mem [299] : 
                            (N353)? \nz.mem [307] : 
                            (N355)? \nz.mem [315] : 
                            (N357)? \nz.mem [323] : 
                            (N359)? \nz.mem [331] : 
                            (N361)? \nz.mem [339] : 
                            (N363)? \nz.mem [347] : 
                            (N365)? \nz.mem [355] : 
                            (N367)? \nz.mem [363] : 
                            (N369)? \nz.mem [371] : 
                            (N371)? \nz.mem [379] : 
                            (N373)? \nz.mem [387] : 
                            (N375)? \nz.mem [395] : 
                            (N377)? \nz.mem [403] : 
                            (N379)? \nz.mem [411] : 
                            (N381)? \nz.mem [419] : 
                            (N383)? \nz.mem [427] : 
                            (N385)? \nz.mem [435] : 
                            (N387)? \nz.mem [443] : 
                            (N389)? \nz.mem [451] : 
                            (N391)? \nz.mem [459] : 
                            (N393)? \nz.mem [467] : 
                            (N395)? \nz.mem [475] : 
                            (N397)? \nz.mem [483] : 
                            (N399)? \nz.mem [491] : 
                            (N401)? \nz.mem [499] : 
                            (N403)? \nz.mem [507] : 
                            (N405)? \nz.mem [515] : 
                            (N407)? \nz.mem [523] : 
                            (N409)? \nz.mem [531] : 
                            (N411)? \nz.mem [539] : 
                            (N413)? \nz.mem [547] : 
                            (N415)? \nz.mem [555] : 
                            (N417)? \nz.mem [563] : 
                            (N419)? \nz.mem [571] : 
                            (N421)? \nz.mem [579] : 
                            (N423)? \nz.mem [587] : 
                            (N425)? \nz.mem [595] : 
                            (N427)? \nz.mem [603] : 
                            (N429)? \nz.mem [611] : 
                            (N431)? \nz.mem [619] : 
                            (N433)? \nz.mem [627] : 
                            (N435)? \nz.mem [635] : 
                            (N437)? \nz.mem [643] : 
                            (N439)? \nz.mem [651] : 
                            (N441)? \nz.mem [659] : 
                            (N443)? \nz.mem [667] : 
                            (N445)? \nz.mem [675] : 
                            (N447)? \nz.mem [683] : 
                            (N449)? \nz.mem [691] : 
                            (N451)? \nz.mem [699] : 
                            (N453)? \nz.mem [707] : 
                            (N455)? \nz.mem [715] : 
                            (N457)? \nz.mem [723] : 
                            (N459)? \nz.mem [731] : 
                            (N461)? \nz.mem [739] : 
                            (N463)? \nz.mem [747] : 
                            (N465)? \nz.mem [755] : 
                            (N467)? \nz.mem [763] : 
                            (N469)? \nz.mem [771] : 
                            (N471)? \nz.mem [779] : 
                            (N473)? \nz.mem [787] : 
                            (N475)? \nz.mem [795] : 
                            (N477)? \nz.mem [803] : 
                            (N479)? \nz.mem [811] : 
                            (N481)? \nz.mem [819] : 
                            (N483)? \nz.mem [827] : 
                            (N485)? \nz.mem [835] : 
                            (N487)? \nz.mem [843] : 
                            (N489)? \nz.mem [851] : 
                            (N491)? \nz.mem [859] : 
                            (N493)? \nz.mem [867] : 
                            (N495)? \nz.mem [875] : 
                            (N497)? \nz.mem [883] : 
                            (N499)? \nz.mem [891] : 
                            (N501)? \nz.mem [899] : 
                            (N503)? \nz.mem [907] : 
                            (N505)? \nz.mem [915] : 
                            (N507)? \nz.mem [923] : 
                            (N509)? \nz.mem [931] : 
                            (N511)? \nz.mem [939] : 
                            (N513)? \nz.mem [947] : 
                            (N515)? \nz.mem [955] : 
                            (N517)? \nz.mem [963] : 
                            (N519)? \nz.mem [971] : 
                            (N521)? \nz.mem [979] : 
                            (N523)? \nz.mem [987] : 
                            (N525)? \nz.mem [995] : 
                            (N527)? \nz.mem [1003] : 
                            (N529)? \nz.mem [1011] : 
                            (N531)? \nz.mem [1019] : 
                            (N278)? \nz.mem [1027] : 
                            (N280)? \nz.mem [1035] : 
                            (N282)? \nz.mem [1043] : 
                            (N284)? \nz.mem [1051] : 
                            (N286)? \nz.mem [1059] : 
                            (N288)? \nz.mem [1067] : 
                            (N290)? \nz.mem [1075] : 
                            (N292)? \nz.mem [1083] : 
                            (N294)? \nz.mem [1091] : 
                            (N296)? \nz.mem [1099] : 
                            (N298)? \nz.mem [1107] : 
                            (N300)? \nz.mem [1115] : 
                            (N302)? \nz.mem [1123] : 
                            (N304)? \nz.mem [1131] : 
                            (N306)? \nz.mem [1139] : 
                            (N308)? \nz.mem [1147] : 
                            (N310)? \nz.mem [1155] : 
                            (N312)? \nz.mem [1163] : 
                            (N314)? \nz.mem [1171] : 
                            (N316)? \nz.mem [1179] : 
                            (N318)? \nz.mem [1187] : 
                            (N320)? \nz.mem [1195] : 
                            (N322)? \nz.mem [1203] : 
                            (N324)? \nz.mem [1211] : 
                            (N326)? \nz.mem [1219] : 
                            (N328)? \nz.mem [1227] : 
                            (N330)? \nz.mem [1235] : 
                            (N332)? \nz.mem [1243] : 
                            (N334)? \nz.mem [1251] : 
                            (N336)? \nz.mem [1259] : 
                            (N338)? \nz.mem [1267] : 
                            (N340)? \nz.mem [1275] : 
                            (N342)? \nz.mem [1283] : 
                            (N344)? \nz.mem [1291] : 
                            (N346)? \nz.mem [1299] : 
                            (N348)? \nz.mem [1307] : 
                            (N350)? \nz.mem [1315] : 
                            (N352)? \nz.mem [1323] : 
                            (N354)? \nz.mem [1331] : 
                            (N356)? \nz.mem [1339] : 
                            (N358)? \nz.mem [1347] : 
                            (N360)? \nz.mem [1355] : 
                            (N362)? \nz.mem [1363] : 
                            (N364)? \nz.mem [1371] : 
                            (N366)? \nz.mem [1379] : 
                            (N368)? \nz.mem [1387] : 
                            (N370)? \nz.mem [1395] : 
                            (N372)? \nz.mem [1403] : 
                            (N374)? \nz.mem [1411] : 
                            (N376)? \nz.mem [1419] : 
                            (N378)? \nz.mem [1427] : 
                            (N380)? \nz.mem [1435] : 
                            (N382)? \nz.mem [1443] : 
                            (N384)? \nz.mem [1451] : 
                            (N386)? \nz.mem [1459] : 
                            (N388)? \nz.mem [1467] : 
                            (N390)? \nz.mem [1475] : 
                            (N392)? \nz.mem [1483] : 
                            (N394)? \nz.mem [1491] : 
                            (N396)? \nz.mem [1499] : 
                            (N398)? \nz.mem [1507] : 
                            (N400)? \nz.mem [1515] : 
                            (N402)? \nz.mem [1523] : 
                            (N404)? \nz.mem [1531] : 
                            (N406)? \nz.mem [1539] : 
                            (N408)? \nz.mem [1547] : 
                            (N410)? \nz.mem [1555] : 
                            (N412)? \nz.mem [1563] : 
                            (N414)? \nz.mem [1571] : 
                            (N416)? \nz.mem [1579] : 
                            (N418)? \nz.mem [1587] : 
                            (N420)? \nz.mem [1595] : 
                            (N422)? \nz.mem [1603] : 
                            (N424)? \nz.mem [1611] : 
                            (N426)? \nz.mem [1619] : 
                            (N428)? \nz.mem [1627] : 
                            (N430)? \nz.mem [1635] : 
                            (N432)? \nz.mem [1643] : 
                            (N434)? \nz.mem [1651] : 
                            (N436)? \nz.mem [1659] : 
                            (N438)? \nz.mem [1667] : 
                            (N440)? \nz.mem [1675] : 
                            (N442)? \nz.mem [1683] : 
                            (N444)? \nz.mem [1691] : 
                            (N446)? \nz.mem [1699] : 
                            (N448)? \nz.mem [1707] : 
                            (N450)? \nz.mem [1715] : 
                            (N452)? \nz.mem [1723] : 
                            (N454)? \nz.mem [1731] : 
                            (N456)? \nz.mem [1739] : 
                            (N458)? \nz.mem [1747] : 
                            (N460)? \nz.mem [1755] : 
                            (N462)? \nz.mem [1763] : 
                            (N464)? \nz.mem [1771] : 
                            (N466)? \nz.mem [1779] : 
                            (N468)? \nz.mem [1787] : 
                            (N470)? \nz.mem [1795] : 
                            (N472)? \nz.mem [1803] : 
                            (N474)? \nz.mem [1811] : 
                            (N476)? \nz.mem [1819] : 
                            (N478)? \nz.mem [1827] : 
                            (N480)? \nz.mem [1835] : 
                            (N482)? \nz.mem [1843] : 
                            (N484)? \nz.mem [1851] : 
                            (N486)? \nz.mem [1859] : 
                            (N488)? \nz.mem [1867] : 
                            (N490)? \nz.mem [1875] : 
                            (N492)? \nz.mem [1883] : 
                            (N494)? \nz.mem [1891] : 
                            (N496)? \nz.mem [1899] : 
                            (N498)? \nz.mem [1907] : 
                            (N500)? \nz.mem [1915] : 
                            (N502)? \nz.mem [1923] : 
                            (N504)? \nz.mem [1931] : 
                            (N506)? \nz.mem [1939] : 
                            (N508)? \nz.mem [1947] : 
                            (N510)? \nz.mem [1955] : 
                            (N512)? \nz.mem [1963] : 
                            (N514)? \nz.mem [1971] : 
                            (N516)? \nz.mem [1979] : 
                            (N518)? \nz.mem [1987] : 
                            (N520)? \nz.mem [1995] : 
                            (N522)? \nz.mem [2003] : 
                            (N524)? \nz.mem [2011] : 
                            (N526)? \nz.mem [2019] : 
                            (N528)? \nz.mem [2027] : 
                            (N530)? \nz.mem [2035] : 
                            (N532)? \nz.mem [2043] : 1'b0;
  assign \nz.data_out [2] = (N277)? \nz.mem [2] : 
                            (N279)? \nz.mem [10] : 
                            (N281)? \nz.mem [18] : 
                            (N283)? \nz.mem [26] : 
                            (N285)? \nz.mem [34] : 
                            (N287)? \nz.mem [42] : 
                            (N289)? \nz.mem [50] : 
                            (N291)? \nz.mem [58] : 
                            (N293)? \nz.mem [66] : 
                            (N295)? \nz.mem [74] : 
                            (N297)? \nz.mem [82] : 
                            (N299)? \nz.mem [90] : 
                            (N301)? \nz.mem [98] : 
                            (N303)? \nz.mem [106] : 
                            (N305)? \nz.mem [114] : 
                            (N307)? \nz.mem [122] : 
                            (N309)? \nz.mem [130] : 
                            (N311)? \nz.mem [138] : 
                            (N313)? \nz.mem [146] : 
                            (N315)? \nz.mem [154] : 
                            (N317)? \nz.mem [162] : 
                            (N319)? \nz.mem [170] : 
                            (N321)? \nz.mem [178] : 
                            (N323)? \nz.mem [186] : 
                            (N325)? \nz.mem [194] : 
                            (N327)? \nz.mem [202] : 
                            (N329)? \nz.mem [210] : 
                            (N331)? \nz.mem [218] : 
                            (N333)? \nz.mem [226] : 
                            (N335)? \nz.mem [234] : 
                            (N337)? \nz.mem [242] : 
                            (N339)? \nz.mem [250] : 
                            (N341)? \nz.mem [258] : 
                            (N343)? \nz.mem [266] : 
                            (N345)? \nz.mem [274] : 
                            (N347)? \nz.mem [282] : 
                            (N349)? \nz.mem [290] : 
                            (N351)? \nz.mem [298] : 
                            (N353)? \nz.mem [306] : 
                            (N355)? \nz.mem [314] : 
                            (N357)? \nz.mem [322] : 
                            (N359)? \nz.mem [330] : 
                            (N361)? \nz.mem [338] : 
                            (N363)? \nz.mem [346] : 
                            (N365)? \nz.mem [354] : 
                            (N367)? \nz.mem [362] : 
                            (N369)? \nz.mem [370] : 
                            (N371)? \nz.mem [378] : 
                            (N373)? \nz.mem [386] : 
                            (N375)? \nz.mem [394] : 
                            (N377)? \nz.mem [402] : 
                            (N379)? \nz.mem [410] : 
                            (N381)? \nz.mem [418] : 
                            (N383)? \nz.mem [426] : 
                            (N385)? \nz.mem [434] : 
                            (N387)? \nz.mem [442] : 
                            (N389)? \nz.mem [450] : 
                            (N391)? \nz.mem [458] : 
                            (N393)? \nz.mem [466] : 
                            (N395)? \nz.mem [474] : 
                            (N397)? \nz.mem [482] : 
                            (N399)? \nz.mem [490] : 
                            (N401)? \nz.mem [498] : 
                            (N403)? \nz.mem [506] : 
                            (N405)? \nz.mem [514] : 
                            (N407)? \nz.mem [522] : 
                            (N409)? \nz.mem [530] : 
                            (N411)? \nz.mem [538] : 
                            (N413)? \nz.mem [546] : 
                            (N415)? \nz.mem [554] : 
                            (N417)? \nz.mem [562] : 
                            (N419)? \nz.mem [570] : 
                            (N421)? \nz.mem [578] : 
                            (N423)? \nz.mem [586] : 
                            (N425)? \nz.mem [594] : 
                            (N427)? \nz.mem [602] : 
                            (N429)? \nz.mem [610] : 
                            (N431)? \nz.mem [618] : 
                            (N433)? \nz.mem [626] : 
                            (N435)? \nz.mem [634] : 
                            (N437)? \nz.mem [642] : 
                            (N439)? \nz.mem [650] : 
                            (N441)? \nz.mem [658] : 
                            (N443)? \nz.mem [666] : 
                            (N445)? \nz.mem [674] : 
                            (N447)? \nz.mem [682] : 
                            (N449)? \nz.mem [690] : 
                            (N451)? \nz.mem [698] : 
                            (N453)? \nz.mem [706] : 
                            (N455)? \nz.mem [714] : 
                            (N457)? \nz.mem [722] : 
                            (N459)? \nz.mem [730] : 
                            (N461)? \nz.mem [738] : 
                            (N463)? \nz.mem [746] : 
                            (N465)? \nz.mem [754] : 
                            (N467)? \nz.mem [762] : 
                            (N469)? \nz.mem [770] : 
                            (N471)? \nz.mem [778] : 
                            (N473)? \nz.mem [786] : 
                            (N475)? \nz.mem [794] : 
                            (N477)? \nz.mem [802] : 
                            (N479)? \nz.mem [810] : 
                            (N481)? \nz.mem [818] : 
                            (N483)? \nz.mem [826] : 
                            (N485)? \nz.mem [834] : 
                            (N487)? \nz.mem [842] : 
                            (N489)? \nz.mem [850] : 
                            (N491)? \nz.mem [858] : 
                            (N493)? \nz.mem [866] : 
                            (N495)? \nz.mem [874] : 
                            (N497)? \nz.mem [882] : 
                            (N499)? \nz.mem [890] : 
                            (N501)? \nz.mem [898] : 
                            (N503)? \nz.mem [906] : 
                            (N505)? \nz.mem [914] : 
                            (N507)? \nz.mem [922] : 
                            (N509)? \nz.mem [930] : 
                            (N511)? \nz.mem [938] : 
                            (N513)? \nz.mem [946] : 
                            (N515)? \nz.mem [954] : 
                            (N517)? \nz.mem [962] : 
                            (N519)? \nz.mem [970] : 
                            (N521)? \nz.mem [978] : 
                            (N523)? \nz.mem [986] : 
                            (N525)? \nz.mem [994] : 
                            (N527)? \nz.mem [1002] : 
                            (N529)? \nz.mem [1010] : 
                            (N531)? \nz.mem [1018] : 
                            (N278)? \nz.mem [1026] : 
                            (N280)? \nz.mem [1034] : 
                            (N282)? \nz.mem [1042] : 
                            (N284)? \nz.mem [1050] : 
                            (N286)? \nz.mem [1058] : 
                            (N288)? \nz.mem [1066] : 
                            (N290)? \nz.mem [1074] : 
                            (N292)? \nz.mem [1082] : 
                            (N294)? \nz.mem [1090] : 
                            (N296)? \nz.mem [1098] : 
                            (N298)? \nz.mem [1106] : 
                            (N300)? \nz.mem [1114] : 
                            (N302)? \nz.mem [1122] : 
                            (N304)? \nz.mem [1130] : 
                            (N306)? \nz.mem [1138] : 
                            (N308)? \nz.mem [1146] : 
                            (N310)? \nz.mem [1154] : 
                            (N312)? \nz.mem [1162] : 
                            (N314)? \nz.mem [1170] : 
                            (N316)? \nz.mem [1178] : 
                            (N318)? \nz.mem [1186] : 
                            (N320)? \nz.mem [1194] : 
                            (N322)? \nz.mem [1202] : 
                            (N324)? \nz.mem [1210] : 
                            (N326)? \nz.mem [1218] : 
                            (N328)? \nz.mem [1226] : 
                            (N330)? \nz.mem [1234] : 
                            (N332)? \nz.mem [1242] : 
                            (N334)? \nz.mem [1250] : 
                            (N336)? \nz.mem [1258] : 
                            (N338)? \nz.mem [1266] : 
                            (N340)? \nz.mem [1274] : 
                            (N342)? \nz.mem [1282] : 
                            (N344)? \nz.mem [1290] : 
                            (N346)? \nz.mem [1298] : 
                            (N348)? \nz.mem [1306] : 
                            (N350)? \nz.mem [1314] : 
                            (N352)? \nz.mem [1322] : 
                            (N354)? \nz.mem [1330] : 
                            (N356)? \nz.mem [1338] : 
                            (N358)? \nz.mem [1346] : 
                            (N360)? \nz.mem [1354] : 
                            (N362)? \nz.mem [1362] : 
                            (N364)? \nz.mem [1370] : 
                            (N366)? \nz.mem [1378] : 
                            (N368)? \nz.mem [1386] : 
                            (N370)? \nz.mem [1394] : 
                            (N372)? \nz.mem [1402] : 
                            (N374)? \nz.mem [1410] : 
                            (N376)? \nz.mem [1418] : 
                            (N378)? \nz.mem [1426] : 
                            (N380)? \nz.mem [1434] : 
                            (N382)? \nz.mem [1442] : 
                            (N384)? \nz.mem [1450] : 
                            (N386)? \nz.mem [1458] : 
                            (N388)? \nz.mem [1466] : 
                            (N390)? \nz.mem [1474] : 
                            (N392)? \nz.mem [1482] : 
                            (N394)? \nz.mem [1490] : 
                            (N396)? \nz.mem [1498] : 
                            (N398)? \nz.mem [1506] : 
                            (N400)? \nz.mem [1514] : 
                            (N402)? \nz.mem [1522] : 
                            (N404)? \nz.mem [1530] : 
                            (N406)? \nz.mem [1538] : 
                            (N408)? \nz.mem [1546] : 
                            (N410)? \nz.mem [1554] : 
                            (N412)? \nz.mem [1562] : 
                            (N414)? \nz.mem [1570] : 
                            (N416)? \nz.mem [1578] : 
                            (N418)? \nz.mem [1586] : 
                            (N420)? \nz.mem [1594] : 
                            (N422)? \nz.mem [1602] : 
                            (N424)? \nz.mem [1610] : 
                            (N426)? \nz.mem [1618] : 
                            (N428)? \nz.mem [1626] : 
                            (N430)? \nz.mem [1634] : 
                            (N432)? \nz.mem [1642] : 
                            (N434)? \nz.mem [1650] : 
                            (N436)? \nz.mem [1658] : 
                            (N438)? \nz.mem [1666] : 
                            (N440)? \nz.mem [1674] : 
                            (N442)? \nz.mem [1682] : 
                            (N444)? \nz.mem [1690] : 
                            (N446)? \nz.mem [1698] : 
                            (N448)? \nz.mem [1706] : 
                            (N450)? \nz.mem [1714] : 
                            (N452)? \nz.mem [1722] : 
                            (N454)? \nz.mem [1730] : 
                            (N456)? \nz.mem [1738] : 
                            (N458)? \nz.mem [1746] : 
                            (N460)? \nz.mem [1754] : 
                            (N462)? \nz.mem [1762] : 
                            (N464)? \nz.mem [1770] : 
                            (N466)? \nz.mem [1778] : 
                            (N468)? \nz.mem [1786] : 
                            (N470)? \nz.mem [1794] : 
                            (N472)? \nz.mem [1802] : 
                            (N474)? \nz.mem [1810] : 
                            (N476)? \nz.mem [1818] : 
                            (N478)? \nz.mem [1826] : 
                            (N480)? \nz.mem [1834] : 
                            (N482)? \nz.mem [1842] : 
                            (N484)? \nz.mem [1850] : 
                            (N486)? \nz.mem [1858] : 
                            (N488)? \nz.mem [1866] : 
                            (N490)? \nz.mem [1874] : 
                            (N492)? \nz.mem [1882] : 
                            (N494)? \nz.mem [1890] : 
                            (N496)? \nz.mem [1898] : 
                            (N498)? \nz.mem [1906] : 
                            (N500)? \nz.mem [1914] : 
                            (N502)? \nz.mem [1922] : 
                            (N504)? \nz.mem [1930] : 
                            (N506)? \nz.mem [1938] : 
                            (N508)? \nz.mem [1946] : 
                            (N510)? \nz.mem [1954] : 
                            (N512)? \nz.mem [1962] : 
                            (N514)? \nz.mem [1970] : 
                            (N516)? \nz.mem [1978] : 
                            (N518)? \nz.mem [1986] : 
                            (N520)? \nz.mem [1994] : 
                            (N522)? \nz.mem [2002] : 
                            (N524)? \nz.mem [2010] : 
                            (N526)? \nz.mem [2018] : 
                            (N528)? \nz.mem [2026] : 
                            (N530)? \nz.mem [2034] : 
                            (N532)? \nz.mem [2042] : 1'b0;
  assign \nz.data_out [1] = (N277)? \nz.mem [1] : 
                            (N279)? \nz.mem [9] : 
                            (N281)? \nz.mem [17] : 
                            (N283)? \nz.mem [25] : 
                            (N285)? \nz.mem [33] : 
                            (N287)? \nz.mem [41] : 
                            (N289)? \nz.mem [49] : 
                            (N291)? \nz.mem [57] : 
                            (N293)? \nz.mem [65] : 
                            (N295)? \nz.mem [73] : 
                            (N297)? \nz.mem [81] : 
                            (N299)? \nz.mem [89] : 
                            (N301)? \nz.mem [97] : 
                            (N303)? \nz.mem [105] : 
                            (N305)? \nz.mem [113] : 
                            (N307)? \nz.mem [121] : 
                            (N309)? \nz.mem [129] : 
                            (N311)? \nz.mem [137] : 
                            (N313)? \nz.mem [145] : 
                            (N315)? \nz.mem [153] : 
                            (N317)? \nz.mem [161] : 
                            (N319)? \nz.mem [169] : 
                            (N321)? \nz.mem [177] : 
                            (N323)? \nz.mem [185] : 
                            (N325)? \nz.mem [193] : 
                            (N327)? \nz.mem [201] : 
                            (N329)? \nz.mem [209] : 
                            (N331)? \nz.mem [217] : 
                            (N333)? \nz.mem [225] : 
                            (N335)? \nz.mem [233] : 
                            (N337)? \nz.mem [241] : 
                            (N339)? \nz.mem [249] : 
                            (N341)? \nz.mem [257] : 
                            (N343)? \nz.mem [265] : 
                            (N345)? \nz.mem [273] : 
                            (N347)? \nz.mem [281] : 
                            (N349)? \nz.mem [289] : 
                            (N351)? \nz.mem [297] : 
                            (N353)? \nz.mem [305] : 
                            (N355)? \nz.mem [313] : 
                            (N357)? \nz.mem [321] : 
                            (N359)? \nz.mem [329] : 
                            (N361)? \nz.mem [337] : 
                            (N363)? \nz.mem [345] : 
                            (N365)? \nz.mem [353] : 
                            (N367)? \nz.mem [361] : 
                            (N369)? \nz.mem [369] : 
                            (N371)? \nz.mem [377] : 
                            (N373)? \nz.mem [385] : 
                            (N375)? \nz.mem [393] : 
                            (N377)? \nz.mem [401] : 
                            (N379)? \nz.mem [409] : 
                            (N381)? \nz.mem [417] : 
                            (N383)? \nz.mem [425] : 
                            (N385)? \nz.mem [433] : 
                            (N387)? \nz.mem [441] : 
                            (N389)? \nz.mem [449] : 
                            (N391)? \nz.mem [457] : 
                            (N393)? \nz.mem [465] : 
                            (N395)? \nz.mem [473] : 
                            (N397)? \nz.mem [481] : 
                            (N399)? \nz.mem [489] : 
                            (N401)? \nz.mem [497] : 
                            (N403)? \nz.mem [505] : 
                            (N405)? \nz.mem [513] : 
                            (N407)? \nz.mem [521] : 
                            (N409)? \nz.mem [529] : 
                            (N411)? \nz.mem [537] : 
                            (N413)? \nz.mem [545] : 
                            (N415)? \nz.mem [553] : 
                            (N417)? \nz.mem [561] : 
                            (N419)? \nz.mem [569] : 
                            (N421)? \nz.mem [577] : 
                            (N423)? \nz.mem [585] : 
                            (N425)? \nz.mem [593] : 
                            (N427)? \nz.mem [601] : 
                            (N429)? \nz.mem [609] : 
                            (N431)? \nz.mem [617] : 
                            (N433)? \nz.mem [625] : 
                            (N435)? \nz.mem [633] : 
                            (N437)? \nz.mem [641] : 
                            (N439)? \nz.mem [649] : 
                            (N441)? \nz.mem [657] : 
                            (N443)? \nz.mem [665] : 
                            (N445)? \nz.mem [673] : 
                            (N447)? \nz.mem [681] : 
                            (N449)? \nz.mem [689] : 
                            (N451)? \nz.mem [697] : 
                            (N453)? \nz.mem [705] : 
                            (N455)? \nz.mem [713] : 
                            (N457)? \nz.mem [721] : 
                            (N459)? \nz.mem [729] : 
                            (N461)? \nz.mem [737] : 
                            (N463)? \nz.mem [745] : 
                            (N465)? \nz.mem [753] : 
                            (N467)? \nz.mem [761] : 
                            (N469)? \nz.mem [769] : 
                            (N471)? \nz.mem [777] : 
                            (N473)? \nz.mem [785] : 
                            (N475)? \nz.mem [793] : 
                            (N477)? \nz.mem [801] : 
                            (N479)? \nz.mem [809] : 
                            (N481)? \nz.mem [817] : 
                            (N483)? \nz.mem [825] : 
                            (N485)? \nz.mem [833] : 
                            (N487)? \nz.mem [841] : 
                            (N489)? \nz.mem [849] : 
                            (N491)? \nz.mem [857] : 
                            (N493)? \nz.mem [865] : 
                            (N495)? \nz.mem [873] : 
                            (N497)? \nz.mem [881] : 
                            (N499)? \nz.mem [889] : 
                            (N501)? \nz.mem [897] : 
                            (N503)? \nz.mem [905] : 
                            (N505)? \nz.mem [913] : 
                            (N507)? \nz.mem [921] : 
                            (N509)? \nz.mem [929] : 
                            (N511)? \nz.mem [937] : 
                            (N513)? \nz.mem [945] : 
                            (N515)? \nz.mem [953] : 
                            (N517)? \nz.mem [961] : 
                            (N519)? \nz.mem [969] : 
                            (N521)? \nz.mem [977] : 
                            (N523)? \nz.mem [985] : 
                            (N525)? \nz.mem [993] : 
                            (N527)? \nz.mem [1001] : 
                            (N529)? \nz.mem [1009] : 
                            (N531)? \nz.mem [1017] : 
                            (N278)? \nz.mem [1025] : 
                            (N280)? \nz.mem [1033] : 
                            (N282)? \nz.mem [1041] : 
                            (N284)? \nz.mem [1049] : 
                            (N286)? \nz.mem [1057] : 
                            (N288)? \nz.mem [1065] : 
                            (N290)? \nz.mem [1073] : 
                            (N292)? \nz.mem [1081] : 
                            (N294)? \nz.mem [1089] : 
                            (N296)? \nz.mem [1097] : 
                            (N298)? \nz.mem [1105] : 
                            (N300)? \nz.mem [1113] : 
                            (N302)? \nz.mem [1121] : 
                            (N304)? \nz.mem [1129] : 
                            (N306)? \nz.mem [1137] : 
                            (N308)? \nz.mem [1145] : 
                            (N310)? \nz.mem [1153] : 
                            (N312)? \nz.mem [1161] : 
                            (N314)? \nz.mem [1169] : 
                            (N316)? \nz.mem [1177] : 
                            (N318)? \nz.mem [1185] : 
                            (N320)? \nz.mem [1193] : 
                            (N322)? \nz.mem [1201] : 
                            (N324)? \nz.mem [1209] : 
                            (N326)? \nz.mem [1217] : 
                            (N328)? \nz.mem [1225] : 
                            (N330)? \nz.mem [1233] : 
                            (N332)? \nz.mem [1241] : 
                            (N334)? \nz.mem [1249] : 
                            (N336)? \nz.mem [1257] : 
                            (N338)? \nz.mem [1265] : 
                            (N340)? \nz.mem [1273] : 
                            (N342)? \nz.mem [1281] : 
                            (N344)? \nz.mem [1289] : 
                            (N346)? \nz.mem [1297] : 
                            (N348)? \nz.mem [1305] : 
                            (N350)? \nz.mem [1313] : 
                            (N352)? \nz.mem [1321] : 
                            (N354)? \nz.mem [1329] : 
                            (N356)? \nz.mem [1337] : 
                            (N358)? \nz.mem [1345] : 
                            (N360)? \nz.mem [1353] : 
                            (N362)? \nz.mem [1361] : 
                            (N364)? \nz.mem [1369] : 
                            (N366)? \nz.mem [1377] : 
                            (N368)? \nz.mem [1385] : 
                            (N370)? \nz.mem [1393] : 
                            (N372)? \nz.mem [1401] : 
                            (N374)? \nz.mem [1409] : 
                            (N376)? \nz.mem [1417] : 
                            (N378)? \nz.mem [1425] : 
                            (N380)? \nz.mem [1433] : 
                            (N382)? \nz.mem [1441] : 
                            (N384)? \nz.mem [1449] : 
                            (N386)? \nz.mem [1457] : 
                            (N388)? \nz.mem [1465] : 
                            (N390)? \nz.mem [1473] : 
                            (N392)? \nz.mem [1481] : 
                            (N394)? \nz.mem [1489] : 
                            (N396)? \nz.mem [1497] : 
                            (N398)? \nz.mem [1505] : 
                            (N400)? \nz.mem [1513] : 
                            (N402)? \nz.mem [1521] : 
                            (N404)? \nz.mem [1529] : 
                            (N406)? \nz.mem [1537] : 
                            (N408)? \nz.mem [1545] : 
                            (N410)? \nz.mem [1553] : 
                            (N412)? \nz.mem [1561] : 
                            (N414)? \nz.mem [1569] : 
                            (N416)? \nz.mem [1577] : 
                            (N418)? \nz.mem [1585] : 
                            (N420)? \nz.mem [1593] : 
                            (N422)? \nz.mem [1601] : 
                            (N424)? \nz.mem [1609] : 
                            (N426)? \nz.mem [1617] : 
                            (N428)? \nz.mem [1625] : 
                            (N430)? \nz.mem [1633] : 
                            (N432)? \nz.mem [1641] : 
                            (N434)? \nz.mem [1649] : 
                            (N436)? \nz.mem [1657] : 
                            (N438)? \nz.mem [1665] : 
                            (N440)? \nz.mem [1673] : 
                            (N442)? \nz.mem [1681] : 
                            (N444)? \nz.mem [1689] : 
                            (N446)? \nz.mem [1697] : 
                            (N448)? \nz.mem [1705] : 
                            (N450)? \nz.mem [1713] : 
                            (N452)? \nz.mem [1721] : 
                            (N454)? \nz.mem [1729] : 
                            (N456)? \nz.mem [1737] : 
                            (N458)? \nz.mem [1745] : 
                            (N460)? \nz.mem [1753] : 
                            (N462)? \nz.mem [1761] : 
                            (N464)? \nz.mem [1769] : 
                            (N466)? \nz.mem [1777] : 
                            (N468)? \nz.mem [1785] : 
                            (N470)? \nz.mem [1793] : 
                            (N472)? \nz.mem [1801] : 
                            (N474)? \nz.mem [1809] : 
                            (N476)? \nz.mem [1817] : 
                            (N478)? \nz.mem [1825] : 
                            (N480)? \nz.mem [1833] : 
                            (N482)? \nz.mem [1841] : 
                            (N484)? \nz.mem [1849] : 
                            (N486)? \nz.mem [1857] : 
                            (N488)? \nz.mem [1865] : 
                            (N490)? \nz.mem [1873] : 
                            (N492)? \nz.mem [1881] : 
                            (N494)? \nz.mem [1889] : 
                            (N496)? \nz.mem [1897] : 
                            (N498)? \nz.mem [1905] : 
                            (N500)? \nz.mem [1913] : 
                            (N502)? \nz.mem [1921] : 
                            (N504)? \nz.mem [1929] : 
                            (N506)? \nz.mem [1937] : 
                            (N508)? \nz.mem [1945] : 
                            (N510)? \nz.mem [1953] : 
                            (N512)? \nz.mem [1961] : 
                            (N514)? \nz.mem [1969] : 
                            (N516)? \nz.mem [1977] : 
                            (N518)? \nz.mem [1985] : 
                            (N520)? \nz.mem [1993] : 
                            (N522)? \nz.mem [2001] : 
                            (N524)? \nz.mem [2009] : 
                            (N526)? \nz.mem [2017] : 
                            (N528)? \nz.mem [2025] : 
                            (N530)? \nz.mem [2033] : 
                            (N532)? \nz.mem [2041] : 1'b0;
  assign \nz.data_out [0] = (N277)? \nz.mem [0] : 
                            (N279)? \nz.mem [8] : 
                            (N281)? \nz.mem [16] : 
                            (N283)? \nz.mem [24] : 
                            (N285)? \nz.mem [32] : 
                            (N287)? \nz.mem [40] : 
                            (N289)? \nz.mem [48] : 
                            (N291)? \nz.mem [56] : 
                            (N293)? \nz.mem [64] : 
                            (N295)? \nz.mem [72] : 
                            (N297)? \nz.mem [80] : 
                            (N299)? \nz.mem [88] : 
                            (N301)? \nz.mem [96] : 
                            (N303)? \nz.mem [104] : 
                            (N305)? \nz.mem [112] : 
                            (N307)? \nz.mem [120] : 
                            (N309)? \nz.mem [128] : 
                            (N311)? \nz.mem [136] : 
                            (N313)? \nz.mem [144] : 
                            (N315)? \nz.mem [152] : 
                            (N317)? \nz.mem [160] : 
                            (N319)? \nz.mem [168] : 
                            (N321)? \nz.mem [176] : 
                            (N323)? \nz.mem [184] : 
                            (N325)? \nz.mem [192] : 
                            (N327)? \nz.mem [200] : 
                            (N329)? \nz.mem [208] : 
                            (N331)? \nz.mem [216] : 
                            (N333)? \nz.mem [224] : 
                            (N335)? \nz.mem [232] : 
                            (N337)? \nz.mem [240] : 
                            (N339)? \nz.mem [248] : 
                            (N341)? \nz.mem [256] : 
                            (N343)? \nz.mem [264] : 
                            (N345)? \nz.mem [272] : 
                            (N347)? \nz.mem [280] : 
                            (N349)? \nz.mem [288] : 
                            (N351)? \nz.mem [296] : 
                            (N353)? \nz.mem [304] : 
                            (N355)? \nz.mem [312] : 
                            (N357)? \nz.mem [320] : 
                            (N359)? \nz.mem [328] : 
                            (N361)? \nz.mem [336] : 
                            (N363)? \nz.mem [344] : 
                            (N365)? \nz.mem [352] : 
                            (N367)? \nz.mem [360] : 
                            (N369)? \nz.mem [368] : 
                            (N371)? \nz.mem [376] : 
                            (N373)? \nz.mem [384] : 
                            (N375)? \nz.mem [392] : 
                            (N377)? \nz.mem [400] : 
                            (N379)? \nz.mem [408] : 
                            (N381)? \nz.mem [416] : 
                            (N383)? \nz.mem [424] : 
                            (N385)? \nz.mem [432] : 
                            (N387)? \nz.mem [440] : 
                            (N389)? \nz.mem [448] : 
                            (N391)? \nz.mem [456] : 
                            (N393)? \nz.mem [464] : 
                            (N395)? \nz.mem [472] : 
                            (N397)? \nz.mem [480] : 
                            (N399)? \nz.mem [488] : 
                            (N401)? \nz.mem [496] : 
                            (N403)? \nz.mem [504] : 
                            (N405)? \nz.mem [512] : 
                            (N407)? \nz.mem [520] : 
                            (N409)? \nz.mem [528] : 
                            (N411)? \nz.mem [536] : 
                            (N413)? \nz.mem [544] : 
                            (N415)? \nz.mem [552] : 
                            (N417)? \nz.mem [560] : 
                            (N419)? \nz.mem [568] : 
                            (N421)? \nz.mem [576] : 
                            (N423)? \nz.mem [584] : 
                            (N425)? \nz.mem [592] : 
                            (N427)? \nz.mem [600] : 
                            (N429)? \nz.mem [608] : 
                            (N431)? \nz.mem [616] : 
                            (N433)? \nz.mem [624] : 
                            (N435)? \nz.mem [632] : 
                            (N437)? \nz.mem [640] : 
                            (N439)? \nz.mem [648] : 
                            (N441)? \nz.mem [656] : 
                            (N443)? \nz.mem [664] : 
                            (N445)? \nz.mem [672] : 
                            (N447)? \nz.mem [680] : 
                            (N449)? \nz.mem [688] : 
                            (N451)? \nz.mem [696] : 
                            (N453)? \nz.mem [704] : 
                            (N455)? \nz.mem [712] : 
                            (N457)? \nz.mem [720] : 
                            (N459)? \nz.mem [728] : 
                            (N461)? \nz.mem [736] : 
                            (N463)? \nz.mem [744] : 
                            (N465)? \nz.mem [752] : 
                            (N467)? \nz.mem [760] : 
                            (N469)? \nz.mem [768] : 
                            (N471)? \nz.mem [776] : 
                            (N473)? \nz.mem [784] : 
                            (N475)? \nz.mem [792] : 
                            (N477)? \nz.mem [800] : 
                            (N479)? \nz.mem [808] : 
                            (N481)? \nz.mem [816] : 
                            (N483)? \nz.mem [824] : 
                            (N485)? \nz.mem [832] : 
                            (N487)? \nz.mem [840] : 
                            (N489)? \nz.mem [848] : 
                            (N491)? \nz.mem [856] : 
                            (N493)? \nz.mem [864] : 
                            (N495)? \nz.mem [872] : 
                            (N497)? \nz.mem [880] : 
                            (N499)? \nz.mem [888] : 
                            (N501)? \nz.mem [896] : 
                            (N503)? \nz.mem [904] : 
                            (N505)? \nz.mem [912] : 
                            (N507)? \nz.mem [920] : 
                            (N509)? \nz.mem [928] : 
                            (N511)? \nz.mem [936] : 
                            (N513)? \nz.mem [944] : 
                            (N515)? \nz.mem [952] : 
                            (N517)? \nz.mem [960] : 
                            (N519)? \nz.mem [968] : 
                            (N521)? \nz.mem [976] : 
                            (N523)? \nz.mem [984] : 
                            (N525)? \nz.mem [992] : 
                            (N527)? \nz.mem [1000] : 
                            (N529)? \nz.mem [1008] : 
                            (N531)? \nz.mem [1016] : 
                            (N278)? \nz.mem [1024] : 
                            (N280)? \nz.mem [1032] : 
                            (N282)? \nz.mem [1040] : 
                            (N284)? \nz.mem [1048] : 
                            (N286)? \nz.mem [1056] : 
                            (N288)? \nz.mem [1064] : 
                            (N290)? \nz.mem [1072] : 
                            (N292)? \nz.mem [1080] : 
                            (N294)? \nz.mem [1088] : 
                            (N296)? \nz.mem [1096] : 
                            (N298)? \nz.mem [1104] : 
                            (N300)? \nz.mem [1112] : 
                            (N302)? \nz.mem [1120] : 
                            (N304)? \nz.mem [1128] : 
                            (N306)? \nz.mem [1136] : 
                            (N308)? \nz.mem [1144] : 
                            (N310)? \nz.mem [1152] : 
                            (N312)? \nz.mem [1160] : 
                            (N314)? \nz.mem [1168] : 
                            (N316)? \nz.mem [1176] : 
                            (N318)? \nz.mem [1184] : 
                            (N320)? \nz.mem [1192] : 
                            (N322)? \nz.mem [1200] : 
                            (N324)? \nz.mem [1208] : 
                            (N326)? \nz.mem [1216] : 
                            (N328)? \nz.mem [1224] : 
                            (N330)? \nz.mem [1232] : 
                            (N332)? \nz.mem [1240] : 
                            (N334)? \nz.mem [1248] : 
                            (N336)? \nz.mem [1256] : 
                            (N338)? \nz.mem [1264] : 
                            (N340)? \nz.mem [1272] : 
                            (N342)? \nz.mem [1280] : 
                            (N344)? \nz.mem [1288] : 
                            (N346)? \nz.mem [1296] : 
                            (N348)? \nz.mem [1304] : 
                            (N350)? \nz.mem [1312] : 
                            (N352)? \nz.mem [1320] : 
                            (N354)? \nz.mem [1328] : 
                            (N356)? \nz.mem [1336] : 
                            (N358)? \nz.mem [1344] : 
                            (N360)? \nz.mem [1352] : 
                            (N362)? \nz.mem [1360] : 
                            (N364)? \nz.mem [1368] : 
                            (N366)? \nz.mem [1376] : 
                            (N368)? \nz.mem [1384] : 
                            (N370)? \nz.mem [1392] : 
                            (N372)? \nz.mem [1400] : 
                            (N374)? \nz.mem [1408] : 
                            (N376)? \nz.mem [1416] : 
                            (N378)? \nz.mem [1424] : 
                            (N380)? \nz.mem [1432] : 
                            (N382)? \nz.mem [1440] : 
                            (N384)? \nz.mem [1448] : 
                            (N386)? \nz.mem [1456] : 
                            (N388)? \nz.mem [1464] : 
                            (N390)? \nz.mem [1472] : 
                            (N392)? \nz.mem [1480] : 
                            (N394)? \nz.mem [1488] : 
                            (N396)? \nz.mem [1496] : 
                            (N398)? \nz.mem [1504] : 
                            (N400)? \nz.mem [1512] : 
                            (N402)? \nz.mem [1520] : 
                            (N404)? \nz.mem [1528] : 
                            (N406)? \nz.mem [1536] : 
                            (N408)? \nz.mem [1544] : 
                            (N410)? \nz.mem [1552] : 
                            (N412)? \nz.mem [1560] : 
                            (N414)? \nz.mem [1568] : 
                            (N416)? \nz.mem [1576] : 
                            (N418)? \nz.mem [1584] : 
                            (N420)? \nz.mem [1592] : 
                            (N422)? \nz.mem [1600] : 
                            (N424)? \nz.mem [1608] : 
                            (N426)? \nz.mem [1616] : 
                            (N428)? \nz.mem [1624] : 
                            (N430)? \nz.mem [1632] : 
                            (N432)? \nz.mem [1640] : 
                            (N434)? \nz.mem [1648] : 
                            (N436)? \nz.mem [1656] : 
                            (N438)? \nz.mem [1664] : 
                            (N440)? \nz.mem [1672] : 
                            (N442)? \nz.mem [1680] : 
                            (N444)? \nz.mem [1688] : 
                            (N446)? \nz.mem [1696] : 
                            (N448)? \nz.mem [1704] : 
                            (N450)? \nz.mem [1712] : 
                            (N452)? \nz.mem [1720] : 
                            (N454)? \nz.mem [1728] : 
                            (N456)? \nz.mem [1736] : 
                            (N458)? \nz.mem [1744] : 
                            (N460)? \nz.mem [1752] : 
                            (N462)? \nz.mem [1760] : 
                            (N464)? \nz.mem [1768] : 
                            (N466)? \nz.mem [1776] : 
                            (N468)? \nz.mem [1784] : 
                            (N470)? \nz.mem [1792] : 
                            (N472)? \nz.mem [1800] : 
                            (N474)? \nz.mem [1808] : 
                            (N476)? \nz.mem [1816] : 
                            (N478)? \nz.mem [1824] : 
                            (N480)? \nz.mem [1832] : 
                            (N482)? \nz.mem [1840] : 
                            (N484)? \nz.mem [1848] : 
                            (N486)? \nz.mem [1856] : 
                            (N488)? \nz.mem [1864] : 
                            (N490)? \nz.mem [1872] : 
                            (N492)? \nz.mem [1880] : 
                            (N494)? \nz.mem [1888] : 
                            (N496)? \nz.mem [1896] : 
                            (N498)? \nz.mem [1904] : 
                            (N500)? \nz.mem [1912] : 
                            (N502)? \nz.mem [1920] : 
                            (N504)? \nz.mem [1928] : 
                            (N506)? \nz.mem [1936] : 
                            (N508)? \nz.mem [1944] : 
                            (N510)? \nz.mem [1952] : 
                            (N512)? \nz.mem [1960] : 
                            (N514)? \nz.mem [1968] : 
                            (N516)? \nz.mem [1976] : 
                            (N518)? \nz.mem [1984] : 
                            (N520)? \nz.mem [1992] : 
                            (N522)? \nz.mem [2000] : 
                            (N524)? \nz.mem [2008] : 
                            (N526)? \nz.mem [2016] : 
                            (N528)? \nz.mem [2024] : 
                            (N530)? \nz.mem [2032] : 
                            (N532)? \nz.mem [2040] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p8
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N1047 = addr_i[6] & addr_i[7];
  assign N1048 = N0 & addr_i[7];
  assign N0 = ~addr_i[6];
  assign N1049 = addr_i[6] & N1;
  assign N1 = ~addr_i[7];
  assign N1050 = N2 & N3;
  assign N2 = ~addr_i[6];
  assign N3 = ~addr_i[7];
  assign N1051 = addr_i[4] & addr_i[5];
  assign N1052 = N4 & addr_i[5];
  assign N4 = ~addr_i[4];
  assign N1053 = addr_i[4] & N5;
  assign N5 = ~addr_i[5];
  assign N1054 = N6 & N7;
  assign N6 = ~addr_i[4];
  assign N7 = ~addr_i[5];
  assign N1055 = N1047 & N1051;
  assign N1056 = N1047 & N1052;
  assign N1057 = N1047 & N1053;
  assign N1058 = N1047 & N1054;
  assign N1059 = N1048 & N1051;
  assign N1060 = N1048 & N1052;
  assign N1061 = N1048 & N1053;
  assign N1062 = N1048 & N1054;
  assign N1063 = N1049 & N1051;
  assign N1064 = N1049 & N1052;
  assign N1065 = N1049 & N1053;
  assign N1066 = N1049 & N1054;
  assign N1067 = N1050 & N1051;
  assign N1068 = N1050 & N1052;
  assign N1069 = N1050 & N1053;
  assign N1070 = N1050 & N1054;
  assign N1071 = addr_i[2] & addr_i[3];
  assign N1072 = N8 & addr_i[3];
  assign N8 = ~addr_i[2];
  assign N1073 = addr_i[2] & N9;
  assign N9 = ~addr_i[3];
  assign N1074 = N10 & N11;
  assign N10 = ~addr_i[2];
  assign N11 = ~addr_i[3];
  assign N1075 = addr_i[0] & addr_i[1];
  assign N1076 = N12 & addr_i[1];
  assign N12 = ~addr_i[0];
  assign N1077 = addr_i[0] & N13;
  assign N13 = ~addr_i[1];
  assign N1078 = N14 & N15;
  assign N14 = ~addr_i[0];
  assign N15 = ~addr_i[1];
  assign N1079 = N1071 & N1075;
  assign N1080 = N1071 & N1076;
  assign N1081 = N1071 & N1077;
  assign N1082 = N1071 & N1078;
  assign N1083 = N1072 & N1075;
  assign N1084 = N1072 & N1076;
  assign N1085 = N1072 & N1077;
  assign N1086 = N1072 & N1078;
  assign N1087 = N1073 & N1075;
  assign N1088 = N1073 & N1076;
  assign N1089 = N1073 & N1077;
  assign N1090 = N1073 & N1078;
  assign N1091 = N1074 & N1075;
  assign N1092 = N1074 & N1076;
  assign N1093 = N1074 & N1077;
  assign N1094 = N1074 & N1078;
  assign N790 = N1055 & N1079;
  assign N789 = N1055 & N1080;
  assign N788 = N1055 & N1081;
  assign N787 = N1055 & N1082;
  assign N786 = N1055 & N1083;
  assign N785 = N1055 & N1084;
  assign N784 = N1055 & N1085;
  assign N783 = N1055 & N1086;
  assign N782 = N1055 & N1087;
  assign N781 = N1055 & N1088;
  assign N780 = N1055 & N1089;
  assign N779 = N1055 & N1090;
  assign N778 = N1055 & N1091;
  assign N777 = N1055 & N1092;
  assign N776 = N1055 & N1093;
  assign N775 = N1055 & N1094;
  assign N774 = N1056 & N1079;
  assign N773 = N1056 & N1080;
  assign N772 = N1056 & N1081;
  assign N771 = N1056 & N1082;
  assign N770 = N1056 & N1083;
  assign N769 = N1056 & N1084;
  assign N768 = N1056 & N1085;
  assign N767 = N1056 & N1086;
  assign N766 = N1056 & N1087;
  assign N765 = N1056 & N1088;
  assign N764 = N1056 & N1089;
  assign N763 = N1056 & N1090;
  assign N762 = N1056 & N1091;
  assign N761 = N1056 & N1092;
  assign N760 = N1056 & N1093;
  assign N759 = N1056 & N1094;
  assign N758 = N1057 & N1079;
  assign N757 = N1057 & N1080;
  assign N756 = N1057 & N1081;
  assign N755 = N1057 & N1082;
  assign N754 = N1057 & N1083;
  assign N753 = N1057 & N1084;
  assign N752 = N1057 & N1085;
  assign N751 = N1057 & N1086;
  assign N750 = N1057 & N1087;
  assign N749 = N1057 & N1088;
  assign N748 = N1057 & N1089;
  assign N747 = N1057 & N1090;
  assign N746 = N1057 & N1091;
  assign N745 = N1057 & N1092;
  assign N744 = N1057 & N1093;
  assign N743 = N1057 & N1094;
  assign N742 = N1058 & N1079;
  assign N741 = N1058 & N1080;
  assign N740 = N1058 & N1081;
  assign N739 = N1058 & N1082;
  assign N738 = N1058 & N1083;
  assign N737 = N1058 & N1084;
  assign N736 = N1058 & N1085;
  assign N735 = N1058 & N1086;
  assign N734 = N1058 & N1087;
  assign N733 = N1058 & N1088;
  assign N732 = N1058 & N1089;
  assign N731 = N1058 & N1090;
  assign N730 = N1058 & N1091;
  assign N729 = N1058 & N1092;
  assign N728 = N1058 & N1093;
  assign N727 = N1058 & N1094;
  assign N726 = N1059 & N1079;
  assign N725 = N1059 & N1080;
  assign N724 = N1059 & N1081;
  assign N723 = N1059 & N1082;
  assign N722 = N1059 & N1083;
  assign N721 = N1059 & N1084;
  assign N720 = N1059 & N1085;
  assign N719 = N1059 & N1086;
  assign N718 = N1059 & N1087;
  assign N717 = N1059 & N1088;
  assign N716 = N1059 & N1089;
  assign N715 = N1059 & N1090;
  assign N714 = N1059 & N1091;
  assign N713 = N1059 & N1092;
  assign N712 = N1059 & N1093;
  assign N711 = N1059 & N1094;
  assign N710 = N1060 & N1079;
  assign N709 = N1060 & N1080;
  assign N708 = N1060 & N1081;
  assign N707 = N1060 & N1082;
  assign N706 = N1060 & N1083;
  assign N705 = N1060 & N1084;
  assign N704 = N1060 & N1085;
  assign N703 = N1060 & N1086;
  assign N702 = N1060 & N1087;
  assign N701 = N1060 & N1088;
  assign N700 = N1060 & N1089;
  assign N699 = N1060 & N1090;
  assign N698 = N1060 & N1091;
  assign N697 = N1060 & N1092;
  assign N696 = N1060 & N1093;
  assign N695 = N1060 & N1094;
  assign N694 = N1061 & N1079;
  assign N693 = N1061 & N1080;
  assign N692 = N1061 & N1081;
  assign N691 = N1061 & N1082;
  assign N690 = N1061 & N1083;
  assign N689 = N1061 & N1084;
  assign N688 = N1061 & N1085;
  assign N687 = N1061 & N1086;
  assign N686 = N1061 & N1087;
  assign N685 = N1061 & N1088;
  assign N684 = N1061 & N1089;
  assign N683 = N1061 & N1090;
  assign N682 = N1061 & N1091;
  assign N681 = N1061 & N1092;
  assign N680 = N1061 & N1093;
  assign N679 = N1061 & N1094;
  assign N678 = N1062 & N1079;
  assign N677 = N1062 & N1080;
  assign N676 = N1062 & N1081;
  assign N675 = N1062 & N1082;
  assign N674 = N1062 & N1083;
  assign N673 = N1062 & N1084;
  assign N672 = N1062 & N1085;
  assign N671 = N1062 & N1086;
  assign N670 = N1062 & N1087;
  assign N669 = N1062 & N1088;
  assign N668 = N1062 & N1089;
  assign N667 = N1062 & N1090;
  assign N666 = N1062 & N1091;
  assign N665 = N1062 & N1092;
  assign N664 = N1062 & N1093;
  assign N663 = N1062 & N1094;
  assign N662 = N1063 & N1079;
  assign N661 = N1063 & N1080;
  assign N660 = N1063 & N1081;
  assign N659 = N1063 & N1082;
  assign N658 = N1063 & N1083;
  assign N657 = N1063 & N1084;
  assign N656 = N1063 & N1085;
  assign N655 = N1063 & N1086;
  assign N654 = N1063 & N1087;
  assign N653 = N1063 & N1088;
  assign N652 = N1063 & N1089;
  assign N651 = N1063 & N1090;
  assign N650 = N1063 & N1091;
  assign N649 = N1063 & N1092;
  assign N648 = N1063 & N1093;
  assign N647 = N1063 & N1094;
  assign N646 = N1064 & N1079;
  assign N645 = N1064 & N1080;
  assign N644 = N1064 & N1081;
  assign N643 = N1064 & N1082;
  assign N642 = N1064 & N1083;
  assign N641 = N1064 & N1084;
  assign N640 = N1064 & N1085;
  assign N639 = N1064 & N1086;
  assign N638 = N1064 & N1087;
  assign N637 = N1064 & N1088;
  assign N636 = N1064 & N1089;
  assign N635 = N1064 & N1090;
  assign N634 = N1064 & N1091;
  assign N633 = N1064 & N1092;
  assign N632 = N1064 & N1093;
  assign N631 = N1064 & N1094;
  assign N630 = N1065 & N1079;
  assign N629 = N1065 & N1080;
  assign N628 = N1065 & N1081;
  assign N627 = N1065 & N1082;
  assign N626 = N1065 & N1083;
  assign N625 = N1065 & N1084;
  assign N624 = N1065 & N1085;
  assign N623 = N1065 & N1086;
  assign N622 = N1065 & N1087;
  assign N621 = N1065 & N1088;
  assign N620 = N1065 & N1089;
  assign N619 = N1065 & N1090;
  assign N618 = N1065 & N1091;
  assign N617 = N1065 & N1092;
  assign N616 = N1065 & N1093;
  assign N615 = N1065 & N1094;
  assign N614 = N1066 & N1079;
  assign N613 = N1066 & N1080;
  assign N612 = N1066 & N1081;
  assign N611 = N1066 & N1082;
  assign N610 = N1066 & N1083;
  assign N609 = N1066 & N1084;
  assign N608 = N1066 & N1085;
  assign N607 = N1066 & N1086;
  assign N606 = N1066 & N1087;
  assign N605 = N1066 & N1088;
  assign N604 = N1066 & N1089;
  assign N603 = N1066 & N1090;
  assign N602 = N1066 & N1091;
  assign N601 = N1066 & N1092;
  assign N600 = N1066 & N1093;
  assign N599 = N1066 & N1094;
  assign N598 = N1067 & N1079;
  assign N597 = N1067 & N1080;
  assign N596 = N1067 & N1081;
  assign N595 = N1067 & N1082;
  assign N594 = N1067 & N1083;
  assign N593 = N1067 & N1084;
  assign N592 = N1067 & N1085;
  assign N591 = N1067 & N1086;
  assign N590 = N1067 & N1087;
  assign N589 = N1067 & N1088;
  assign N588 = N1067 & N1089;
  assign N587 = N1067 & N1090;
  assign N586 = N1067 & N1091;
  assign N585 = N1067 & N1092;
  assign N584 = N1067 & N1093;
  assign N583 = N1067 & N1094;
  assign N582 = N1068 & N1079;
  assign N581 = N1068 & N1080;
  assign N580 = N1068 & N1081;
  assign N579 = N1068 & N1082;
  assign N578 = N1068 & N1083;
  assign N577 = N1068 & N1084;
  assign N576 = N1068 & N1085;
  assign N575 = N1068 & N1086;
  assign N574 = N1068 & N1087;
  assign N573 = N1068 & N1088;
  assign N572 = N1068 & N1089;
  assign N571 = N1068 & N1090;
  assign N570 = N1068 & N1091;
  assign N569 = N1068 & N1092;
  assign N568 = N1068 & N1093;
  assign N567 = N1068 & N1094;
  assign N566 = N1069 & N1079;
  assign N565 = N1069 & N1080;
  assign N564 = N1069 & N1081;
  assign N563 = N1069 & N1082;
  assign N562 = N1069 & N1083;
  assign N561 = N1069 & N1084;
  assign N560 = N1069 & N1085;
  assign N559 = N1069 & N1086;
  assign N558 = N1069 & N1087;
  assign N557 = N1069 & N1088;
  assign N556 = N1069 & N1089;
  assign N555 = N1069 & N1090;
  assign N554 = N1069 & N1091;
  assign N553 = N1069 & N1092;
  assign N552 = N1069 & N1093;
  assign N551 = N1069 & N1094;
  assign N550 = N1070 & N1079;
  assign N549 = N1070 & N1080;
  assign N548 = N1070 & N1081;
  assign N547 = N1070 & N1082;
  assign N546 = N1070 & N1083;
  assign N545 = N1070 & N1084;
  assign N544 = N1070 & N1085;
  assign N543 = N1070 & N1086;
  assign N542 = N1070 & N1087;
  assign N541 = N1070 & N1088;
  assign N540 = N1070 & N1089;
  assign N539 = N1070 & N1090;
  assign N538 = N1070 & N1091;
  assign N537 = N1070 & N1092;
  assign N536 = N1070 & N1093;
  assign N535 = N1070 & N1094;
  assign { N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791 } = (N16)? { N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N533;
  assign \nz.read_en  = v_i & N1095;
  assign N1095 = ~w_i;
  assign N17 = ~\nz.addr_r [0];
  assign N18 = ~\nz.addr_r [1];
  assign N19 = N17 & N18;
  assign N20 = N17 & \nz.addr_r [1];
  assign N21 = \nz.addr_r [0] & N18;
  assign N22 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N23 = ~\nz.addr_r [2];
  assign N24 = N19 & N23;
  assign N25 = N19 & \nz.addr_r [2];
  assign N26 = N21 & N23;
  assign N27 = N21 & \nz.addr_r [2];
  assign N28 = N20 & N23;
  assign N29 = N20 & \nz.addr_r [2];
  assign N30 = N22 & N23;
  assign N31 = N22 & \nz.addr_r [2];
  assign N32 = ~\nz.addr_r [3];
  assign N33 = N24 & N32;
  assign N34 = N24 & \nz.addr_r [3];
  assign N35 = N26 & N32;
  assign N36 = N26 & \nz.addr_r [3];
  assign N37 = N28 & N32;
  assign N38 = N28 & \nz.addr_r [3];
  assign N39 = N30 & N32;
  assign N40 = N30 & \nz.addr_r [3];
  assign N41 = N25 & N32;
  assign N42 = N25 & \nz.addr_r [3];
  assign N43 = N27 & N32;
  assign N44 = N27 & \nz.addr_r [3];
  assign N45 = N29 & N32;
  assign N46 = N29 & \nz.addr_r [3];
  assign N47 = N31 & N32;
  assign N48 = N31 & \nz.addr_r [3];
  assign N49 = ~\nz.addr_r [4];
  assign N50 = N33 & N49;
  assign N51 = N33 & \nz.addr_r [4];
  assign N52 = N35 & N49;
  assign N53 = N35 & \nz.addr_r [4];
  assign N54 = N37 & N49;
  assign N55 = N37 & \nz.addr_r [4];
  assign N56 = N39 & N49;
  assign N57 = N39 & \nz.addr_r [4];
  assign N58 = N41 & N49;
  assign N59 = N41 & \nz.addr_r [4];
  assign N60 = N43 & N49;
  assign N61 = N43 & \nz.addr_r [4];
  assign N62 = N45 & N49;
  assign N63 = N45 & \nz.addr_r [4];
  assign N64 = N47 & N49;
  assign N65 = N47 & \nz.addr_r [4];
  assign N66 = N34 & N49;
  assign N67 = N34 & \nz.addr_r [4];
  assign N68 = N36 & N49;
  assign N69 = N36 & \nz.addr_r [4];
  assign N70 = N38 & N49;
  assign N71 = N38 & \nz.addr_r [4];
  assign N72 = N40 & N49;
  assign N73 = N40 & \nz.addr_r [4];
  assign N74 = N42 & N49;
  assign N75 = N42 & \nz.addr_r [4];
  assign N76 = N44 & N49;
  assign N77 = N44 & \nz.addr_r [4];
  assign N78 = N46 & N49;
  assign N79 = N46 & \nz.addr_r [4];
  assign N80 = N48 & N49;
  assign N81 = N48 & \nz.addr_r [4];
  assign N82 = ~\nz.addr_r [5];
  assign N83 = N50 & N82;
  assign N84 = N50 & \nz.addr_r [5];
  assign N85 = N52 & N82;
  assign N86 = N52 & \nz.addr_r [5];
  assign N87 = N54 & N82;
  assign N88 = N54 & \nz.addr_r [5];
  assign N89 = N56 & N82;
  assign N90 = N56 & \nz.addr_r [5];
  assign N91 = N58 & N82;
  assign N92 = N58 & \nz.addr_r [5];
  assign N93 = N60 & N82;
  assign N94 = N60 & \nz.addr_r [5];
  assign N95 = N62 & N82;
  assign N96 = N62 & \nz.addr_r [5];
  assign N97 = N64 & N82;
  assign N98 = N64 & \nz.addr_r [5];
  assign N99 = N66 & N82;
  assign N100 = N66 & \nz.addr_r [5];
  assign N101 = N68 & N82;
  assign N102 = N68 & \nz.addr_r [5];
  assign N103 = N70 & N82;
  assign N104 = N70 & \nz.addr_r [5];
  assign N105 = N72 & N82;
  assign N106 = N72 & \nz.addr_r [5];
  assign N107 = N74 & N82;
  assign N108 = N74 & \nz.addr_r [5];
  assign N109 = N76 & N82;
  assign N110 = N76 & \nz.addr_r [5];
  assign N111 = N78 & N82;
  assign N112 = N78 & \nz.addr_r [5];
  assign N113 = N80 & N82;
  assign N114 = N80 & \nz.addr_r [5];
  assign N115 = N51 & N82;
  assign N116 = N51 & \nz.addr_r [5];
  assign N117 = N53 & N82;
  assign N118 = N53 & \nz.addr_r [5];
  assign N119 = N55 & N82;
  assign N120 = N55 & \nz.addr_r [5];
  assign N121 = N57 & N82;
  assign N122 = N57 & \nz.addr_r [5];
  assign N123 = N59 & N82;
  assign N124 = N59 & \nz.addr_r [5];
  assign N125 = N61 & N82;
  assign N126 = N61 & \nz.addr_r [5];
  assign N127 = N63 & N82;
  assign N128 = N63 & \nz.addr_r [5];
  assign N129 = N65 & N82;
  assign N130 = N65 & \nz.addr_r [5];
  assign N131 = N67 & N82;
  assign N132 = N67 & \nz.addr_r [5];
  assign N133 = N69 & N82;
  assign N134 = N69 & \nz.addr_r [5];
  assign N135 = N71 & N82;
  assign N136 = N71 & \nz.addr_r [5];
  assign N137 = N73 & N82;
  assign N138 = N73 & \nz.addr_r [5];
  assign N139 = N75 & N82;
  assign N140 = N75 & \nz.addr_r [5];
  assign N141 = N77 & N82;
  assign N142 = N77 & \nz.addr_r [5];
  assign N143 = N79 & N82;
  assign N144 = N79 & \nz.addr_r [5];
  assign N145 = N81 & N82;
  assign N146 = N81 & \nz.addr_r [5];
  assign N147 = ~\nz.addr_r [6];
  assign N148 = N83 & N147;
  assign N149 = N83 & \nz.addr_r [6];
  assign N150 = N85 & N147;
  assign N151 = N85 & \nz.addr_r [6];
  assign N152 = N87 & N147;
  assign N153 = N87 & \nz.addr_r [6];
  assign N154 = N89 & N147;
  assign N155 = N89 & \nz.addr_r [6];
  assign N156 = N91 & N147;
  assign N157 = N91 & \nz.addr_r [6];
  assign N158 = N93 & N147;
  assign N159 = N93 & \nz.addr_r [6];
  assign N160 = N95 & N147;
  assign N161 = N95 & \nz.addr_r [6];
  assign N162 = N97 & N147;
  assign N163 = N97 & \nz.addr_r [6];
  assign N164 = N99 & N147;
  assign N165 = N99 & \nz.addr_r [6];
  assign N166 = N101 & N147;
  assign N167 = N101 & \nz.addr_r [6];
  assign N168 = N103 & N147;
  assign N169 = N103 & \nz.addr_r [6];
  assign N170 = N105 & N147;
  assign N171 = N105 & \nz.addr_r [6];
  assign N172 = N107 & N147;
  assign N173 = N107 & \nz.addr_r [6];
  assign N174 = N109 & N147;
  assign N175 = N109 & \nz.addr_r [6];
  assign N176 = N111 & N147;
  assign N177 = N111 & \nz.addr_r [6];
  assign N178 = N113 & N147;
  assign N179 = N113 & \nz.addr_r [6];
  assign N180 = N115 & N147;
  assign N181 = N115 & \nz.addr_r [6];
  assign N182 = N117 & N147;
  assign N183 = N117 & \nz.addr_r [6];
  assign N184 = N119 & N147;
  assign N185 = N119 & \nz.addr_r [6];
  assign N186 = N121 & N147;
  assign N187 = N121 & \nz.addr_r [6];
  assign N188 = N123 & N147;
  assign N189 = N123 & \nz.addr_r [6];
  assign N190 = N125 & N147;
  assign N191 = N125 & \nz.addr_r [6];
  assign N192 = N127 & N147;
  assign N193 = N127 & \nz.addr_r [6];
  assign N194 = N129 & N147;
  assign N195 = N129 & \nz.addr_r [6];
  assign N196 = N131 & N147;
  assign N197 = N131 & \nz.addr_r [6];
  assign N198 = N133 & N147;
  assign N199 = N133 & \nz.addr_r [6];
  assign N200 = N135 & N147;
  assign N201 = N135 & \nz.addr_r [6];
  assign N202 = N137 & N147;
  assign N203 = N137 & \nz.addr_r [6];
  assign N204 = N139 & N147;
  assign N205 = N139 & \nz.addr_r [6];
  assign N206 = N141 & N147;
  assign N207 = N141 & \nz.addr_r [6];
  assign N208 = N143 & N147;
  assign N209 = N143 & \nz.addr_r [6];
  assign N210 = N145 & N147;
  assign N211 = N145 & \nz.addr_r [6];
  assign N212 = N84 & N147;
  assign N213 = N84 & \nz.addr_r [6];
  assign N214 = N86 & N147;
  assign N215 = N86 & \nz.addr_r [6];
  assign N216 = N88 & N147;
  assign N217 = N88 & \nz.addr_r [6];
  assign N218 = N90 & N147;
  assign N219 = N90 & \nz.addr_r [6];
  assign N220 = N92 & N147;
  assign N221 = N92 & \nz.addr_r [6];
  assign N222 = N94 & N147;
  assign N223 = N94 & \nz.addr_r [6];
  assign N224 = N96 & N147;
  assign N225 = N96 & \nz.addr_r [6];
  assign N226 = N98 & N147;
  assign N227 = N98 & \nz.addr_r [6];
  assign N228 = N100 & N147;
  assign N229 = N100 & \nz.addr_r [6];
  assign N230 = N102 & N147;
  assign N231 = N102 & \nz.addr_r [6];
  assign N232 = N104 & N147;
  assign N233 = N104 & \nz.addr_r [6];
  assign N234 = N106 & N147;
  assign N235 = N106 & \nz.addr_r [6];
  assign N236 = N108 & N147;
  assign N237 = N108 & \nz.addr_r [6];
  assign N238 = N110 & N147;
  assign N239 = N110 & \nz.addr_r [6];
  assign N240 = N112 & N147;
  assign N241 = N112 & \nz.addr_r [6];
  assign N242 = N114 & N147;
  assign N243 = N114 & \nz.addr_r [6];
  assign N244 = N116 & N147;
  assign N245 = N116 & \nz.addr_r [6];
  assign N246 = N118 & N147;
  assign N247 = N118 & \nz.addr_r [6];
  assign N248 = N120 & N147;
  assign N249 = N120 & \nz.addr_r [6];
  assign N250 = N122 & N147;
  assign N251 = N122 & \nz.addr_r [6];
  assign N252 = N124 & N147;
  assign N253 = N124 & \nz.addr_r [6];
  assign N254 = N126 & N147;
  assign N255 = N126 & \nz.addr_r [6];
  assign N256 = N128 & N147;
  assign N257 = N128 & \nz.addr_r [6];
  assign N258 = N130 & N147;
  assign N259 = N130 & \nz.addr_r [6];
  assign N260 = N132 & N147;
  assign N261 = N132 & \nz.addr_r [6];
  assign N262 = N134 & N147;
  assign N263 = N134 & \nz.addr_r [6];
  assign N264 = N136 & N147;
  assign N265 = N136 & \nz.addr_r [6];
  assign N266 = N138 & N147;
  assign N267 = N138 & \nz.addr_r [6];
  assign N268 = N140 & N147;
  assign N269 = N140 & \nz.addr_r [6];
  assign N270 = N142 & N147;
  assign N271 = N142 & \nz.addr_r [6];
  assign N272 = N144 & N147;
  assign N273 = N144 & \nz.addr_r [6];
  assign N274 = N146 & N147;
  assign N275 = N146 & \nz.addr_r [6];
  assign N276 = ~\nz.addr_r [7];
  assign N277 = N148 & N276;
  assign N278 = N148 & \nz.addr_r [7];
  assign N279 = N150 & N276;
  assign N280 = N150 & \nz.addr_r [7];
  assign N281 = N152 & N276;
  assign N282 = N152 & \nz.addr_r [7];
  assign N283 = N154 & N276;
  assign N284 = N154 & \nz.addr_r [7];
  assign N285 = N156 & N276;
  assign N286 = N156 & \nz.addr_r [7];
  assign N287 = N158 & N276;
  assign N288 = N158 & \nz.addr_r [7];
  assign N289 = N160 & N276;
  assign N290 = N160 & \nz.addr_r [7];
  assign N291 = N162 & N276;
  assign N292 = N162 & \nz.addr_r [7];
  assign N293 = N164 & N276;
  assign N294 = N164 & \nz.addr_r [7];
  assign N295 = N166 & N276;
  assign N296 = N166 & \nz.addr_r [7];
  assign N297 = N168 & N276;
  assign N298 = N168 & \nz.addr_r [7];
  assign N299 = N170 & N276;
  assign N300 = N170 & \nz.addr_r [7];
  assign N301 = N172 & N276;
  assign N302 = N172 & \nz.addr_r [7];
  assign N303 = N174 & N276;
  assign N304 = N174 & \nz.addr_r [7];
  assign N305 = N176 & N276;
  assign N306 = N176 & \nz.addr_r [7];
  assign N307 = N178 & N276;
  assign N308 = N178 & \nz.addr_r [7];
  assign N309 = N180 & N276;
  assign N310 = N180 & \nz.addr_r [7];
  assign N311 = N182 & N276;
  assign N312 = N182 & \nz.addr_r [7];
  assign N313 = N184 & N276;
  assign N314 = N184 & \nz.addr_r [7];
  assign N315 = N186 & N276;
  assign N316 = N186 & \nz.addr_r [7];
  assign N317 = N188 & N276;
  assign N318 = N188 & \nz.addr_r [7];
  assign N319 = N190 & N276;
  assign N320 = N190 & \nz.addr_r [7];
  assign N321 = N192 & N276;
  assign N322 = N192 & \nz.addr_r [7];
  assign N323 = N194 & N276;
  assign N324 = N194 & \nz.addr_r [7];
  assign N325 = N196 & N276;
  assign N326 = N196 & \nz.addr_r [7];
  assign N327 = N198 & N276;
  assign N328 = N198 & \nz.addr_r [7];
  assign N329 = N200 & N276;
  assign N330 = N200 & \nz.addr_r [7];
  assign N331 = N202 & N276;
  assign N332 = N202 & \nz.addr_r [7];
  assign N333 = N204 & N276;
  assign N334 = N204 & \nz.addr_r [7];
  assign N335 = N206 & N276;
  assign N336 = N206 & \nz.addr_r [7];
  assign N337 = N208 & N276;
  assign N338 = N208 & \nz.addr_r [7];
  assign N339 = N210 & N276;
  assign N340 = N210 & \nz.addr_r [7];
  assign N341 = N212 & N276;
  assign N342 = N212 & \nz.addr_r [7];
  assign N343 = N214 & N276;
  assign N344 = N214 & \nz.addr_r [7];
  assign N345 = N216 & N276;
  assign N346 = N216 & \nz.addr_r [7];
  assign N347 = N218 & N276;
  assign N348 = N218 & \nz.addr_r [7];
  assign N349 = N220 & N276;
  assign N350 = N220 & \nz.addr_r [7];
  assign N351 = N222 & N276;
  assign N352 = N222 & \nz.addr_r [7];
  assign N353 = N224 & N276;
  assign N354 = N224 & \nz.addr_r [7];
  assign N355 = N226 & N276;
  assign N356 = N226 & \nz.addr_r [7];
  assign N357 = N228 & N276;
  assign N358 = N228 & \nz.addr_r [7];
  assign N359 = N230 & N276;
  assign N360 = N230 & \nz.addr_r [7];
  assign N361 = N232 & N276;
  assign N362 = N232 & \nz.addr_r [7];
  assign N363 = N234 & N276;
  assign N364 = N234 & \nz.addr_r [7];
  assign N365 = N236 & N276;
  assign N366 = N236 & \nz.addr_r [7];
  assign N367 = N238 & N276;
  assign N368 = N238 & \nz.addr_r [7];
  assign N369 = N240 & N276;
  assign N370 = N240 & \nz.addr_r [7];
  assign N371 = N242 & N276;
  assign N372 = N242 & \nz.addr_r [7];
  assign N373 = N244 & N276;
  assign N374 = N244 & \nz.addr_r [7];
  assign N375 = N246 & N276;
  assign N376 = N246 & \nz.addr_r [7];
  assign N377 = N248 & N276;
  assign N378 = N248 & \nz.addr_r [7];
  assign N379 = N250 & N276;
  assign N380 = N250 & \nz.addr_r [7];
  assign N381 = N252 & N276;
  assign N382 = N252 & \nz.addr_r [7];
  assign N383 = N254 & N276;
  assign N384 = N254 & \nz.addr_r [7];
  assign N385 = N256 & N276;
  assign N386 = N256 & \nz.addr_r [7];
  assign N387 = N258 & N276;
  assign N388 = N258 & \nz.addr_r [7];
  assign N389 = N260 & N276;
  assign N390 = N260 & \nz.addr_r [7];
  assign N391 = N262 & N276;
  assign N392 = N262 & \nz.addr_r [7];
  assign N393 = N264 & N276;
  assign N394 = N264 & \nz.addr_r [7];
  assign N395 = N266 & N276;
  assign N396 = N266 & \nz.addr_r [7];
  assign N397 = N268 & N276;
  assign N398 = N268 & \nz.addr_r [7];
  assign N399 = N270 & N276;
  assign N400 = N270 & \nz.addr_r [7];
  assign N401 = N272 & N276;
  assign N402 = N272 & \nz.addr_r [7];
  assign N403 = N274 & N276;
  assign N404 = N274 & \nz.addr_r [7];
  assign N405 = N149 & N276;
  assign N406 = N149 & \nz.addr_r [7];
  assign N407 = N151 & N276;
  assign N408 = N151 & \nz.addr_r [7];
  assign N409 = N153 & N276;
  assign N410 = N153 & \nz.addr_r [7];
  assign N411 = N155 & N276;
  assign N412 = N155 & \nz.addr_r [7];
  assign N413 = N157 & N276;
  assign N414 = N157 & \nz.addr_r [7];
  assign N415 = N159 & N276;
  assign N416 = N159 & \nz.addr_r [7];
  assign N417 = N161 & N276;
  assign N418 = N161 & \nz.addr_r [7];
  assign N419 = N163 & N276;
  assign N420 = N163 & \nz.addr_r [7];
  assign N421 = N165 & N276;
  assign N422 = N165 & \nz.addr_r [7];
  assign N423 = N167 & N276;
  assign N424 = N167 & \nz.addr_r [7];
  assign N425 = N169 & N276;
  assign N426 = N169 & \nz.addr_r [7];
  assign N427 = N171 & N276;
  assign N428 = N171 & \nz.addr_r [7];
  assign N429 = N173 & N276;
  assign N430 = N173 & \nz.addr_r [7];
  assign N431 = N175 & N276;
  assign N432 = N175 & \nz.addr_r [7];
  assign N433 = N177 & N276;
  assign N434 = N177 & \nz.addr_r [7];
  assign N435 = N179 & N276;
  assign N436 = N179 & \nz.addr_r [7];
  assign N437 = N181 & N276;
  assign N438 = N181 & \nz.addr_r [7];
  assign N439 = N183 & N276;
  assign N440 = N183 & \nz.addr_r [7];
  assign N441 = N185 & N276;
  assign N442 = N185 & \nz.addr_r [7];
  assign N443 = N187 & N276;
  assign N444 = N187 & \nz.addr_r [7];
  assign N445 = N189 & N276;
  assign N446 = N189 & \nz.addr_r [7];
  assign N447 = N191 & N276;
  assign N448 = N191 & \nz.addr_r [7];
  assign N449 = N193 & N276;
  assign N450 = N193 & \nz.addr_r [7];
  assign N451 = N195 & N276;
  assign N452 = N195 & \nz.addr_r [7];
  assign N453 = N197 & N276;
  assign N454 = N197 & \nz.addr_r [7];
  assign N455 = N199 & N276;
  assign N456 = N199 & \nz.addr_r [7];
  assign N457 = N201 & N276;
  assign N458 = N201 & \nz.addr_r [7];
  assign N459 = N203 & N276;
  assign N460 = N203 & \nz.addr_r [7];
  assign N461 = N205 & N276;
  assign N462 = N205 & \nz.addr_r [7];
  assign N463 = N207 & N276;
  assign N464 = N207 & \nz.addr_r [7];
  assign N465 = N209 & N276;
  assign N466 = N209 & \nz.addr_r [7];
  assign N467 = N211 & N276;
  assign N468 = N211 & \nz.addr_r [7];
  assign N469 = N213 & N276;
  assign N470 = N213 & \nz.addr_r [7];
  assign N471 = N215 & N276;
  assign N472 = N215 & \nz.addr_r [7];
  assign N473 = N217 & N276;
  assign N474 = N217 & \nz.addr_r [7];
  assign N475 = N219 & N276;
  assign N476 = N219 & \nz.addr_r [7];
  assign N477 = N221 & N276;
  assign N478 = N221 & \nz.addr_r [7];
  assign N479 = N223 & N276;
  assign N480 = N223 & \nz.addr_r [7];
  assign N481 = N225 & N276;
  assign N482 = N225 & \nz.addr_r [7];
  assign N483 = N227 & N276;
  assign N484 = N227 & \nz.addr_r [7];
  assign N485 = N229 & N276;
  assign N486 = N229 & \nz.addr_r [7];
  assign N487 = N231 & N276;
  assign N488 = N231 & \nz.addr_r [7];
  assign N489 = N233 & N276;
  assign N490 = N233 & \nz.addr_r [7];
  assign N491 = N235 & N276;
  assign N492 = N235 & \nz.addr_r [7];
  assign N493 = N237 & N276;
  assign N494 = N237 & \nz.addr_r [7];
  assign N495 = N239 & N276;
  assign N496 = N239 & \nz.addr_r [7];
  assign N497 = N241 & N276;
  assign N498 = N241 & \nz.addr_r [7];
  assign N499 = N243 & N276;
  assign N500 = N243 & \nz.addr_r [7];
  assign N501 = N245 & N276;
  assign N502 = N245 & \nz.addr_r [7];
  assign N503 = N247 & N276;
  assign N504 = N247 & \nz.addr_r [7];
  assign N505 = N249 & N276;
  assign N506 = N249 & \nz.addr_r [7];
  assign N507 = N251 & N276;
  assign N508 = N251 & \nz.addr_r [7];
  assign N509 = N253 & N276;
  assign N510 = N253 & \nz.addr_r [7];
  assign N511 = N255 & N276;
  assign N512 = N255 & \nz.addr_r [7];
  assign N513 = N257 & N276;
  assign N514 = N257 & \nz.addr_r [7];
  assign N515 = N259 & N276;
  assign N516 = N259 & \nz.addr_r [7];
  assign N517 = N261 & N276;
  assign N518 = N261 & \nz.addr_r [7];
  assign N519 = N263 & N276;
  assign N520 = N263 & \nz.addr_r [7];
  assign N521 = N265 & N276;
  assign N522 = N265 & \nz.addr_r [7];
  assign N523 = N267 & N276;
  assign N524 = N267 & \nz.addr_r [7];
  assign N525 = N269 & N276;
  assign N526 = N269 & \nz.addr_r [7];
  assign N527 = N271 & N276;
  assign N528 = N271 & \nz.addr_r [7];
  assign N529 = N273 & N276;
  assign N530 = N273 & \nz.addr_r [7];
  assign N531 = N275 & N276;
  assign N532 = N275 & \nz.addr_r [7];
  assign N533 = v_i & w_i;
  assign N534 = ~N533;

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_7_sv2v_reg  <= addr_i[7];
      \nz.addr_r_6_sv2v_reg  <= addr_i[6];
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N1046) begin
      \nz.mem_2047_sv2v_reg  <= data_i[7];
      \nz.mem_2046_sv2v_reg  <= data_i[6];
      \nz.mem_2045_sv2v_reg  <= data_i[5];
      \nz.mem_2044_sv2v_reg  <= data_i[4];
      \nz.mem_2043_sv2v_reg  <= data_i[3];
      \nz.mem_2042_sv2v_reg  <= data_i[2];
      \nz.mem_2041_sv2v_reg  <= data_i[1];
      \nz.mem_2040_sv2v_reg  <= data_i[0];
    end 
    if(N1045) begin
      \nz.mem_2039_sv2v_reg  <= data_i[7];
      \nz.mem_2038_sv2v_reg  <= data_i[6];
      \nz.mem_2037_sv2v_reg  <= data_i[5];
      \nz.mem_2036_sv2v_reg  <= data_i[4];
      \nz.mem_2035_sv2v_reg  <= data_i[3];
      \nz.mem_2034_sv2v_reg  <= data_i[2];
      \nz.mem_2033_sv2v_reg  <= data_i[1];
      \nz.mem_2032_sv2v_reg  <= data_i[0];
    end 
    if(N1044) begin
      \nz.mem_2031_sv2v_reg  <= data_i[7];
      \nz.mem_2030_sv2v_reg  <= data_i[6];
      \nz.mem_2029_sv2v_reg  <= data_i[5];
      \nz.mem_2028_sv2v_reg  <= data_i[4];
      \nz.mem_2027_sv2v_reg  <= data_i[3];
      \nz.mem_2026_sv2v_reg  <= data_i[2];
      \nz.mem_2025_sv2v_reg  <= data_i[1];
      \nz.mem_2024_sv2v_reg  <= data_i[0];
    end 
    if(N1043) begin
      \nz.mem_2023_sv2v_reg  <= data_i[7];
      \nz.mem_2022_sv2v_reg  <= data_i[6];
      \nz.mem_2021_sv2v_reg  <= data_i[5];
      \nz.mem_2020_sv2v_reg  <= data_i[4];
      \nz.mem_2019_sv2v_reg  <= data_i[3];
      \nz.mem_2018_sv2v_reg  <= data_i[2];
      \nz.mem_2017_sv2v_reg  <= data_i[1];
      \nz.mem_2016_sv2v_reg  <= data_i[0];
    end 
    if(N1042) begin
      \nz.mem_2015_sv2v_reg  <= data_i[7];
      \nz.mem_2014_sv2v_reg  <= data_i[6];
      \nz.mem_2013_sv2v_reg  <= data_i[5];
      \nz.mem_2012_sv2v_reg  <= data_i[4];
      \nz.mem_2011_sv2v_reg  <= data_i[3];
      \nz.mem_2010_sv2v_reg  <= data_i[2];
      \nz.mem_2009_sv2v_reg  <= data_i[1];
      \nz.mem_2008_sv2v_reg  <= data_i[0];
    end 
    if(N1041) begin
      \nz.mem_2007_sv2v_reg  <= data_i[7];
      \nz.mem_2006_sv2v_reg  <= data_i[6];
      \nz.mem_2005_sv2v_reg  <= data_i[5];
      \nz.mem_2004_sv2v_reg  <= data_i[4];
      \nz.mem_2003_sv2v_reg  <= data_i[3];
      \nz.mem_2002_sv2v_reg  <= data_i[2];
      \nz.mem_2001_sv2v_reg  <= data_i[1];
      \nz.mem_2000_sv2v_reg  <= data_i[0];
    end 
    if(N1040) begin
      \nz.mem_1999_sv2v_reg  <= data_i[7];
      \nz.mem_1998_sv2v_reg  <= data_i[6];
      \nz.mem_1997_sv2v_reg  <= data_i[5];
      \nz.mem_1996_sv2v_reg  <= data_i[4];
      \nz.mem_1995_sv2v_reg  <= data_i[3];
      \nz.mem_1994_sv2v_reg  <= data_i[2];
      \nz.mem_1993_sv2v_reg  <= data_i[1];
      \nz.mem_1992_sv2v_reg  <= data_i[0];
    end 
    if(N1039) begin
      \nz.mem_1991_sv2v_reg  <= data_i[7];
      \nz.mem_1990_sv2v_reg  <= data_i[6];
      \nz.mem_1989_sv2v_reg  <= data_i[5];
      \nz.mem_1988_sv2v_reg  <= data_i[4];
      \nz.mem_1987_sv2v_reg  <= data_i[3];
      \nz.mem_1986_sv2v_reg  <= data_i[2];
      \nz.mem_1985_sv2v_reg  <= data_i[1];
      \nz.mem_1984_sv2v_reg  <= data_i[0];
    end 
    if(N1038) begin
      \nz.mem_1983_sv2v_reg  <= data_i[7];
      \nz.mem_1982_sv2v_reg  <= data_i[6];
      \nz.mem_1981_sv2v_reg  <= data_i[5];
      \nz.mem_1980_sv2v_reg  <= data_i[4];
      \nz.mem_1979_sv2v_reg  <= data_i[3];
      \nz.mem_1978_sv2v_reg  <= data_i[2];
      \nz.mem_1977_sv2v_reg  <= data_i[1];
      \nz.mem_1976_sv2v_reg  <= data_i[0];
    end 
    if(N1037) begin
      \nz.mem_1975_sv2v_reg  <= data_i[7];
      \nz.mem_1974_sv2v_reg  <= data_i[6];
      \nz.mem_1973_sv2v_reg  <= data_i[5];
      \nz.mem_1972_sv2v_reg  <= data_i[4];
      \nz.mem_1971_sv2v_reg  <= data_i[3];
      \nz.mem_1970_sv2v_reg  <= data_i[2];
      \nz.mem_1969_sv2v_reg  <= data_i[1];
      \nz.mem_1968_sv2v_reg  <= data_i[0];
    end 
    if(N1036) begin
      \nz.mem_1967_sv2v_reg  <= data_i[7];
      \nz.mem_1966_sv2v_reg  <= data_i[6];
      \nz.mem_1965_sv2v_reg  <= data_i[5];
      \nz.mem_1964_sv2v_reg  <= data_i[4];
      \nz.mem_1963_sv2v_reg  <= data_i[3];
      \nz.mem_1962_sv2v_reg  <= data_i[2];
      \nz.mem_1961_sv2v_reg  <= data_i[1];
      \nz.mem_1960_sv2v_reg  <= data_i[0];
    end 
    if(N1035) begin
      \nz.mem_1959_sv2v_reg  <= data_i[7];
      \nz.mem_1958_sv2v_reg  <= data_i[6];
      \nz.mem_1957_sv2v_reg  <= data_i[5];
      \nz.mem_1956_sv2v_reg  <= data_i[4];
      \nz.mem_1955_sv2v_reg  <= data_i[3];
      \nz.mem_1954_sv2v_reg  <= data_i[2];
      \nz.mem_1953_sv2v_reg  <= data_i[1];
      \nz.mem_1952_sv2v_reg  <= data_i[0];
    end 
    if(N1034) begin
      \nz.mem_1951_sv2v_reg  <= data_i[7];
      \nz.mem_1950_sv2v_reg  <= data_i[6];
      \nz.mem_1949_sv2v_reg  <= data_i[5];
      \nz.mem_1948_sv2v_reg  <= data_i[4];
      \nz.mem_1947_sv2v_reg  <= data_i[3];
      \nz.mem_1946_sv2v_reg  <= data_i[2];
      \nz.mem_1945_sv2v_reg  <= data_i[1];
      \nz.mem_1944_sv2v_reg  <= data_i[0];
    end 
    if(N1033) begin
      \nz.mem_1943_sv2v_reg  <= data_i[7];
      \nz.mem_1942_sv2v_reg  <= data_i[6];
      \nz.mem_1941_sv2v_reg  <= data_i[5];
      \nz.mem_1940_sv2v_reg  <= data_i[4];
      \nz.mem_1939_sv2v_reg  <= data_i[3];
      \nz.mem_1938_sv2v_reg  <= data_i[2];
      \nz.mem_1937_sv2v_reg  <= data_i[1];
      \nz.mem_1936_sv2v_reg  <= data_i[0];
    end 
    if(N1032) begin
      \nz.mem_1935_sv2v_reg  <= data_i[7];
      \nz.mem_1934_sv2v_reg  <= data_i[6];
      \nz.mem_1933_sv2v_reg  <= data_i[5];
      \nz.mem_1932_sv2v_reg  <= data_i[4];
      \nz.mem_1931_sv2v_reg  <= data_i[3];
      \nz.mem_1930_sv2v_reg  <= data_i[2];
      \nz.mem_1929_sv2v_reg  <= data_i[1];
      \nz.mem_1928_sv2v_reg  <= data_i[0];
    end 
    if(N1031) begin
      \nz.mem_1927_sv2v_reg  <= data_i[7];
      \nz.mem_1926_sv2v_reg  <= data_i[6];
      \nz.mem_1925_sv2v_reg  <= data_i[5];
      \nz.mem_1924_sv2v_reg  <= data_i[4];
      \nz.mem_1923_sv2v_reg  <= data_i[3];
      \nz.mem_1922_sv2v_reg  <= data_i[2];
      \nz.mem_1921_sv2v_reg  <= data_i[1];
      \nz.mem_1920_sv2v_reg  <= data_i[0];
    end 
    if(N1030) begin
      \nz.mem_1919_sv2v_reg  <= data_i[7];
      \nz.mem_1918_sv2v_reg  <= data_i[6];
      \nz.mem_1917_sv2v_reg  <= data_i[5];
      \nz.mem_1916_sv2v_reg  <= data_i[4];
      \nz.mem_1915_sv2v_reg  <= data_i[3];
      \nz.mem_1914_sv2v_reg  <= data_i[2];
      \nz.mem_1913_sv2v_reg  <= data_i[1];
      \nz.mem_1912_sv2v_reg  <= data_i[0];
    end 
    if(N1029) begin
      \nz.mem_1911_sv2v_reg  <= data_i[7];
      \nz.mem_1910_sv2v_reg  <= data_i[6];
      \nz.mem_1909_sv2v_reg  <= data_i[5];
      \nz.mem_1908_sv2v_reg  <= data_i[4];
      \nz.mem_1907_sv2v_reg  <= data_i[3];
      \nz.mem_1906_sv2v_reg  <= data_i[2];
      \nz.mem_1905_sv2v_reg  <= data_i[1];
      \nz.mem_1904_sv2v_reg  <= data_i[0];
    end 
    if(N1028) begin
      \nz.mem_1903_sv2v_reg  <= data_i[7];
      \nz.mem_1902_sv2v_reg  <= data_i[6];
      \nz.mem_1901_sv2v_reg  <= data_i[5];
      \nz.mem_1900_sv2v_reg  <= data_i[4];
      \nz.mem_1899_sv2v_reg  <= data_i[3];
      \nz.mem_1898_sv2v_reg  <= data_i[2];
      \nz.mem_1897_sv2v_reg  <= data_i[1];
      \nz.mem_1896_sv2v_reg  <= data_i[0];
    end 
    if(N1027) begin
      \nz.mem_1895_sv2v_reg  <= data_i[7];
      \nz.mem_1894_sv2v_reg  <= data_i[6];
      \nz.mem_1893_sv2v_reg  <= data_i[5];
      \nz.mem_1892_sv2v_reg  <= data_i[4];
      \nz.mem_1891_sv2v_reg  <= data_i[3];
      \nz.mem_1890_sv2v_reg  <= data_i[2];
      \nz.mem_1889_sv2v_reg  <= data_i[1];
      \nz.mem_1888_sv2v_reg  <= data_i[0];
    end 
    if(N1026) begin
      \nz.mem_1887_sv2v_reg  <= data_i[7];
      \nz.mem_1886_sv2v_reg  <= data_i[6];
      \nz.mem_1885_sv2v_reg  <= data_i[5];
      \nz.mem_1884_sv2v_reg  <= data_i[4];
      \nz.mem_1883_sv2v_reg  <= data_i[3];
      \nz.mem_1882_sv2v_reg  <= data_i[2];
      \nz.mem_1881_sv2v_reg  <= data_i[1];
      \nz.mem_1880_sv2v_reg  <= data_i[0];
    end 
    if(N1025) begin
      \nz.mem_1879_sv2v_reg  <= data_i[7];
      \nz.mem_1878_sv2v_reg  <= data_i[6];
      \nz.mem_1877_sv2v_reg  <= data_i[5];
      \nz.mem_1876_sv2v_reg  <= data_i[4];
      \nz.mem_1875_sv2v_reg  <= data_i[3];
      \nz.mem_1874_sv2v_reg  <= data_i[2];
      \nz.mem_1873_sv2v_reg  <= data_i[1];
      \nz.mem_1872_sv2v_reg  <= data_i[0];
    end 
    if(N1024) begin
      \nz.mem_1871_sv2v_reg  <= data_i[7];
      \nz.mem_1870_sv2v_reg  <= data_i[6];
      \nz.mem_1869_sv2v_reg  <= data_i[5];
      \nz.mem_1868_sv2v_reg  <= data_i[4];
      \nz.mem_1867_sv2v_reg  <= data_i[3];
      \nz.mem_1866_sv2v_reg  <= data_i[2];
      \nz.mem_1865_sv2v_reg  <= data_i[1];
      \nz.mem_1864_sv2v_reg  <= data_i[0];
    end 
    if(N1023) begin
      \nz.mem_1863_sv2v_reg  <= data_i[7];
      \nz.mem_1862_sv2v_reg  <= data_i[6];
      \nz.mem_1861_sv2v_reg  <= data_i[5];
      \nz.mem_1860_sv2v_reg  <= data_i[4];
      \nz.mem_1859_sv2v_reg  <= data_i[3];
      \nz.mem_1858_sv2v_reg  <= data_i[2];
      \nz.mem_1857_sv2v_reg  <= data_i[1];
      \nz.mem_1856_sv2v_reg  <= data_i[0];
    end 
    if(N1022) begin
      \nz.mem_1855_sv2v_reg  <= data_i[7];
      \nz.mem_1854_sv2v_reg  <= data_i[6];
      \nz.mem_1853_sv2v_reg  <= data_i[5];
      \nz.mem_1852_sv2v_reg  <= data_i[4];
      \nz.mem_1851_sv2v_reg  <= data_i[3];
      \nz.mem_1850_sv2v_reg  <= data_i[2];
      \nz.mem_1849_sv2v_reg  <= data_i[1];
      \nz.mem_1848_sv2v_reg  <= data_i[0];
    end 
    if(N1021) begin
      \nz.mem_1847_sv2v_reg  <= data_i[7];
      \nz.mem_1846_sv2v_reg  <= data_i[6];
      \nz.mem_1845_sv2v_reg  <= data_i[5];
      \nz.mem_1844_sv2v_reg  <= data_i[4];
      \nz.mem_1843_sv2v_reg  <= data_i[3];
      \nz.mem_1842_sv2v_reg  <= data_i[2];
      \nz.mem_1841_sv2v_reg  <= data_i[1];
      \nz.mem_1840_sv2v_reg  <= data_i[0];
    end 
    if(N1020) begin
      \nz.mem_1839_sv2v_reg  <= data_i[7];
      \nz.mem_1838_sv2v_reg  <= data_i[6];
      \nz.mem_1837_sv2v_reg  <= data_i[5];
      \nz.mem_1836_sv2v_reg  <= data_i[4];
      \nz.mem_1835_sv2v_reg  <= data_i[3];
      \nz.mem_1834_sv2v_reg  <= data_i[2];
      \nz.mem_1833_sv2v_reg  <= data_i[1];
      \nz.mem_1832_sv2v_reg  <= data_i[0];
    end 
    if(N1019) begin
      \nz.mem_1831_sv2v_reg  <= data_i[7];
      \nz.mem_1830_sv2v_reg  <= data_i[6];
      \nz.mem_1829_sv2v_reg  <= data_i[5];
      \nz.mem_1828_sv2v_reg  <= data_i[4];
      \nz.mem_1827_sv2v_reg  <= data_i[3];
      \nz.mem_1826_sv2v_reg  <= data_i[2];
      \nz.mem_1825_sv2v_reg  <= data_i[1];
      \nz.mem_1824_sv2v_reg  <= data_i[0];
    end 
    if(N1018) begin
      \nz.mem_1823_sv2v_reg  <= data_i[7];
      \nz.mem_1822_sv2v_reg  <= data_i[6];
      \nz.mem_1821_sv2v_reg  <= data_i[5];
      \nz.mem_1820_sv2v_reg  <= data_i[4];
      \nz.mem_1819_sv2v_reg  <= data_i[3];
      \nz.mem_1818_sv2v_reg  <= data_i[2];
      \nz.mem_1817_sv2v_reg  <= data_i[1];
      \nz.mem_1816_sv2v_reg  <= data_i[0];
    end 
    if(N1017) begin
      \nz.mem_1815_sv2v_reg  <= data_i[7];
      \nz.mem_1814_sv2v_reg  <= data_i[6];
      \nz.mem_1813_sv2v_reg  <= data_i[5];
      \nz.mem_1812_sv2v_reg  <= data_i[4];
      \nz.mem_1811_sv2v_reg  <= data_i[3];
      \nz.mem_1810_sv2v_reg  <= data_i[2];
      \nz.mem_1809_sv2v_reg  <= data_i[1];
      \nz.mem_1808_sv2v_reg  <= data_i[0];
    end 
    if(N1016) begin
      \nz.mem_1807_sv2v_reg  <= data_i[7];
      \nz.mem_1806_sv2v_reg  <= data_i[6];
      \nz.mem_1805_sv2v_reg  <= data_i[5];
      \nz.mem_1804_sv2v_reg  <= data_i[4];
      \nz.mem_1803_sv2v_reg  <= data_i[3];
      \nz.mem_1802_sv2v_reg  <= data_i[2];
      \nz.mem_1801_sv2v_reg  <= data_i[1];
      \nz.mem_1800_sv2v_reg  <= data_i[0];
    end 
    if(N1015) begin
      \nz.mem_1799_sv2v_reg  <= data_i[7];
      \nz.mem_1798_sv2v_reg  <= data_i[6];
      \nz.mem_1797_sv2v_reg  <= data_i[5];
      \nz.mem_1796_sv2v_reg  <= data_i[4];
      \nz.mem_1795_sv2v_reg  <= data_i[3];
      \nz.mem_1794_sv2v_reg  <= data_i[2];
      \nz.mem_1793_sv2v_reg  <= data_i[1];
      \nz.mem_1792_sv2v_reg  <= data_i[0];
    end 
    if(N1014) begin
      \nz.mem_1791_sv2v_reg  <= data_i[7];
      \nz.mem_1790_sv2v_reg  <= data_i[6];
      \nz.mem_1789_sv2v_reg  <= data_i[5];
      \nz.mem_1788_sv2v_reg  <= data_i[4];
      \nz.mem_1787_sv2v_reg  <= data_i[3];
      \nz.mem_1786_sv2v_reg  <= data_i[2];
      \nz.mem_1785_sv2v_reg  <= data_i[1];
      \nz.mem_1784_sv2v_reg  <= data_i[0];
    end 
    if(N1013) begin
      \nz.mem_1783_sv2v_reg  <= data_i[7];
      \nz.mem_1782_sv2v_reg  <= data_i[6];
      \nz.mem_1781_sv2v_reg  <= data_i[5];
      \nz.mem_1780_sv2v_reg  <= data_i[4];
      \nz.mem_1779_sv2v_reg  <= data_i[3];
      \nz.mem_1778_sv2v_reg  <= data_i[2];
      \nz.mem_1777_sv2v_reg  <= data_i[1];
      \nz.mem_1776_sv2v_reg  <= data_i[0];
    end 
    if(N1012) begin
      \nz.mem_1775_sv2v_reg  <= data_i[7];
      \nz.mem_1774_sv2v_reg  <= data_i[6];
      \nz.mem_1773_sv2v_reg  <= data_i[5];
      \nz.mem_1772_sv2v_reg  <= data_i[4];
      \nz.mem_1771_sv2v_reg  <= data_i[3];
      \nz.mem_1770_sv2v_reg  <= data_i[2];
      \nz.mem_1769_sv2v_reg  <= data_i[1];
      \nz.mem_1768_sv2v_reg  <= data_i[0];
    end 
    if(N1011) begin
      \nz.mem_1767_sv2v_reg  <= data_i[7];
      \nz.mem_1766_sv2v_reg  <= data_i[6];
      \nz.mem_1765_sv2v_reg  <= data_i[5];
      \nz.mem_1764_sv2v_reg  <= data_i[4];
      \nz.mem_1763_sv2v_reg  <= data_i[3];
      \nz.mem_1762_sv2v_reg  <= data_i[2];
      \nz.mem_1761_sv2v_reg  <= data_i[1];
      \nz.mem_1760_sv2v_reg  <= data_i[0];
    end 
    if(N1010) begin
      \nz.mem_1759_sv2v_reg  <= data_i[7];
      \nz.mem_1758_sv2v_reg  <= data_i[6];
      \nz.mem_1757_sv2v_reg  <= data_i[5];
      \nz.mem_1756_sv2v_reg  <= data_i[4];
      \nz.mem_1755_sv2v_reg  <= data_i[3];
      \nz.mem_1754_sv2v_reg  <= data_i[2];
      \nz.mem_1753_sv2v_reg  <= data_i[1];
      \nz.mem_1752_sv2v_reg  <= data_i[0];
    end 
    if(N1009) begin
      \nz.mem_1751_sv2v_reg  <= data_i[7];
      \nz.mem_1750_sv2v_reg  <= data_i[6];
      \nz.mem_1749_sv2v_reg  <= data_i[5];
      \nz.mem_1748_sv2v_reg  <= data_i[4];
      \nz.mem_1747_sv2v_reg  <= data_i[3];
      \nz.mem_1746_sv2v_reg  <= data_i[2];
      \nz.mem_1745_sv2v_reg  <= data_i[1];
      \nz.mem_1744_sv2v_reg  <= data_i[0];
    end 
    if(N1008) begin
      \nz.mem_1743_sv2v_reg  <= data_i[7];
      \nz.mem_1742_sv2v_reg  <= data_i[6];
      \nz.mem_1741_sv2v_reg  <= data_i[5];
      \nz.mem_1740_sv2v_reg  <= data_i[4];
      \nz.mem_1739_sv2v_reg  <= data_i[3];
      \nz.mem_1738_sv2v_reg  <= data_i[2];
      \nz.mem_1737_sv2v_reg  <= data_i[1];
      \nz.mem_1736_sv2v_reg  <= data_i[0];
    end 
    if(N1007) begin
      \nz.mem_1735_sv2v_reg  <= data_i[7];
      \nz.mem_1734_sv2v_reg  <= data_i[6];
      \nz.mem_1733_sv2v_reg  <= data_i[5];
      \nz.mem_1732_sv2v_reg  <= data_i[4];
      \nz.mem_1731_sv2v_reg  <= data_i[3];
      \nz.mem_1730_sv2v_reg  <= data_i[2];
      \nz.mem_1729_sv2v_reg  <= data_i[1];
      \nz.mem_1728_sv2v_reg  <= data_i[0];
    end 
    if(N1006) begin
      \nz.mem_1727_sv2v_reg  <= data_i[7];
      \nz.mem_1726_sv2v_reg  <= data_i[6];
      \nz.mem_1725_sv2v_reg  <= data_i[5];
      \nz.mem_1724_sv2v_reg  <= data_i[4];
      \nz.mem_1723_sv2v_reg  <= data_i[3];
      \nz.mem_1722_sv2v_reg  <= data_i[2];
      \nz.mem_1721_sv2v_reg  <= data_i[1];
      \nz.mem_1720_sv2v_reg  <= data_i[0];
    end 
    if(N1005) begin
      \nz.mem_1719_sv2v_reg  <= data_i[7];
      \nz.mem_1718_sv2v_reg  <= data_i[6];
      \nz.mem_1717_sv2v_reg  <= data_i[5];
      \nz.mem_1716_sv2v_reg  <= data_i[4];
      \nz.mem_1715_sv2v_reg  <= data_i[3];
      \nz.mem_1714_sv2v_reg  <= data_i[2];
      \nz.mem_1713_sv2v_reg  <= data_i[1];
      \nz.mem_1712_sv2v_reg  <= data_i[0];
    end 
    if(N1004) begin
      \nz.mem_1711_sv2v_reg  <= data_i[7];
      \nz.mem_1710_sv2v_reg  <= data_i[6];
      \nz.mem_1709_sv2v_reg  <= data_i[5];
      \nz.mem_1708_sv2v_reg  <= data_i[4];
      \nz.mem_1707_sv2v_reg  <= data_i[3];
      \nz.mem_1706_sv2v_reg  <= data_i[2];
      \nz.mem_1705_sv2v_reg  <= data_i[1];
      \nz.mem_1704_sv2v_reg  <= data_i[0];
    end 
    if(N1003) begin
      \nz.mem_1703_sv2v_reg  <= data_i[7];
      \nz.mem_1702_sv2v_reg  <= data_i[6];
      \nz.mem_1701_sv2v_reg  <= data_i[5];
      \nz.mem_1700_sv2v_reg  <= data_i[4];
      \nz.mem_1699_sv2v_reg  <= data_i[3];
      \nz.mem_1698_sv2v_reg  <= data_i[2];
      \nz.mem_1697_sv2v_reg  <= data_i[1];
      \nz.mem_1696_sv2v_reg  <= data_i[0];
    end 
    if(N1002) begin
      \nz.mem_1695_sv2v_reg  <= data_i[7];
      \nz.mem_1694_sv2v_reg  <= data_i[6];
      \nz.mem_1693_sv2v_reg  <= data_i[5];
      \nz.mem_1692_sv2v_reg  <= data_i[4];
      \nz.mem_1691_sv2v_reg  <= data_i[3];
      \nz.mem_1690_sv2v_reg  <= data_i[2];
      \nz.mem_1689_sv2v_reg  <= data_i[1];
      \nz.mem_1688_sv2v_reg  <= data_i[0];
    end 
    if(N1001) begin
      \nz.mem_1687_sv2v_reg  <= data_i[7];
      \nz.mem_1686_sv2v_reg  <= data_i[6];
      \nz.mem_1685_sv2v_reg  <= data_i[5];
      \nz.mem_1684_sv2v_reg  <= data_i[4];
      \nz.mem_1683_sv2v_reg  <= data_i[3];
      \nz.mem_1682_sv2v_reg  <= data_i[2];
      \nz.mem_1681_sv2v_reg  <= data_i[1];
      \nz.mem_1680_sv2v_reg  <= data_i[0];
    end 
    if(N1000) begin
      \nz.mem_1679_sv2v_reg  <= data_i[7];
      \nz.mem_1678_sv2v_reg  <= data_i[6];
      \nz.mem_1677_sv2v_reg  <= data_i[5];
      \nz.mem_1676_sv2v_reg  <= data_i[4];
      \nz.mem_1675_sv2v_reg  <= data_i[3];
      \nz.mem_1674_sv2v_reg  <= data_i[2];
      \nz.mem_1673_sv2v_reg  <= data_i[1];
      \nz.mem_1672_sv2v_reg  <= data_i[0];
    end 
    if(N999) begin
      \nz.mem_1671_sv2v_reg  <= data_i[7];
      \nz.mem_1670_sv2v_reg  <= data_i[6];
      \nz.mem_1669_sv2v_reg  <= data_i[5];
      \nz.mem_1668_sv2v_reg  <= data_i[4];
      \nz.mem_1667_sv2v_reg  <= data_i[3];
      \nz.mem_1666_sv2v_reg  <= data_i[2];
      \nz.mem_1665_sv2v_reg  <= data_i[1];
      \nz.mem_1664_sv2v_reg  <= data_i[0];
    end 
    if(N998) begin
      \nz.mem_1663_sv2v_reg  <= data_i[7];
      \nz.mem_1662_sv2v_reg  <= data_i[6];
      \nz.mem_1661_sv2v_reg  <= data_i[5];
      \nz.mem_1660_sv2v_reg  <= data_i[4];
      \nz.mem_1659_sv2v_reg  <= data_i[3];
      \nz.mem_1658_sv2v_reg  <= data_i[2];
      \nz.mem_1657_sv2v_reg  <= data_i[1];
      \nz.mem_1656_sv2v_reg  <= data_i[0];
    end 
    if(N997) begin
      \nz.mem_1655_sv2v_reg  <= data_i[7];
      \nz.mem_1654_sv2v_reg  <= data_i[6];
      \nz.mem_1653_sv2v_reg  <= data_i[5];
      \nz.mem_1652_sv2v_reg  <= data_i[4];
      \nz.mem_1651_sv2v_reg  <= data_i[3];
      \nz.mem_1650_sv2v_reg  <= data_i[2];
      \nz.mem_1649_sv2v_reg  <= data_i[1];
      \nz.mem_1648_sv2v_reg  <= data_i[0];
    end 
    if(N996) begin
      \nz.mem_1647_sv2v_reg  <= data_i[7];
      \nz.mem_1646_sv2v_reg  <= data_i[6];
      \nz.mem_1645_sv2v_reg  <= data_i[5];
      \nz.mem_1644_sv2v_reg  <= data_i[4];
      \nz.mem_1643_sv2v_reg  <= data_i[3];
      \nz.mem_1642_sv2v_reg  <= data_i[2];
      \nz.mem_1641_sv2v_reg  <= data_i[1];
      \nz.mem_1640_sv2v_reg  <= data_i[0];
    end 
    if(N995) begin
      \nz.mem_1639_sv2v_reg  <= data_i[7];
      \nz.mem_1638_sv2v_reg  <= data_i[6];
      \nz.mem_1637_sv2v_reg  <= data_i[5];
      \nz.mem_1636_sv2v_reg  <= data_i[4];
      \nz.mem_1635_sv2v_reg  <= data_i[3];
      \nz.mem_1634_sv2v_reg  <= data_i[2];
      \nz.mem_1633_sv2v_reg  <= data_i[1];
      \nz.mem_1632_sv2v_reg  <= data_i[0];
    end 
    if(N994) begin
      \nz.mem_1631_sv2v_reg  <= data_i[7];
      \nz.mem_1630_sv2v_reg  <= data_i[6];
      \nz.mem_1629_sv2v_reg  <= data_i[5];
      \nz.mem_1628_sv2v_reg  <= data_i[4];
      \nz.mem_1627_sv2v_reg  <= data_i[3];
      \nz.mem_1626_sv2v_reg  <= data_i[2];
      \nz.mem_1625_sv2v_reg  <= data_i[1];
      \nz.mem_1624_sv2v_reg  <= data_i[0];
    end 
    if(N993) begin
      \nz.mem_1623_sv2v_reg  <= data_i[7];
      \nz.mem_1622_sv2v_reg  <= data_i[6];
      \nz.mem_1621_sv2v_reg  <= data_i[5];
      \nz.mem_1620_sv2v_reg  <= data_i[4];
      \nz.mem_1619_sv2v_reg  <= data_i[3];
      \nz.mem_1618_sv2v_reg  <= data_i[2];
      \nz.mem_1617_sv2v_reg  <= data_i[1];
      \nz.mem_1616_sv2v_reg  <= data_i[0];
    end 
    if(N992) begin
      \nz.mem_1615_sv2v_reg  <= data_i[7];
      \nz.mem_1614_sv2v_reg  <= data_i[6];
      \nz.mem_1613_sv2v_reg  <= data_i[5];
      \nz.mem_1612_sv2v_reg  <= data_i[4];
      \nz.mem_1611_sv2v_reg  <= data_i[3];
      \nz.mem_1610_sv2v_reg  <= data_i[2];
      \nz.mem_1609_sv2v_reg  <= data_i[1];
      \nz.mem_1608_sv2v_reg  <= data_i[0];
    end 
    if(N991) begin
      \nz.mem_1607_sv2v_reg  <= data_i[7];
      \nz.mem_1606_sv2v_reg  <= data_i[6];
      \nz.mem_1605_sv2v_reg  <= data_i[5];
      \nz.mem_1604_sv2v_reg  <= data_i[4];
      \nz.mem_1603_sv2v_reg  <= data_i[3];
      \nz.mem_1602_sv2v_reg  <= data_i[2];
      \nz.mem_1601_sv2v_reg  <= data_i[1];
      \nz.mem_1600_sv2v_reg  <= data_i[0];
    end 
    if(N990) begin
      \nz.mem_1599_sv2v_reg  <= data_i[7];
      \nz.mem_1598_sv2v_reg  <= data_i[6];
      \nz.mem_1597_sv2v_reg  <= data_i[5];
      \nz.mem_1596_sv2v_reg  <= data_i[4];
      \nz.mem_1595_sv2v_reg  <= data_i[3];
      \nz.mem_1594_sv2v_reg  <= data_i[2];
      \nz.mem_1593_sv2v_reg  <= data_i[1];
      \nz.mem_1592_sv2v_reg  <= data_i[0];
    end 
    if(N989) begin
      \nz.mem_1591_sv2v_reg  <= data_i[7];
      \nz.mem_1590_sv2v_reg  <= data_i[6];
      \nz.mem_1589_sv2v_reg  <= data_i[5];
      \nz.mem_1588_sv2v_reg  <= data_i[4];
      \nz.mem_1587_sv2v_reg  <= data_i[3];
      \nz.mem_1586_sv2v_reg  <= data_i[2];
      \nz.mem_1585_sv2v_reg  <= data_i[1];
      \nz.mem_1584_sv2v_reg  <= data_i[0];
    end 
    if(N988) begin
      \nz.mem_1583_sv2v_reg  <= data_i[7];
      \nz.mem_1582_sv2v_reg  <= data_i[6];
      \nz.mem_1581_sv2v_reg  <= data_i[5];
      \nz.mem_1580_sv2v_reg  <= data_i[4];
      \nz.mem_1579_sv2v_reg  <= data_i[3];
      \nz.mem_1578_sv2v_reg  <= data_i[2];
      \nz.mem_1577_sv2v_reg  <= data_i[1];
      \nz.mem_1576_sv2v_reg  <= data_i[0];
    end 
    if(N987) begin
      \nz.mem_1575_sv2v_reg  <= data_i[7];
      \nz.mem_1574_sv2v_reg  <= data_i[6];
      \nz.mem_1573_sv2v_reg  <= data_i[5];
      \nz.mem_1572_sv2v_reg  <= data_i[4];
      \nz.mem_1571_sv2v_reg  <= data_i[3];
      \nz.mem_1570_sv2v_reg  <= data_i[2];
      \nz.mem_1569_sv2v_reg  <= data_i[1];
      \nz.mem_1568_sv2v_reg  <= data_i[0];
    end 
    if(N986) begin
      \nz.mem_1567_sv2v_reg  <= data_i[7];
      \nz.mem_1566_sv2v_reg  <= data_i[6];
      \nz.mem_1565_sv2v_reg  <= data_i[5];
      \nz.mem_1564_sv2v_reg  <= data_i[4];
      \nz.mem_1563_sv2v_reg  <= data_i[3];
      \nz.mem_1562_sv2v_reg  <= data_i[2];
      \nz.mem_1561_sv2v_reg  <= data_i[1];
      \nz.mem_1560_sv2v_reg  <= data_i[0];
    end 
    if(N985) begin
      \nz.mem_1559_sv2v_reg  <= data_i[7];
      \nz.mem_1558_sv2v_reg  <= data_i[6];
      \nz.mem_1557_sv2v_reg  <= data_i[5];
      \nz.mem_1556_sv2v_reg  <= data_i[4];
      \nz.mem_1555_sv2v_reg  <= data_i[3];
      \nz.mem_1554_sv2v_reg  <= data_i[2];
      \nz.mem_1553_sv2v_reg  <= data_i[1];
      \nz.mem_1552_sv2v_reg  <= data_i[0];
    end 
    if(N984) begin
      \nz.mem_1551_sv2v_reg  <= data_i[7];
      \nz.mem_1550_sv2v_reg  <= data_i[6];
      \nz.mem_1549_sv2v_reg  <= data_i[5];
      \nz.mem_1548_sv2v_reg  <= data_i[4];
      \nz.mem_1547_sv2v_reg  <= data_i[3];
      \nz.mem_1546_sv2v_reg  <= data_i[2];
      \nz.mem_1545_sv2v_reg  <= data_i[1];
      \nz.mem_1544_sv2v_reg  <= data_i[0];
    end 
    if(N983) begin
      \nz.mem_1543_sv2v_reg  <= data_i[7];
      \nz.mem_1542_sv2v_reg  <= data_i[6];
      \nz.mem_1541_sv2v_reg  <= data_i[5];
      \nz.mem_1540_sv2v_reg  <= data_i[4];
      \nz.mem_1539_sv2v_reg  <= data_i[3];
      \nz.mem_1538_sv2v_reg  <= data_i[2];
      \nz.mem_1537_sv2v_reg  <= data_i[1];
      \nz.mem_1536_sv2v_reg  <= data_i[0];
    end 
    if(N982) begin
      \nz.mem_1535_sv2v_reg  <= data_i[7];
      \nz.mem_1534_sv2v_reg  <= data_i[6];
      \nz.mem_1533_sv2v_reg  <= data_i[5];
      \nz.mem_1532_sv2v_reg  <= data_i[4];
      \nz.mem_1531_sv2v_reg  <= data_i[3];
      \nz.mem_1530_sv2v_reg  <= data_i[2];
      \nz.mem_1529_sv2v_reg  <= data_i[1];
      \nz.mem_1528_sv2v_reg  <= data_i[0];
    end 
    if(N981) begin
      \nz.mem_1527_sv2v_reg  <= data_i[7];
      \nz.mem_1526_sv2v_reg  <= data_i[6];
      \nz.mem_1525_sv2v_reg  <= data_i[5];
      \nz.mem_1524_sv2v_reg  <= data_i[4];
      \nz.mem_1523_sv2v_reg  <= data_i[3];
      \nz.mem_1522_sv2v_reg  <= data_i[2];
      \nz.mem_1521_sv2v_reg  <= data_i[1];
      \nz.mem_1520_sv2v_reg  <= data_i[0];
    end 
    if(N980) begin
      \nz.mem_1519_sv2v_reg  <= data_i[7];
      \nz.mem_1518_sv2v_reg  <= data_i[6];
      \nz.mem_1517_sv2v_reg  <= data_i[5];
      \nz.mem_1516_sv2v_reg  <= data_i[4];
      \nz.mem_1515_sv2v_reg  <= data_i[3];
      \nz.mem_1514_sv2v_reg  <= data_i[2];
      \nz.mem_1513_sv2v_reg  <= data_i[1];
      \nz.mem_1512_sv2v_reg  <= data_i[0];
    end 
    if(N979) begin
      \nz.mem_1511_sv2v_reg  <= data_i[7];
      \nz.mem_1510_sv2v_reg  <= data_i[6];
      \nz.mem_1509_sv2v_reg  <= data_i[5];
      \nz.mem_1508_sv2v_reg  <= data_i[4];
      \nz.mem_1507_sv2v_reg  <= data_i[3];
      \nz.mem_1506_sv2v_reg  <= data_i[2];
      \nz.mem_1505_sv2v_reg  <= data_i[1];
      \nz.mem_1504_sv2v_reg  <= data_i[0];
    end 
    if(N978) begin
      \nz.mem_1503_sv2v_reg  <= data_i[7];
      \nz.mem_1502_sv2v_reg  <= data_i[6];
      \nz.mem_1501_sv2v_reg  <= data_i[5];
      \nz.mem_1500_sv2v_reg  <= data_i[4];
      \nz.mem_1499_sv2v_reg  <= data_i[3];
      \nz.mem_1498_sv2v_reg  <= data_i[2];
      \nz.mem_1497_sv2v_reg  <= data_i[1];
      \nz.mem_1496_sv2v_reg  <= data_i[0];
    end 
    if(N977) begin
      \nz.mem_1495_sv2v_reg  <= data_i[7];
      \nz.mem_1494_sv2v_reg  <= data_i[6];
      \nz.mem_1493_sv2v_reg  <= data_i[5];
      \nz.mem_1492_sv2v_reg  <= data_i[4];
      \nz.mem_1491_sv2v_reg  <= data_i[3];
      \nz.mem_1490_sv2v_reg  <= data_i[2];
      \nz.mem_1489_sv2v_reg  <= data_i[1];
      \nz.mem_1488_sv2v_reg  <= data_i[0];
    end 
    if(N976) begin
      \nz.mem_1487_sv2v_reg  <= data_i[7];
      \nz.mem_1486_sv2v_reg  <= data_i[6];
      \nz.mem_1485_sv2v_reg  <= data_i[5];
      \nz.mem_1484_sv2v_reg  <= data_i[4];
      \nz.mem_1483_sv2v_reg  <= data_i[3];
      \nz.mem_1482_sv2v_reg  <= data_i[2];
      \nz.mem_1481_sv2v_reg  <= data_i[1];
      \nz.mem_1480_sv2v_reg  <= data_i[0];
    end 
    if(N975) begin
      \nz.mem_1479_sv2v_reg  <= data_i[7];
      \nz.mem_1478_sv2v_reg  <= data_i[6];
      \nz.mem_1477_sv2v_reg  <= data_i[5];
      \nz.mem_1476_sv2v_reg  <= data_i[4];
      \nz.mem_1475_sv2v_reg  <= data_i[3];
      \nz.mem_1474_sv2v_reg  <= data_i[2];
      \nz.mem_1473_sv2v_reg  <= data_i[1];
      \nz.mem_1472_sv2v_reg  <= data_i[0];
    end 
    if(N974) begin
      \nz.mem_1471_sv2v_reg  <= data_i[7];
      \nz.mem_1470_sv2v_reg  <= data_i[6];
      \nz.mem_1469_sv2v_reg  <= data_i[5];
      \nz.mem_1468_sv2v_reg  <= data_i[4];
      \nz.mem_1467_sv2v_reg  <= data_i[3];
      \nz.mem_1466_sv2v_reg  <= data_i[2];
      \nz.mem_1465_sv2v_reg  <= data_i[1];
      \nz.mem_1464_sv2v_reg  <= data_i[0];
    end 
    if(N973) begin
      \nz.mem_1463_sv2v_reg  <= data_i[7];
      \nz.mem_1462_sv2v_reg  <= data_i[6];
      \nz.mem_1461_sv2v_reg  <= data_i[5];
      \nz.mem_1460_sv2v_reg  <= data_i[4];
      \nz.mem_1459_sv2v_reg  <= data_i[3];
      \nz.mem_1458_sv2v_reg  <= data_i[2];
      \nz.mem_1457_sv2v_reg  <= data_i[1];
      \nz.mem_1456_sv2v_reg  <= data_i[0];
    end 
    if(N972) begin
      \nz.mem_1455_sv2v_reg  <= data_i[7];
      \nz.mem_1454_sv2v_reg  <= data_i[6];
      \nz.mem_1453_sv2v_reg  <= data_i[5];
      \nz.mem_1452_sv2v_reg  <= data_i[4];
      \nz.mem_1451_sv2v_reg  <= data_i[3];
      \nz.mem_1450_sv2v_reg  <= data_i[2];
      \nz.mem_1449_sv2v_reg  <= data_i[1];
      \nz.mem_1448_sv2v_reg  <= data_i[0];
    end 
    if(N971) begin
      \nz.mem_1447_sv2v_reg  <= data_i[7];
      \nz.mem_1446_sv2v_reg  <= data_i[6];
      \nz.mem_1445_sv2v_reg  <= data_i[5];
      \nz.mem_1444_sv2v_reg  <= data_i[4];
      \nz.mem_1443_sv2v_reg  <= data_i[3];
      \nz.mem_1442_sv2v_reg  <= data_i[2];
      \nz.mem_1441_sv2v_reg  <= data_i[1];
      \nz.mem_1440_sv2v_reg  <= data_i[0];
    end 
    if(N970) begin
      \nz.mem_1439_sv2v_reg  <= data_i[7];
      \nz.mem_1438_sv2v_reg  <= data_i[6];
      \nz.mem_1437_sv2v_reg  <= data_i[5];
      \nz.mem_1436_sv2v_reg  <= data_i[4];
      \nz.mem_1435_sv2v_reg  <= data_i[3];
      \nz.mem_1434_sv2v_reg  <= data_i[2];
      \nz.mem_1433_sv2v_reg  <= data_i[1];
      \nz.mem_1432_sv2v_reg  <= data_i[0];
    end 
    if(N969) begin
      \nz.mem_1431_sv2v_reg  <= data_i[7];
      \nz.mem_1430_sv2v_reg  <= data_i[6];
      \nz.mem_1429_sv2v_reg  <= data_i[5];
      \nz.mem_1428_sv2v_reg  <= data_i[4];
      \nz.mem_1427_sv2v_reg  <= data_i[3];
      \nz.mem_1426_sv2v_reg  <= data_i[2];
      \nz.mem_1425_sv2v_reg  <= data_i[1];
      \nz.mem_1424_sv2v_reg  <= data_i[0];
    end 
    if(N968) begin
      \nz.mem_1423_sv2v_reg  <= data_i[7];
      \nz.mem_1422_sv2v_reg  <= data_i[6];
      \nz.mem_1421_sv2v_reg  <= data_i[5];
      \nz.mem_1420_sv2v_reg  <= data_i[4];
      \nz.mem_1419_sv2v_reg  <= data_i[3];
      \nz.mem_1418_sv2v_reg  <= data_i[2];
      \nz.mem_1417_sv2v_reg  <= data_i[1];
      \nz.mem_1416_sv2v_reg  <= data_i[0];
    end 
    if(N967) begin
      \nz.mem_1415_sv2v_reg  <= data_i[7];
      \nz.mem_1414_sv2v_reg  <= data_i[6];
      \nz.mem_1413_sv2v_reg  <= data_i[5];
      \nz.mem_1412_sv2v_reg  <= data_i[4];
      \nz.mem_1411_sv2v_reg  <= data_i[3];
      \nz.mem_1410_sv2v_reg  <= data_i[2];
      \nz.mem_1409_sv2v_reg  <= data_i[1];
      \nz.mem_1408_sv2v_reg  <= data_i[0];
    end 
    if(N966) begin
      \nz.mem_1407_sv2v_reg  <= data_i[7];
      \nz.mem_1406_sv2v_reg  <= data_i[6];
      \nz.mem_1405_sv2v_reg  <= data_i[5];
      \nz.mem_1404_sv2v_reg  <= data_i[4];
      \nz.mem_1403_sv2v_reg  <= data_i[3];
      \nz.mem_1402_sv2v_reg  <= data_i[2];
      \nz.mem_1401_sv2v_reg  <= data_i[1];
      \nz.mem_1400_sv2v_reg  <= data_i[0];
    end 
    if(N965) begin
      \nz.mem_1399_sv2v_reg  <= data_i[7];
      \nz.mem_1398_sv2v_reg  <= data_i[6];
      \nz.mem_1397_sv2v_reg  <= data_i[5];
      \nz.mem_1396_sv2v_reg  <= data_i[4];
      \nz.mem_1395_sv2v_reg  <= data_i[3];
      \nz.mem_1394_sv2v_reg  <= data_i[2];
      \nz.mem_1393_sv2v_reg  <= data_i[1];
      \nz.mem_1392_sv2v_reg  <= data_i[0];
    end 
    if(N964) begin
      \nz.mem_1391_sv2v_reg  <= data_i[7];
      \nz.mem_1390_sv2v_reg  <= data_i[6];
      \nz.mem_1389_sv2v_reg  <= data_i[5];
      \nz.mem_1388_sv2v_reg  <= data_i[4];
      \nz.mem_1387_sv2v_reg  <= data_i[3];
      \nz.mem_1386_sv2v_reg  <= data_i[2];
      \nz.mem_1385_sv2v_reg  <= data_i[1];
      \nz.mem_1384_sv2v_reg  <= data_i[0];
    end 
    if(N963) begin
      \nz.mem_1383_sv2v_reg  <= data_i[7];
      \nz.mem_1382_sv2v_reg  <= data_i[6];
      \nz.mem_1381_sv2v_reg  <= data_i[5];
      \nz.mem_1380_sv2v_reg  <= data_i[4];
      \nz.mem_1379_sv2v_reg  <= data_i[3];
      \nz.mem_1378_sv2v_reg  <= data_i[2];
      \nz.mem_1377_sv2v_reg  <= data_i[1];
      \nz.mem_1376_sv2v_reg  <= data_i[0];
    end 
    if(N962) begin
      \nz.mem_1375_sv2v_reg  <= data_i[7];
      \nz.mem_1374_sv2v_reg  <= data_i[6];
      \nz.mem_1373_sv2v_reg  <= data_i[5];
      \nz.mem_1372_sv2v_reg  <= data_i[4];
      \nz.mem_1371_sv2v_reg  <= data_i[3];
      \nz.mem_1370_sv2v_reg  <= data_i[2];
      \nz.mem_1369_sv2v_reg  <= data_i[1];
      \nz.mem_1368_sv2v_reg  <= data_i[0];
    end 
    if(N961) begin
      \nz.mem_1367_sv2v_reg  <= data_i[7];
      \nz.mem_1366_sv2v_reg  <= data_i[6];
      \nz.mem_1365_sv2v_reg  <= data_i[5];
      \nz.mem_1364_sv2v_reg  <= data_i[4];
      \nz.mem_1363_sv2v_reg  <= data_i[3];
      \nz.mem_1362_sv2v_reg  <= data_i[2];
      \nz.mem_1361_sv2v_reg  <= data_i[1];
      \nz.mem_1360_sv2v_reg  <= data_i[0];
    end 
    if(N960) begin
      \nz.mem_1359_sv2v_reg  <= data_i[7];
      \nz.mem_1358_sv2v_reg  <= data_i[6];
      \nz.mem_1357_sv2v_reg  <= data_i[5];
      \nz.mem_1356_sv2v_reg  <= data_i[4];
      \nz.mem_1355_sv2v_reg  <= data_i[3];
      \nz.mem_1354_sv2v_reg  <= data_i[2];
      \nz.mem_1353_sv2v_reg  <= data_i[1];
      \nz.mem_1352_sv2v_reg  <= data_i[0];
    end 
    if(N959) begin
      \nz.mem_1351_sv2v_reg  <= data_i[7];
      \nz.mem_1350_sv2v_reg  <= data_i[6];
      \nz.mem_1349_sv2v_reg  <= data_i[5];
      \nz.mem_1348_sv2v_reg  <= data_i[4];
      \nz.mem_1347_sv2v_reg  <= data_i[3];
      \nz.mem_1346_sv2v_reg  <= data_i[2];
      \nz.mem_1345_sv2v_reg  <= data_i[1];
      \nz.mem_1344_sv2v_reg  <= data_i[0];
    end 
    if(N958) begin
      \nz.mem_1343_sv2v_reg  <= data_i[7];
      \nz.mem_1342_sv2v_reg  <= data_i[6];
      \nz.mem_1341_sv2v_reg  <= data_i[5];
      \nz.mem_1340_sv2v_reg  <= data_i[4];
      \nz.mem_1339_sv2v_reg  <= data_i[3];
      \nz.mem_1338_sv2v_reg  <= data_i[2];
      \nz.mem_1337_sv2v_reg  <= data_i[1];
      \nz.mem_1336_sv2v_reg  <= data_i[0];
    end 
    if(N957) begin
      \nz.mem_1335_sv2v_reg  <= data_i[7];
      \nz.mem_1334_sv2v_reg  <= data_i[6];
      \nz.mem_1333_sv2v_reg  <= data_i[5];
      \nz.mem_1332_sv2v_reg  <= data_i[4];
      \nz.mem_1331_sv2v_reg  <= data_i[3];
      \nz.mem_1330_sv2v_reg  <= data_i[2];
      \nz.mem_1329_sv2v_reg  <= data_i[1];
      \nz.mem_1328_sv2v_reg  <= data_i[0];
    end 
    if(N956) begin
      \nz.mem_1327_sv2v_reg  <= data_i[7];
      \nz.mem_1326_sv2v_reg  <= data_i[6];
      \nz.mem_1325_sv2v_reg  <= data_i[5];
      \nz.mem_1324_sv2v_reg  <= data_i[4];
      \nz.mem_1323_sv2v_reg  <= data_i[3];
      \nz.mem_1322_sv2v_reg  <= data_i[2];
      \nz.mem_1321_sv2v_reg  <= data_i[1];
      \nz.mem_1320_sv2v_reg  <= data_i[0];
    end 
    if(N955) begin
      \nz.mem_1319_sv2v_reg  <= data_i[7];
      \nz.mem_1318_sv2v_reg  <= data_i[6];
      \nz.mem_1317_sv2v_reg  <= data_i[5];
      \nz.mem_1316_sv2v_reg  <= data_i[4];
      \nz.mem_1315_sv2v_reg  <= data_i[3];
      \nz.mem_1314_sv2v_reg  <= data_i[2];
      \nz.mem_1313_sv2v_reg  <= data_i[1];
      \nz.mem_1312_sv2v_reg  <= data_i[0];
    end 
    if(N954) begin
      \nz.mem_1311_sv2v_reg  <= data_i[7];
      \nz.mem_1310_sv2v_reg  <= data_i[6];
      \nz.mem_1309_sv2v_reg  <= data_i[5];
      \nz.mem_1308_sv2v_reg  <= data_i[4];
      \nz.mem_1307_sv2v_reg  <= data_i[3];
      \nz.mem_1306_sv2v_reg  <= data_i[2];
      \nz.mem_1305_sv2v_reg  <= data_i[1];
      \nz.mem_1304_sv2v_reg  <= data_i[0];
    end 
    if(N953) begin
      \nz.mem_1303_sv2v_reg  <= data_i[7];
      \nz.mem_1302_sv2v_reg  <= data_i[6];
      \nz.mem_1301_sv2v_reg  <= data_i[5];
      \nz.mem_1300_sv2v_reg  <= data_i[4];
      \nz.mem_1299_sv2v_reg  <= data_i[3];
      \nz.mem_1298_sv2v_reg  <= data_i[2];
      \nz.mem_1297_sv2v_reg  <= data_i[1];
      \nz.mem_1296_sv2v_reg  <= data_i[0];
    end 
    if(N952) begin
      \nz.mem_1295_sv2v_reg  <= data_i[7];
      \nz.mem_1294_sv2v_reg  <= data_i[6];
      \nz.mem_1293_sv2v_reg  <= data_i[5];
      \nz.mem_1292_sv2v_reg  <= data_i[4];
      \nz.mem_1291_sv2v_reg  <= data_i[3];
      \nz.mem_1290_sv2v_reg  <= data_i[2];
      \nz.mem_1289_sv2v_reg  <= data_i[1];
      \nz.mem_1288_sv2v_reg  <= data_i[0];
    end 
    if(N951) begin
      \nz.mem_1287_sv2v_reg  <= data_i[7];
      \nz.mem_1286_sv2v_reg  <= data_i[6];
      \nz.mem_1285_sv2v_reg  <= data_i[5];
      \nz.mem_1284_sv2v_reg  <= data_i[4];
      \nz.mem_1283_sv2v_reg  <= data_i[3];
      \nz.mem_1282_sv2v_reg  <= data_i[2];
      \nz.mem_1281_sv2v_reg  <= data_i[1];
      \nz.mem_1280_sv2v_reg  <= data_i[0];
    end 
    if(N950) begin
      \nz.mem_1279_sv2v_reg  <= data_i[7];
      \nz.mem_1278_sv2v_reg  <= data_i[6];
      \nz.mem_1277_sv2v_reg  <= data_i[5];
      \nz.mem_1276_sv2v_reg  <= data_i[4];
      \nz.mem_1275_sv2v_reg  <= data_i[3];
      \nz.mem_1274_sv2v_reg  <= data_i[2];
      \nz.mem_1273_sv2v_reg  <= data_i[1];
      \nz.mem_1272_sv2v_reg  <= data_i[0];
    end 
    if(N949) begin
      \nz.mem_1271_sv2v_reg  <= data_i[7];
      \nz.mem_1270_sv2v_reg  <= data_i[6];
      \nz.mem_1269_sv2v_reg  <= data_i[5];
      \nz.mem_1268_sv2v_reg  <= data_i[4];
      \nz.mem_1267_sv2v_reg  <= data_i[3];
      \nz.mem_1266_sv2v_reg  <= data_i[2];
      \nz.mem_1265_sv2v_reg  <= data_i[1];
      \nz.mem_1264_sv2v_reg  <= data_i[0];
    end 
    if(N948) begin
      \nz.mem_1263_sv2v_reg  <= data_i[7];
      \nz.mem_1262_sv2v_reg  <= data_i[6];
      \nz.mem_1261_sv2v_reg  <= data_i[5];
      \nz.mem_1260_sv2v_reg  <= data_i[4];
      \nz.mem_1259_sv2v_reg  <= data_i[3];
      \nz.mem_1258_sv2v_reg  <= data_i[2];
      \nz.mem_1257_sv2v_reg  <= data_i[1];
      \nz.mem_1256_sv2v_reg  <= data_i[0];
    end 
    if(N947) begin
      \nz.mem_1255_sv2v_reg  <= data_i[7];
      \nz.mem_1254_sv2v_reg  <= data_i[6];
      \nz.mem_1253_sv2v_reg  <= data_i[5];
      \nz.mem_1252_sv2v_reg  <= data_i[4];
      \nz.mem_1251_sv2v_reg  <= data_i[3];
      \nz.mem_1250_sv2v_reg  <= data_i[2];
      \nz.mem_1249_sv2v_reg  <= data_i[1];
      \nz.mem_1248_sv2v_reg  <= data_i[0];
    end 
    if(N946) begin
      \nz.mem_1247_sv2v_reg  <= data_i[7];
      \nz.mem_1246_sv2v_reg  <= data_i[6];
      \nz.mem_1245_sv2v_reg  <= data_i[5];
      \nz.mem_1244_sv2v_reg  <= data_i[4];
      \nz.mem_1243_sv2v_reg  <= data_i[3];
      \nz.mem_1242_sv2v_reg  <= data_i[2];
      \nz.mem_1241_sv2v_reg  <= data_i[1];
      \nz.mem_1240_sv2v_reg  <= data_i[0];
    end 
    if(N945) begin
      \nz.mem_1239_sv2v_reg  <= data_i[7];
      \nz.mem_1238_sv2v_reg  <= data_i[6];
      \nz.mem_1237_sv2v_reg  <= data_i[5];
      \nz.mem_1236_sv2v_reg  <= data_i[4];
      \nz.mem_1235_sv2v_reg  <= data_i[3];
      \nz.mem_1234_sv2v_reg  <= data_i[2];
      \nz.mem_1233_sv2v_reg  <= data_i[1];
      \nz.mem_1232_sv2v_reg  <= data_i[0];
    end 
    if(N944) begin
      \nz.mem_1231_sv2v_reg  <= data_i[7];
      \nz.mem_1230_sv2v_reg  <= data_i[6];
      \nz.mem_1229_sv2v_reg  <= data_i[5];
      \nz.mem_1228_sv2v_reg  <= data_i[4];
      \nz.mem_1227_sv2v_reg  <= data_i[3];
      \nz.mem_1226_sv2v_reg  <= data_i[2];
      \nz.mem_1225_sv2v_reg  <= data_i[1];
      \nz.mem_1224_sv2v_reg  <= data_i[0];
    end 
    if(N943) begin
      \nz.mem_1223_sv2v_reg  <= data_i[7];
      \nz.mem_1222_sv2v_reg  <= data_i[6];
      \nz.mem_1221_sv2v_reg  <= data_i[5];
      \nz.mem_1220_sv2v_reg  <= data_i[4];
      \nz.mem_1219_sv2v_reg  <= data_i[3];
      \nz.mem_1218_sv2v_reg  <= data_i[2];
      \nz.mem_1217_sv2v_reg  <= data_i[1];
      \nz.mem_1216_sv2v_reg  <= data_i[0];
    end 
    if(N942) begin
      \nz.mem_1215_sv2v_reg  <= data_i[7];
      \nz.mem_1214_sv2v_reg  <= data_i[6];
      \nz.mem_1213_sv2v_reg  <= data_i[5];
      \nz.mem_1212_sv2v_reg  <= data_i[4];
      \nz.mem_1211_sv2v_reg  <= data_i[3];
      \nz.mem_1210_sv2v_reg  <= data_i[2];
      \nz.mem_1209_sv2v_reg  <= data_i[1];
      \nz.mem_1208_sv2v_reg  <= data_i[0];
    end 
    if(N941) begin
      \nz.mem_1207_sv2v_reg  <= data_i[7];
      \nz.mem_1206_sv2v_reg  <= data_i[6];
      \nz.mem_1205_sv2v_reg  <= data_i[5];
      \nz.mem_1204_sv2v_reg  <= data_i[4];
      \nz.mem_1203_sv2v_reg  <= data_i[3];
      \nz.mem_1202_sv2v_reg  <= data_i[2];
      \nz.mem_1201_sv2v_reg  <= data_i[1];
      \nz.mem_1200_sv2v_reg  <= data_i[0];
    end 
    if(N940) begin
      \nz.mem_1199_sv2v_reg  <= data_i[7];
      \nz.mem_1198_sv2v_reg  <= data_i[6];
      \nz.mem_1197_sv2v_reg  <= data_i[5];
      \nz.mem_1196_sv2v_reg  <= data_i[4];
      \nz.mem_1195_sv2v_reg  <= data_i[3];
      \nz.mem_1194_sv2v_reg  <= data_i[2];
      \nz.mem_1193_sv2v_reg  <= data_i[1];
      \nz.mem_1192_sv2v_reg  <= data_i[0];
    end 
    if(N939) begin
      \nz.mem_1191_sv2v_reg  <= data_i[7];
      \nz.mem_1190_sv2v_reg  <= data_i[6];
      \nz.mem_1189_sv2v_reg  <= data_i[5];
      \nz.mem_1188_sv2v_reg  <= data_i[4];
      \nz.mem_1187_sv2v_reg  <= data_i[3];
      \nz.mem_1186_sv2v_reg  <= data_i[2];
      \nz.mem_1185_sv2v_reg  <= data_i[1];
      \nz.mem_1184_sv2v_reg  <= data_i[0];
    end 
    if(N938) begin
      \nz.mem_1183_sv2v_reg  <= data_i[7];
      \nz.mem_1182_sv2v_reg  <= data_i[6];
      \nz.mem_1181_sv2v_reg  <= data_i[5];
      \nz.mem_1180_sv2v_reg  <= data_i[4];
      \nz.mem_1179_sv2v_reg  <= data_i[3];
      \nz.mem_1178_sv2v_reg  <= data_i[2];
      \nz.mem_1177_sv2v_reg  <= data_i[1];
      \nz.mem_1176_sv2v_reg  <= data_i[0];
    end 
    if(N937) begin
      \nz.mem_1175_sv2v_reg  <= data_i[7];
      \nz.mem_1174_sv2v_reg  <= data_i[6];
      \nz.mem_1173_sv2v_reg  <= data_i[5];
      \nz.mem_1172_sv2v_reg  <= data_i[4];
      \nz.mem_1171_sv2v_reg  <= data_i[3];
      \nz.mem_1170_sv2v_reg  <= data_i[2];
      \nz.mem_1169_sv2v_reg  <= data_i[1];
      \nz.mem_1168_sv2v_reg  <= data_i[0];
    end 
    if(N936) begin
      \nz.mem_1167_sv2v_reg  <= data_i[7];
      \nz.mem_1166_sv2v_reg  <= data_i[6];
      \nz.mem_1165_sv2v_reg  <= data_i[5];
      \nz.mem_1164_sv2v_reg  <= data_i[4];
      \nz.mem_1163_sv2v_reg  <= data_i[3];
      \nz.mem_1162_sv2v_reg  <= data_i[2];
      \nz.mem_1161_sv2v_reg  <= data_i[1];
      \nz.mem_1160_sv2v_reg  <= data_i[0];
    end 
    if(N935) begin
      \nz.mem_1159_sv2v_reg  <= data_i[7];
      \nz.mem_1158_sv2v_reg  <= data_i[6];
      \nz.mem_1157_sv2v_reg  <= data_i[5];
      \nz.mem_1156_sv2v_reg  <= data_i[4];
      \nz.mem_1155_sv2v_reg  <= data_i[3];
      \nz.mem_1154_sv2v_reg  <= data_i[2];
      \nz.mem_1153_sv2v_reg  <= data_i[1];
      \nz.mem_1152_sv2v_reg  <= data_i[0];
    end 
    if(N934) begin
      \nz.mem_1151_sv2v_reg  <= data_i[7];
      \nz.mem_1150_sv2v_reg  <= data_i[6];
      \nz.mem_1149_sv2v_reg  <= data_i[5];
      \nz.mem_1148_sv2v_reg  <= data_i[4];
      \nz.mem_1147_sv2v_reg  <= data_i[3];
      \nz.mem_1146_sv2v_reg  <= data_i[2];
      \nz.mem_1145_sv2v_reg  <= data_i[1];
      \nz.mem_1144_sv2v_reg  <= data_i[0];
    end 
    if(N933) begin
      \nz.mem_1143_sv2v_reg  <= data_i[7];
      \nz.mem_1142_sv2v_reg  <= data_i[6];
      \nz.mem_1141_sv2v_reg  <= data_i[5];
      \nz.mem_1140_sv2v_reg  <= data_i[4];
      \nz.mem_1139_sv2v_reg  <= data_i[3];
      \nz.mem_1138_sv2v_reg  <= data_i[2];
      \nz.mem_1137_sv2v_reg  <= data_i[1];
      \nz.mem_1136_sv2v_reg  <= data_i[0];
    end 
    if(N932) begin
      \nz.mem_1135_sv2v_reg  <= data_i[7];
      \nz.mem_1134_sv2v_reg  <= data_i[6];
      \nz.mem_1133_sv2v_reg  <= data_i[5];
      \nz.mem_1132_sv2v_reg  <= data_i[4];
      \nz.mem_1131_sv2v_reg  <= data_i[3];
      \nz.mem_1130_sv2v_reg  <= data_i[2];
      \nz.mem_1129_sv2v_reg  <= data_i[1];
      \nz.mem_1128_sv2v_reg  <= data_i[0];
    end 
    if(N931) begin
      \nz.mem_1127_sv2v_reg  <= data_i[7];
      \nz.mem_1126_sv2v_reg  <= data_i[6];
      \nz.mem_1125_sv2v_reg  <= data_i[5];
      \nz.mem_1124_sv2v_reg  <= data_i[4];
      \nz.mem_1123_sv2v_reg  <= data_i[3];
      \nz.mem_1122_sv2v_reg  <= data_i[2];
      \nz.mem_1121_sv2v_reg  <= data_i[1];
      \nz.mem_1120_sv2v_reg  <= data_i[0];
    end 
    if(N930) begin
      \nz.mem_1119_sv2v_reg  <= data_i[7];
      \nz.mem_1118_sv2v_reg  <= data_i[6];
      \nz.mem_1117_sv2v_reg  <= data_i[5];
      \nz.mem_1116_sv2v_reg  <= data_i[4];
      \nz.mem_1115_sv2v_reg  <= data_i[3];
      \nz.mem_1114_sv2v_reg  <= data_i[2];
      \nz.mem_1113_sv2v_reg  <= data_i[1];
      \nz.mem_1112_sv2v_reg  <= data_i[0];
    end 
    if(N929) begin
      \nz.mem_1111_sv2v_reg  <= data_i[7];
      \nz.mem_1110_sv2v_reg  <= data_i[6];
      \nz.mem_1109_sv2v_reg  <= data_i[5];
      \nz.mem_1108_sv2v_reg  <= data_i[4];
      \nz.mem_1107_sv2v_reg  <= data_i[3];
      \nz.mem_1106_sv2v_reg  <= data_i[2];
      \nz.mem_1105_sv2v_reg  <= data_i[1];
      \nz.mem_1104_sv2v_reg  <= data_i[0];
    end 
    if(N928) begin
      \nz.mem_1103_sv2v_reg  <= data_i[7];
      \nz.mem_1102_sv2v_reg  <= data_i[6];
      \nz.mem_1101_sv2v_reg  <= data_i[5];
      \nz.mem_1100_sv2v_reg  <= data_i[4];
      \nz.mem_1099_sv2v_reg  <= data_i[3];
      \nz.mem_1098_sv2v_reg  <= data_i[2];
      \nz.mem_1097_sv2v_reg  <= data_i[1];
      \nz.mem_1096_sv2v_reg  <= data_i[0];
    end 
    if(N927) begin
      \nz.mem_1095_sv2v_reg  <= data_i[7];
      \nz.mem_1094_sv2v_reg  <= data_i[6];
      \nz.mem_1093_sv2v_reg  <= data_i[5];
      \nz.mem_1092_sv2v_reg  <= data_i[4];
      \nz.mem_1091_sv2v_reg  <= data_i[3];
      \nz.mem_1090_sv2v_reg  <= data_i[2];
      \nz.mem_1089_sv2v_reg  <= data_i[1];
      \nz.mem_1088_sv2v_reg  <= data_i[0];
    end 
    if(N926) begin
      \nz.mem_1087_sv2v_reg  <= data_i[7];
      \nz.mem_1086_sv2v_reg  <= data_i[6];
      \nz.mem_1085_sv2v_reg  <= data_i[5];
      \nz.mem_1084_sv2v_reg  <= data_i[4];
      \nz.mem_1083_sv2v_reg  <= data_i[3];
      \nz.mem_1082_sv2v_reg  <= data_i[2];
      \nz.mem_1081_sv2v_reg  <= data_i[1];
      \nz.mem_1080_sv2v_reg  <= data_i[0];
    end 
    if(N925) begin
      \nz.mem_1079_sv2v_reg  <= data_i[7];
      \nz.mem_1078_sv2v_reg  <= data_i[6];
      \nz.mem_1077_sv2v_reg  <= data_i[5];
      \nz.mem_1076_sv2v_reg  <= data_i[4];
      \nz.mem_1075_sv2v_reg  <= data_i[3];
      \nz.mem_1074_sv2v_reg  <= data_i[2];
      \nz.mem_1073_sv2v_reg  <= data_i[1];
      \nz.mem_1072_sv2v_reg  <= data_i[0];
    end 
    if(N924) begin
      \nz.mem_1071_sv2v_reg  <= data_i[7];
      \nz.mem_1070_sv2v_reg  <= data_i[6];
      \nz.mem_1069_sv2v_reg  <= data_i[5];
      \nz.mem_1068_sv2v_reg  <= data_i[4];
      \nz.mem_1067_sv2v_reg  <= data_i[3];
      \nz.mem_1066_sv2v_reg  <= data_i[2];
      \nz.mem_1065_sv2v_reg  <= data_i[1];
      \nz.mem_1064_sv2v_reg  <= data_i[0];
    end 
    if(N923) begin
      \nz.mem_1063_sv2v_reg  <= data_i[7];
      \nz.mem_1062_sv2v_reg  <= data_i[6];
      \nz.mem_1061_sv2v_reg  <= data_i[5];
      \nz.mem_1060_sv2v_reg  <= data_i[4];
      \nz.mem_1059_sv2v_reg  <= data_i[3];
      \nz.mem_1058_sv2v_reg  <= data_i[2];
      \nz.mem_1057_sv2v_reg  <= data_i[1];
      \nz.mem_1056_sv2v_reg  <= data_i[0];
    end 
    if(N922) begin
      \nz.mem_1055_sv2v_reg  <= data_i[7];
      \nz.mem_1054_sv2v_reg  <= data_i[6];
      \nz.mem_1053_sv2v_reg  <= data_i[5];
      \nz.mem_1052_sv2v_reg  <= data_i[4];
      \nz.mem_1051_sv2v_reg  <= data_i[3];
      \nz.mem_1050_sv2v_reg  <= data_i[2];
      \nz.mem_1049_sv2v_reg  <= data_i[1];
      \nz.mem_1048_sv2v_reg  <= data_i[0];
    end 
    if(N921) begin
      \nz.mem_1047_sv2v_reg  <= data_i[7];
      \nz.mem_1046_sv2v_reg  <= data_i[6];
      \nz.mem_1045_sv2v_reg  <= data_i[5];
      \nz.mem_1044_sv2v_reg  <= data_i[4];
      \nz.mem_1043_sv2v_reg  <= data_i[3];
      \nz.mem_1042_sv2v_reg  <= data_i[2];
      \nz.mem_1041_sv2v_reg  <= data_i[1];
      \nz.mem_1040_sv2v_reg  <= data_i[0];
    end 
    if(N920) begin
      \nz.mem_1039_sv2v_reg  <= data_i[7];
      \nz.mem_1038_sv2v_reg  <= data_i[6];
      \nz.mem_1037_sv2v_reg  <= data_i[5];
      \nz.mem_1036_sv2v_reg  <= data_i[4];
      \nz.mem_1035_sv2v_reg  <= data_i[3];
      \nz.mem_1034_sv2v_reg  <= data_i[2];
      \nz.mem_1033_sv2v_reg  <= data_i[1];
      \nz.mem_1032_sv2v_reg  <= data_i[0];
    end 
    if(N919) begin
      \nz.mem_1031_sv2v_reg  <= data_i[7];
      \nz.mem_1030_sv2v_reg  <= data_i[6];
      \nz.mem_1029_sv2v_reg  <= data_i[5];
      \nz.mem_1028_sv2v_reg  <= data_i[4];
      \nz.mem_1027_sv2v_reg  <= data_i[3];
      \nz.mem_1026_sv2v_reg  <= data_i[2];
      \nz.mem_1025_sv2v_reg  <= data_i[1];
      \nz.mem_1024_sv2v_reg  <= data_i[0];
    end 
    if(N918) begin
      \nz.mem_1023_sv2v_reg  <= data_i[7];
      \nz.mem_1022_sv2v_reg  <= data_i[6];
      \nz.mem_1021_sv2v_reg  <= data_i[5];
      \nz.mem_1020_sv2v_reg  <= data_i[4];
      \nz.mem_1019_sv2v_reg  <= data_i[3];
      \nz.mem_1018_sv2v_reg  <= data_i[2];
      \nz.mem_1017_sv2v_reg  <= data_i[1];
      \nz.mem_1016_sv2v_reg  <= data_i[0];
    end 
    if(N917) begin
      \nz.mem_1015_sv2v_reg  <= data_i[7];
      \nz.mem_1014_sv2v_reg  <= data_i[6];
      \nz.mem_1013_sv2v_reg  <= data_i[5];
      \nz.mem_1012_sv2v_reg  <= data_i[4];
      \nz.mem_1011_sv2v_reg  <= data_i[3];
      \nz.mem_1010_sv2v_reg  <= data_i[2];
      \nz.mem_1009_sv2v_reg  <= data_i[1];
      \nz.mem_1008_sv2v_reg  <= data_i[0];
    end 
    if(N916) begin
      \nz.mem_1007_sv2v_reg  <= data_i[7];
      \nz.mem_1006_sv2v_reg  <= data_i[6];
      \nz.mem_1005_sv2v_reg  <= data_i[5];
      \nz.mem_1004_sv2v_reg  <= data_i[4];
      \nz.mem_1003_sv2v_reg  <= data_i[3];
      \nz.mem_1002_sv2v_reg  <= data_i[2];
      \nz.mem_1001_sv2v_reg  <= data_i[1];
      \nz.mem_1000_sv2v_reg  <= data_i[0];
    end 
    if(N915) begin
      \nz.mem_999_sv2v_reg  <= data_i[7];
      \nz.mem_998_sv2v_reg  <= data_i[6];
      \nz.mem_997_sv2v_reg  <= data_i[5];
      \nz.mem_996_sv2v_reg  <= data_i[4];
      \nz.mem_995_sv2v_reg  <= data_i[3];
      \nz.mem_994_sv2v_reg  <= data_i[2];
      \nz.mem_993_sv2v_reg  <= data_i[1];
      \nz.mem_992_sv2v_reg  <= data_i[0];
    end 
    if(N914) begin
      \nz.mem_991_sv2v_reg  <= data_i[7];
      \nz.mem_990_sv2v_reg  <= data_i[6];
      \nz.mem_989_sv2v_reg  <= data_i[5];
      \nz.mem_988_sv2v_reg  <= data_i[4];
      \nz.mem_987_sv2v_reg  <= data_i[3];
      \nz.mem_986_sv2v_reg  <= data_i[2];
      \nz.mem_985_sv2v_reg  <= data_i[1];
      \nz.mem_984_sv2v_reg  <= data_i[0];
    end 
    if(N913) begin
      \nz.mem_983_sv2v_reg  <= data_i[7];
      \nz.mem_982_sv2v_reg  <= data_i[6];
      \nz.mem_981_sv2v_reg  <= data_i[5];
      \nz.mem_980_sv2v_reg  <= data_i[4];
      \nz.mem_979_sv2v_reg  <= data_i[3];
      \nz.mem_978_sv2v_reg  <= data_i[2];
      \nz.mem_977_sv2v_reg  <= data_i[1];
      \nz.mem_976_sv2v_reg  <= data_i[0];
    end 
    if(N912) begin
      \nz.mem_975_sv2v_reg  <= data_i[7];
      \nz.mem_974_sv2v_reg  <= data_i[6];
      \nz.mem_973_sv2v_reg  <= data_i[5];
      \nz.mem_972_sv2v_reg  <= data_i[4];
      \nz.mem_971_sv2v_reg  <= data_i[3];
      \nz.mem_970_sv2v_reg  <= data_i[2];
      \nz.mem_969_sv2v_reg  <= data_i[1];
      \nz.mem_968_sv2v_reg  <= data_i[0];
    end 
    if(N911) begin
      \nz.mem_967_sv2v_reg  <= data_i[7];
      \nz.mem_966_sv2v_reg  <= data_i[6];
      \nz.mem_965_sv2v_reg  <= data_i[5];
      \nz.mem_964_sv2v_reg  <= data_i[4];
      \nz.mem_963_sv2v_reg  <= data_i[3];
      \nz.mem_962_sv2v_reg  <= data_i[2];
      \nz.mem_961_sv2v_reg  <= data_i[1];
      \nz.mem_960_sv2v_reg  <= data_i[0];
    end 
    if(N910) begin
      \nz.mem_959_sv2v_reg  <= data_i[7];
      \nz.mem_958_sv2v_reg  <= data_i[6];
      \nz.mem_957_sv2v_reg  <= data_i[5];
      \nz.mem_956_sv2v_reg  <= data_i[4];
      \nz.mem_955_sv2v_reg  <= data_i[3];
      \nz.mem_954_sv2v_reg  <= data_i[2];
      \nz.mem_953_sv2v_reg  <= data_i[1];
      \nz.mem_952_sv2v_reg  <= data_i[0];
    end 
    if(N909) begin
      \nz.mem_951_sv2v_reg  <= data_i[7];
      \nz.mem_950_sv2v_reg  <= data_i[6];
      \nz.mem_949_sv2v_reg  <= data_i[5];
      \nz.mem_948_sv2v_reg  <= data_i[4];
      \nz.mem_947_sv2v_reg  <= data_i[3];
      \nz.mem_946_sv2v_reg  <= data_i[2];
      \nz.mem_945_sv2v_reg  <= data_i[1];
      \nz.mem_944_sv2v_reg  <= data_i[0];
    end 
    if(N908) begin
      \nz.mem_943_sv2v_reg  <= data_i[7];
      \nz.mem_942_sv2v_reg  <= data_i[6];
      \nz.mem_941_sv2v_reg  <= data_i[5];
      \nz.mem_940_sv2v_reg  <= data_i[4];
      \nz.mem_939_sv2v_reg  <= data_i[3];
      \nz.mem_938_sv2v_reg  <= data_i[2];
      \nz.mem_937_sv2v_reg  <= data_i[1];
      \nz.mem_936_sv2v_reg  <= data_i[0];
    end 
    if(N907) begin
      \nz.mem_935_sv2v_reg  <= data_i[7];
      \nz.mem_934_sv2v_reg  <= data_i[6];
      \nz.mem_933_sv2v_reg  <= data_i[5];
      \nz.mem_932_sv2v_reg  <= data_i[4];
      \nz.mem_931_sv2v_reg  <= data_i[3];
      \nz.mem_930_sv2v_reg  <= data_i[2];
      \nz.mem_929_sv2v_reg  <= data_i[1];
      \nz.mem_928_sv2v_reg  <= data_i[0];
    end 
    if(N906) begin
      \nz.mem_927_sv2v_reg  <= data_i[7];
      \nz.mem_926_sv2v_reg  <= data_i[6];
      \nz.mem_925_sv2v_reg  <= data_i[5];
      \nz.mem_924_sv2v_reg  <= data_i[4];
      \nz.mem_923_sv2v_reg  <= data_i[3];
      \nz.mem_922_sv2v_reg  <= data_i[2];
      \nz.mem_921_sv2v_reg  <= data_i[1];
      \nz.mem_920_sv2v_reg  <= data_i[0];
    end 
    if(N905) begin
      \nz.mem_919_sv2v_reg  <= data_i[7];
      \nz.mem_918_sv2v_reg  <= data_i[6];
      \nz.mem_917_sv2v_reg  <= data_i[5];
      \nz.mem_916_sv2v_reg  <= data_i[4];
      \nz.mem_915_sv2v_reg  <= data_i[3];
      \nz.mem_914_sv2v_reg  <= data_i[2];
      \nz.mem_913_sv2v_reg  <= data_i[1];
      \nz.mem_912_sv2v_reg  <= data_i[0];
    end 
    if(N904) begin
      \nz.mem_911_sv2v_reg  <= data_i[7];
      \nz.mem_910_sv2v_reg  <= data_i[6];
      \nz.mem_909_sv2v_reg  <= data_i[5];
      \nz.mem_908_sv2v_reg  <= data_i[4];
      \nz.mem_907_sv2v_reg  <= data_i[3];
      \nz.mem_906_sv2v_reg  <= data_i[2];
      \nz.mem_905_sv2v_reg  <= data_i[1];
      \nz.mem_904_sv2v_reg  <= data_i[0];
    end 
    if(N903) begin
      \nz.mem_903_sv2v_reg  <= data_i[7];
      \nz.mem_902_sv2v_reg  <= data_i[6];
      \nz.mem_901_sv2v_reg  <= data_i[5];
      \nz.mem_900_sv2v_reg  <= data_i[4];
      \nz.mem_899_sv2v_reg  <= data_i[3];
      \nz.mem_898_sv2v_reg  <= data_i[2];
      \nz.mem_897_sv2v_reg  <= data_i[1];
      \nz.mem_896_sv2v_reg  <= data_i[0];
    end 
    if(N902) begin
      \nz.mem_895_sv2v_reg  <= data_i[7];
      \nz.mem_894_sv2v_reg  <= data_i[6];
      \nz.mem_893_sv2v_reg  <= data_i[5];
      \nz.mem_892_sv2v_reg  <= data_i[4];
      \nz.mem_891_sv2v_reg  <= data_i[3];
      \nz.mem_890_sv2v_reg  <= data_i[2];
      \nz.mem_889_sv2v_reg  <= data_i[1];
      \nz.mem_888_sv2v_reg  <= data_i[0];
    end 
    if(N901) begin
      \nz.mem_887_sv2v_reg  <= data_i[7];
      \nz.mem_886_sv2v_reg  <= data_i[6];
      \nz.mem_885_sv2v_reg  <= data_i[5];
      \nz.mem_884_sv2v_reg  <= data_i[4];
      \nz.mem_883_sv2v_reg  <= data_i[3];
      \nz.mem_882_sv2v_reg  <= data_i[2];
      \nz.mem_881_sv2v_reg  <= data_i[1];
      \nz.mem_880_sv2v_reg  <= data_i[0];
    end 
    if(N900) begin
      \nz.mem_879_sv2v_reg  <= data_i[7];
      \nz.mem_878_sv2v_reg  <= data_i[6];
      \nz.mem_877_sv2v_reg  <= data_i[5];
      \nz.mem_876_sv2v_reg  <= data_i[4];
      \nz.mem_875_sv2v_reg  <= data_i[3];
      \nz.mem_874_sv2v_reg  <= data_i[2];
      \nz.mem_873_sv2v_reg  <= data_i[1];
      \nz.mem_872_sv2v_reg  <= data_i[0];
    end 
    if(N899) begin
      \nz.mem_871_sv2v_reg  <= data_i[7];
      \nz.mem_870_sv2v_reg  <= data_i[6];
      \nz.mem_869_sv2v_reg  <= data_i[5];
      \nz.mem_868_sv2v_reg  <= data_i[4];
      \nz.mem_867_sv2v_reg  <= data_i[3];
      \nz.mem_866_sv2v_reg  <= data_i[2];
      \nz.mem_865_sv2v_reg  <= data_i[1];
      \nz.mem_864_sv2v_reg  <= data_i[0];
    end 
    if(N898) begin
      \nz.mem_863_sv2v_reg  <= data_i[7];
      \nz.mem_862_sv2v_reg  <= data_i[6];
      \nz.mem_861_sv2v_reg  <= data_i[5];
      \nz.mem_860_sv2v_reg  <= data_i[4];
      \nz.mem_859_sv2v_reg  <= data_i[3];
      \nz.mem_858_sv2v_reg  <= data_i[2];
      \nz.mem_857_sv2v_reg  <= data_i[1];
      \nz.mem_856_sv2v_reg  <= data_i[0];
    end 
    if(N897) begin
      \nz.mem_855_sv2v_reg  <= data_i[7];
      \nz.mem_854_sv2v_reg  <= data_i[6];
      \nz.mem_853_sv2v_reg  <= data_i[5];
      \nz.mem_852_sv2v_reg  <= data_i[4];
      \nz.mem_851_sv2v_reg  <= data_i[3];
      \nz.mem_850_sv2v_reg  <= data_i[2];
      \nz.mem_849_sv2v_reg  <= data_i[1];
      \nz.mem_848_sv2v_reg  <= data_i[0];
    end 
    if(N896) begin
      \nz.mem_847_sv2v_reg  <= data_i[7];
      \nz.mem_846_sv2v_reg  <= data_i[6];
      \nz.mem_845_sv2v_reg  <= data_i[5];
      \nz.mem_844_sv2v_reg  <= data_i[4];
      \nz.mem_843_sv2v_reg  <= data_i[3];
      \nz.mem_842_sv2v_reg  <= data_i[2];
      \nz.mem_841_sv2v_reg  <= data_i[1];
      \nz.mem_840_sv2v_reg  <= data_i[0];
    end 
    if(N895) begin
      \nz.mem_839_sv2v_reg  <= data_i[7];
      \nz.mem_838_sv2v_reg  <= data_i[6];
      \nz.mem_837_sv2v_reg  <= data_i[5];
      \nz.mem_836_sv2v_reg  <= data_i[4];
      \nz.mem_835_sv2v_reg  <= data_i[3];
      \nz.mem_834_sv2v_reg  <= data_i[2];
      \nz.mem_833_sv2v_reg  <= data_i[1];
      \nz.mem_832_sv2v_reg  <= data_i[0];
    end 
    if(N894) begin
      \nz.mem_831_sv2v_reg  <= data_i[7];
      \nz.mem_830_sv2v_reg  <= data_i[6];
      \nz.mem_829_sv2v_reg  <= data_i[5];
      \nz.mem_828_sv2v_reg  <= data_i[4];
      \nz.mem_827_sv2v_reg  <= data_i[3];
      \nz.mem_826_sv2v_reg  <= data_i[2];
      \nz.mem_825_sv2v_reg  <= data_i[1];
      \nz.mem_824_sv2v_reg  <= data_i[0];
    end 
    if(N893) begin
      \nz.mem_823_sv2v_reg  <= data_i[7];
      \nz.mem_822_sv2v_reg  <= data_i[6];
      \nz.mem_821_sv2v_reg  <= data_i[5];
      \nz.mem_820_sv2v_reg  <= data_i[4];
      \nz.mem_819_sv2v_reg  <= data_i[3];
      \nz.mem_818_sv2v_reg  <= data_i[2];
      \nz.mem_817_sv2v_reg  <= data_i[1];
      \nz.mem_816_sv2v_reg  <= data_i[0];
    end 
    if(N892) begin
      \nz.mem_815_sv2v_reg  <= data_i[7];
      \nz.mem_814_sv2v_reg  <= data_i[6];
      \nz.mem_813_sv2v_reg  <= data_i[5];
      \nz.mem_812_sv2v_reg  <= data_i[4];
      \nz.mem_811_sv2v_reg  <= data_i[3];
      \nz.mem_810_sv2v_reg  <= data_i[2];
      \nz.mem_809_sv2v_reg  <= data_i[1];
      \nz.mem_808_sv2v_reg  <= data_i[0];
    end 
    if(N891) begin
      \nz.mem_807_sv2v_reg  <= data_i[7];
      \nz.mem_806_sv2v_reg  <= data_i[6];
      \nz.mem_805_sv2v_reg  <= data_i[5];
      \nz.mem_804_sv2v_reg  <= data_i[4];
      \nz.mem_803_sv2v_reg  <= data_i[3];
      \nz.mem_802_sv2v_reg  <= data_i[2];
      \nz.mem_801_sv2v_reg  <= data_i[1];
      \nz.mem_800_sv2v_reg  <= data_i[0];
    end 
    if(N890) begin
      \nz.mem_799_sv2v_reg  <= data_i[7];
      \nz.mem_798_sv2v_reg  <= data_i[6];
      \nz.mem_797_sv2v_reg  <= data_i[5];
      \nz.mem_796_sv2v_reg  <= data_i[4];
      \nz.mem_795_sv2v_reg  <= data_i[3];
      \nz.mem_794_sv2v_reg  <= data_i[2];
      \nz.mem_793_sv2v_reg  <= data_i[1];
      \nz.mem_792_sv2v_reg  <= data_i[0];
    end 
    if(N889) begin
      \nz.mem_791_sv2v_reg  <= data_i[7];
      \nz.mem_790_sv2v_reg  <= data_i[6];
      \nz.mem_789_sv2v_reg  <= data_i[5];
      \nz.mem_788_sv2v_reg  <= data_i[4];
      \nz.mem_787_sv2v_reg  <= data_i[3];
      \nz.mem_786_sv2v_reg  <= data_i[2];
      \nz.mem_785_sv2v_reg  <= data_i[1];
      \nz.mem_784_sv2v_reg  <= data_i[0];
    end 
    if(N888) begin
      \nz.mem_783_sv2v_reg  <= data_i[7];
      \nz.mem_782_sv2v_reg  <= data_i[6];
      \nz.mem_781_sv2v_reg  <= data_i[5];
      \nz.mem_780_sv2v_reg  <= data_i[4];
      \nz.mem_779_sv2v_reg  <= data_i[3];
      \nz.mem_778_sv2v_reg  <= data_i[2];
      \nz.mem_777_sv2v_reg  <= data_i[1];
      \nz.mem_776_sv2v_reg  <= data_i[0];
    end 
    if(N887) begin
      \nz.mem_775_sv2v_reg  <= data_i[7];
      \nz.mem_774_sv2v_reg  <= data_i[6];
      \nz.mem_773_sv2v_reg  <= data_i[5];
      \nz.mem_772_sv2v_reg  <= data_i[4];
      \nz.mem_771_sv2v_reg  <= data_i[3];
      \nz.mem_770_sv2v_reg  <= data_i[2];
      \nz.mem_769_sv2v_reg  <= data_i[1];
      \nz.mem_768_sv2v_reg  <= data_i[0];
    end 
    if(N886) begin
      \nz.mem_767_sv2v_reg  <= data_i[7];
      \nz.mem_766_sv2v_reg  <= data_i[6];
      \nz.mem_765_sv2v_reg  <= data_i[5];
      \nz.mem_764_sv2v_reg  <= data_i[4];
      \nz.mem_763_sv2v_reg  <= data_i[3];
      \nz.mem_762_sv2v_reg  <= data_i[2];
      \nz.mem_761_sv2v_reg  <= data_i[1];
      \nz.mem_760_sv2v_reg  <= data_i[0];
    end 
    if(N885) begin
      \nz.mem_759_sv2v_reg  <= data_i[7];
      \nz.mem_758_sv2v_reg  <= data_i[6];
      \nz.mem_757_sv2v_reg  <= data_i[5];
      \nz.mem_756_sv2v_reg  <= data_i[4];
      \nz.mem_755_sv2v_reg  <= data_i[3];
      \nz.mem_754_sv2v_reg  <= data_i[2];
      \nz.mem_753_sv2v_reg  <= data_i[1];
      \nz.mem_752_sv2v_reg  <= data_i[0];
    end 
    if(N884) begin
      \nz.mem_751_sv2v_reg  <= data_i[7];
      \nz.mem_750_sv2v_reg  <= data_i[6];
      \nz.mem_749_sv2v_reg  <= data_i[5];
      \nz.mem_748_sv2v_reg  <= data_i[4];
      \nz.mem_747_sv2v_reg  <= data_i[3];
      \nz.mem_746_sv2v_reg  <= data_i[2];
      \nz.mem_745_sv2v_reg  <= data_i[1];
      \nz.mem_744_sv2v_reg  <= data_i[0];
    end 
    if(N883) begin
      \nz.mem_743_sv2v_reg  <= data_i[7];
      \nz.mem_742_sv2v_reg  <= data_i[6];
      \nz.mem_741_sv2v_reg  <= data_i[5];
      \nz.mem_740_sv2v_reg  <= data_i[4];
      \nz.mem_739_sv2v_reg  <= data_i[3];
      \nz.mem_738_sv2v_reg  <= data_i[2];
      \nz.mem_737_sv2v_reg  <= data_i[1];
      \nz.mem_736_sv2v_reg  <= data_i[0];
    end 
    if(N882) begin
      \nz.mem_735_sv2v_reg  <= data_i[7];
      \nz.mem_734_sv2v_reg  <= data_i[6];
      \nz.mem_733_sv2v_reg  <= data_i[5];
      \nz.mem_732_sv2v_reg  <= data_i[4];
      \nz.mem_731_sv2v_reg  <= data_i[3];
      \nz.mem_730_sv2v_reg  <= data_i[2];
      \nz.mem_729_sv2v_reg  <= data_i[1];
      \nz.mem_728_sv2v_reg  <= data_i[0];
    end 
    if(N881) begin
      \nz.mem_727_sv2v_reg  <= data_i[7];
      \nz.mem_726_sv2v_reg  <= data_i[6];
      \nz.mem_725_sv2v_reg  <= data_i[5];
      \nz.mem_724_sv2v_reg  <= data_i[4];
      \nz.mem_723_sv2v_reg  <= data_i[3];
      \nz.mem_722_sv2v_reg  <= data_i[2];
      \nz.mem_721_sv2v_reg  <= data_i[1];
      \nz.mem_720_sv2v_reg  <= data_i[0];
    end 
    if(N880) begin
      \nz.mem_719_sv2v_reg  <= data_i[7];
      \nz.mem_718_sv2v_reg  <= data_i[6];
      \nz.mem_717_sv2v_reg  <= data_i[5];
      \nz.mem_716_sv2v_reg  <= data_i[4];
      \nz.mem_715_sv2v_reg  <= data_i[3];
      \nz.mem_714_sv2v_reg  <= data_i[2];
      \nz.mem_713_sv2v_reg  <= data_i[1];
      \nz.mem_712_sv2v_reg  <= data_i[0];
    end 
    if(N879) begin
      \nz.mem_711_sv2v_reg  <= data_i[7];
      \nz.mem_710_sv2v_reg  <= data_i[6];
      \nz.mem_709_sv2v_reg  <= data_i[5];
      \nz.mem_708_sv2v_reg  <= data_i[4];
      \nz.mem_707_sv2v_reg  <= data_i[3];
      \nz.mem_706_sv2v_reg  <= data_i[2];
      \nz.mem_705_sv2v_reg  <= data_i[1];
      \nz.mem_704_sv2v_reg  <= data_i[0];
    end 
    if(N878) begin
      \nz.mem_703_sv2v_reg  <= data_i[7];
      \nz.mem_702_sv2v_reg  <= data_i[6];
      \nz.mem_701_sv2v_reg  <= data_i[5];
      \nz.mem_700_sv2v_reg  <= data_i[4];
      \nz.mem_699_sv2v_reg  <= data_i[3];
      \nz.mem_698_sv2v_reg  <= data_i[2];
      \nz.mem_697_sv2v_reg  <= data_i[1];
      \nz.mem_696_sv2v_reg  <= data_i[0];
    end 
    if(N877) begin
      \nz.mem_695_sv2v_reg  <= data_i[7];
      \nz.mem_694_sv2v_reg  <= data_i[6];
      \nz.mem_693_sv2v_reg  <= data_i[5];
      \nz.mem_692_sv2v_reg  <= data_i[4];
      \nz.mem_691_sv2v_reg  <= data_i[3];
      \nz.mem_690_sv2v_reg  <= data_i[2];
      \nz.mem_689_sv2v_reg  <= data_i[1];
      \nz.mem_688_sv2v_reg  <= data_i[0];
    end 
    if(N876) begin
      \nz.mem_687_sv2v_reg  <= data_i[7];
      \nz.mem_686_sv2v_reg  <= data_i[6];
      \nz.mem_685_sv2v_reg  <= data_i[5];
      \nz.mem_684_sv2v_reg  <= data_i[4];
      \nz.mem_683_sv2v_reg  <= data_i[3];
      \nz.mem_682_sv2v_reg  <= data_i[2];
      \nz.mem_681_sv2v_reg  <= data_i[1];
      \nz.mem_680_sv2v_reg  <= data_i[0];
    end 
    if(N875) begin
      \nz.mem_679_sv2v_reg  <= data_i[7];
      \nz.mem_678_sv2v_reg  <= data_i[6];
      \nz.mem_677_sv2v_reg  <= data_i[5];
      \nz.mem_676_sv2v_reg  <= data_i[4];
      \nz.mem_675_sv2v_reg  <= data_i[3];
      \nz.mem_674_sv2v_reg  <= data_i[2];
      \nz.mem_673_sv2v_reg  <= data_i[1];
      \nz.mem_672_sv2v_reg  <= data_i[0];
    end 
    if(N874) begin
      \nz.mem_671_sv2v_reg  <= data_i[7];
      \nz.mem_670_sv2v_reg  <= data_i[6];
      \nz.mem_669_sv2v_reg  <= data_i[5];
      \nz.mem_668_sv2v_reg  <= data_i[4];
      \nz.mem_667_sv2v_reg  <= data_i[3];
      \nz.mem_666_sv2v_reg  <= data_i[2];
      \nz.mem_665_sv2v_reg  <= data_i[1];
      \nz.mem_664_sv2v_reg  <= data_i[0];
    end 
    if(N873) begin
      \nz.mem_663_sv2v_reg  <= data_i[7];
      \nz.mem_662_sv2v_reg  <= data_i[6];
      \nz.mem_661_sv2v_reg  <= data_i[5];
      \nz.mem_660_sv2v_reg  <= data_i[4];
      \nz.mem_659_sv2v_reg  <= data_i[3];
      \nz.mem_658_sv2v_reg  <= data_i[2];
      \nz.mem_657_sv2v_reg  <= data_i[1];
      \nz.mem_656_sv2v_reg  <= data_i[0];
    end 
    if(N872) begin
      \nz.mem_655_sv2v_reg  <= data_i[7];
      \nz.mem_654_sv2v_reg  <= data_i[6];
      \nz.mem_653_sv2v_reg  <= data_i[5];
      \nz.mem_652_sv2v_reg  <= data_i[4];
      \nz.mem_651_sv2v_reg  <= data_i[3];
      \nz.mem_650_sv2v_reg  <= data_i[2];
      \nz.mem_649_sv2v_reg  <= data_i[1];
      \nz.mem_648_sv2v_reg  <= data_i[0];
    end 
    if(N871) begin
      \nz.mem_647_sv2v_reg  <= data_i[7];
      \nz.mem_646_sv2v_reg  <= data_i[6];
      \nz.mem_645_sv2v_reg  <= data_i[5];
      \nz.mem_644_sv2v_reg  <= data_i[4];
      \nz.mem_643_sv2v_reg  <= data_i[3];
      \nz.mem_642_sv2v_reg  <= data_i[2];
      \nz.mem_641_sv2v_reg  <= data_i[1];
      \nz.mem_640_sv2v_reg  <= data_i[0];
    end 
    if(N870) begin
      \nz.mem_639_sv2v_reg  <= data_i[7];
      \nz.mem_638_sv2v_reg  <= data_i[6];
      \nz.mem_637_sv2v_reg  <= data_i[5];
      \nz.mem_636_sv2v_reg  <= data_i[4];
      \nz.mem_635_sv2v_reg  <= data_i[3];
      \nz.mem_634_sv2v_reg  <= data_i[2];
      \nz.mem_633_sv2v_reg  <= data_i[1];
      \nz.mem_632_sv2v_reg  <= data_i[0];
    end 
    if(N869) begin
      \nz.mem_631_sv2v_reg  <= data_i[7];
      \nz.mem_630_sv2v_reg  <= data_i[6];
      \nz.mem_629_sv2v_reg  <= data_i[5];
      \nz.mem_628_sv2v_reg  <= data_i[4];
      \nz.mem_627_sv2v_reg  <= data_i[3];
      \nz.mem_626_sv2v_reg  <= data_i[2];
      \nz.mem_625_sv2v_reg  <= data_i[1];
      \nz.mem_624_sv2v_reg  <= data_i[0];
    end 
    if(N868) begin
      \nz.mem_623_sv2v_reg  <= data_i[7];
      \nz.mem_622_sv2v_reg  <= data_i[6];
      \nz.mem_621_sv2v_reg  <= data_i[5];
      \nz.mem_620_sv2v_reg  <= data_i[4];
      \nz.mem_619_sv2v_reg  <= data_i[3];
      \nz.mem_618_sv2v_reg  <= data_i[2];
      \nz.mem_617_sv2v_reg  <= data_i[1];
      \nz.mem_616_sv2v_reg  <= data_i[0];
    end 
    if(N867) begin
      \nz.mem_615_sv2v_reg  <= data_i[7];
      \nz.mem_614_sv2v_reg  <= data_i[6];
      \nz.mem_613_sv2v_reg  <= data_i[5];
      \nz.mem_612_sv2v_reg  <= data_i[4];
      \nz.mem_611_sv2v_reg  <= data_i[3];
      \nz.mem_610_sv2v_reg  <= data_i[2];
      \nz.mem_609_sv2v_reg  <= data_i[1];
      \nz.mem_608_sv2v_reg  <= data_i[0];
    end 
    if(N866) begin
      \nz.mem_607_sv2v_reg  <= data_i[7];
      \nz.mem_606_sv2v_reg  <= data_i[6];
      \nz.mem_605_sv2v_reg  <= data_i[5];
      \nz.mem_604_sv2v_reg  <= data_i[4];
      \nz.mem_603_sv2v_reg  <= data_i[3];
      \nz.mem_602_sv2v_reg  <= data_i[2];
      \nz.mem_601_sv2v_reg  <= data_i[1];
      \nz.mem_600_sv2v_reg  <= data_i[0];
    end 
    if(N865) begin
      \nz.mem_599_sv2v_reg  <= data_i[7];
      \nz.mem_598_sv2v_reg  <= data_i[6];
      \nz.mem_597_sv2v_reg  <= data_i[5];
      \nz.mem_596_sv2v_reg  <= data_i[4];
      \nz.mem_595_sv2v_reg  <= data_i[3];
      \nz.mem_594_sv2v_reg  <= data_i[2];
      \nz.mem_593_sv2v_reg  <= data_i[1];
      \nz.mem_592_sv2v_reg  <= data_i[0];
    end 
    if(N864) begin
      \nz.mem_591_sv2v_reg  <= data_i[7];
      \nz.mem_590_sv2v_reg  <= data_i[6];
      \nz.mem_589_sv2v_reg  <= data_i[5];
      \nz.mem_588_sv2v_reg  <= data_i[4];
      \nz.mem_587_sv2v_reg  <= data_i[3];
      \nz.mem_586_sv2v_reg  <= data_i[2];
      \nz.mem_585_sv2v_reg  <= data_i[1];
      \nz.mem_584_sv2v_reg  <= data_i[0];
    end 
    if(N863) begin
      \nz.mem_583_sv2v_reg  <= data_i[7];
      \nz.mem_582_sv2v_reg  <= data_i[6];
      \nz.mem_581_sv2v_reg  <= data_i[5];
      \nz.mem_580_sv2v_reg  <= data_i[4];
      \nz.mem_579_sv2v_reg  <= data_i[3];
      \nz.mem_578_sv2v_reg  <= data_i[2];
      \nz.mem_577_sv2v_reg  <= data_i[1];
      \nz.mem_576_sv2v_reg  <= data_i[0];
    end 
    if(N862) begin
      \nz.mem_575_sv2v_reg  <= data_i[7];
      \nz.mem_574_sv2v_reg  <= data_i[6];
      \nz.mem_573_sv2v_reg  <= data_i[5];
      \nz.mem_572_sv2v_reg  <= data_i[4];
      \nz.mem_571_sv2v_reg  <= data_i[3];
      \nz.mem_570_sv2v_reg  <= data_i[2];
      \nz.mem_569_sv2v_reg  <= data_i[1];
      \nz.mem_568_sv2v_reg  <= data_i[0];
    end 
    if(N861) begin
      \nz.mem_567_sv2v_reg  <= data_i[7];
      \nz.mem_566_sv2v_reg  <= data_i[6];
      \nz.mem_565_sv2v_reg  <= data_i[5];
      \nz.mem_564_sv2v_reg  <= data_i[4];
      \nz.mem_563_sv2v_reg  <= data_i[3];
      \nz.mem_562_sv2v_reg  <= data_i[2];
      \nz.mem_561_sv2v_reg  <= data_i[1];
      \nz.mem_560_sv2v_reg  <= data_i[0];
    end 
    if(N860) begin
      \nz.mem_559_sv2v_reg  <= data_i[7];
      \nz.mem_558_sv2v_reg  <= data_i[6];
      \nz.mem_557_sv2v_reg  <= data_i[5];
      \nz.mem_556_sv2v_reg  <= data_i[4];
      \nz.mem_555_sv2v_reg  <= data_i[3];
      \nz.mem_554_sv2v_reg  <= data_i[2];
      \nz.mem_553_sv2v_reg  <= data_i[1];
      \nz.mem_552_sv2v_reg  <= data_i[0];
    end 
    if(N859) begin
      \nz.mem_551_sv2v_reg  <= data_i[7];
      \nz.mem_550_sv2v_reg  <= data_i[6];
      \nz.mem_549_sv2v_reg  <= data_i[5];
      \nz.mem_548_sv2v_reg  <= data_i[4];
      \nz.mem_547_sv2v_reg  <= data_i[3];
      \nz.mem_546_sv2v_reg  <= data_i[2];
      \nz.mem_545_sv2v_reg  <= data_i[1];
      \nz.mem_544_sv2v_reg  <= data_i[0];
    end 
    if(N858) begin
      \nz.mem_543_sv2v_reg  <= data_i[7];
      \nz.mem_542_sv2v_reg  <= data_i[6];
      \nz.mem_541_sv2v_reg  <= data_i[5];
      \nz.mem_540_sv2v_reg  <= data_i[4];
      \nz.mem_539_sv2v_reg  <= data_i[3];
      \nz.mem_538_sv2v_reg  <= data_i[2];
      \nz.mem_537_sv2v_reg  <= data_i[1];
      \nz.mem_536_sv2v_reg  <= data_i[0];
    end 
    if(N857) begin
      \nz.mem_535_sv2v_reg  <= data_i[7];
      \nz.mem_534_sv2v_reg  <= data_i[6];
      \nz.mem_533_sv2v_reg  <= data_i[5];
      \nz.mem_532_sv2v_reg  <= data_i[4];
      \nz.mem_531_sv2v_reg  <= data_i[3];
      \nz.mem_530_sv2v_reg  <= data_i[2];
      \nz.mem_529_sv2v_reg  <= data_i[1];
      \nz.mem_528_sv2v_reg  <= data_i[0];
    end 
    if(N856) begin
      \nz.mem_527_sv2v_reg  <= data_i[7];
      \nz.mem_526_sv2v_reg  <= data_i[6];
      \nz.mem_525_sv2v_reg  <= data_i[5];
      \nz.mem_524_sv2v_reg  <= data_i[4];
      \nz.mem_523_sv2v_reg  <= data_i[3];
      \nz.mem_522_sv2v_reg  <= data_i[2];
      \nz.mem_521_sv2v_reg  <= data_i[1];
      \nz.mem_520_sv2v_reg  <= data_i[0];
    end 
    if(N855) begin
      \nz.mem_519_sv2v_reg  <= data_i[7];
      \nz.mem_518_sv2v_reg  <= data_i[6];
      \nz.mem_517_sv2v_reg  <= data_i[5];
      \nz.mem_516_sv2v_reg  <= data_i[4];
      \nz.mem_515_sv2v_reg  <= data_i[3];
      \nz.mem_514_sv2v_reg  <= data_i[2];
      \nz.mem_513_sv2v_reg  <= data_i[1];
      \nz.mem_512_sv2v_reg  <= data_i[0];
    end 
    if(N854) begin
      \nz.mem_511_sv2v_reg  <= data_i[7];
      \nz.mem_510_sv2v_reg  <= data_i[6];
      \nz.mem_509_sv2v_reg  <= data_i[5];
      \nz.mem_508_sv2v_reg  <= data_i[4];
      \nz.mem_507_sv2v_reg  <= data_i[3];
      \nz.mem_506_sv2v_reg  <= data_i[2];
      \nz.mem_505_sv2v_reg  <= data_i[1];
      \nz.mem_504_sv2v_reg  <= data_i[0];
    end 
    if(N853) begin
      \nz.mem_503_sv2v_reg  <= data_i[7];
      \nz.mem_502_sv2v_reg  <= data_i[6];
      \nz.mem_501_sv2v_reg  <= data_i[5];
      \nz.mem_500_sv2v_reg  <= data_i[4];
      \nz.mem_499_sv2v_reg  <= data_i[3];
      \nz.mem_498_sv2v_reg  <= data_i[2];
      \nz.mem_497_sv2v_reg  <= data_i[1];
      \nz.mem_496_sv2v_reg  <= data_i[0];
    end 
    if(N852) begin
      \nz.mem_495_sv2v_reg  <= data_i[7];
      \nz.mem_494_sv2v_reg  <= data_i[6];
      \nz.mem_493_sv2v_reg  <= data_i[5];
      \nz.mem_492_sv2v_reg  <= data_i[4];
      \nz.mem_491_sv2v_reg  <= data_i[3];
      \nz.mem_490_sv2v_reg  <= data_i[2];
      \nz.mem_489_sv2v_reg  <= data_i[1];
      \nz.mem_488_sv2v_reg  <= data_i[0];
    end 
    if(N851) begin
      \nz.mem_487_sv2v_reg  <= data_i[7];
      \nz.mem_486_sv2v_reg  <= data_i[6];
      \nz.mem_485_sv2v_reg  <= data_i[5];
      \nz.mem_484_sv2v_reg  <= data_i[4];
      \nz.mem_483_sv2v_reg  <= data_i[3];
      \nz.mem_482_sv2v_reg  <= data_i[2];
      \nz.mem_481_sv2v_reg  <= data_i[1];
      \nz.mem_480_sv2v_reg  <= data_i[0];
    end 
    if(N850) begin
      \nz.mem_479_sv2v_reg  <= data_i[7];
      \nz.mem_478_sv2v_reg  <= data_i[6];
      \nz.mem_477_sv2v_reg  <= data_i[5];
      \nz.mem_476_sv2v_reg  <= data_i[4];
      \nz.mem_475_sv2v_reg  <= data_i[3];
      \nz.mem_474_sv2v_reg  <= data_i[2];
      \nz.mem_473_sv2v_reg  <= data_i[1];
      \nz.mem_472_sv2v_reg  <= data_i[0];
    end 
    if(N849) begin
      \nz.mem_471_sv2v_reg  <= data_i[7];
      \nz.mem_470_sv2v_reg  <= data_i[6];
      \nz.mem_469_sv2v_reg  <= data_i[5];
      \nz.mem_468_sv2v_reg  <= data_i[4];
      \nz.mem_467_sv2v_reg  <= data_i[3];
      \nz.mem_466_sv2v_reg  <= data_i[2];
      \nz.mem_465_sv2v_reg  <= data_i[1];
      \nz.mem_464_sv2v_reg  <= data_i[0];
    end 
    if(N848) begin
      \nz.mem_463_sv2v_reg  <= data_i[7];
      \nz.mem_462_sv2v_reg  <= data_i[6];
      \nz.mem_461_sv2v_reg  <= data_i[5];
      \nz.mem_460_sv2v_reg  <= data_i[4];
      \nz.mem_459_sv2v_reg  <= data_i[3];
      \nz.mem_458_sv2v_reg  <= data_i[2];
      \nz.mem_457_sv2v_reg  <= data_i[1];
      \nz.mem_456_sv2v_reg  <= data_i[0];
    end 
    if(N847) begin
      \nz.mem_455_sv2v_reg  <= data_i[7];
      \nz.mem_454_sv2v_reg  <= data_i[6];
      \nz.mem_453_sv2v_reg  <= data_i[5];
      \nz.mem_452_sv2v_reg  <= data_i[4];
      \nz.mem_451_sv2v_reg  <= data_i[3];
      \nz.mem_450_sv2v_reg  <= data_i[2];
      \nz.mem_449_sv2v_reg  <= data_i[1];
      \nz.mem_448_sv2v_reg  <= data_i[0];
    end 
    if(N846) begin
      \nz.mem_447_sv2v_reg  <= data_i[7];
      \nz.mem_446_sv2v_reg  <= data_i[6];
      \nz.mem_445_sv2v_reg  <= data_i[5];
      \nz.mem_444_sv2v_reg  <= data_i[4];
      \nz.mem_443_sv2v_reg  <= data_i[3];
      \nz.mem_442_sv2v_reg  <= data_i[2];
      \nz.mem_441_sv2v_reg  <= data_i[1];
      \nz.mem_440_sv2v_reg  <= data_i[0];
    end 
    if(N845) begin
      \nz.mem_439_sv2v_reg  <= data_i[7];
      \nz.mem_438_sv2v_reg  <= data_i[6];
      \nz.mem_437_sv2v_reg  <= data_i[5];
      \nz.mem_436_sv2v_reg  <= data_i[4];
      \nz.mem_435_sv2v_reg  <= data_i[3];
      \nz.mem_434_sv2v_reg  <= data_i[2];
      \nz.mem_433_sv2v_reg  <= data_i[1];
      \nz.mem_432_sv2v_reg  <= data_i[0];
    end 
    if(N844) begin
      \nz.mem_431_sv2v_reg  <= data_i[7];
      \nz.mem_430_sv2v_reg  <= data_i[6];
      \nz.mem_429_sv2v_reg  <= data_i[5];
      \nz.mem_428_sv2v_reg  <= data_i[4];
      \nz.mem_427_sv2v_reg  <= data_i[3];
      \nz.mem_426_sv2v_reg  <= data_i[2];
      \nz.mem_425_sv2v_reg  <= data_i[1];
      \nz.mem_424_sv2v_reg  <= data_i[0];
    end 
    if(N843) begin
      \nz.mem_423_sv2v_reg  <= data_i[7];
      \nz.mem_422_sv2v_reg  <= data_i[6];
      \nz.mem_421_sv2v_reg  <= data_i[5];
      \nz.mem_420_sv2v_reg  <= data_i[4];
      \nz.mem_419_sv2v_reg  <= data_i[3];
      \nz.mem_418_sv2v_reg  <= data_i[2];
      \nz.mem_417_sv2v_reg  <= data_i[1];
      \nz.mem_416_sv2v_reg  <= data_i[0];
    end 
    if(N842) begin
      \nz.mem_415_sv2v_reg  <= data_i[7];
      \nz.mem_414_sv2v_reg  <= data_i[6];
      \nz.mem_413_sv2v_reg  <= data_i[5];
      \nz.mem_412_sv2v_reg  <= data_i[4];
      \nz.mem_411_sv2v_reg  <= data_i[3];
      \nz.mem_410_sv2v_reg  <= data_i[2];
      \nz.mem_409_sv2v_reg  <= data_i[1];
      \nz.mem_408_sv2v_reg  <= data_i[0];
    end 
    if(N841) begin
      \nz.mem_407_sv2v_reg  <= data_i[7];
      \nz.mem_406_sv2v_reg  <= data_i[6];
      \nz.mem_405_sv2v_reg  <= data_i[5];
      \nz.mem_404_sv2v_reg  <= data_i[4];
      \nz.mem_403_sv2v_reg  <= data_i[3];
      \nz.mem_402_sv2v_reg  <= data_i[2];
      \nz.mem_401_sv2v_reg  <= data_i[1];
      \nz.mem_400_sv2v_reg  <= data_i[0];
    end 
    if(N840) begin
      \nz.mem_399_sv2v_reg  <= data_i[7];
      \nz.mem_398_sv2v_reg  <= data_i[6];
      \nz.mem_397_sv2v_reg  <= data_i[5];
      \nz.mem_396_sv2v_reg  <= data_i[4];
      \nz.mem_395_sv2v_reg  <= data_i[3];
      \nz.mem_394_sv2v_reg  <= data_i[2];
      \nz.mem_393_sv2v_reg  <= data_i[1];
      \nz.mem_392_sv2v_reg  <= data_i[0];
    end 
    if(N839) begin
      \nz.mem_391_sv2v_reg  <= data_i[7];
      \nz.mem_390_sv2v_reg  <= data_i[6];
      \nz.mem_389_sv2v_reg  <= data_i[5];
      \nz.mem_388_sv2v_reg  <= data_i[4];
      \nz.mem_387_sv2v_reg  <= data_i[3];
      \nz.mem_386_sv2v_reg  <= data_i[2];
      \nz.mem_385_sv2v_reg  <= data_i[1];
      \nz.mem_384_sv2v_reg  <= data_i[0];
    end 
    if(N838) begin
      \nz.mem_383_sv2v_reg  <= data_i[7];
      \nz.mem_382_sv2v_reg  <= data_i[6];
      \nz.mem_381_sv2v_reg  <= data_i[5];
      \nz.mem_380_sv2v_reg  <= data_i[4];
      \nz.mem_379_sv2v_reg  <= data_i[3];
      \nz.mem_378_sv2v_reg  <= data_i[2];
      \nz.mem_377_sv2v_reg  <= data_i[1];
      \nz.mem_376_sv2v_reg  <= data_i[0];
    end 
    if(N837) begin
      \nz.mem_375_sv2v_reg  <= data_i[7];
      \nz.mem_374_sv2v_reg  <= data_i[6];
      \nz.mem_373_sv2v_reg  <= data_i[5];
      \nz.mem_372_sv2v_reg  <= data_i[4];
      \nz.mem_371_sv2v_reg  <= data_i[3];
      \nz.mem_370_sv2v_reg  <= data_i[2];
      \nz.mem_369_sv2v_reg  <= data_i[1];
      \nz.mem_368_sv2v_reg  <= data_i[0];
    end 
    if(N836) begin
      \nz.mem_367_sv2v_reg  <= data_i[7];
      \nz.mem_366_sv2v_reg  <= data_i[6];
      \nz.mem_365_sv2v_reg  <= data_i[5];
      \nz.mem_364_sv2v_reg  <= data_i[4];
      \nz.mem_363_sv2v_reg  <= data_i[3];
      \nz.mem_362_sv2v_reg  <= data_i[2];
      \nz.mem_361_sv2v_reg  <= data_i[1];
      \nz.mem_360_sv2v_reg  <= data_i[0];
    end 
    if(N835) begin
      \nz.mem_359_sv2v_reg  <= data_i[7];
      \nz.mem_358_sv2v_reg  <= data_i[6];
      \nz.mem_357_sv2v_reg  <= data_i[5];
      \nz.mem_356_sv2v_reg  <= data_i[4];
      \nz.mem_355_sv2v_reg  <= data_i[3];
      \nz.mem_354_sv2v_reg  <= data_i[2];
      \nz.mem_353_sv2v_reg  <= data_i[1];
      \nz.mem_352_sv2v_reg  <= data_i[0];
    end 
    if(N834) begin
      \nz.mem_351_sv2v_reg  <= data_i[7];
      \nz.mem_350_sv2v_reg  <= data_i[6];
      \nz.mem_349_sv2v_reg  <= data_i[5];
      \nz.mem_348_sv2v_reg  <= data_i[4];
      \nz.mem_347_sv2v_reg  <= data_i[3];
      \nz.mem_346_sv2v_reg  <= data_i[2];
      \nz.mem_345_sv2v_reg  <= data_i[1];
      \nz.mem_344_sv2v_reg  <= data_i[0];
    end 
    if(N833) begin
      \nz.mem_343_sv2v_reg  <= data_i[7];
      \nz.mem_342_sv2v_reg  <= data_i[6];
      \nz.mem_341_sv2v_reg  <= data_i[5];
      \nz.mem_340_sv2v_reg  <= data_i[4];
      \nz.mem_339_sv2v_reg  <= data_i[3];
      \nz.mem_338_sv2v_reg  <= data_i[2];
      \nz.mem_337_sv2v_reg  <= data_i[1];
      \nz.mem_336_sv2v_reg  <= data_i[0];
    end 
    if(N832) begin
      \nz.mem_335_sv2v_reg  <= data_i[7];
      \nz.mem_334_sv2v_reg  <= data_i[6];
      \nz.mem_333_sv2v_reg  <= data_i[5];
      \nz.mem_332_sv2v_reg  <= data_i[4];
      \nz.mem_331_sv2v_reg  <= data_i[3];
      \nz.mem_330_sv2v_reg  <= data_i[2];
      \nz.mem_329_sv2v_reg  <= data_i[1];
      \nz.mem_328_sv2v_reg  <= data_i[0];
    end 
    if(N831) begin
      \nz.mem_327_sv2v_reg  <= data_i[7];
      \nz.mem_326_sv2v_reg  <= data_i[6];
      \nz.mem_325_sv2v_reg  <= data_i[5];
      \nz.mem_324_sv2v_reg  <= data_i[4];
      \nz.mem_323_sv2v_reg  <= data_i[3];
      \nz.mem_322_sv2v_reg  <= data_i[2];
      \nz.mem_321_sv2v_reg  <= data_i[1];
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N830) begin
      \nz.mem_319_sv2v_reg  <= data_i[7];
      \nz.mem_318_sv2v_reg  <= data_i[6];
      \nz.mem_317_sv2v_reg  <= data_i[5];
      \nz.mem_316_sv2v_reg  <= data_i[4];
      \nz.mem_315_sv2v_reg  <= data_i[3];
      \nz.mem_314_sv2v_reg  <= data_i[2];
      \nz.mem_313_sv2v_reg  <= data_i[1];
      \nz.mem_312_sv2v_reg  <= data_i[0];
    end 
    if(N829) begin
      \nz.mem_311_sv2v_reg  <= data_i[7];
      \nz.mem_310_sv2v_reg  <= data_i[6];
      \nz.mem_309_sv2v_reg  <= data_i[5];
      \nz.mem_308_sv2v_reg  <= data_i[4];
      \nz.mem_307_sv2v_reg  <= data_i[3];
      \nz.mem_306_sv2v_reg  <= data_i[2];
      \nz.mem_305_sv2v_reg  <= data_i[1];
      \nz.mem_304_sv2v_reg  <= data_i[0];
    end 
    if(N828) begin
      \nz.mem_303_sv2v_reg  <= data_i[7];
      \nz.mem_302_sv2v_reg  <= data_i[6];
      \nz.mem_301_sv2v_reg  <= data_i[5];
      \nz.mem_300_sv2v_reg  <= data_i[4];
      \nz.mem_299_sv2v_reg  <= data_i[3];
      \nz.mem_298_sv2v_reg  <= data_i[2];
      \nz.mem_297_sv2v_reg  <= data_i[1];
      \nz.mem_296_sv2v_reg  <= data_i[0];
    end 
    if(N827) begin
      \nz.mem_295_sv2v_reg  <= data_i[7];
      \nz.mem_294_sv2v_reg  <= data_i[6];
      \nz.mem_293_sv2v_reg  <= data_i[5];
      \nz.mem_292_sv2v_reg  <= data_i[4];
      \nz.mem_291_sv2v_reg  <= data_i[3];
      \nz.mem_290_sv2v_reg  <= data_i[2];
      \nz.mem_289_sv2v_reg  <= data_i[1];
      \nz.mem_288_sv2v_reg  <= data_i[0];
    end 
    if(N826) begin
      \nz.mem_287_sv2v_reg  <= data_i[7];
      \nz.mem_286_sv2v_reg  <= data_i[6];
      \nz.mem_285_sv2v_reg  <= data_i[5];
      \nz.mem_284_sv2v_reg  <= data_i[4];
      \nz.mem_283_sv2v_reg  <= data_i[3];
      \nz.mem_282_sv2v_reg  <= data_i[2];
      \nz.mem_281_sv2v_reg  <= data_i[1];
      \nz.mem_280_sv2v_reg  <= data_i[0];
    end 
    if(N825) begin
      \nz.mem_279_sv2v_reg  <= data_i[7];
      \nz.mem_278_sv2v_reg  <= data_i[6];
      \nz.mem_277_sv2v_reg  <= data_i[5];
      \nz.mem_276_sv2v_reg  <= data_i[4];
      \nz.mem_275_sv2v_reg  <= data_i[3];
      \nz.mem_274_sv2v_reg  <= data_i[2];
      \nz.mem_273_sv2v_reg  <= data_i[1];
      \nz.mem_272_sv2v_reg  <= data_i[0];
    end 
    if(N824) begin
      \nz.mem_271_sv2v_reg  <= data_i[7];
      \nz.mem_270_sv2v_reg  <= data_i[6];
      \nz.mem_269_sv2v_reg  <= data_i[5];
      \nz.mem_268_sv2v_reg  <= data_i[4];
      \nz.mem_267_sv2v_reg  <= data_i[3];
      \nz.mem_266_sv2v_reg  <= data_i[2];
      \nz.mem_265_sv2v_reg  <= data_i[1];
      \nz.mem_264_sv2v_reg  <= data_i[0];
    end 
    if(N823) begin
      \nz.mem_263_sv2v_reg  <= data_i[7];
      \nz.mem_262_sv2v_reg  <= data_i[6];
      \nz.mem_261_sv2v_reg  <= data_i[5];
      \nz.mem_260_sv2v_reg  <= data_i[4];
      \nz.mem_259_sv2v_reg  <= data_i[3];
      \nz.mem_258_sv2v_reg  <= data_i[2];
      \nz.mem_257_sv2v_reg  <= data_i[1];
      \nz.mem_256_sv2v_reg  <= data_i[0];
    end 
    if(N822) begin
      \nz.mem_255_sv2v_reg  <= data_i[7];
      \nz.mem_254_sv2v_reg  <= data_i[6];
      \nz.mem_253_sv2v_reg  <= data_i[5];
      \nz.mem_252_sv2v_reg  <= data_i[4];
      \nz.mem_251_sv2v_reg  <= data_i[3];
      \nz.mem_250_sv2v_reg  <= data_i[2];
      \nz.mem_249_sv2v_reg  <= data_i[1];
      \nz.mem_248_sv2v_reg  <= data_i[0];
    end 
    if(N821) begin
      \nz.mem_247_sv2v_reg  <= data_i[7];
      \nz.mem_246_sv2v_reg  <= data_i[6];
      \nz.mem_245_sv2v_reg  <= data_i[5];
      \nz.mem_244_sv2v_reg  <= data_i[4];
      \nz.mem_243_sv2v_reg  <= data_i[3];
      \nz.mem_242_sv2v_reg  <= data_i[2];
      \nz.mem_241_sv2v_reg  <= data_i[1];
      \nz.mem_240_sv2v_reg  <= data_i[0];
    end 
    if(N820) begin
      \nz.mem_239_sv2v_reg  <= data_i[7];
      \nz.mem_238_sv2v_reg  <= data_i[6];
      \nz.mem_237_sv2v_reg  <= data_i[5];
      \nz.mem_236_sv2v_reg  <= data_i[4];
      \nz.mem_235_sv2v_reg  <= data_i[3];
      \nz.mem_234_sv2v_reg  <= data_i[2];
      \nz.mem_233_sv2v_reg  <= data_i[1];
      \nz.mem_232_sv2v_reg  <= data_i[0];
    end 
    if(N819) begin
      \nz.mem_231_sv2v_reg  <= data_i[7];
      \nz.mem_230_sv2v_reg  <= data_i[6];
      \nz.mem_229_sv2v_reg  <= data_i[5];
      \nz.mem_228_sv2v_reg  <= data_i[4];
      \nz.mem_227_sv2v_reg  <= data_i[3];
      \nz.mem_226_sv2v_reg  <= data_i[2];
      \nz.mem_225_sv2v_reg  <= data_i[1];
      \nz.mem_224_sv2v_reg  <= data_i[0];
    end 
    if(N818) begin
      \nz.mem_223_sv2v_reg  <= data_i[7];
      \nz.mem_222_sv2v_reg  <= data_i[6];
      \nz.mem_221_sv2v_reg  <= data_i[5];
      \nz.mem_220_sv2v_reg  <= data_i[4];
      \nz.mem_219_sv2v_reg  <= data_i[3];
      \nz.mem_218_sv2v_reg  <= data_i[2];
      \nz.mem_217_sv2v_reg  <= data_i[1];
      \nz.mem_216_sv2v_reg  <= data_i[0];
    end 
    if(N817) begin
      \nz.mem_215_sv2v_reg  <= data_i[7];
      \nz.mem_214_sv2v_reg  <= data_i[6];
      \nz.mem_213_sv2v_reg  <= data_i[5];
      \nz.mem_212_sv2v_reg  <= data_i[4];
      \nz.mem_211_sv2v_reg  <= data_i[3];
      \nz.mem_210_sv2v_reg  <= data_i[2];
      \nz.mem_209_sv2v_reg  <= data_i[1];
      \nz.mem_208_sv2v_reg  <= data_i[0];
    end 
    if(N816) begin
      \nz.mem_207_sv2v_reg  <= data_i[7];
      \nz.mem_206_sv2v_reg  <= data_i[6];
      \nz.mem_205_sv2v_reg  <= data_i[5];
      \nz.mem_204_sv2v_reg  <= data_i[4];
      \nz.mem_203_sv2v_reg  <= data_i[3];
      \nz.mem_202_sv2v_reg  <= data_i[2];
      \nz.mem_201_sv2v_reg  <= data_i[1];
      \nz.mem_200_sv2v_reg  <= data_i[0];
    end 
    if(N815) begin
      \nz.mem_199_sv2v_reg  <= data_i[7];
      \nz.mem_198_sv2v_reg  <= data_i[6];
      \nz.mem_197_sv2v_reg  <= data_i[5];
      \nz.mem_196_sv2v_reg  <= data_i[4];
      \nz.mem_195_sv2v_reg  <= data_i[3];
      \nz.mem_194_sv2v_reg  <= data_i[2];
      \nz.mem_193_sv2v_reg  <= data_i[1];
      \nz.mem_192_sv2v_reg  <= data_i[0];
    end 
    if(N814) begin
      \nz.mem_191_sv2v_reg  <= data_i[7];
      \nz.mem_190_sv2v_reg  <= data_i[6];
      \nz.mem_189_sv2v_reg  <= data_i[5];
      \nz.mem_188_sv2v_reg  <= data_i[4];
      \nz.mem_187_sv2v_reg  <= data_i[3];
      \nz.mem_186_sv2v_reg  <= data_i[2];
      \nz.mem_185_sv2v_reg  <= data_i[1];
      \nz.mem_184_sv2v_reg  <= data_i[0];
    end 
    if(N813) begin
      \nz.mem_183_sv2v_reg  <= data_i[7];
      \nz.mem_182_sv2v_reg  <= data_i[6];
      \nz.mem_181_sv2v_reg  <= data_i[5];
      \nz.mem_180_sv2v_reg  <= data_i[4];
      \nz.mem_179_sv2v_reg  <= data_i[3];
      \nz.mem_178_sv2v_reg  <= data_i[2];
      \nz.mem_177_sv2v_reg  <= data_i[1];
      \nz.mem_176_sv2v_reg  <= data_i[0];
    end 
    if(N812) begin
      \nz.mem_175_sv2v_reg  <= data_i[7];
      \nz.mem_174_sv2v_reg  <= data_i[6];
      \nz.mem_173_sv2v_reg  <= data_i[5];
      \nz.mem_172_sv2v_reg  <= data_i[4];
      \nz.mem_171_sv2v_reg  <= data_i[3];
      \nz.mem_170_sv2v_reg  <= data_i[2];
      \nz.mem_169_sv2v_reg  <= data_i[1];
      \nz.mem_168_sv2v_reg  <= data_i[0];
    end 
    if(N811) begin
      \nz.mem_167_sv2v_reg  <= data_i[7];
      \nz.mem_166_sv2v_reg  <= data_i[6];
      \nz.mem_165_sv2v_reg  <= data_i[5];
      \nz.mem_164_sv2v_reg  <= data_i[4];
      \nz.mem_163_sv2v_reg  <= data_i[3];
      \nz.mem_162_sv2v_reg  <= data_i[2];
      \nz.mem_161_sv2v_reg  <= data_i[1];
      \nz.mem_160_sv2v_reg  <= data_i[0];
    end 
    if(N810) begin
      \nz.mem_159_sv2v_reg  <= data_i[7];
      \nz.mem_158_sv2v_reg  <= data_i[6];
      \nz.mem_157_sv2v_reg  <= data_i[5];
      \nz.mem_156_sv2v_reg  <= data_i[4];
      \nz.mem_155_sv2v_reg  <= data_i[3];
      \nz.mem_154_sv2v_reg  <= data_i[2];
      \nz.mem_153_sv2v_reg  <= data_i[1];
      \nz.mem_152_sv2v_reg  <= data_i[0];
    end 
    if(N809) begin
      \nz.mem_151_sv2v_reg  <= data_i[7];
      \nz.mem_150_sv2v_reg  <= data_i[6];
      \nz.mem_149_sv2v_reg  <= data_i[5];
      \nz.mem_148_sv2v_reg  <= data_i[4];
      \nz.mem_147_sv2v_reg  <= data_i[3];
      \nz.mem_146_sv2v_reg  <= data_i[2];
      \nz.mem_145_sv2v_reg  <= data_i[1];
      \nz.mem_144_sv2v_reg  <= data_i[0];
    end 
    if(N808) begin
      \nz.mem_143_sv2v_reg  <= data_i[7];
      \nz.mem_142_sv2v_reg  <= data_i[6];
      \nz.mem_141_sv2v_reg  <= data_i[5];
      \nz.mem_140_sv2v_reg  <= data_i[4];
      \nz.mem_139_sv2v_reg  <= data_i[3];
      \nz.mem_138_sv2v_reg  <= data_i[2];
      \nz.mem_137_sv2v_reg  <= data_i[1];
      \nz.mem_136_sv2v_reg  <= data_i[0];
    end 
    if(N807) begin
      \nz.mem_135_sv2v_reg  <= data_i[7];
      \nz.mem_134_sv2v_reg  <= data_i[6];
      \nz.mem_133_sv2v_reg  <= data_i[5];
      \nz.mem_132_sv2v_reg  <= data_i[4];
      \nz.mem_131_sv2v_reg  <= data_i[3];
      \nz.mem_130_sv2v_reg  <= data_i[2];
      \nz.mem_129_sv2v_reg  <= data_i[1];
      \nz.mem_128_sv2v_reg  <= data_i[0];
    end 
    if(N806) begin
      \nz.mem_127_sv2v_reg  <= data_i[7];
      \nz.mem_126_sv2v_reg  <= data_i[6];
      \nz.mem_125_sv2v_reg  <= data_i[5];
      \nz.mem_124_sv2v_reg  <= data_i[4];
      \nz.mem_123_sv2v_reg  <= data_i[3];
      \nz.mem_122_sv2v_reg  <= data_i[2];
      \nz.mem_121_sv2v_reg  <= data_i[1];
      \nz.mem_120_sv2v_reg  <= data_i[0];
    end 
    if(N805) begin
      \nz.mem_119_sv2v_reg  <= data_i[7];
      \nz.mem_118_sv2v_reg  <= data_i[6];
      \nz.mem_117_sv2v_reg  <= data_i[5];
      \nz.mem_116_sv2v_reg  <= data_i[4];
      \nz.mem_115_sv2v_reg  <= data_i[3];
      \nz.mem_114_sv2v_reg  <= data_i[2];
      \nz.mem_113_sv2v_reg  <= data_i[1];
      \nz.mem_112_sv2v_reg  <= data_i[0];
    end 
    if(N804) begin
      \nz.mem_111_sv2v_reg  <= data_i[7];
      \nz.mem_110_sv2v_reg  <= data_i[6];
      \nz.mem_109_sv2v_reg  <= data_i[5];
      \nz.mem_108_sv2v_reg  <= data_i[4];
      \nz.mem_107_sv2v_reg  <= data_i[3];
      \nz.mem_106_sv2v_reg  <= data_i[2];
      \nz.mem_105_sv2v_reg  <= data_i[1];
      \nz.mem_104_sv2v_reg  <= data_i[0];
    end 
    if(N803) begin
      \nz.mem_103_sv2v_reg  <= data_i[7];
      \nz.mem_102_sv2v_reg  <= data_i[6];
      \nz.mem_101_sv2v_reg  <= data_i[5];
      \nz.mem_100_sv2v_reg  <= data_i[4];
      \nz.mem_99_sv2v_reg  <= data_i[3];
      \nz.mem_98_sv2v_reg  <= data_i[2];
      \nz.mem_97_sv2v_reg  <= data_i[1];
      \nz.mem_96_sv2v_reg  <= data_i[0];
    end 
    if(N802) begin
      \nz.mem_95_sv2v_reg  <= data_i[7];
      \nz.mem_94_sv2v_reg  <= data_i[6];
      \nz.mem_93_sv2v_reg  <= data_i[5];
      \nz.mem_92_sv2v_reg  <= data_i[4];
      \nz.mem_91_sv2v_reg  <= data_i[3];
      \nz.mem_90_sv2v_reg  <= data_i[2];
      \nz.mem_89_sv2v_reg  <= data_i[1];
      \nz.mem_88_sv2v_reg  <= data_i[0];
    end 
    if(N801) begin
      \nz.mem_87_sv2v_reg  <= data_i[7];
      \nz.mem_86_sv2v_reg  <= data_i[6];
      \nz.mem_85_sv2v_reg  <= data_i[5];
      \nz.mem_84_sv2v_reg  <= data_i[4];
      \nz.mem_83_sv2v_reg  <= data_i[3];
      \nz.mem_82_sv2v_reg  <= data_i[2];
      \nz.mem_81_sv2v_reg  <= data_i[1];
      \nz.mem_80_sv2v_reg  <= data_i[0];
    end 
    if(N800) begin
      \nz.mem_79_sv2v_reg  <= data_i[7];
      \nz.mem_78_sv2v_reg  <= data_i[6];
      \nz.mem_77_sv2v_reg  <= data_i[5];
      \nz.mem_76_sv2v_reg  <= data_i[4];
      \nz.mem_75_sv2v_reg  <= data_i[3];
      \nz.mem_74_sv2v_reg  <= data_i[2];
      \nz.mem_73_sv2v_reg  <= data_i[1];
      \nz.mem_72_sv2v_reg  <= data_i[0];
    end 
    if(N799) begin
      \nz.mem_71_sv2v_reg  <= data_i[7];
      \nz.mem_70_sv2v_reg  <= data_i[6];
      \nz.mem_69_sv2v_reg  <= data_i[5];
      \nz.mem_68_sv2v_reg  <= data_i[4];
      \nz.mem_67_sv2v_reg  <= data_i[3];
      \nz.mem_66_sv2v_reg  <= data_i[2];
      \nz.mem_65_sv2v_reg  <= data_i[1];
      \nz.mem_64_sv2v_reg  <= data_i[0];
    end 
    if(N798) begin
      \nz.mem_63_sv2v_reg  <= data_i[7];
      \nz.mem_62_sv2v_reg  <= data_i[6];
      \nz.mem_61_sv2v_reg  <= data_i[5];
      \nz.mem_60_sv2v_reg  <= data_i[4];
      \nz.mem_59_sv2v_reg  <= data_i[3];
      \nz.mem_58_sv2v_reg  <= data_i[2];
      \nz.mem_57_sv2v_reg  <= data_i[1];
      \nz.mem_56_sv2v_reg  <= data_i[0];
    end 
    if(N797) begin
      \nz.mem_55_sv2v_reg  <= data_i[7];
      \nz.mem_54_sv2v_reg  <= data_i[6];
      \nz.mem_53_sv2v_reg  <= data_i[5];
      \nz.mem_52_sv2v_reg  <= data_i[4];
      \nz.mem_51_sv2v_reg  <= data_i[3];
      \nz.mem_50_sv2v_reg  <= data_i[2];
      \nz.mem_49_sv2v_reg  <= data_i[1];
      \nz.mem_48_sv2v_reg  <= data_i[0];
    end 
    if(N796) begin
      \nz.mem_47_sv2v_reg  <= data_i[7];
      \nz.mem_46_sv2v_reg  <= data_i[6];
      \nz.mem_45_sv2v_reg  <= data_i[5];
      \nz.mem_44_sv2v_reg  <= data_i[4];
      \nz.mem_43_sv2v_reg  <= data_i[3];
      \nz.mem_42_sv2v_reg  <= data_i[2];
      \nz.mem_41_sv2v_reg  <= data_i[1];
      \nz.mem_40_sv2v_reg  <= data_i[0];
    end 
    if(N795) begin
      \nz.mem_39_sv2v_reg  <= data_i[7];
      \nz.mem_38_sv2v_reg  <= data_i[6];
      \nz.mem_37_sv2v_reg  <= data_i[5];
      \nz.mem_36_sv2v_reg  <= data_i[4];
      \nz.mem_35_sv2v_reg  <= data_i[3];
      \nz.mem_34_sv2v_reg  <= data_i[2];
      \nz.mem_33_sv2v_reg  <= data_i[1];
      \nz.mem_32_sv2v_reg  <= data_i[0];
    end 
    if(N794) begin
      \nz.mem_31_sv2v_reg  <= data_i[7];
      \nz.mem_30_sv2v_reg  <= data_i[6];
      \nz.mem_29_sv2v_reg  <= data_i[5];
      \nz.mem_28_sv2v_reg  <= data_i[4];
      \nz.mem_27_sv2v_reg  <= data_i[3];
      \nz.mem_26_sv2v_reg  <= data_i[2];
      \nz.mem_25_sv2v_reg  <= data_i[1];
      \nz.mem_24_sv2v_reg  <= data_i[0];
    end 
    if(N793) begin
      \nz.mem_23_sv2v_reg  <= data_i[7];
      \nz.mem_22_sv2v_reg  <= data_i[6];
      \nz.mem_21_sv2v_reg  <= data_i[5];
      \nz.mem_20_sv2v_reg  <= data_i[4];
      \nz.mem_19_sv2v_reg  <= data_i[3];
      \nz.mem_18_sv2v_reg  <= data_i[2];
      \nz.mem_17_sv2v_reg  <= data_i[1];
      \nz.mem_16_sv2v_reg  <= data_i[0];
    end 
    if(N792) begin
      \nz.mem_15_sv2v_reg  <= data_i[7];
      \nz.mem_14_sv2v_reg  <= data_i[6];
      \nz.mem_13_sv2v_reg  <= data_i[5];
      \nz.mem_12_sv2v_reg  <= data_i[4];
      \nz.mem_11_sv2v_reg  <= data_i[3];
      \nz.mem_10_sv2v_reg  <= data_i[2];
      \nz.mem_9_sv2v_reg  <= data_i[1];
      \nz.mem_8_sv2v_reg  <= data_i[0];
    end 
    if(N791) begin
      \nz.mem_7_sv2v_reg  <= data_i[7];
      \nz.mem_6_sv2v_reg  <= data_i[6];
      \nz.mem_5_sv2v_reg  <= data_i[5];
      \nz.mem_4_sv2v_reg  <= data_i[4];
      \nz.mem_3_sv2v_reg  <= data_i[3];
      \nz.mem_2_sv2v_reg  <= data_i[2];
      \nz.mem_1_sv2v_reg  <= data_i[1];
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [7:0] addr_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [7:0] data_o;

  bsg_mem_1rw_sync_synth_width_p8_els_p256_latch_last_read_p1_verbose_p0
  synth
  (
    .clk_i(clk_i),
    .v_i(v_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p64
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;
  wire N0,N1,_0_net__0_,_1_net_,N2,N3,_2_net__0_,_3_net_,N4,_4_net__0_,_5_net_,N5,
  _6_net__0_,_7_net_,N6,_8_net__0_,_9_net_,N7,_10_net__0_,_11_net_,N8,_12_net__0_,
  _13_net_,N9,_14_net__0_,_15_net_,N10;

  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_0_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[7:0]),
    .addr_i(addr_i),
    .v_i(_0_net__0_),
    .w_i(_1_net_),
    .data_o(data_o[7:0])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_1_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[15:8]),
    .addr_i(addr_i),
    .v_i(_2_net__0_),
    .w_i(_3_net_),
    .data_o(data_o[15:8])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_2_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[23:16]),
    .addr_i(addr_i),
    .v_i(_4_net__0_),
    .w_i(_5_net_),
    .data_o(data_o[23:16])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_3_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[31:24]),
    .addr_i(addr_i),
    .v_i(_6_net__0_),
    .w_i(_7_net_),
    .data_o(data_o[31:24])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_4_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[39:32]),
    .addr_i(addr_i),
    .v_i(_8_net__0_),
    .w_i(_9_net_),
    .data_o(data_o[39:32])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_5_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[47:40]),
    .addr_i(addr_i),
    .v_i(_10_net__0_),
    .w_i(_11_net_),
    .data_o(data_o[47:40])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_6_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[55:48]),
    .addr_i(addr_i),
    .v_i(_12_net__0_),
    .w_i(_13_net_),
    .data_o(data_o[55:48])
  );


  bsg_mem_1rw_sync_width_p8_els_p256_latch_last_read_p1_addr_width_lp8_verbose_if_synth_p0
  \nz.bk_7_.mem_1rw_sync 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i[63:56]),
    .addr_i(addr_i),
    .v_i(_14_net__0_),
    .w_i(_15_net_),
    .data_o(data_o[63:56])
  );

  assign N3 = (N0)? write_mask_i[0] : 
              (N1)? 1'b1 : 1'b0;
  assign N0 = w_i;
  assign N1 = N2;
  assign N4 = (N0)? write_mask_i[1] : 
              (N1)? 1'b1 : 1'b0;
  assign N5 = (N0)? write_mask_i[2] : 
              (N1)? 1'b1 : 1'b0;
  assign N6 = (N0)? write_mask_i[3] : 
              (N1)? 1'b1 : 1'b0;
  assign N7 = (N0)? write_mask_i[4] : 
              (N1)? 1'b1 : 1'b0;
  assign N8 = (N0)? write_mask_i[5] : 
              (N1)? 1'b1 : 1'b0;
  assign N9 = (N0)? write_mask_i[6] : 
              (N1)? 1'b1 : 1'b0;
  assign N10 = (N0)? write_mask_i[7] : 
               (N1)? 1'b1 : 1'b0;
  assign _1_net_ = w_i & write_mask_i[0];
  assign N2 = ~w_i;
  assign _0_net__0_ = v_i & N3;
  assign _3_net_ = w_i & write_mask_i[1];
  assign _2_net__0_ = v_i & N4;
  assign _5_net_ = w_i & write_mask_i[2];
  assign _4_net__0_ = v_i & N5;
  assign _7_net_ = w_i & write_mask_i[3];
  assign _6_net__0_ = v_i & N6;
  assign _9_net_ = w_i & write_mask_i[4];
  assign _8_net__0_ = v_i & N7;
  assign _11_net_ = w_i & write_mask_i[5];
  assign _10_net__0_ = v_i & N8;
  assign _13_net_ = w_i & write_mask_i[6];
  assign _12_net__0_ = v_i & N9;
  assign _15_net_ = w_i & write_mask_i[7];
  assign _14_net__0_ = v_i & N10;

endmodule



module bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  v_i,
  w_i,
  addr_i,
  data_i,
  write_mask_i,
  data_o
);

  input [7:0] addr_i;
  input [63:0] data_i;
  input [7:0] write_mask_i;
  output [63:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [63:0] data_o;

  bsg_mem_1rw_sync_mask_write_byte_synth_els_p256_latch_last_read_p1_data_width_p64
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .w_i(w_i),
    .addr_i(addr_i),
    .data_i(data_i),
    .write_mask_i(write_mask_i),
    .data_o(data_o)
  );


endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p8_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [5:0] addr_i;
  input [7:0] w_mask_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [7:0] data_o,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,\nz.read_en ,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,
  \nz.llr.read_en_r ,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271;
  wire [5:0] \nz.addr_r ;
  wire [511:0] \nz.mem ;
  reg \nz.addr_r_5_sv2v_reg ,\nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,
  \nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,\nz.mem_511_sv2v_reg ,
  \nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,
  \nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,
  \nz.mem_500_sv2v_reg ,\nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,
  \nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,
  \nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,
  \nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,
  \nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,
  \nz.mem_460_sv2v_reg ,\nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,
  \nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,
  \nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,
  \nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,
  \nz.mem_420_sv2v_reg ,\nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,
  \nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,
  \nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,
  \nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,
  \nz.mem_380_sv2v_reg ,\nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,
  \nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,
  \nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,
  \nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,
  \nz.mem_340_sv2v_reg ,\nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,
  \nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,
  \nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,
  \nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,
  \nz.mem_300_sv2v_reg ,\nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,
  \nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,
  \nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,
  \nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,
  \nz.mem_260_sv2v_reg ,\nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,
  \nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,
  \nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,
  \nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,
  \nz.mem_220_sv2v_reg ,\nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,
  \nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,
  \nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [7] = (N83)? \nz.mem [7] : 
                            (N85)? \nz.mem [15] : 
                            (N87)? \nz.mem [23] : 
                            (N89)? \nz.mem [31] : 
                            (N91)? \nz.mem [39] : 
                            (N93)? \nz.mem [47] : 
                            (N95)? \nz.mem [55] : 
                            (N97)? \nz.mem [63] : 
                            (N99)? \nz.mem [71] : 
                            (N101)? \nz.mem [79] : 
                            (N103)? \nz.mem [87] : 
                            (N105)? \nz.mem [95] : 
                            (N107)? \nz.mem [103] : 
                            (N109)? \nz.mem [111] : 
                            (N111)? \nz.mem [119] : 
                            (N113)? \nz.mem [127] : 
                            (N115)? \nz.mem [135] : 
                            (N117)? \nz.mem [143] : 
                            (N119)? \nz.mem [151] : 
                            (N121)? \nz.mem [159] : 
                            (N123)? \nz.mem [167] : 
                            (N125)? \nz.mem [175] : 
                            (N127)? \nz.mem [183] : 
                            (N129)? \nz.mem [191] : 
                            (N131)? \nz.mem [199] : 
                            (N133)? \nz.mem [207] : 
                            (N135)? \nz.mem [215] : 
                            (N137)? \nz.mem [223] : 
                            (N139)? \nz.mem [231] : 
                            (N141)? \nz.mem [239] : 
                            (N143)? \nz.mem [247] : 
                            (N145)? \nz.mem [255] : 
                            (N84)? \nz.mem [263] : 
                            (N86)? \nz.mem [271] : 
                            (N88)? \nz.mem [279] : 
                            (N90)? \nz.mem [287] : 
                            (N92)? \nz.mem [295] : 
                            (N94)? \nz.mem [303] : 
                            (N96)? \nz.mem [311] : 
                            (N98)? \nz.mem [319] : 
                            (N100)? \nz.mem [327] : 
                            (N102)? \nz.mem [335] : 
                            (N104)? \nz.mem [343] : 
                            (N106)? \nz.mem [351] : 
                            (N108)? \nz.mem [359] : 
                            (N110)? \nz.mem [367] : 
                            (N112)? \nz.mem [375] : 
                            (N114)? \nz.mem [383] : 
                            (N116)? \nz.mem [391] : 
                            (N118)? \nz.mem [399] : 
                            (N120)? \nz.mem [407] : 
                            (N122)? \nz.mem [415] : 
                            (N124)? \nz.mem [423] : 
                            (N126)? \nz.mem [431] : 
                            (N128)? \nz.mem [439] : 
                            (N130)? \nz.mem [447] : 
                            (N132)? \nz.mem [455] : 
                            (N134)? \nz.mem [463] : 
                            (N136)? \nz.mem [471] : 
                            (N138)? \nz.mem [479] : 
                            (N140)? \nz.mem [487] : 
                            (N142)? \nz.mem [495] : 
                            (N144)? \nz.mem [503] : 
                            (N146)? \nz.mem [511] : 1'b0;
  assign \nz.data_out [6] = (N83)? \nz.mem [6] : 
                            (N85)? \nz.mem [14] : 
                            (N87)? \nz.mem [22] : 
                            (N89)? \nz.mem [30] : 
                            (N91)? \nz.mem [38] : 
                            (N93)? \nz.mem [46] : 
                            (N95)? \nz.mem [54] : 
                            (N97)? \nz.mem [62] : 
                            (N99)? \nz.mem [70] : 
                            (N101)? \nz.mem [78] : 
                            (N103)? \nz.mem [86] : 
                            (N105)? \nz.mem [94] : 
                            (N107)? \nz.mem [102] : 
                            (N109)? \nz.mem [110] : 
                            (N111)? \nz.mem [118] : 
                            (N113)? \nz.mem [126] : 
                            (N115)? \nz.mem [134] : 
                            (N117)? \nz.mem [142] : 
                            (N119)? \nz.mem [150] : 
                            (N121)? \nz.mem [158] : 
                            (N123)? \nz.mem [166] : 
                            (N125)? \nz.mem [174] : 
                            (N127)? \nz.mem [182] : 
                            (N129)? \nz.mem [190] : 
                            (N131)? \nz.mem [198] : 
                            (N133)? \nz.mem [206] : 
                            (N135)? \nz.mem [214] : 
                            (N137)? \nz.mem [222] : 
                            (N139)? \nz.mem [230] : 
                            (N141)? \nz.mem [238] : 
                            (N143)? \nz.mem [246] : 
                            (N145)? \nz.mem [254] : 
                            (N84)? \nz.mem [262] : 
                            (N86)? \nz.mem [270] : 
                            (N88)? \nz.mem [278] : 
                            (N90)? \nz.mem [286] : 
                            (N92)? \nz.mem [294] : 
                            (N94)? \nz.mem [302] : 
                            (N96)? \nz.mem [310] : 
                            (N98)? \nz.mem [318] : 
                            (N100)? \nz.mem [326] : 
                            (N102)? \nz.mem [334] : 
                            (N104)? \nz.mem [342] : 
                            (N106)? \nz.mem [350] : 
                            (N108)? \nz.mem [358] : 
                            (N110)? \nz.mem [366] : 
                            (N112)? \nz.mem [374] : 
                            (N114)? \nz.mem [382] : 
                            (N116)? \nz.mem [390] : 
                            (N118)? \nz.mem [398] : 
                            (N120)? \nz.mem [406] : 
                            (N122)? \nz.mem [414] : 
                            (N124)? \nz.mem [422] : 
                            (N126)? \nz.mem [430] : 
                            (N128)? \nz.mem [438] : 
                            (N130)? \nz.mem [446] : 
                            (N132)? \nz.mem [454] : 
                            (N134)? \nz.mem [462] : 
                            (N136)? \nz.mem [470] : 
                            (N138)? \nz.mem [478] : 
                            (N140)? \nz.mem [486] : 
                            (N142)? \nz.mem [494] : 
                            (N144)? \nz.mem [502] : 
                            (N146)? \nz.mem [510] : 1'b0;
  assign \nz.data_out [5] = (N83)? \nz.mem [5] : 
                            (N85)? \nz.mem [13] : 
                            (N87)? \nz.mem [21] : 
                            (N89)? \nz.mem [29] : 
                            (N91)? \nz.mem [37] : 
                            (N93)? \nz.mem [45] : 
                            (N95)? \nz.mem [53] : 
                            (N97)? \nz.mem [61] : 
                            (N99)? \nz.mem [69] : 
                            (N101)? \nz.mem [77] : 
                            (N103)? \nz.mem [85] : 
                            (N105)? \nz.mem [93] : 
                            (N107)? \nz.mem [101] : 
                            (N109)? \nz.mem [109] : 
                            (N111)? \nz.mem [117] : 
                            (N113)? \nz.mem [125] : 
                            (N115)? \nz.mem [133] : 
                            (N117)? \nz.mem [141] : 
                            (N119)? \nz.mem [149] : 
                            (N121)? \nz.mem [157] : 
                            (N123)? \nz.mem [165] : 
                            (N125)? \nz.mem [173] : 
                            (N127)? \nz.mem [181] : 
                            (N129)? \nz.mem [189] : 
                            (N131)? \nz.mem [197] : 
                            (N133)? \nz.mem [205] : 
                            (N135)? \nz.mem [213] : 
                            (N137)? \nz.mem [221] : 
                            (N139)? \nz.mem [229] : 
                            (N141)? \nz.mem [237] : 
                            (N143)? \nz.mem [245] : 
                            (N145)? \nz.mem [253] : 
                            (N84)? \nz.mem [261] : 
                            (N86)? \nz.mem [269] : 
                            (N88)? \nz.mem [277] : 
                            (N90)? \nz.mem [285] : 
                            (N92)? \nz.mem [293] : 
                            (N94)? \nz.mem [301] : 
                            (N96)? \nz.mem [309] : 
                            (N98)? \nz.mem [317] : 
                            (N100)? \nz.mem [325] : 
                            (N102)? \nz.mem [333] : 
                            (N104)? \nz.mem [341] : 
                            (N106)? \nz.mem [349] : 
                            (N108)? \nz.mem [357] : 
                            (N110)? \nz.mem [365] : 
                            (N112)? \nz.mem [373] : 
                            (N114)? \nz.mem [381] : 
                            (N116)? \nz.mem [389] : 
                            (N118)? \nz.mem [397] : 
                            (N120)? \nz.mem [405] : 
                            (N122)? \nz.mem [413] : 
                            (N124)? \nz.mem [421] : 
                            (N126)? \nz.mem [429] : 
                            (N128)? \nz.mem [437] : 
                            (N130)? \nz.mem [445] : 
                            (N132)? \nz.mem [453] : 
                            (N134)? \nz.mem [461] : 
                            (N136)? \nz.mem [469] : 
                            (N138)? \nz.mem [477] : 
                            (N140)? \nz.mem [485] : 
                            (N142)? \nz.mem [493] : 
                            (N144)? \nz.mem [501] : 
                            (N146)? \nz.mem [509] : 1'b0;
  assign \nz.data_out [4] = (N83)? \nz.mem [4] : 
                            (N85)? \nz.mem [12] : 
                            (N87)? \nz.mem [20] : 
                            (N89)? \nz.mem [28] : 
                            (N91)? \nz.mem [36] : 
                            (N93)? \nz.mem [44] : 
                            (N95)? \nz.mem [52] : 
                            (N97)? \nz.mem [60] : 
                            (N99)? \nz.mem [68] : 
                            (N101)? \nz.mem [76] : 
                            (N103)? \nz.mem [84] : 
                            (N105)? \nz.mem [92] : 
                            (N107)? \nz.mem [100] : 
                            (N109)? \nz.mem [108] : 
                            (N111)? \nz.mem [116] : 
                            (N113)? \nz.mem [124] : 
                            (N115)? \nz.mem [132] : 
                            (N117)? \nz.mem [140] : 
                            (N119)? \nz.mem [148] : 
                            (N121)? \nz.mem [156] : 
                            (N123)? \nz.mem [164] : 
                            (N125)? \nz.mem [172] : 
                            (N127)? \nz.mem [180] : 
                            (N129)? \nz.mem [188] : 
                            (N131)? \nz.mem [196] : 
                            (N133)? \nz.mem [204] : 
                            (N135)? \nz.mem [212] : 
                            (N137)? \nz.mem [220] : 
                            (N139)? \nz.mem [228] : 
                            (N141)? \nz.mem [236] : 
                            (N143)? \nz.mem [244] : 
                            (N145)? \nz.mem [252] : 
                            (N84)? \nz.mem [260] : 
                            (N86)? \nz.mem [268] : 
                            (N88)? \nz.mem [276] : 
                            (N90)? \nz.mem [284] : 
                            (N92)? \nz.mem [292] : 
                            (N94)? \nz.mem [300] : 
                            (N96)? \nz.mem [308] : 
                            (N98)? \nz.mem [316] : 
                            (N100)? \nz.mem [324] : 
                            (N102)? \nz.mem [332] : 
                            (N104)? \nz.mem [340] : 
                            (N106)? \nz.mem [348] : 
                            (N108)? \nz.mem [356] : 
                            (N110)? \nz.mem [364] : 
                            (N112)? \nz.mem [372] : 
                            (N114)? \nz.mem [380] : 
                            (N116)? \nz.mem [388] : 
                            (N118)? \nz.mem [396] : 
                            (N120)? \nz.mem [404] : 
                            (N122)? \nz.mem [412] : 
                            (N124)? \nz.mem [420] : 
                            (N126)? \nz.mem [428] : 
                            (N128)? \nz.mem [436] : 
                            (N130)? \nz.mem [444] : 
                            (N132)? \nz.mem [452] : 
                            (N134)? \nz.mem [460] : 
                            (N136)? \nz.mem [468] : 
                            (N138)? \nz.mem [476] : 
                            (N140)? \nz.mem [484] : 
                            (N142)? \nz.mem [492] : 
                            (N144)? \nz.mem [500] : 
                            (N146)? \nz.mem [508] : 1'b0;
  assign \nz.data_out [3] = (N83)? \nz.mem [3] : 
                            (N85)? \nz.mem [11] : 
                            (N87)? \nz.mem [19] : 
                            (N89)? \nz.mem [27] : 
                            (N91)? \nz.mem [35] : 
                            (N93)? \nz.mem [43] : 
                            (N95)? \nz.mem [51] : 
                            (N97)? \nz.mem [59] : 
                            (N99)? \nz.mem [67] : 
                            (N101)? \nz.mem [75] : 
                            (N103)? \nz.mem [83] : 
                            (N105)? \nz.mem [91] : 
                            (N107)? \nz.mem [99] : 
                            (N109)? \nz.mem [107] : 
                            (N111)? \nz.mem [115] : 
                            (N113)? \nz.mem [123] : 
                            (N115)? \nz.mem [131] : 
                            (N117)? \nz.mem [139] : 
                            (N119)? \nz.mem [147] : 
                            (N121)? \nz.mem [155] : 
                            (N123)? \nz.mem [163] : 
                            (N125)? \nz.mem [171] : 
                            (N127)? \nz.mem [179] : 
                            (N129)? \nz.mem [187] : 
                            (N131)? \nz.mem [195] : 
                            (N133)? \nz.mem [203] : 
                            (N135)? \nz.mem [211] : 
                            (N137)? \nz.mem [219] : 
                            (N139)? \nz.mem [227] : 
                            (N141)? \nz.mem [235] : 
                            (N143)? \nz.mem [243] : 
                            (N145)? \nz.mem [251] : 
                            (N84)? \nz.mem [259] : 
                            (N86)? \nz.mem [267] : 
                            (N88)? \nz.mem [275] : 
                            (N90)? \nz.mem [283] : 
                            (N92)? \nz.mem [291] : 
                            (N94)? \nz.mem [299] : 
                            (N96)? \nz.mem [307] : 
                            (N98)? \nz.mem [315] : 
                            (N100)? \nz.mem [323] : 
                            (N102)? \nz.mem [331] : 
                            (N104)? \nz.mem [339] : 
                            (N106)? \nz.mem [347] : 
                            (N108)? \nz.mem [355] : 
                            (N110)? \nz.mem [363] : 
                            (N112)? \nz.mem [371] : 
                            (N114)? \nz.mem [379] : 
                            (N116)? \nz.mem [387] : 
                            (N118)? \nz.mem [395] : 
                            (N120)? \nz.mem [403] : 
                            (N122)? \nz.mem [411] : 
                            (N124)? \nz.mem [419] : 
                            (N126)? \nz.mem [427] : 
                            (N128)? \nz.mem [435] : 
                            (N130)? \nz.mem [443] : 
                            (N132)? \nz.mem [451] : 
                            (N134)? \nz.mem [459] : 
                            (N136)? \nz.mem [467] : 
                            (N138)? \nz.mem [475] : 
                            (N140)? \nz.mem [483] : 
                            (N142)? \nz.mem [491] : 
                            (N144)? \nz.mem [499] : 
                            (N146)? \nz.mem [507] : 1'b0;
  assign \nz.data_out [2] = (N83)? \nz.mem [2] : 
                            (N85)? \nz.mem [10] : 
                            (N87)? \nz.mem [18] : 
                            (N89)? \nz.mem [26] : 
                            (N91)? \nz.mem [34] : 
                            (N93)? \nz.mem [42] : 
                            (N95)? \nz.mem [50] : 
                            (N97)? \nz.mem [58] : 
                            (N99)? \nz.mem [66] : 
                            (N101)? \nz.mem [74] : 
                            (N103)? \nz.mem [82] : 
                            (N105)? \nz.mem [90] : 
                            (N107)? \nz.mem [98] : 
                            (N109)? \nz.mem [106] : 
                            (N111)? \nz.mem [114] : 
                            (N113)? \nz.mem [122] : 
                            (N115)? \nz.mem [130] : 
                            (N117)? \nz.mem [138] : 
                            (N119)? \nz.mem [146] : 
                            (N121)? \nz.mem [154] : 
                            (N123)? \nz.mem [162] : 
                            (N125)? \nz.mem [170] : 
                            (N127)? \nz.mem [178] : 
                            (N129)? \nz.mem [186] : 
                            (N131)? \nz.mem [194] : 
                            (N133)? \nz.mem [202] : 
                            (N135)? \nz.mem [210] : 
                            (N137)? \nz.mem [218] : 
                            (N139)? \nz.mem [226] : 
                            (N141)? \nz.mem [234] : 
                            (N143)? \nz.mem [242] : 
                            (N145)? \nz.mem [250] : 
                            (N84)? \nz.mem [258] : 
                            (N86)? \nz.mem [266] : 
                            (N88)? \nz.mem [274] : 
                            (N90)? \nz.mem [282] : 
                            (N92)? \nz.mem [290] : 
                            (N94)? \nz.mem [298] : 
                            (N96)? \nz.mem [306] : 
                            (N98)? \nz.mem [314] : 
                            (N100)? \nz.mem [322] : 
                            (N102)? \nz.mem [330] : 
                            (N104)? \nz.mem [338] : 
                            (N106)? \nz.mem [346] : 
                            (N108)? \nz.mem [354] : 
                            (N110)? \nz.mem [362] : 
                            (N112)? \nz.mem [370] : 
                            (N114)? \nz.mem [378] : 
                            (N116)? \nz.mem [386] : 
                            (N118)? \nz.mem [394] : 
                            (N120)? \nz.mem [402] : 
                            (N122)? \nz.mem [410] : 
                            (N124)? \nz.mem [418] : 
                            (N126)? \nz.mem [426] : 
                            (N128)? \nz.mem [434] : 
                            (N130)? \nz.mem [442] : 
                            (N132)? \nz.mem [450] : 
                            (N134)? \nz.mem [458] : 
                            (N136)? \nz.mem [466] : 
                            (N138)? \nz.mem [474] : 
                            (N140)? \nz.mem [482] : 
                            (N142)? \nz.mem [490] : 
                            (N144)? \nz.mem [498] : 
                            (N146)? \nz.mem [506] : 1'b0;
  assign \nz.data_out [1] = (N83)? \nz.mem [1] : 
                            (N85)? \nz.mem [9] : 
                            (N87)? \nz.mem [17] : 
                            (N89)? \nz.mem [25] : 
                            (N91)? \nz.mem [33] : 
                            (N93)? \nz.mem [41] : 
                            (N95)? \nz.mem [49] : 
                            (N97)? \nz.mem [57] : 
                            (N99)? \nz.mem [65] : 
                            (N101)? \nz.mem [73] : 
                            (N103)? \nz.mem [81] : 
                            (N105)? \nz.mem [89] : 
                            (N107)? \nz.mem [97] : 
                            (N109)? \nz.mem [105] : 
                            (N111)? \nz.mem [113] : 
                            (N113)? \nz.mem [121] : 
                            (N115)? \nz.mem [129] : 
                            (N117)? \nz.mem [137] : 
                            (N119)? \nz.mem [145] : 
                            (N121)? \nz.mem [153] : 
                            (N123)? \nz.mem [161] : 
                            (N125)? \nz.mem [169] : 
                            (N127)? \nz.mem [177] : 
                            (N129)? \nz.mem [185] : 
                            (N131)? \nz.mem [193] : 
                            (N133)? \nz.mem [201] : 
                            (N135)? \nz.mem [209] : 
                            (N137)? \nz.mem [217] : 
                            (N139)? \nz.mem [225] : 
                            (N141)? \nz.mem [233] : 
                            (N143)? \nz.mem [241] : 
                            (N145)? \nz.mem [249] : 
                            (N84)? \nz.mem [257] : 
                            (N86)? \nz.mem [265] : 
                            (N88)? \nz.mem [273] : 
                            (N90)? \nz.mem [281] : 
                            (N92)? \nz.mem [289] : 
                            (N94)? \nz.mem [297] : 
                            (N96)? \nz.mem [305] : 
                            (N98)? \nz.mem [313] : 
                            (N100)? \nz.mem [321] : 
                            (N102)? \nz.mem [329] : 
                            (N104)? \nz.mem [337] : 
                            (N106)? \nz.mem [345] : 
                            (N108)? \nz.mem [353] : 
                            (N110)? \nz.mem [361] : 
                            (N112)? \nz.mem [369] : 
                            (N114)? \nz.mem [377] : 
                            (N116)? \nz.mem [385] : 
                            (N118)? \nz.mem [393] : 
                            (N120)? \nz.mem [401] : 
                            (N122)? \nz.mem [409] : 
                            (N124)? \nz.mem [417] : 
                            (N126)? \nz.mem [425] : 
                            (N128)? \nz.mem [433] : 
                            (N130)? \nz.mem [441] : 
                            (N132)? \nz.mem [449] : 
                            (N134)? \nz.mem [457] : 
                            (N136)? \nz.mem [465] : 
                            (N138)? \nz.mem [473] : 
                            (N140)? \nz.mem [481] : 
                            (N142)? \nz.mem [489] : 
                            (N144)? \nz.mem [497] : 
                            (N146)? \nz.mem [505] : 1'b0;
  assign \nz.data_out [0] = (N83)? \nz.mem [0] : 
                            (N85)? \nz.mem [8] : 
                            (N87)? \nz.mem [16] : 
                            (N89)? \nz.mem [24] : 
                            (N91)? \nz.mem [32] : 
                            (N93)? \nz.mem [40] : 
                            (N95)? \nz.mem [48] : 
                            (N97)? \nz.mem [56] : 
                            (N99)? \nz.mem [64] : 
                            (N101)? \nz.mem [72] : 
                            (N103)? \nz.mem [80] : 
                            (N105)? \nz.mem [88] : 
                            (N107)? \nz.mem [96] : 
                            (N109)? \nz.mem [104] : 
                            (N111)? \nz.mem [112] : 
                            (N113)? \nz.mem [120] : 
                            (N115)? \nz.mem [128] : 
                            (N117)? \nz.mem [136] : 
                            (N119)? \nz.mem [144] : 
                            (N121)? \nz.mem [152] : 
                            (N123)? \nz.mem [160] : 
                            (N125)? \nz.mem [168] : 
                            (N127)? \nz.mem [176] : 
                            (N129)? \nz.mem [184] : 
                            (N131)? \nz.mem [192] : 
                            (N133)? \nz.mem [200] : 
                            (N135)? \nz.mem [208] : 
                            (N137)? \nz.mem [216] : 
                            (N139)? \nz.mem [224] : 
                            (N141)? \nz.mem [232] : 
                            (N143)? \nz.mem [240] : 
                            (N145)? \nz.mem [248] : 
                            (N84)? \nz.mem [256] : 
                            (N86)? \nz.mem [264] : 
                            (N88)? \nz.mem [272] : 
                            (N90)? \nz.mem [280] : 
                            (N92)? \nz.mem [288] : 
                            (N94)? \nz.mem [296] : 
                            (N96)? \nz.mem [304] : 
                            (N98)? \nz.mem [312] : 
                            (N100)? \nz.mem [320] : 
                            (N102)? \nz.mem [328] : 
                            (N104)? \nz.mem [336] : 
                            (N106)? \nz.mem [344] : 
                            (N108)? \nz.mem [352] : 
                            (N110)? \nz.mem [360] : 
                            (N112)? \nz.mem [368] : 
                            (N114)? \nz.mem [376] : 
                            (N116)? \nz.mem [384] : 
                            (N118)? \nz.mem [392] : 
                            (N120)? \nz.mem [400] : 
                            (N122)? \nz.mem [408] : 
                            (N124)? \nz.mem [416] : 
                            (N126)? \nz.mem [424] : 
                            (N128)? \nz.mem [432] : 
                            (N130)? \nz.mem [440] : 
                            (N132)? \nz.mem [448] : 
                            (N134)? \nz.mem [456] : 
                            (N136)? \nz.mem [464] : 
                            (N138)? \nz.mem [472] : 
                            (N140)? \nz.mem [480] : 
                            (N142)? \nz.mem [488] : 
                            (N144)? \nz.mem [496] : 
                            (N146)? \nz.mem [504] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p8
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N1245 = ~addr_i[5];
  assign N1246 = addr_i[3] & addr_i[4];
  assign N1247 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N1248 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N1249 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N1250 = addr_i[5] & N1246;
  assign N1251 = addr_i[5] & N1247;
  assign N1252 = addr_i[5] & N1248;
  assign N1253 = addr_i[5] & N1249;
  assign N1254 = N1245 & N1246;
  assign N1255 = N1245 & N1247;
  assign N1256 = N1245 & N1248;
  assign N1257 = N1245 & N1249;
  assign N1258 = ~addr_i[2];
  assign N1259 = addr_i[0] & addr_i[1];
  assign N1260 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N1261 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N1262 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N1263 = addr_i[2] & N1259;
  assign N1264 = addr_i[2] & N1260;
  assign N1265 = addr_i[2] & N1261;
  assign N1266 = addr_i[2] & N1262;
  assign N1267 = N1258 & N1259;
  assign N1268 = N1258 & N1260;
  assign N1269 = N1258 & N1261;
  assign N1270 = N1258 & N1262;
  assign N668 = N1250 & N1263;
  assign N667 = N1250 & N1264;
  assign N666 = N1250 & N1265;
  assign N665 = N1250 & N1266;
  assign N664 = N1250 & N1267;
  assign N663 = N1250 & N1268;
  assign N662 = N1250 & N1269;
  assign N661 = N1250 & N1270;
  assign N660 = N1251 & N1263;
  assign N659 = N1251 & N1264;
  assign N658 = N1251 & N1265;
  assign N657 = N1251 & N1266;
  assign N656 = N1251 & N1267;
  assign N655 = N1251 & N1268;
  assign N654 = N1251 & N1269;
  assign N653 = N1251 & N1270;
  assign N652 = N1252 & N1263;
  assign N651 = N1252 & N1264;
  assign N650 = N1252 & N1265;
  assign N649 = N1252 & N1266;
  assign N648 = N1252 & N1267;
  assign N647 = N1252 & N1268;
  assign N646 = N1252 & N1269;
  assign N645 = N1252 & N1270;
  assign N644 = N1253 & N1263;
  assign N643 = N1253 & N1264;
  assign N642 = N1253 & N1265;
  assign N641 = N1253 & N1266;
  assign N640 = N1253 & N1267;
  assign N639 = N1253 & N1268;
  assign N638 = N1253 & N1269;
  assign N637 = N1253 & N1270;
  assign N636 = N1254 & N1263;
  assign N635 = N1254 & N1264;
  assign N634 = N1254 & N1265;
  assign N633 = N1254 & N1266;
  assign N632 = N1254 & N1267;
  assign N631 = N1254 & N1268;
  assign N630 = N1254 & N1269;
  assign N629 = N1254 & N1270;
  assign N628 = N1255 & N1263;
  assign N627 = N1255 & N1264;
  assign N626 = N1255 & N1265;
  assign N625 = N1255 & N1266;
  assign N624 = N1255 & N1267;
  assign N623 = N1255 & N1268;
  assign N622 = N1255 & N1269;
  assign N621 = N1255 & N1270;
  assign N620 = N1256 & N1263;
  assign N619 = N1256 & N1264;
  assign N618 = N1256 & N1265;
  assign N617 = N1256 & N1266;
  assign N616 = N1256 & N1267;
  assign N615 = N1256 & N1268;
  assign N614 = N1256 & N1269;
  assign N613 = N1256 & N1270;
  assign N612 = N1257 & N1263;
  assign N611 = N1257 & N1264;
  assign N610 = N1257 & N1265;
  assign N609 = N1257 & N1266;
  assign N608 = N1257 & N1267;
  assign N607 = N1257 & N1268;
  assign N606 = N1257 & N1269;
  assign N605 = N1257 & N1270;
  assign { N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150 } = (N8)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N149)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215 } = (N9)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N214)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280 } = (N10)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N279)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345 } = (N11)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N344)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410 } = (N12)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N409)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475 } = (N13)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N474)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540 } = (N14)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N539)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669 } = (N15)? { N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N604)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = w_mask_i[7];
  assign { N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733 } = (N16)? { N732, N603, N538, N473, N408, N343, N278, N213, N731, N602, N537, N472, N407, N342, N277, N212, N730, N601, N536, N471, N406, N341, N276, N211, N729, N600, N535, N470, N405, N340, N275, N210, N728, N599, N534, N469, N404, N339, N274, N209, N727, N598, N533, N468, N403, N338, N273, N208, N726, N597, N532, N467, N402, N337, N272, N207, N725, N596, N531, N466, N401, N336, N271, N206, N724, N595, N530, N465, N400, N335, N270, N205, N723, N594, N529, N464, N399, N334, N269, N204, N722, N593, N528, N463, N398, N333, N268, N203, N721, N592, N527, N462, N397, N332, N267, N202, N720, N591, N526, N461, N396, N331, N266, N201, N719, N590, N525, N460, N395, N330, N265, N200, N718, N589, N524, N459, N394, N329, N264, N199, N717, N588, N523, N458, N393, N328, N263, N198, N716, N587, N522, N457, N392, N327, N262, N197, N715, N586, N521, N456, N391, N326, N261, N196, N714, N585, N520, N455, N390, N325, N260, N195, N713, N584, N519, N454, N389, N324, N259, N194, N712, N583, N518, N453, N388, N323, N258, N193, N711, N582, N517, N452, N387, N322, N257, N192, N710, N581, N516, N451, N386, N321, N256, N191, N709, N580, N515, N450, N385, N320, N255, N190, N708, N579, N514, N449, N384, N319, N254, N189, N707, N578, N513, N448, N383, N318, N253, N188, N706, N577, N512, N447, N382, N317, N252, N187, N705, N576, N511, N446, N381, N316, N251, N186, N704, N575, N510, N445, N380, N315, N250, N185, N703, N574, N509, N444, N379, N314, N249, N184, N702, N573, N508, N443, N378, N313, N248, N183, N701, N572, N507, N442, N377, N312, N247, N182, N700, N571, N506, N441, N376, N311, N246, N181, N699, N570, N505, N440, N375, N310, N245, N180, N698, N569, N504, N439, N374, N309, N244, N179, N697, N568, N503, N438, N373, N308, N243, N178, N696, N567, N502, N437, N372, N307, N242, N177, N695, N566, N501, N436, N371, N306, N241, N176, N694, N565, N500, N435, N370, N305, N240, N175, N693, N564, N499, N434, N369, N304, N239, N174, N692, N563, N498, N433, N368, N303, N238, N173, N691, N562, N497, N432, N367, N302, N237, N172, N690, N561, N496, N431, N366, N301, N236, N171, N689, N560, N495, N430, N365, N300, N235, N170, N688, N559, N494, N429, N364, N299, N234, N169, N687, N558, N493, N428, N363, N298, N233, N168, N686, N557, N492, N427, N362, N297, N232, N167, N685, N556, N491, N426, N361, N296, N231, N166, N684, N555, N490, N425, N360, N295, N230, N165, N683, N554, N489, N424, N359, N294, N229, N164, N682, N553, N488, N423, N358, N293, N228, N163, N681, N552, N487, N422, N357, N292, N227, N162, N680, N551, N486, N421, N356, N291, N226, N161, N679, N550, N485, N420, N355, N290, N225, N160, N678, N549, N484, N419, N354, N289, N224, N159, N677, N548, N483, N418, N353, N288, N223, N158, N676, N547, N482, N417, N352, N287, N222, N157, N675, N546, N481, N416, N351, N286, N221, N156, N674, N545, N480, N415, N350, N285, N220, N155, N673, N544, N479, N414, N349, N284, N219, N154, N672, N543, N478, N413, N348, N283, N218, N153, N671, N542, N477, N412, N347, N282, N217, N152, N670, N541, N476, N411, N346, N281, N216, N151, N669, N540, N475, N410, N345, N280, N215, N150 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   (N148)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = N147;
  assign \nz.read_en  = v_i & N1271;
  assign N1271 = ~w_i;
  assign N17 = ~\nz.addr_r [0];
  assign N18 = ~\nz.addr_r [1];
  assign N19 = N17 & N18;
  assign N20 = N17 & \nz.addr_r [1];
  assign N21 = \nz.addr_r [0] & N18;
  assign N22 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N23 = ~\nz.addr_r [2];
  assign N24 = N19 & N23;
  assign N25 = N19 & \nz.addr_r [2];
  assign N26 = N21 & N23;
  assign N27 = N21 & \nz.addr_r [2];
  assign N28 = N20 & N23;
  assign N29 = N20 & \nz.addr_r [2];
  assign N30 = N22 & N23;
  assign N31 = N22 & \nz.addr_r [2];
  assign N32 = ~\nz.addr_r [3];
  assign N33 = N24 & N32;
  assign N34 = N24 & \nz.addr_r [3];
  assign N35 = N26 & N32;
  assign N36 = N26 & \nz.addr_r [3];
  assign N37 = N28 & N32;
  assign N38 = N28 & \nz.addr_r [3];
  assign N39 = N30 & N32;
  assign N40 = N30 & \nz.addr_r [3];
  assign N41 = N25 & N32;
  assign N42 = N25 & \nz.addr_r [3];
  assign N43 = N27 & N32;
  assign N44 = N27 & \nz.addr_r [3];
  assign N45 = N29 & N32;
  assign N46 = N29 & \nz.addr_r [3];
  assign N47 = N31 & N32;
  assign N48 = N31 & \nz.addr_r [3];
  assign N49 = ~\nz.addr_r [4];
  assign N50 = N33 & N49;
  assign N51 = N33 & \nz.addr_r [4];
  assign N52 = N35 & N49;
  assign N53 = N35 & \nz.addr_r [4];
  assign N54 = N37 & N49;
  assign N55 = N37 & \nz.addr_r [4];
  assign N56 = N39 & N49;
  assign N57 = N39 & \nz.addr_r [4];
  assign N58 = N41 & N49;
  assign N59 = N41 & \nz.addr_r [4];
  assign N60 = N43 & N49;
  assign N61 = N43 & \nz.addr_r [4];
  assign N62 = N45 & N49;
  assign N63 = N45 & \nz.addr_r [4];
  assign N64 = N47 & N49;
  assign N65 = N47 & \nz.addr_r [4];
  assign N66 = N34 & N49;
  assign N67 = N34 & \nz.addr_r [4];
  assign N68 = N36 & N49;
  assign N69 = N36 & \nz.addr_r [4];
  assign N70 = N38 & N49;
  assign N71 = N38 & \nz.addr_r [4];
  assign N72 = N40 & N49;
  assign N73 = N40 & \nz.addr_r [4];
  assign N74 = N42 & N49;
  assign N75 = N42 & \nz.addr_r [4];
  assign N76 = N44 & N49;
  assign N77 = N44 & \nz.addr_r [4];
  assign N78 = N46 & N49;
  assign N79 = N46 & \nz.addr_r [4];
  assign N80 = N48 & N49;
  assign N81 = N48 & \nz.addr_r [4];
  assign N82 = ~\nz.addr_r [5];
  assign N83 = N50 & N82;
  assign N84 = N50 & \nz.addr_r [5];
  assign N85 = N52 & N82;
  assign N86 = N52 & \nz.addr_r [5];
  assign N87 = N54 & N82;
  assign N88 = N54 & \nz.addr_r [5];
  assign N89 = N56 & N82;
  assign N90 = N56 & \nz.addr_r [5];
  assign N91 = N58 & N82;
  assign N92 = N58 & \nz.addr_r [5];
  assign N93 = N60 & N82;
  assign N94 = N60 & \nz.addr_r [5];
  assign N95 = N62 & N82;
  assign N96 = N62 & \nz.addr_r [5];
  assign N97 = N64 & N82;
  assign N98 = N64 & \nz.addr_r [5];
  assign N99 = N66 & N82;
  assign N100 = N66 & \nz.addr_r [5];
  assign N101 = N68 & N82;
  assign N102 = N68 & \nz.addr_r [5];
  assign N103 = N70 & N82;
  assign N104 = N70 & \nz.addr_r [5];
  assign N105 = N72 & N82;
  assign N106 = N72 & \nz.addr_r [5];
  assign N107 = N74 & N82;
  assign N108 = N74 & \nz.addr_r [5];
  assign N109 = N76 & N82;
  assign N110 = N76 & \nz.addr_r [5];
  assign N111 = N78 & N82;
  assign N112 = N78 & \nz.addr_r [5];
  assign N113 = N80 & N82;
  assign N114 = N80 & \nz.addr_r [5];
  assign N115 = N51 & N82;
  assign N116 = N51 & \nz.addr_r [5];
  assign N117 = N53 & N82;
  assign N118 = N53 & \nz.addr_r [5];
  assign N119 = N55 & N82;
  assign N120 = N55 & \nz.addr_r [5];
  assign N121 = N57 & N82;
  assign N122 = N57 & \nz.addr_r [5];
  assign N123 = N59 & N82;
  assign N124 = N59 & \nz.addr_r [5];
  assign N125 = N61 & N82;
  assign N126 = N61 & \nz.addr_r [5];
  assign N127 = N63 & N82;
  assign N128 = N63 & \nz.addr_r [5];
  assign N129 = N65 & N82;
  assign N130 = N65 & \nz.addr_r [5];
  assign N131 = N67 & N82;
  assign N132 = N67 & \nz.addr_r [5];
  assign N133 = N69 & N82;
  assign N134 = N69 & \nz.addr_r [5];
  assign N135 = N71 & N82;
  assign N136 = N71 & \nz.addr_r [5];
  assign N137 = N73 & N82;
  assign N138 = N73 & \nz.addr_r [5];
  assign N139 = N75 & N82;
  assign N140 = N75 & \nz.addr_r [5];
  assign N141 = N77 & N82;
  assign N142 = N77 & \nz.addr_r [5];
  assign N143 = N79 & N82;
  assign N144 = N79 & \nz.addr_r [5];
  assign N145 = N81 & N82;
  assign N146 = N81 & \nz.addr_r [5];
  assign N147 = v_i & w_i;
  assign N148 = ~N147;
  assign N149 = ~w_mask_i[0];
  assign N214 = ~w_mask_i[1];
  assign N279 = ~w_mask_i[2];
  assign N344 = ~w_mask_i[3];
  assign N409 = ~w_mask_i[4];
  assign N474 = ~w_mask_i[5];
  assign N539 = ~w_mask_i[6];
  assign N604 = ~w_mask_i[7];

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N1244) begin
      \nz.mem_511_sv2v_reg  <= data_i[7];
    end 
    if(N1243) begin
      \nz.mem_510_sv2v_reg  <= data_i[6];
    end 
    if(N1242) begin
      \nz.mem_509_sv2v_reg  <= data_i[5];
    end 
    if(N1241) begin
      \nz.mem_508_sv2v_reg  <= data_i[4];
    end 
    if(N1240) begin
      \nz.mem_507_sv2v_reg  <= data_i[3];
    end 
    if(N1239) begin
      \nz.mem_506_sv2v_reg  <= data_i[2];
    end 
    if(N1238) begin
      \nz.mem_505_sv2v_reg  <= data_i[1];
    end 
    if(N1237) begin
      \nz.mem_504_sv2v_reg  <= data_i[0];
    end 
    if(N1236) begin
      \nz.mem_503_sv2v_reg  <= data_i[7];
    end 
    if(N1235) begin
      \nz.mem_502_sv2v_reg  <= data_i[6];
    end 
    if(N1234) begin
      \nz.mem_501_sv2v_reg  <= data_i[5];
    end 
    if(N1233) begin
      \nz.mem_500_sv2v_reg  <= data_i[4];
    end 
    if(N1232) begin
      \nz.mem_499_sv2v_reg  <= data_i[3];
    end 
    if(N1231) begin
      \nz.mem_498_sv2v_reg  <= data_i[2];
    end 
    if(N1230) begin
      \nz.mem_497_sv2v_reg  <= data_i[1];
    end 
    if(N1229) begin
      \nz.mem_496_sv2v_reg  <= data_i[0];
    end 
    if(N1228) begin
      \nz.mem_495_sv2v_reg  <= data_i[7];
    end 
    if(N1227) begin
      \nz.mem_494_sv2v_reg  <= data_i[6];
    end 
    if(N1226) begin
      \nz.mem_493_sv2v_reg  <= data_i[5];
    end 
    if(N1225) begin
      \nz.mem_492_sv2v_reg  <= data_i[4];
    end 
    if(N1224) begin
      \nz.mem_491_sv2v_reg  <= data_i[3];
    end 
    if(N1223) begin
      \nz.mem_490_sv2v_reg  <= data_i[2];
    end 
    if(N1222) begin
      \nz.mem_489_sv2v_reg  <= data_i[1];
    end 
    if(N1221) begin
      \nz.mem_488_sv2v_reg  <= data_i[0];
    end 
    if(N1220) begin
      \nz.mem_487_sv2v_reg  <= data_i[7];
    end 
    if(N1219) begin
      \nz.mem_486_sv2v_reg  <= data_i[6];
    end 
    if(N1218) begin
      \nz.mem_485_sv2v_reg  <= data_i[5];
    end 
    if(N1217) begin
      \nz.mem_484_sv2v_reg  <= data_i[4];
    end 
    if(N1216) begin
      \nz.mem_483_sv2v_reg  <= data_i[3];
    end 
    if(N1215) begin
      \nz.mem_482_sv2v_reg  <= data_i[2];
    end 
    if(N1214) begin
      \nz.mem_481_sv2v_reg  <= data_i[1];
    end 
    if(N1213) begin
      \nz.mem_480_sv2v_reg  <= data_i[0];
    end 
    if(N1212) begin
      \nz.mem_479_sv2v_reg  <= data_i[7];
    end 
    if(N1211) begin
      \nz.mem_478_sv2v_reg  <= data_i[6];
    end 
    if(N1210) begin
      \nz.mem_477_sv2v_reg  <= data_i[5];
    end 
    if(N1209) begin
      \nz.mem_476_sv2v_reg  <= data_i[4];
    end 
    if(N1208) begin
      \nz.mem_475_sv2v_reg  <= data_i[3];
    end 
    if(N1207) begin
      \nz.mem_474_sv2v_reg  <= data_i[2];
    end 
    if(N1206) begin
      \nz.mem_473_sv2v_reg  <= data_i[1];
    end 
    if(N1205) begin
      \nz.mem_472_sv2v_reg  <= data_i[0];
    end 
    if(N1204) begin
      \nz.mem_471_sv2v_reg  <= data_i[7];
    end 
    if(N1203) begin
      \nz.mem_470_sv2v_reg  <= data_i[6];
    end 
    if(N1202) begin
      \nz.mem_469_sv2v_reg  <= data_i[5];
    end 
    if(N1201) begin
      \nz.mem_468_sv2v_reg  <= data_i[4];
    end 
    if(N1200) begin
      \nz.mem_467_sv2v_reg  <= data_i[3];
    end 
    if(N1199) begin
      \nz.mem_466_sv2v_reg  <= data_i[2];
    end 
    if(N1198) begin
      \nz.mem_465_sv2v_reg  <= data_i[1];
    end 
    if(N1197) begin
      \nz.mem_464_sv2v_reg  <= data_i[0];
    end 
    if(N1196) begin
      \nz.mem_463_sv2v_reg  <= data_i[7];
    end 
    if(N1195) begin
      \nz.mem_462_sv2v_reg  <= data_i[6];
    end 
    if(N1194) begin
      \nz.mem_461_sv2v_reg  <= data_i[5];
    end 
    if(N1193) begin
      \nz.mem_460_sv2v_reg  <= data_i[4];
    end 
    if(N1192) begin
      \nz.mem_459_sv2v_reg  <= data_i[3];
    end 
    if(N1191) begin
      \nz.mem_458_sv2v_reg  <= data_i[2];
    end 
    if(N1190) begin
      \nz.mem_457_sv2v_reg  <= data_i[1];
    end 
    if(N1189) begin
      \nz.mem_456_sv2v_reg  <= data_i[0];
    end 
    if(N1188) begin
      \nz.mem_455_sv2v_reg  <= data_i[7];
    end 
    if(N1187) begin
      \nz.mem_454_sv2v_reg  <= data_i[6];
    end 
    if(N1186) begin
      \nz.mem_453_sv2v_reg  <= data_i[5];
    end 
    if(N1185) begin
      \nz.mem_452_sv2v_reg  <= data_i[4];
    end 
    if(N1184) begin
      \nz.mem_451_sv2v_reg  <= data_i[3];
    end 
    if(N1183) begin
      \nz.mem_450_sv2v_reg  <= data_i[2];
    end 
    if(N1182) begin
      \nz.mem_449_sv2v_reg  <= data_i[1];
    end 
    if(N1181) begin
      \nz.mem_448_sv2v_reg  <= data_i[0];
    end 
    if(N1180) begin
      \nz.mem_447_sv2v_reg  <= data_i[7];
    end 
    if(N1179) begin
      \nz.mem_446_sv2v_reg  <= data_i[6];
    end 
    if(N1178) begin
      \nz.mem_445_sv2v_reg  <= data_i[5];
    end 
    if(N1177) begin
      \nz.mem_444_sv2v_reg  <= data_i[4];
    end 
    if(N1176) begin
      \nz.mem_443_sv2v_reg  <= data_i[3];
    end 
    if(N1175) begin
      \nz.mem_442_sv2v_reg  <= data_i[2];
    end 
    if(N1174) begin
      \nz.mem_441_sv2v_reg  <= data_i[1];
    end 
    if(N1173) begin
      \nz.mem_440_sv2v_reg  <= data_i[0];
    end 
    if(N1172) begin
      \nz.mem_439_sv2v_reg  <= data_i[7];
    end 
    if(N1171) begin
      \nz.mem_438_sv2v_reg  <= data_i[6];
    end 
    if(N1170) begin
      \nz.mem_437_sv2v_reg  <= data_i[5];
    end 
    if(N1169) begin
      \nz.mem_436_sv2v_reg  <= data_i[4];
    end 
    if(N1168) begin
      \nz.mem_435_sv2v_reg  <= data_i[3];
    end 
    if(N1167) begin
      \nz.mem_434_sv2v_reg  <= data_i[2];
    end 
    if(N1166) begin
      \nz.mem_433_sv2v_reg  <= data_i[1];
    end 
    if(N1165) begin
      \nz.mem_432_sv2v_reg  <= data_i[0];
    end 
    if(N1164) begin
      \nz.mem_431_sv2v_reg  <= data_i[7];
    end 
    if(N1163) begin
      \nz.mem_430_sv2v_reg  <= data_i[6];
    end 
    if(N1162) begin
      \nz.mem_429_sv2v_reg  <= data_i[5];
    end 
    if(N1161) begin
      \nz.mem_428_sv2v_reg  <= data_i[4];
    end 
    if(N1160) begin
      \nz.mem_427_sv2v_reg  <= data_i[3];
    end 
    if(N1159) begin
      \nz.mem_426_sv2v_reg  <= data_i[2];
    end 
    if(N1158) begin
      \nz.mem_425_sv2v_reg  <= data_i[1];
    end 
    if(N1157) begin
      \nz.mem_424_sv2v_reg  <= data_i[0];
    end 
    if(N1156) begin
      \nz.mem_423_sv2v_reg  <= data_i[7];
    end 
    if(N1155) begin
      \nz.mem_422_sv2v_reg  <= data_i[6];
    end 
    if(N1154) begin
      \nz.mem_421_sv2v_reg  <= data_i[5];
    end 
    if(N1153) begin
      \nz.mem_420_sv2v_reg  <= data_i[4];
    end 
    if(N1152) begin
      \nz.mem_419_sv2v_reg  <= data_i[3];
    end 
    if(N1151) begin
      \nz.mem_418_sv2v_reg  <= data_i[2];
    end 
    if(N1150) begin
      \nz.mem_417_sv2v_reg  <= data_i[1];
    end 
    if(N1149) begin
      \nz.mem_416_sv2v_reg  <= data_i[0];
    end 
    if(N1148) begin
      \nz.mem_415_sv2v_reg  <= data_i[7];
    end 
    if(N1147) begin
      \nz.mem_414_sv2v_reg  <= data_i[6];
    end 
    if(N1146) begin
      \nz.mem_413_sv2v_reg  <= data_i[5];
    end 
    if(N1145) begin
      \nz.mem_412_sv2v_reg  <= data_i[4];
    end 
    if(N1144) begin
      \nz.mem_411_sv2v_reg  <= data_i[3];
    end 
    if(N1143) begin
      \nz.mem_410_sv2v_reg  <= data_i[2];
    end 
    if(N1142) begin
      \nz.mem_409_sv2v_reg  <= data_i[1];
    end 
    if(N1141) begin
      \nz.mem_408_sv2v_reg  <= data_i[0];
    end 
    if(N1140) begin
      \nz.mem_407_sv2v_reg  <= data_i[7];
    end 
    if(N1139) begin
      \nz.mem_406_sv2v_reg  <= data_i[6];
    end 
    if(N1138) begin
      \nz.mem_405_sv2v_reg  <= data_i[5];
    end 
    if(N1137) begin
      \nz.mem_404_sv2v_reg  <= data_i[4];
    end 
    if(N1136) begin
      \nz.mem_403_sv2v_reg  <= data_i[3];
    end 
    if(N1135) begin
      \nz.mem_402_sv2v_reg  <= data_i[2];
    end 
    if(N1134) begin
      \nz.mem_401_sv2v_reg  <= data_i[1];
    end 
    if(N1133) begin
      \nz.mem_400_sv2v_reg  <= data_i[0];
    end 
    if(N1132) begin
      \nz.mem_399_sv2v_reg  <= data_i[7];
    end 
    if(N1131) begin
      \nz.mem_398_sv2v_reg  <= data_i[6];
    end 
    if(N1130) begin
      \nz.mem_397_sv2v_reg  <= data_i[5];
    end 
    if(N1129) begin
      \nz.mem_396_sv2v_reg  <= data_i[4];
    end 
    if(N1128) begin
      \nz.mem_395_sv2v_reg  <= data_i[3];
    end 
    if(N1127) begin
      \nz.mem_394_sv2v_reg  <= data_i[2];
    end 
    if(N1126) begin
      \nz.mem_393_sv2v_reg  <= data_i[1];
    end 
    if(N1125) begin
      \nz.mem_392_sv2v_reg  <= data_i[0];
    end 
    if(N1124) begin
      \nz.mem_391_sv2v_reg  <= data_i[7];
    end 
    if(N1123) begin
      \nz.mem_390_sv2v_reg  <= data_i[6];
    end 
    if(N1122) begin
      \nz.mem_389_sv2v_reg  <= data_i[5];
    end 
    if(N1121) begin
      \nz.mem_388_sv2v_reg  <= data_i[4];
    end 
    if(N1120) begin
      \nz.mem_387_sv2v_reg  <= data_i[3];
    end 
    if(N1119) begin
      \nz.mem_386_sv2v_reg  <= data_i[2];
    end 
    if(N1118) begin
      \nz.mem_385_sv2v_reg  <= data_i[1];
    end 
    if(N1117) begin
      \nz.mem_384_sv2v_reg  <= data_i[0];
    end 
    if(N1116) begin
      \nz.mem_383_sv2v_reg  <= data_i[7];
    end 
    if(N1115) begin
      \nz.mem_382_sv2v_reg  <= data_i[6];
    end 
    if(N1114) begin
      \nz.mem_381_sv2v_reg  <= data_i[5];
    end 
    if(N1113) begin
      \nz.mem_380_sv2v_reg  <= data_i[4];
    end 
    if(N1112) begin
      \nz.mem_379_sv2v_reg  <= data_i[3];
    end 
    if(N1111) begin
      \nz.mem_378_sv2v_reg  <= data_i[2];
    end 
    if(N1110) begin
      \nz.mem_377_sv2v_reg  <= data_i[1];
    end 
    if(N1109) begin
      \nz.mem_376_sv2v_reg  <= data_i[0];
    end 
    if(N1108) begin
      \nz.mem_375_sv2v_reg  <= data_i[7];
    end 
    if(N1107) begin
      \nz.mem_374_sv2v_reg  <= data_i[6];
    end 
    if(N1106) begin
      \nz.mem_373_sv2v_reg  <= data_i[5];
    end 
    if(N1105) begin
      \nz.mem_372_sv2v_reg  <= data_i[4];
    end 
    if(N1104) begin
      \nz.mem_371_sv2v_reg  <= data_i[3];
    end 
    if(N1103) begin
      \nz.mem_370_sv2v_reg  <= data_i[2];
    end 
    if(N1102) begin
      \nz.mem_369_sv2v_reg  <= data_i[1];
    end 
    if(N1101) begin
      \nz.mem_368_sv2v_reg  <= data_i[0];
    end 
    if(N1100) begin
      \nz.mem_367_sv2v_reg  <= data_i[7];
    end 
    if(N1099) begin
      \nz.mem_366_sv2v_reg  <= data_i[6];
    end 
    if(N1098) begin
      \nz.mem_365_sv2v_reg  <= data_i[5];
    end 
    if(N1097) begin
      \nz.mem_364_sv2v_reg  <= data_i[4];
    end 
    if(N1096) begin
      \nz.mem_363_sv2v_reg  <= data_i[3];
    end 
    if(N1095) begin
      \nz.mem_362_sv2v_reg  <= data_i[2];
    end 
    if(N1094) begin
      \nz.mem_361_sv2v_reg  <= data_i[1];
    end 
    if(N1093) begin
      \nz.mem_360_sv2v_reg  <= data_i[0];
    end 
    if(N1092) begin
      \nz.mem_359_sv2v_reg  <= data_i[7];
    end 
    if(N1091) begin
      \nz.mem_358_sv2v_reg  <= data_i[6];
    end 
    if(N1090) begin
      \nz.mem_357_sv2v_reg  <= data_i[5];
    end 
    if(N1089) begin
      \nz.mem_356_sv2v_reg  <= data_i[4];
    end 
    if(N1088) begin
      \nz.mem_355_sv2v_reg  <= data_i[3];
    end 
    if(N1087) begin
      \nz.mem_354_sv2v_reg  <= data_i[2];
    end 
    if(N1086) begin
      \nz.mem_353_sv2v_reg  <= data_i[1];
    end 
    if(N1085) begin
      \nz.mem_352_sv2v_reg  <= data_i[0];
    end 
    if(N1084) begin
      \nz.mem_351_sv2v_reg  <= data_i[7];
    end 
    if(N1083) begin
      \nz.mem_350_sv2v_reg  <= data_i[6];
    end 
    if(N1082) begin
      \nz.mem_349_sv2v_reg  <= data_i[5];
    end 
    if(N1081) begin
      \nz.mem_348_sv2v_reg  <= data_i[4];
    end 
    if(N1080) begin
      \nz.mem_347_sv2v_reg  <= data_i[3];
    end 
    if(N1079) begin
      \nz.mem_346_sv2v_reg  <= data_i[2];
    end 
    if(N1078) begin
      \nz.mem_345_sv2v_reg  <= data_i[1];
    end 
    if(N1077) begin
      \nz.mem_344_sv2v_reg  <= data_i[0];
    end 
    if(N1076) begin
      \nz.mem_343_sv2v_reg  <= data_i[7];
    end 
    if(N1075) begin
      \nz.mem_342_sv2v_reg  <= data_i[6];
    end 
    if(N1074) begin
      \nz.mem_341_sv2v_reg  <= data_i[5];
    end 
    if(N1073) begin
      \nz.mem_340_sv2v_reg  <= data_i[4];
    end 
    if(N1072) begin
      \nz.mem_339_sv2v_reg  <= data_i[3];
    end 
    if(N1071) begin
      \nz.mem_338_sv2v_reg  <= data_i[2];
    end 
    if(N1070) begin
      \nz.mem_337_sv2v_reg  <= data_i[1];
    end 
    if(N1069) begin
      \nz.mem_336_sv2v_reg  <= data_i[0];
    end 
    if(N1068) begin
      \nz.mem_335_sv2v_reg  <= data_i[7];
    end 
    if(N1067) begin
      \nz.mem_334_sv2v_reg  <= data_i[6];
    end 
    if(N1066) begin
      \nz.mem_333_sv2v_reg  <= data_i[5];
    end 
    if(N1065) begin
      \nz.mem_332_sv2v_reg  <= data_i[4];
    end 
    if(N1064) begin
      \nz.mem_331_sv2v_reg  <= data_i[3];
    end 
    if(N1063) begin
      \nz.mem_330_sv2v_reg  <= data_i[2];
    end 
    if(N1062) begin
      \nz.mem_329_sv2v_reg  <= data_i[1];
    end 
    if(N1061) begin
      \nz.mem_328_sv2v_reg  <= data_i[0];
    end 
    if(N1060) begin
      \nz.mem_327_sv2v_reg  <= data_i[7];
    end 
    if(N1059) begin
      \nz.mem_326_sv2v_reg  <= data_i[6];
    end 
    if(N1058) begin
      \nz.mem_325_sv2v_reg  <= data_i[5];
    end 
    if(N1057) begin
      \nz.mem_324_sv2v_reg  <= data_i[4];
    end 
    if(N1056) begin
      \nz.mem_323_sv2v_reg  <= data_i[3];
    end 
    if(N1055) begin
      \nz.mem_322_sv2v_reg  <= data_i[2];
    end 
    if(N1054) begin
      \nz.mem_321_sv2v_reg  <= data_i[1];
    end 
    if(N1053) begin
      \nz.mem_320_sv2v_reg  <= data_i[0];
    end 
    if(N1052) begin
      \nz.mem_319_sv2v_reg  <= data_i[7];
    end 
    if(N1051) begin
      \nz.mem_318_sv2v_reg  <= data_i[6];
    end 
    if(N1050) begin
      \nz.mem_317_sv2v_reg  <= data_i[5];
    end 
    if(N1049) begin
      \nz.mem_316_sv2v_reg  <= data_i[4];
    end 
    if(N1048) begin
      \nz.mem_315_sv2v_reg  <= data_i[3];
    end 
    if(N1047) begin
      \nz.mem_314_sv2v_reg  <= data_i[2];
    end 
    if(N1046) begin
      \nz.mem_313_sv2v_reg  <= data_i[1];
    end 
    if(N1045) begin
      \nz.mem_312_sv2v_reg  <= data_i[0];
    end 
    if(N1044) begin
      \nz.mem_311_sv2v_reg  <= data_i[7];
    end 
    if(N1043) begin
      \nz.mem_310_sv2v_reg  <= data_i[6];
    end 
    if(N1042) begin
      \nz.mem_309_sv2v_reg  <= data_i[5];
    end 
    if(N1041) begin
      \nz.mem_308_sv2v_reg  <= data_i[4];
    end 
    if(N1040) begin
      \nz.mem_307_sv2v_reg  <= data_i[3];
    end 
    if(N1039) begin
      \nz.mem_306_sv2v_reg  <= data_i[2];
    end 
    if(N1038) begin
      \nz.mem_305_sv2v_reg  <= data_i[1];
    end 
    if(N1037) begin
      \nz.mem_304_sv2v_reg  <= data_i[0];
    end 
    if(N1036) begin
      \nz.mem_303_sv2v_reg  <= data_i[7];
    end 
    if(N1035) begin
      \nz.mem_302_sv2v_reg  <= data_i[6];
    end 
    if(N1034) begin
      \nz.mem_301_sv2v_reg  <= data_i[5];
    end 
    if(N1033) begin
      \nz.mem_300_sv2v_reg  <= data_i[4];
    end 
    if(N1032) begin
      \nz.mem_299_sv2v_reg  <= data_i[3];
    end 
    if(N1031) begin
      \nz.mem_298_sv2v_reg  <= data_i[2];
    end 
    if(N1030) begin
      \nz.mem_297_sv2v_reg  <= data_i[1];
    end 
    if(N1029) begin
      \nz.mem_296_sv2v_reg  <= data_i[0];
    end 
    if(N1028) begin
      \nz.mem_295_sv2v_reg  <= data_i[7];
    end 
    if(N1027) begin
      \nz.mem_294_sv2v_reg  <= data_i[6];
    end 
    if(N1026) begin
      \nz.mem_293_sv2v_reg  <= data_i[5];
    end 
    if(N1025) begin
      \nz.mem_292_sv2v_reg  <= data_i[4];
    end 
    if(N1024) begin
      \nz.mem_291_sv2v_reg  <= data_i[3];
    end 
    if(N1023) begin
      \nz.mem_290_sv2v_reg  <= data_i[2];
    end 
    if(N1022) begin
      \nz.mem_289_sv2v_reg  <= data_i[1];
    end 
    if(N1021) begin
      \nz.mem_288_sv2v_reg  <= data_i[0];
    end 
    if(N1020) begin
      \nz.mem_287_sv2v_reg  <= data_i[7];
    end 
    if(N1019) begin
      \nz.mem_286_sv2v_reg  <= data_i[6];
    end 
    if(N1018) begin
      \nz.mem_285_sv2v_reg  <= data_i[5];
    end 
    if(N1017) begin
      \nz.mem_284_sv2v_reg  <= data_i[4];
    end 
    if(N1016) begin
      \nz.mem_283_sv2v_reg  <= data_i[3];
    end 
    if(N1015) begin
      \nz.mem_282_sv2v_reg  <= data_i[2];
    end 
    if(N1014) begin
      \nz.mem_281_sv2v_reg  <= data_i[1];
    end 
    if(N1013) begin
      \nz.mem_280_sv2v_reg  <= data_i[0];
    end 
    if(N1012) begin
      \nz.mem_279_sv2v_reg  <= data_i[7];
    end 
    if(N1011) begin
      \nz.mem_278_sv2v_reg  <= data_i[6];
    end 
    if(N1010) begin
      \nz.mem_277_sv2v_reg  <= data_i[5];
    end 
    if(N1009) begin
      \nz.mem_276_sv2v_reg  <= data_i[4];
    end 
    if(N1008) begin
      \nz.mem_275_sv2v_reg  <= data_i[3];
    end 
    if(N1007) begin
      \nz.mem_274_sv2v_reg  <= data_i[2];
    end 
    if(N1006) begin
      \nz.mem_273_sv2v_reg  <= data_i[1];
    end 
    if(N1005) begin
      \nz.mem_272_sv2v_reg  <= data_i[0];
    end 
    if(N1004) begin
      \nz.mem_271_sv2v_reg  <= data_i[7];
    end 
    if(N1003) begin
      \nz.mem_270_sv2v_reg  <= data_i[6];
    end 
    if(N1002) begin
      \nz.mem_269_sv2v_reg  <= data_i[5];
    end 
    if(N1001) begin
      \nz.mem_268_sv2v_reg  <= data_i[4];
    end 
    if(N1000) begin
      \nz.mem_267_sv2v_reg  <= data_i[3];
    end 
    if(N999) begin
      \nz.mem_266_sv2v_reg  <= data_i[2];
    end 
    if(N998) begin
      \nz.mem_265_sv2v_reg  <= data_i[1];
    end 
    if(N997) begin
      \nz.mem_264_sv2v_reg  <= data_i[0];
    end 
    if(N996) begin
      \nz.mem_263_sv2v_reg  <= data_i[7];
    end 
    if(N995) begin
      \nz.mem_262_sv2v_reg  <= data_i[6];
    end 
    if(N994) begin
      \nz.mem_261_sv2v_reg  <= data_i[5];
    end 
    if(N993) begin
      \nz.mem_260_sv2v_reg  <= data_i[4];
    end 
    if(N992) begin
      \nz.mem_259_sv2v_reg  <= data_i[3];
    end 
    if(N991) begin
      \nz.mem_258_sv2v_reg  <= data_i[2];
    end 
    if(N990) begin
      \nz.mem_257_sv2v_reg  <= data_i[1];
    end 
    if(N989) begin
      \nz.mem_256_sv2v_reg  <= data_i[0];
    end 
    if(N988) begin
      \nz.mem_255_sv2v_reg  <= data_i[7];
    end 
    if(N987) begin
      \nz.mem_254_sv2v_reg  <= data_i[6];
    end 
    if(N986) begin
      \nz.mem_253_sv2v_reg  <= data_i[5];
    end 
    if(N985) begin
      \nz.mem_252_sv2v_reg  <= data_i[4];
    end 
    if(N984) begin
      \nz.mem_251_sv2v_reg  <= data_i[3];
    end 
    if(N983) begin
      \nz.mem_250_sv2v_reg  <= data_i[2];
    end 
    if(N982) begin
      \nz.mem_249_sv2v_reg  <= data_i[1];
    end 
    if(N981) begin
      \nz.mem_248_sv2v_reg  <= data_i[0];
    end 
    if(N980) begin
      \nz.mem_247_sv2v_reg  <= data_i[7];
    end 
    if(N979) begin
      \nz.mem_246_sv2v_reg  <= data_i[6];
    end 
    if(N978) begin
      \nz.mem_245_sv2v_reg  <= data_i[5];
    end 
    if(N977) begin
      \nz.mem_244_sv2v_reg  <= data_i[4];
    end 
    if(N976) begin
      \nz.mem_243_sv2v_reg  <= data_i[3];
    end 
    if(N975) begin
      \nz.mem_242_sv2v_reg  <= data_i[2];
    end 
    if(N974) begin
      \nz.mem_241_sv2v_reg  <= data_i[1];
    end 
    if(N973) begin
      \nz.mem_240_sv2v_reg  <= data_i[0];
    end 
    if(N972) begin
      \nz.mem_239_sv2v_reg  <= data_i[7];
    end 
    if(N971) begin
      \nz.mem_238_sv2v_reg  <= data_i[6];
    end 
    if(N970) begin
      \nz.mem_237_sv2v_reg  <= data_i[5];
    end 
    if(N969) begin
      \nz.mem_236_sv2v_reg  <= data_i[4];
    end 
    if(N968) begin
      \nz.mem_235_sv2v_reg  <= data_i[3];
    end 
    if(N967) begin
      \nz.mem_234_sv2v_reg  <= data_i[2];
    end 
    if(N966) begin
      \nz.mem_233_sv2v_reg  <= data_i[1];
    end 
    if(N965) begin
      \nz.mem_232_sv2v_reg  <= data_i[0];
    end 
    if(N964) begin
      \nz.mem_231_sv2v_reg  <= data_i[7];
    end 
    if(N963) begin
      \nz.mem_230_sv2v_reg  <= data_i[6];
    end 
    if(N962) begin
      \nz.mem_229_sv2v_reg  <= data_i[5];
    end 
    if(N961) begin
      \nz.mem_228_sv2v_reg  <= data_i[4];
    end 
    if(N960) begin
      \nz.mem_227_sv2v_reg  <= data_i[3];
    end 
    if(N959) begin
      \nz.mem_226_sv2v_reg  <= data_i[2];
    end 
    if(N958) begin
      \nz.mem_225_sv2v_reg  <= data_i[1];
    end 
    if(N957) begin
      \nz.mem_224_sv2v_reg  <= data_i[0];
    end 
    if(N956) begin
      \nz.mem_223_sv2v_reg  <= data_i[7];
    end 
    if(N955) begin
      \nz.mem_222_sv2v_reg  <= data_i[6];
    end 
    if(N954) begin
      \nz.mem_221_sv2v_reg  <= data_i[5];
    end 
    if(N953) begin
      \nz.mem_220_sv2v_reg  <= data_i[4];
    end 
    if(N952) begin
      \nz.mem_219_sv2v_reg  <= data_i[3];
    end 
    if(N951) begin
      \nz.mem_218_sv2v_reg  <= data_i[2];
    end 
    if(N950) begin
      \nz.mem_217_sv2v_reg  <= data_i[1];
    end 
    if(N949) begin
      \nz.mem_216_sv2v_reg  <= data_i[0];
    end 
    if(N948) begin
      \nz.mem_215_sv2v_reg  <= data_i[7];
    end 
    if(N947) begin
      \nz.mem_214_sv2v_reg  <= data_i[6];
    end 
    if(N946) begin
      \nz.mem_213_sv2v_reg  <= data_i[5];
    end 
    if(N945) begin
      \nz.mem_212_sv2v_reg  <= data_i[4];
    end 
    if(N944) begin
      \nz.mem_211_sv2v_reg  <= data_i[3];
    end 
    if(N943) begin
      \nz.mem_210_sv2v_reg  <= data_i[2];
    end 
    if(N942) begin
      \nz.mem_209_sv2v_reg  <= data_i[1];
    end 
    if(N941) begin
      \nz.mem_208_sv2v_reg  <= data_i[0];
    end 
    if(N940) begin
      \nz.mem_207_sv2v_reg  <= data_i[7];
    end 
    if(N939) begin
      \nz.mem_206_sv2v_reg  <= data_i[6];
    end 
    if(N938) begin
      \nz.mem_205_sv2v_reg  <= data_i[5];
    end 
    if(N937) begin
      \nz.mem_204_sv2v_reg  <= data_i[4];
    end 
    if(N936) begin
      \nz.mem_203_sv2v_reg  <= data_i[3];
    end 
    if(N935) begin
      \nz.mem_202_sv2v_reg  <= data_i[2];
    end 
    if(N934) begin
      \nz.mem_201_sv2v_reg  <= data_i[1];
    end 
    if(N933) begin
      \nz.mem_200_sv2v_reg  <= data_i[0];
    end 
    if(N932) begin
      \nz.mem_199_sv2v_reg  <= data_i[7];
    end 
    if(N931) begin
      \nz.mem_198_sv2v_reg  <= data_i[6];
    end 
    if(N930) begin
      \nz.mem_197_sv2v_reg  <= data_i[5];
    end 
    if(N929) begin
      \nz.mem_196_sv2v_reg  <= data_i[4];
    end 
    if(N928) begin
      \nz.mem_195_sv2v_reg  <= data_i[3];
    end 
    if(N927) begin
      \nz.mem_194_sv2v_reg  <= data_i[2];
    end 
    if(N926) begin
      \nz.mem_193_sv2v_reg  <= data_i[1];
    end 
    if(N925) begin
      \nz.mem_192_sv2v_reg  <= data_i[0];
    end 
    if(N924) begin
      \nz.mem_191_sv2v_reg  <= data_i[7];
    end 
    if(N923) begin
      \nz.mem_190_sv2v_reg  <= data_i[6];
    end 
    if(N922) begin
      \nz.mem_189_sv2v_reg  <= data_i[5];
    end 
    if(N921) begin
      \nz.mem_188_sv2v_reg  <= data_i[4];
    end 
    if(N920) begin
      \nz.mem_187_sv2v_reg  <= data_i[3];
    end 
    if(N919) begin
      \nz.mem_186_sv2v_reg  <= data_i[2];
    end 
    if(N918) begin
      \nz.mem_185_sv2v_reg  <= data_i[1];
    end 
    if(N917) begin
      \nz.mem_184_sv2v_reg  <= data_i[0];
    end 
    if(N916) begin
      \nz.mem_183_sv2v_reg  <= data_i[7];
    end 
    if(N915) begin
      \nz.mem_182_sv2v_reg  <= data_i[6];
    end 
    if(N914) begin
      \nz.mem_181_sv2v_reg  <= data_i[5];
    end 
    if(N913) begin
      \nz.mem_180_sv2v_reg  <= data_i[4];
    end 
    if(N912) begin
      \nz.mem_179_sv2v_reg  <= data_i[3];
    end 
    if(N911) begin
      \nz.mem_178_sv2v_reg  <= data_i[2];
    end 
    if(N910) begin
      \nz.mem_177_sv2v_reg  <= data_i[1];
    end 
    if(N909) begin
      \nz.mem_176_sv2v_reg  <= data_i[0];
    end 
    if(N908) begin
      \nz.mem_175_sv2v_reg  <= data_i[7];
    end 
    if(N907) begin
      \nz.mem_174_sv2v_reg  <= data_i[6];
    end 
    if(N906) begin
      \nz.mem_173_sv2v_reg  <= data_i[5];
    end 
    if(N905) begin
      \nz.mem_172_sv2v_reg  <= data_i[4];
    end 
    if(N904) begin
      \nz.mem_171_sv2v_reg  <= data_i[3];
    end 
    if(N903) begin
      \nz.mem_170_sv2v_reg  <= data_i[2];
    end 
    if(N902) begin
      \nz.mem_169_sv2v_reg  <= data_i[1];
    end 
    if(N901) begin
      \nz.mem_168_sv2v_reg  <= data_i[0];
    end 
    if(N900) begin
      \nz.mem_167_sv2v_reg  <= data_i[7];
    end 
    if(N899) begin
      \nz.mem_166_sv2v_reg  <= data_i[6];
    end 
    if(N898) begin
      \nz.mem_165_sv2v_reg  <= data_i[5];
    end 
    if(N897) begin
      \nz.mem_164_sv2v_reg  <= data_i[4];
    end 
    if(N896) begin
      \nz.mem_163_sv2v_reg  <= data_i[3];
    end 
    if(N895) begin
      \nz.mem_162_sv2v_reg  <= data_i[2];
    end 
    if(N894) begin
      \nz.mem_161_sv2v_reg  <= data_i[1];
    end 
    if(N893) begin
      \nz.mem_160_sv2v_reg  <= data_i[0];
    end 
    if(N892) begin
      \nz.mem_159_sv2v_reg  <= data_i[7];
    end 
    if(N891) begin
      \nz.mem_158_sv2v_reg  <= data_i[6];
    end 
    if(N890) begin
      \nz.mem_157_sv2v_reg  <= data_i[5];
    end 
    if(N889) begin
      \nz.mem_156_sv2v_reg  <= data_i[4];
    end 
    if(N888) begin
      \nz.mem_155_sv2v_reg  <= data_i[3];
    end 
    if(N887) begin
      \nz.mem_154_sv2v_reg  <= data_i[2];
    end 
    if(N886) begin
      \nz.mem_153_sv2v_reg  <= data_i[1];
    end 
    if(N885) begin
      \nz.mem_152_sv2v_reg  <= data_i[0];
    end 
    if(N884) begin
      \nz.mem_151_sv2v_reg  <= data_i[7];
    end 
    if(N883) begin
      \nz.mem_150_sv2v_reg  <= data_i[6];
    end 
    if(N882) begin
      \nz.mem_149_sv2v_reg  <= data_i[5];
    end 
    if(N881) begin
      \nz.mem_148_sv2v_reg  <= data_i[4];
    end 
    if(N880) begin
      \nz.mem_147_sv2v_reg  <= data_i[3];
    end 
    if(N879) begin
      \nz.mem_146_sv2v_reg  <= data_i[2];
    end 
    if(N878) begin
      \nz.mem_145_sv2v_reg  <= data_i[1];
    end 
    if(N877) begin
      \nz.mem_144_sv2v_reg  <= data_i[0];
    end 
    if(N876) begin
      \nz.mem_143_sv2v_reg  <= data_i[7];
    end 
    if(N875) begin
      \nz.mem_142_sv2v_reg  <= data_i[6];
    end 
    if(N874) begin
      \nz.mem_141_sv2v_reg  <= data_i[5];
    end 
    if(N873) begin
      \nz.mem_140_sv2v_reg  <= data_i[4];
    end 
    if(N872) begin
      \nz.mem_139_sv2v_reg  <= data_i[3];
    end 
    if(N871) begin
      \nz.mem_138_sv2v_reg  <= data_i[2];
    end 
    if(N870) begin
      \nz.mem_137_sv2v_reg  <= data_i[1];
    end 
    if(N869) begin
      \nz.mem_136_sv2v_reg  <= data_i[0];
    end 
    if(N868) begin
      \nz.mem_135_sv2v_reg  <= data_i[7];
    end 
    if(N867) begin
      \nz.mem_134_sv2v_reg  <= data_i[6];
    end 
    if(N866) begin
      \nz.mem_133_sv2v_reg  <= data_i[5];
    end 
    if(N865) begin
      \nz.mem_132_sv2v_reg  <= data_i[4];
    end 
    if(N864) begin
      \nz.mem_131_sv2v_reg  <= data_i[3];
    end 
    if(N863) begin
      \nz.mem_130_sv2v_reg  <= data_i[2];
    end 
    if(N862) begin
      \nz.mem_129_sv2v_reg  <= data_i[1];
    end 
    if(N861) begin
      \nz.mem_128_sv2v_reg  <= data_i[0];
    end 
    if(N860) begin
      \nz.mem_127_sv2v_reg  <= data_i[7];
    end 
    if(N859) begin
      \nz.mem_126_sv2v_reg  <= data_i[6];
    end 
    if(N858) begin
      \nz.mem_125_sv2v_reg  <= data_i[5];
    end 
    if(N857) begin
      \nz.mem_124_sv2v_reg  <= data_i[4];
    end 
    if(N856) begin
      \nz.mem_123_sv2v_reg  <= data_i[3];
    end 
    if(N855) begin
      \nz.mem_122_sv2v_reg  <= data_i[2];
    end 
    if(N854) begin
      \nz.mem_121_sv2v_reg  <= data_i[1];
    end 
    if(N853) begin
      \nz.mem_120_sv2v_reg  <= data_i[0];
    end 
    if(N852) begin
      \nz.mem_119_sv2v_reg  <= data_i[7];
    end 
    if(N851) begin
      \nz.mem_118_sv2v_reg  <= data_i[6];
    end 
    if(N850) begin
      \nz.mem_117_sv2v_reg  <= data_i[5];
    end 
    if(N849) begin
      \nz.mem_116_sv2v_reg  <= data_i[4];
    end 
    if(N848) begin
      \nz.mem_115_sv2v_reg  <= data_i[3];
    end 
    if(N847) begin
      \nz.mem_114_sv2v_reg  <= data_i[2];
    end 
    if(N846) begin
      \nz.mem_113_sv2v_reg  <= data_i[1];
    end 
    if(N845) begin
      \nz.mem_112_sv2v_reg  <= data_i[0];
    end 
    if(N844) begin
      \nz.mem_111_sv2v_reg  <= data_i[7];
    end 
    if(N843) begin
      \nz.mem_110_sv2v_reg  <= data_i[6];
    end 
    if(N842) begin
      \nz.mem_109_sv2v_reg  <= data_i[5];
    end 
    if(N841) begin
      \nz.mem_108_sv2v_reg  <= data_i[4];
    end 
    if(N840) begin
      \nz.mem_107_sv2v_reg  <= data_i[3];
    end 
    if(N839) begin
      \nz.mem_106_sv2v_reg  <= data_i[2];
    end 
    if(N838) begin
      \nz.mem_105_sv2v_reg  <= data_i[1];
    end 
    if(N837) begin
      \nz.mem_104_sv2v_reg  <= data_i[0];
    end 
    if(N836) begin
      \nz.mem_103_sv2v_reg  <= data_i[7];
    end 
    if(N835) begin
      \nz.mem_102_sv2v_reg  <= data_i[6];
    end 
    if(N834) begin
      \nz.mem_101_sv2v_reg  <= data_i[5];
    end 
    if(N833) begin
      \nz.mem_100_sv2v_reg  <= data_i[4];
    end 
    if(N832) begin
      \nz.mem_99_sv2v_reg  <= data_i[3];
    end 
    if(N831) begin
      \nz.mem_98_sv2v_reg  <= data_i[2];
    end 
    if(N830) begin
      \nz.mem_97_sv2v_reg  <= data_i[1];
    end 
    if(N829) begin
      \nz.mem_96_sv2v_reg  <= data_i[0];
    end 
    if(N828) begin
      \nz.mem_95_sv2v_reg  <= data_i[7];
    end 
    if(N827) begin
      \nz.mem_94_sv2v_reg  <= data_i[6];
    end 
    if(N826) begin
      \nz.mem_93_sv2v_reg  <= data_i[5];
    end 
    if(N825) begin
      \nz.mem_92_sv2v_reg  <= data_i[4];
    end 
    if(N824) begin
      \nz.mem_91_sv2v_reg  <= data_i[3];
    end 
    if(N823) begin
      \nz.mem_90_sv2v_reg  <= data_i[2];
    end 
    if(N822) begin
      \nz.mem_89_sv2v_reg  <= data_i[1];
    end 
    if(N821) begin
      \nz.mem_88_sv2v_reg  <= data_i[0];
    end 
    if(N820) begin
      \nz.mem_87_sv2v_reg  <= data_i[7];
    end 
    if(N819) begin
      \nz.mem_86_sv2v_reg  <= data_i[6];
    end 
    if(N818) begin
      \nz.mem_85_sv2v_reg  <= data_i[5];
    end 
    if(N817) begin
      \nz.mem_84_sv2v_reg  <= data_i[4];
    end 
    if(N816) begin
      \nz.mem_83_sv2v_reg  <= data_i[3];
    end 
    if(N815) begin
      \nz.mem_82_sv2v_reg  <= data_i[2];
    end 
    if(N814) begin
      \nz.mem_81_sv2v_reg  <= data_i[1];
    end 
    if(N813) begin
      \nz.mem_80_sv2v_reg  <= data_i[0];
    end 
    if(N812) begin
      \nz.mem_79_sv2v_reg  <= data_i[7];
    end 
    if(N811) begin
      \nz.mem_78_sv2v_reg  <= data_i[6];
    end 
    if(N810) begin
      \nz.mem_77_sv2v_reg  <= data_i[5];
    end 
    if(N809) begin
      \nz.mem_76_sv2v_reg  <= data_i[4];
    end 
    if(N808) begin
      \nz.mem_75_sv2v_reg  <= data_i[3];
    end 
    if(N807) begin
      \nz.mem_74_sv2v_reg  <= data_i[2];
    end 
    if(N806) begin
      \nz.mem_73_sv2v_reg  <= data_i[1];
    end 
    if(N805) begin
      \nz.mem_72_sv2v_reg  <= data_i[0];
    end 
    if(N804) begin
      \nz.mem_71_sv2v_reg  <= data_i[7];
    end 
    if(N803) begin
      \nz.mem_70_sv2v_reg  <= data_i[6];
    end 
    if(N802) begin
      \nz.mem_69_sv2v_reg  <= data_i[5];
    end 
    if(N801) begin
      \nz.mem_68_sv2v_reg  <= data_i[4];
    end 
    if(N800) begin
      \nz.mem_67_sv2v_reg  <= data_i[3];
    end 
    if(N799) begin
      \nz.mem_66_sv2v_reg  <= data_i[2];
    end 
    if(N798) begin
      \nz.mem_65_sv2v_reg  <= data_i[1];
    end 
    if(N797) begin
      \nz.mem_64_sv2v_reg  <= data_i[0];
    end 
    if(N796) begin
      \nz.mem_63_sv2v_reg  <= data_i[7];
    end 
    if(N795) begin
      \nz.mem_62_sv2v_reg  <= data_i[6];
    end 
    if(N794) begin
      \nz.mem_61_sv2v_reg  <= data_i[5];
    end 
    if(N793) begin
      \nz.mem_60_sv2v_reg  <= data_i[4];
    end 
    if(N792) begin
      \nz.mem_59_sv2v_reg  <= data_i[3];
    end 
    if(N791) begin
      \nz.mem_58_sv2v_reg  <= data_i[2];
    end 
    if(N790) begin
      \nz.mem_57_sv2v_reg  <= data_i[1];
    end 
    if(N789) begin
      \nz.mem_56_sv2v_reg  <= data_i[0];
    end 
    if(N788) begin
      \nz.mem_55_sv2v_reg  <= data_i[7];
    end 
    if(N787) begin
      \nz.mem_54_sv2v_reg  <= data_i[6];
    end 
    if(N786) begin
      \nz.mem_53_sv2v_reg  <= data_i[5];
    end 
    if(N785) begin
      \nz.mem_52_sv2v_reg  <= data_i[4];
    end 
    if(N784) begin
      \nz.mem_51_sv2v_reg  <= data_i[3];
    end 
    if(N783) begin
      \nz.mem_50_sv2v_reg  <= data_i[2];
    end 
    if(N782) begin
      \nz.mem_49_sv2v_reg  <= data_i[1];
    end 
    if(N781) begin
      \nz.mem_48_sv2v_reg  <= data_i[0];
    end 
    if(N780) begin
      \nz.mem_47_sv2v_reg  <= data_i[7];
    end 
    if(N779) begin
      \nz.mem_46_sv2v_reg  <= data_i[6];
    end 
    if(N778) begin
      \nz.mem_45_sv2v_reg  <= data_i[5];
    end 
    if(N777) begin
      \nz.mem_44_sv2v_reg  <= data_i[4];
    end 
    if(N776) begin
      \nz.mem_43_sv2v_reg  <= data_i[3];
    end 
    if(N775) begin
      \nz.mem_42_sv2v_reg  <= data_i[2];
    end 
    if(N774) begin
      \nz.mem_41_sv2v_reg  <= data_i[1];
    end 
    if(N773) begin
      \nz.mem_40_sv2v_reg  <= data_i[0];
    end 
    if(N772) begin
      \nz.mem_39_sv2v_reg  <= data_i[7];
    end 
    if(N771) begin
      \nz.mem_38_sv2v_reg  <= data_i[6];
    end 
    if(N770) begin
      \nz.mem_37_sv2v_reg  <= data_i[5];
    end 
    if(N769) begin
      \nz.mem_36_sv2v_reg  <= data_i[4];
    end 
    if(N768) begin
      \nz.mem_35_sv2v_reg  <= data_i[3];
    end 
    if(N767) begin
      \nz.mem_34_sv2v_reg  <= data_i[2];
    end 
    if(N766) begin
      \nz.mem_33_sv2v_reg  <= data_i[1];
    end 
    if(N765) begin
      \nz.mem_32_sv2v_reg  <= data_i[0];
    end 
    if(N764) begin
      \nz.mem_31_sv2v_reg  <= data_i[7];
    end 
    if(N763) begin
      \nz.mem_30_sv2v_reg  <= data_i[6];
    end 
    if(N762) begin
      \nz.mem_29_sv2v_reg  <= data_i[5];
    end 
    if(N761) begin
      \nz.mem_28_sv2v_reg  <= data_i[4];
    end 
    if(N760) begin
      \nz.mem_27_sv2v_reg  <= data_i[3];
    end 
    if(N759) begin
      \nz.mem_26_sv2v_reg  <= data_i[2];
    end 
    if(N758) begin
      \nz.mem_25_sv2v_reg  <= data_i[1];
    end 
    if(N757) begin
      \nz.mem_24_sv2v_reg  <= data_i[0];
    end 
    if(N756) begin
      \nz.mem_23_sv2v_reg  <= data_i[7];
    end 
    if(N755) begin
      \nz.mem_22_sv2v_reg  <= data_i[6];
    end 
    if(N754) begin
      \nz.mem_21_sv2v_reg  <= data_i[5];
    end 
    if(N753) begin
      \nz.mem_20_sv2v_reg  <= data_i[4];
    end 
    if(N752) begin
      \nz.mem_19_sv2v_reg  <= data_i[3];
    end 
    if(N751) begin
      \nz.mem_18_sv2v_reg  <= data_i[2];
    end 
    if(N750) begin
      \nz.mem_17_sv2v_reg  <= data_i[1];
    end 
    if(N749) begin
      \nz.mem_16_sv2v_reg  <= data_i[0];
    end 
    if(N748) begin
      \nz.mem_15_sv2v_reg  <= data_i[7];
    end 
    if(N747) begin
      \nz.mem_14_sv2v_reg  <= data_i[6];
    end 
    if(N746) begin
      \nz.mem_13_sv2v_reg  <= data_i[5];
    end 
    if(N745) begin
      \nz.mem_12_sv2v_reg  <= data_i[4];
    end 
    if(N744) begin
      \nz.mem_11_sv2v_reg  <= data_i[3];
    end 
    if(N743) begin
      \nz.mem_10_sv2v_reg  <= data_i[2];
    end 
    if(N742) begin
      \nz.mem_9_sv2v_reg  <= data_i[1];
    end 
    if(N741) begin
      \nz.mem_8_sv2v_reg  <= data_i[0];
    end 
    if(N740) begin
      \nz.mem_7_sv2v_reg  <= data_i[7];
    end 
    if(N739) begin
      \nz.mem_6_sv2v_reg  <= data_i[6];
    end 
    if(N738) begin
      \nz.mem_5_sv2v_reg  <= data_i[5];
    end 
    if(N737) begin
      \nz.mem_4_sv2v_reg  <= data_i[4];
    end 
    if(N736) begin
      \nz.mem_3_sv2v_reg  <= data_i[3];
    end 
    if(N735) begin
      \nz.mem_2_sv2v_reg  <= data_i[2];
    end 
    if(N734) begin
      \nz.mem_1_sv2v_reg  <= data_i[1];
    end 
    if(N733) begin
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p8_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [7:0] data_i;
  input [5:0] addr_i;
  input [7:0] w_mask_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [7:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p8_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_scan_width_p2_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [1:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o[0] = i[0] | 1'b0;
  assign o[1] = i[1] | i[0];

endmodule



module bsg_priority_encode_one_hot_out_width_p2_lo_to_hi_p1
(
  i,
  o,
  v_o
);

  input [1:0] i;
  output [1:0] o;
  output v_o;
  wire [1:0] o;
  wire v_o,N0;

  bsg_scan_width_p2_or_p1_lo_to_hi_p1
  \nw1.scan 
  (
    .i(i),
    .o({ v_o, o[0:0] })
  );

  assign o[1] = v_o & N0;
  assign N0 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p2_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign addr_o[0] = i[1];
  assign v_o = addr_o[0] | i[0];

endmodule



module bsg_priority_encode_width_p2_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  wire [1:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p2_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo),
    .v_o(v_o)
  );


  bsg_encode_one_hot_width_p2_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o[0])
  );


endmodule



module bsg_dff_en_width_p3_harden_p0_strength_p0
(
  clk_i,
  data_i,
  en_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input en_i;
  wire [2:0] data_o;
  reg data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(en_i) begin
      data_o_2_sv2v_reg <= data_i[2];
      data_o_1_sv2v_reg <= data_i[1];
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule



module bsg_dff_en_bypass_width_p3
(
  clk_i,
  en_i,
  data_i,
  data_o
);

  input [2:0] data_i;
  output [2:0] data_o;
  input clk_i;
  input en_i;
  wire [2:0] data_o,data_r;
  wire N0,N1,N2,N3;

  bsg_dff_en_width_p3_harden_p0_strength_p0
  dff
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .en_i(en_i),
    .data_o(data_r)
  );

  assign data_o = (N0)? data_i : 
                  (N1)? data_r : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N2 = ~en_i;
  assign N3 = en_i;

endmodule



module bsg_mem_1rw_sync_mask_write_bit_synth_width_p3_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [2:0] data_i;
  input [5:0] addr_i;
  input [2:0] w_mask_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [2:0] data_o,\nz.data_out ;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,\nz.read_en ,N12,N13,N14,N15,N16,N17,N18,
  N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,
  N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,
  N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,
  N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,
  N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,
  N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,
  N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,\nz.llr.read_en_r ,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621;
  wire [5:0] \nz.addr_r ;
  wire [191:0] \nz.mem ;
  reg \nz.addr_r_5_sv2v_reg ,\nz.addr_r_4_sv2v_reg ,\nz.addr_r_3_sv2v_reg ,
  \nz.addr_r_2_sv2v_reg ,\nz.addr_r_1_sv2v_reg ,\nz.addr_r_0_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,
  \nz.mem_180_sv2v_reg ,\nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,
  \nz.mem_140_sv2v_reg ,\nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,
  \nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,
  \nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,
  \nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.addr_r [5] = \nz.addr_r_5_sv2v_reg ;
  assign \nz.addr_r [4] = \nz.addr_r_4_sv2v_reg ;
  assign \nz.addr_r [3] = \nz.addr_r_3_sv2v_reg ;
  assign \nz.addr_r [2] = \nz.addr_r_2_sv2v_reg ;
  assign \nz.addr_r [1] = \nz.addr_r_1_sv2v_reg ;
  assign \nz.addr_r [0] = \nz.addr_r_0_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign \nz.data_out [2] = (N78)? \nz.mem [2] : 
                            (N80)? \nz.mem [5] : 
                            (N82)? \nz.mem [8] : 
                            (N84)? \nz.mem [11] : 
                            (N86)? \nz.mem [14] : 
                            (N88)? \nz.mem [17] : 
                            (N90)? \nz.mem [20] : 
                            (N92)? \nz.mem [23] : 
                            (N94)? \nz.mem [26] : 
                            (N96)? \nz.mem [29] : 
                            (N98)? \nz.mem [32] : 
                            (N100)? \nz.mem [35] : 
                            (N102)? \nz.mem [38] : 
                            (N104)? \nz.mem [41] : 
                            (N106)? \nz.mem [44] : 
                            (N108)? \nz.mem [47] : 
                            (N110)? \nz.mem [50] : 
                            (N112)? \nz.mem [53] : 
                            (N114)? \nz.mem [56] : 
                            (N116)? \nz.mem [59] : 
                            (N118)? \nz.mem [62] : 
                            (N120)? \nz.mem [65] : 
                            (N122)? \nz.mem [68] : 
                            (N124)? \nz.mem [71] : 
                            (N126)? \nz.mem [74] : 
                            (N128)? \nz.mem [77] : 
                            (N130)? \nz.mem [80] : 
                            (N132)? \nz.mem [83] : 
                            (N134)? \nz.mem [86] : 
                            (N136)? \nz.mem [89] : 
                            (N138)? \nz.mem [92] : 
                            (N140)? \nz.mem [95] : 
                            (N79)? \nz.mem [98] : 
                            (N81)? \nz.mem [101] : 
                            (N83)? \nz.mem [104] : 
                            (N85)? \nz.mem [107] : 
                            (N87)? \nz.mem [110] : 
                            (N89)? \nz.mem [113] : 
                            (N91)? \nz.mem [116] : 
                            (N93)? \nz.mem [119] : 
                            (N95)? \nz.mem [122] : 
                            (N97)? \nz.mem [125] : 
                            (N99)? \nz.mem [128] : 
                            (N101)? \nz.mem [131] : 
                            (N103)? \nz.mem [134] : 
                            (N105)? \nz.mem [137] : 
                            (N107)? \nz.mem [140] : 
                            (N109)? \nz.mem [143] : 
                            (N111)? \nz.mem [146] : 
                            (N113)? \nz.mem [149] : 
                            (N115)? \nz.mem [152] : 
                            (N117)? \nz.mem [155] : 
                            (N119)? \nz.mem [158] : 
                            (N121)? \nz.mem [161] : 
                            (N123)? \nz.mem [164] : 
                            (N125)? \nz.mem [167] : 
                            (N127)? \nz.mem [170] : 
                            (N129)? \nz.mem [173] : 
                            (N131)? \nz.mem [176] : 
                            (N133)? \nz.mem [179] : 
                            (N135)? \nz.mem [182] : 
                            (N137)? \nz.mem [185] : 
                            (N139)? \nz.mem [188] : 
                            (N141)? \nz.mem [191] : 1'b0;
  assign \nz.data_out [1] = (N78)? \nz.mem [1] : 
                            (N80)? \nz.mem [4] : 
                            (N82)? \nz.mem [7] : 
                            (N84)? \nz.mem [10] : 
                            (N86)? \nz.mem [13] : 
                            (N88)? \nz.mem [16] : 
                            (N90)? \nz.mem [19] : 
                            (N92)? \nz.mem [22] : 
                            (N94)? \nz.mem [25] : 
                            (N96)? \nz.mem [28] : 
                            (N98)? \nz.mem [31] : 
                            (N100)? \nz.mem [34] : 
                            (N102)? \nz.mem [37] : 
                            (N104)? \nz.mem [40] : 
                            (N106)? \nz.mem [43] : 
                            (N108)? \nz.mem [46] : 
                            (N110)? \nz.mem [49] : 
                            (N112)? \nz.mem [52] : 
                            (N114)? \nz.mem [55] : 
                            (N116)? \nz.mem [58] : 
                            (N118)? \nz.mem [61] : 
                            (N120)? \nz.mem [64] : 
                            (N122)? \nz.mem [67] : 
                            (N124)? \nz.mem [70] : 
                            (N126)? \nz.mem [73] : 
                            (N128)? \nz.mem [76] : 
                            (N130)? \nz.mem [79] : 
                            (N132)? \nz.mem [82] : 
                            (N134)? \nz.mem [85] : 
                            (N136)? \nz.mem [88] : 
                            (N138)? \nz.mem [91] : 
                            (N140)? \nz.mem [94] : 
                            (N79)? \nz.mem [97] : 
                            (N81)? \nz.mem [100] : 
                            (N83)? \nz.mem [103] : 
                            (N85)? \nz.mem [106] : 
                            (N87)? \nz.mem [109] : 
                            (N89)? \nz.mem [112] : 
                            (N91)? \nz.mem [115] : 
                            (N93)? \nz.mem [118] : 
                            (N95)? \nz.mem [121] : 
                            (N97)? \nz.mem [124] : 
                            (N99)? \nz.mem [127] : 
                            (N101)? \nz.mem [130] : 
                            (N103)? \nz.mem [133] : 
                            (N105)? \nz.mem [136] : 
                            (N107)? \nz.mem [139] : 
                            (N109)? \nz.mem [142] : 
                            (N111)? \nz.mem [145] : 
                            (N113)? \nz.mem [148] : 
                            (N115)? \nz.mem [151] : 
                            (N117)? \nz.mem [154] : 
                            (N119)? \nz.mem [157] : 
                            (N121)? \nz.mem [160] : 
                            (N123)? \nz.mem [163] : 
                            (N125)? \nz.mem [166] : 
                            (N127)? \nz.mem [169] : 
                            (N129)? \nz.mem [172] : 
                            (N131)? \nz.mem [175] : 
                            (N133)? \nz.mem [178] : 
                            (N135)? \nz.mem [181] : 
                            (N137)? \nz.mem [184] : 
                            (N139)? \nz.mem [187] : 
                            (N141)? \nz.mem [190] : 1'b0;
  assign \nz.data_out [0] = (N78)? \nz.mem [0] : 
                            (N80)? \nz.mem [3] : 
                            (N82)? \nz.mem [6] : 
                            (N84)? \nz.mem [9] : 
                            (N86)? \nz.mem [12] : 
                            (N88)? \nz.mem [15] : 
                            (N90)? \nz.mem [18] : 
                            (N92)? \nz.mem [21] : 
                            (N94)? \nz.mem [24] : 
                            (N96)? \nz.mem [27] : 
                            (N98)? \nz.mem [30] : 
                            (N100)? \nz.mem [33] : 
                            (N102)? \nz.mem [36] : 
                            (N104)? \nz.mem [39] : 
                            (N106)? \nz.mem [42] : 
                            (N108)? \nz.mem [45] : 
                            (N110)? \nz.mem [48] : 
                            (N112)? \nz.mem [51] : 
                            (N114)? \nz.mem [54] : 
                            (N116)? \nz.mem [57] : 
                            (N118)? \nz.mem [60] : 
                            (N120)? \nz.mem [63] : 
                            (N122)? \nz.mem [66] : 
                            (N124)? \nz.mem [69] : 
                            (N126)? \nz.mem [72] : 
                            (N128)? \nz.mem [75] : 
                            (N130)? \nz.mem [78] : 
                            (N132)? \nz.mem [81] : 
                            (N134)? \nz.mem [84] : 
                            (N136)? \nz.mem [87] : 
                            (N138)? \nz.mem [90] : 
                            (N140)? \nz.mem [93] : 
                            (N79)? \nz.mem [96] : 
                            (N81)? \nz.mem [99] : 
                            (N83)? \nz.mem [102] : 
                            (N85)? \nz.mem [105] : 
                            (N87)? \nz.mem [108] : 
                            (N89)? \nz.mem [111] : 
                            (N91)? \nz.mem [114] : 
                            (N93)? \nz.mem [117] : 
                            (N95)? \nz.mem [120] : 
                            (N97)? \nz.mem [123] : 
                            (N99)? \nz.mem [126] : 
                            (N101)? \nz.mem [129] : 
                            (N103)? \nz.mem [132] : 
                            (N105)? \nz.mem [135] : 
                            (N107)? \nz.mem [138] : 
                            (N109)? \nz.mem [141] : 
                            (N111)? \nz.mem [144] : 
                            (N113)? \nz.mem [147] : 
                            (N115)? \nz.mem [150] : 
                            (N117)? \nz.mem [153] : 
                            (N119)? \nz.mem [156] : 
                            (N121)? \nz.mem [159] : 
                            (N123)? \nz.mem [162] : 
                            (N125)? \nz.mem [165] : 
                            (N127)? \nz.mem [168] : 
                            (N129)? \nz.mem [171] : 
                            (N131)? \nz.mem [174] : 
                            (N133)? \nz.mem [177] : 
                            (N135)? \nz.mem [180] : 
                            (N137)? \nz.mem [183] : 
                            (N139)? \nz.mem [186] : 
                            (N141)? \nz.mem [189] : 1'b0;

  bsg_dff_width_p1
  \nz.llr.read_en_dff 
  (
    .clk_i(clk_i),
    .data_i(\nz.read_en ),
    .data_o(\nz.llr.read_en_r )
  );


  bsg_dff_en_bypass_width_p3
  \nz.llr.dff_bypass 
  (
    .clk_i(clk_i),
    .en_i(\nz.llr.read_en_r ),
    .data_i(\nz.data_out ),
    .data_o(data_o)
  );

  assign N595 = ~addr_i[5];
  assign N596 = addr_i[3] & addr_i[4];
  assign N597 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N598 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N599 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N600 = addr_i[5] & N596;
  assign N601 = addr_i[5] & N597;
  assign N602 = addr_i[5] & N598;
  assign N603 = addr_i[5] & N599;
  assign N604 = N595 & N596;
  assign N605 = N595 & N597;
  assign N606 = N595 & N598;
  assign N607 = N595 & N599;
  assign N608 = ~addr_i[2];
  assign N609 = addr_i[0] & addr_i[1];
  assign N610 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N611 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N612 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N613 = addr_i[2] & N609;
  assign N614 = addr_i[2] & N610;
  assign N615 = addr_i[2] & N611;
  assign N616 = addr_i[2] & N612;
  assign N617 = N608 & N609;
  assign N618 = N608 & N610;
  assign N619 = N608 & N611;
  assign N620 = N608 & N612;
  assign N338 = N600 & N613;
  assign N337 = N600 & N614;
  assign N336 = N600 & N615;
  assign N335 = N600 & N616;
  assign N334 = N600 & N617;
  assign N333 = N600 & N618;
  assign N332 = N600 & N619;
  assign N331 = N600 & N620;
  assign N330 = N601 & N613;
  assign N329 = N601 & N614;
  assign N328 = N601 & N615;
  assign N327 = N601 & N616;
  assign N326 = N601 & N617;
  assign N325 = N601 & N618;
  assign N324 = N601 & N619;
  assign N323 = N601 & N620;
  assign N322 = N602 & N613;
  assign N321 = N602 & N614;
  assign N320 = N602 & N615;
  assign N319 = N602 & N616;
  assign N318 = N602 & N617;
  assign N317 = N602 & N618;
  assign N316 = N602 & N619;
  assign N315 = N602 & N620;
  assign N314 = N603 & N613;
  assign N313 = N603 & N614;
  assign N312 = N603 & N615;
  assign N311 = N603 & N616;
  assign N310 = N603 & N617;
  assign N309 = N603 & N618;
  assign N308 = N603 & N619;
  assign N307 = N603 & N620;
  assign N306 = N604 & N613;
  assign N305 = N604 & N614;
  assign N304 = N604 & N615;
  assign N303 = N604 & N616;
  assign N302 = N604 & N617;
  assign N301 = N604 & N618;
  assign N300 = N604 & N619;
  assign N299 = N604 & N620;
  assign N298 = N605 & N613;
  assign N297 = N605 & N614;
  assign N296 = N605 & N615;
  assign N295 = N605 & N616;
  assign N294 = N605 & N617;
  assign N293 = N605 & N618;
  assign N292 = N605 & N619;
  assign N291 = N605 & N620;
  assign N290 = N606 & N613;
  assign N289 = N606 & N614;
  assign N288 = N606 & N615;
  assign N287 = N606 & N616;
  assign N286 = N606 & N617;
  assign N285 = N606 & N618;
  assign N284 = N606 & N619;
  assign N283 = N606 & N620;
  assign N282 = N607 & N613;
  assign N281 = N607 & N614;
  assign N280 = N607 & N615;
  assign N279 = N607 & N616;
  assign N278 = N607 & N617;
  assign N277 = N607 & N618;
  assign N276 = N607 & N619;
  assign N275 = N607 & N620;
  assign { N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145 } = (N8)? { N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N144)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210 } = (N9)? { N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N209)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339 } = (N10)? { N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N274)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403 } = (N11)? { N402, N273, N208, N401, N272, N207, N400, N271, N206, N399, N270, N205, N398, N269, N204, N397, N268, N203, N396, N267, N202, N395, N266, N201, N394, N265, N200, N393, N264, N199, N392, N263, N198, N391, N262, N197, N390, N261, N196, N389, N260, N195, N388, N259, N194, N387, N258, N193, N386, N257, N192, N385, N256, N191, N384, N255, N190, N383, N254, N189, N382, N253, N188, N381, N252, N187, N380, N251, N186, N379, N250, N185, N378, N249, N184, N377, N248, N183, N376, N247, N182, N375, N246, N181, N374, N245, N180, N373, N244, N179, N372, N243, N178, N371, N242, N177, N370, N241, N176, N369, N240, N175, N368, N239, N174, N367, N238, N173, N366, N237, N172, N365, N236, N171, N364, N235, N170, N363, N234, N169, N362, N233, N168, N361, N232, N167, N360, N231, N166, N359, N230, N165, N358, N229, N164, N357, N228, N163, N356, N227, N162, N355, N226, N161, N354, N225, N160, N353, N224, N159, N352, N223, N158, N351, N222, N157, N350, N221, N156, N349, N220, N155, N348, N219, N154, N347, N218, N153, N346, N217, N152, N345, N216, N151, N344, N215, N150, N343, N214, N149, N342, N213, N148, N341, N212, N147, N340, N211, N146, N339, N210, N145 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N143)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = N142;
  assign \nz.read_en  = v_i & N621;
  assign N621 = ~w_i;
  assign N12 = ~\nz.addr_r [0];
  assign N13 = ~\nz.addr_r [1];
  assign N14 = N12 & N13;
  assign N15 = N12 & \nz.addr_r [1];
  assign N16 = \nz.addr_r [0] & N13;
  assign N17 = \nz.addr_r [0] & \nz.addr_r [1];
  assign N18 = ~\nz.addr_r [2];
  assign N19 = N14 & N18;
  assign N20 = N14 & \nz.addr_r [2];
  assign N21 = N16 & N18;
  assign N22 = N16 & \nz.addr_r [2];
  assign N23 = N15 & N18;
  assign N24 = N15 & \nz.addr_r [2];
  assign N25 = N17 & N18;
  assign N26 = N17 & \nz.addr_r [2];
  assign N27 = ~\nz.addr_r [3];
  assign N28 = N19 & N27;
  assign N29 = N19 & \nz.addr_r [3];
  assign N30 = N21 & N27;
  assign N31 = N21 & \nz.addr_r [3];
  assign N32 = N23 & N27;
  assign N33 = N23 & \nz.addr_r [3];
  assign N34 = N25 & N27;
  assign N35 = N25 & \nz.addr_r [3];
  assign N36 = N20 & N27;
  assign N37 = N20 & \nz.addr_r [3];
  assign N38 = N22 & N27;
  assign N39 = N22 & \nz.addr_r [3];
  assign N40 = N24 & N27;
  assign N41 = N24 & \nz.addr_r [3];
  assign N42 = N26 & N27;
  assign N43 = N26 & \nz.addr_r [3];
  assign N44 = ~\nz.addr_r [4];
  assign N45 = N28 & N44;
  assign N46 = N28 & \nz.addr_r [4];
  assign N47 = N30 & N44;
  assign N48 = N30 & \nz.addr_r [4];
  assign N49 = N32 & N44;
  assign N50 = N32 & \nz.addr_r [4];
  assign N51 = N34 & N44;
  assign N52 = N34 & \nz.addr_r [4];
  assign N53 = N36 & N44;
  assign N54 = N36 & \nz.addr_r [4];
  assign N55 = N38 & N44;
  assign N56 = N38 & \nz.addr_r [4];
  assign N57 = N40 & N44;
  assign N58 = N40 & \nz.addr_r [4];
  assign N59 = N42 & N44;
  assign N60 = N42 & \nz.addr_r [4];
  assign N61 = N29 & N44;
  assign N62 = N29 & \nz.addr_r [4];
  assign N63 = N31 & N44;
  assign N64 = N31 & \nz.addr_r [4];
  assign N65 = N33 & N44;
  assign N66 = N33 & \nz.addr_r [4];
  assign N67 = N35 & N44;
  assign N68 = N35 & \nz.addr_r [4];
  assign N69 = N37 & N44;
  assign N70 = N37 & \nz.addr_r [4];
  assign N71 = N39 & N44;
  assign N72 = N39 & \nz.addr_r [4];
  assign N73 = N41 & N44;
  assign N74 = N41 & \nz.addr_r [4];
  assign N75 = N43 & N44;
  assign N76 = N43 & \nz.addr_r [4];
  assign N77 = ~\nz.addr_r [5];
  assign N78 = N45 & N77;
  assign N79 = N45 & \nz.addr_r [5];
  assign N80 = N47 & N77;
  assign N81 = N47 & \nz.addr_r [5];
  assign N82 = N49 & N77;
  assign N83 = N49 & \nz.addr_r [5];
  assign N84 = N51 & N77;
  assign N85 = N51 & \nz.addr_r [5];
  assign N86 = N53 & N77;
  assign N87 = N53 & \nz.addr_r [5];
  assign N88 = N55 & N77;
  assign N89 = N55 & \nz.addr_r [5];
  assign N90 = N57 & N77;
  assign N91 = N57 & \nz.addr_r [5];
  assign N92 = N59 & N77;
  assign N93 = N59 & \nz.addr_r [5];
  assign N94 = N61 & N77;
  assign N95 = N61 & \nz.addr_r [5];
  assign N96 = N63 & N77;
  assign N97 = N63 & \nz.addr_r [5];
  assign N98 = N65 & N77;
  assign N99 = N65 & \nz.addr_r [5];
  assign N100 = N67 & N77;
  assign N101 = N67 & \nz.addr_r [5];
  assign N102 = N69 & N77;
  assign N103 = N69 & \nz.addr_r [5];
  assign N104 = N71 & N77;
  assign N105 = N71 & \nz.addr_r [5];
  assign N106 = N73 & N77;
  assign N107 = N73 & \nz.addr_r [5];
  assign N108 = N75 & N77;
  assign N109 = N75 & \nz.addr_r [5];
  assign N110 = N46 & N77;
  assign N111 = N46 & \nz.addr_r [5];
  assign N112 = N48 & N77;
  assign N113 = N48 & \nz.addr_r [5];
  assign N114 = N50 & N77;
  assign N115 = N50 & \nz.addr_r [5];
  assign N116 = N52 & N77;
  assign N117 = N52 & \nz.addr_r [5];
  assign N118 = N54 & N77;
  assign N119 = N54 & \nz.addr_r [5];
  assign N120 = N56 & N77;
  assign N121 = N56 & \nz.addr_r [5];
  assign N122 = N58 & N77;
  assign N123 = N58 & \nz.addr_r [5];
  assign N124 = N60 & N77;
  assign N125 = N60 & \nz.addr_r [5];
  assign N126 = N62 & N77;
  assign N127 = N62 & \nz.addr_r [5];
  assign N128 = N64 & N77;
  assign N129 = N64 & \nz.addr_r [5];
  assign N130 = N66 & N77;
  assign N131 = N66 & \nz.addr_r [5];
  assign N132 = N68 & N77;
  assign N133 = N68 & \nz.addr_r [5];
  assign N134 = N70 & N77;
  assign N135 = N70 & \nz.addr_r [5];
  assign N136 = N72 & N77;
  assign N137 = N72 & \nz.addr_r [5];
  assign N138 = N74 & N77;
  assign N139 = N74 & \nz.addr_r [5];
  assign N140 = N76 & N77;
  assign N141 = N76 & \nz.addr_r [5];
  assign N142 = v_i & w_i;
  assign N143 = ~N142;
  assign N144 = ~w_mask_i[0];
  assign N209 = ~w_mask_i[1];
  assign N274 = ~w_mask_i[2];

  always @(posedge clk_i) begin
    if(1'b1) begin
      \nz.addr_r_5_sv2v_reg  <= addr_i[5];
      \nz.addr_r_4_sv2v_reg  <= addr_i[4];
      \nz.addr_r_3_sv2v_reg  <= addr_i[3];
      \nz.addr_r_2_sv2v_reg  <= addr_i[2];
      \nz.addr_r_1_sv2v_reg  <= addr_i[1];
      \nz.addr_r_0_sv2v_reg  <= addr_i[0];
    end 
    if(N594) begin
      \nz.mem_191_sv2v_reg  <= data_i[2];
    end 
    if(N593) begin
      \nz.mem_190_sv2v_reg  <= data_i[1];
    end 
    if(N592) begin
      \nz.mem_189_sv2v_reg  <= data_i[0];
    end 
    if(N591) begin
      \nz.mem_188_sv2v_reg  <= data_i[2];
    end 
    if(N590) begin
      \nz.mem_187_sv2v_reg  <= data_i[1];
    end 
    if(N589) begin
      \nz.mem_186_sv2v_reg  <= data_i[0];
    end 
    if(N588) begin
      \nz.mem_185_sv2v_reg  <= data_i[2];
    end 
    if(N587) begin
      \nz.mem_184_sv2v_reg  <= data_i[1];
    end 
    if(N586) begin
      \nz.mem_183_sv2v_reg  <= data_i[0];
    end 
    if(N585) begin
      \nz.mem_182_sv2v_reg  <= data_i[2];
    end 
    if(N584) begin
      \nz.mem_181_sv2v_reg  <= data_i[1];
    end 
    if(N583) begin
      \nz.mem_180_sv2v_reg  <= data_i[0];
    end 
    if(N582) begin
      \nz.mem_179_sv2v_reg  <= data_i[2];
    end 
    if(N581) begin
      \nz.mem_178_sv2v_reg  <= data_i[1];
    end 
    if(N580) begin
      \nz.mem_177_sv2v_reg  <= data_i[0];
    end 
    if(N579) begin
      \nz.mem_176_sv2v_reg  <= data_i[2];
    end 
    if(N578) begin
      \nz.mem_175_sv2v_reg  <= data_i[1];
    end 
    if(N577) begin
      \nz.mem_174_sv2v_reg  <= data_i[0];
    end 
    if(N576) begin
      \nz.mem_173_sv2v_reg  <= data_i[2];
    end 
    if(N575) begin
      \nz.mem_172_sv2v_reg  <= data_i[1];
    end 
    if(N574) begin
      \nz.mem_171_sv2v_reg  <= data_i[0];
    end 
    if(N573) begin
      \nz.mem_170_sv2v_reg  <= data_i[2];
    end 
    if(N572) begin
      \nz.mem_169_sv2v_reg  <= data_i[1];
    end 
    if(N571) begin
      \nz.mem_168_sv2v_reg  <= data_i[0];
    end 
    if(N570) begin
      \nz.mem_167_sv2v_reg  <= data_i[2];
    end 
    if(N569) begin
      \nz.mem_166_sv2v_reg  <= data_i[1];
    end 
    if(N568) begin
      \nz.mem_165_sv2v_reg  <= data_i[0];
    end 
    if(N567) begin
      \nz.mem_164_sv2v_reg  <= data_i[2];
    end 
    if(N566) begin
      \nz.mem_163_sv2v_reg  <= data_i[1];
    end 
    if(N565) begin
      \nz.mem_162_sv2v_reg  <= data_i[0];
    end 
    if(N564) begin
      \nz.mem_161_sv2v_reg  <= data_i[2];
    end 
    if(N563) begin
      \nz.mem_160_sv2v_reg  <= data_i[1];
    end 
    if(N562) begin
      \nz.mem_159_sv2v_reg  <= data_i[0];
    end 
    if(N561) begin
      \nz.mem_158_sv2v_reg  <= data_i[2];
    end 
    if(N560) begin
      \nz.mem_157_sv2v_reg  <= data_i[1];
    end 
    if(N559) begin
      \nz.mem_156_sv2v_reg  <= data_i[0];
    end 
    if(N558) begin
      \nz.mem_155_sv2v_reg  <= data_i[2];
    end 
    if(N557) begin
      \nz.mem_154_sv2v_reg  <= data_i[1];
    end 
    if(N556) begin
      \nz.mem_153_sv2v_reg  <= data_i[0];
    end 
    if(N555) begin
      \nz.mem_152_sv2v_reg  <= data_i[2];
    end 
    if(N554) begin
      \nz.mem_151_sv2v_reg  <= data_i[1];
    end 
    if(N553) begin
      \nz.mem_150_sv2v_reg  <= data_i[0];
    end 
    if(N552) begin
      \nz.mem_149_sv2v_reg  <= data_i[2];
    end 
    if(N551) begin
      \nz.mem_148_sv2v_reg  <= data_i[1];
    end 
    if(N550) begin
      \nz.mem_147_sv2v_reg  <= data_i[0];
    end 
    if(N549) begin
      \nz.mem_146_sv2v_reg  <= data_i[2];
    end 
    if(N548) begin
      \nz.mem_145_sv2v_reg  <= data_i[1];
    end 
    if(N547) begin
      \nz.mem_144_sv2v_reg  <= data_i[0];
    end 
    if(N546) begin
      \nz.mem_143_sv2v_reg  <= data_i[2];
    end 
    if(N545) begin
      \nz.mem_142_sv2v_reg  <= data_i[1];
    end 
    if(N544) begin
      \nz.mem_141_sv2v_reg  <= data_i[0];
    end 
    if(N543) begin
      \nz.mem_140_sv2v_reg  <= data_i[2];
    end 
    if(N542) begin
      \nz.mem_139_sv2v_reg  <= data_i[1];
    end 
    if(N541) begin
      \nz.mem_138_sv2v_reg  <= data_i[0];
    end 
    if(N540) begin
      \nz.mem_137_sv2v_reg  <= data_i[2];
    end 
    if(N539) begin
      \nz.mem_136_sv2v_reg  <= data_i[1];
    end 
    if(N538) begin
      \nz.mem_135_sv2v_reg  <= data_i[0];
    end 
    if(N537) begin
      \nz.mem_134_sv2v_reg  <= data_i[2];
    end 
    if(N536) begin
      \nz.mem_133_sv2v_reg  <= data_i[1];
    end 
    if(N535) begin
      \nz.mem_132_sv2v_reg  <= data_i[0];
    end 
    if(N534) begin
      \nz.mem_131_sv2v_reg  <= data_i[2];
    end 
    if(N533) begin
      \nz.mem_130_sv2v_reg  <= data_i[1];
    end 
    if(N532) begin
      \nz.mem_129_sv2v_reg  <= data_i[0];
    end 
    if(N531) begin
      \nz.mem_128_sv2v_reg  <= data_i[2];
    end 
    if(N530) begin
      \nz.mem_127_sv2v_reg  <= data_i[1];
    end 
    if(N529) begin
      \nz.mem_126_sv2v_reg  <= data_i[0];
    end 
    if(N528) begin
      \nz.mem_125_sv2v_reg  <= data_i[2];
    end 
    if(N527) begin
      \nz.mem_124_sv2v_reg  <= data_i[1];
    end 
    if(N526) begin
      \nz.mem_123_sv2v_reg  <= data_i[0];
    end 
    if(N525) begin
      \nz.mem_122_sv2v_reg  <= data_i[2];
    end 
    if(N524) begin
      \nz.mem_121_sv2v_reg  <= data_i[1];
    end 
    if(N523) begin
      \nz.mem_120_sv2v_reg  <= data_i[0];
    end 
    if(N522) begin
      \nz.mem_119_sv2v_reg  <= data_i[2];
    end 
    if(N521) begin
      \nz.mem_118_sv2v_reg  <= data_i[1];
    end 
    if(N520) begin
      \nz.mem_117_sv2v_reg  <= data_i[0];
    end 
    if(N519) begin
      \nz.mem_116_sv2v_reg  <= data_i[2];
    end 
    if(N518) begin
      \nz.mem_115_sv2v_reg  <= data_i[1];
    end 
    if(N517) begin
      \nz.mem_114_sv2v_reg  <= data_i[0];
    end 
    if(N516) begin
      \nz.mem_113_sv2v_reg  <= data_i[2];
    end 
    if(N515) begin
      \nz.mem_112_sv2v_reg  <= data_i[1];
    end 
    if(N514) begin
      \nz.mem_111_sv2v_reg  <= data_i[0];
    end 
    if(N513) begin
      \nz.mem_110_sv2v_reg  <= data_i[2];
    end 
    if(N512) begin
      \nz.mem_109_sv2v_reg  <= data_i[1];
    end 
    if(N511) begin
      \nz.mem_108_sv2v_reg  <= data_i[0];
    end 
    if(N510) begin
      \nz.mem_107_sv2v_reg  <= data_i[2];
    end 
    if(N509) begin
      \nz.mem_106_sv2v_reg  <= data_i[1];
    end 
    if(N508) begin
      \nz.mem_105_sv2v_reg  <= data_i[0];
    end 
    if(N507) begin
      \nz.mem_104_sv2v_reg  <= data_i[2];
    end 
    if(N506) begin
      \nz.mem_103_sv2v_reg  <= data_i[1];
    end 
    if(N505) begin
      \nz.mem_102_sv2v_reg  <= data_i[0];
    end 
    if(N504) begin
      \nz.mem_101_sv2v_reg  <= data_i[2];
    end 
    if(N503) begin
      \nz.mem_100_sv2v_reg  <= data_i[1];
    end 
    if(N502) begin
      \nz.mem_99_sv2v_reg  <= data_i[0];
    end 
    if(N501) begin
      \nz.mem_98_sv2v_reg  <= data_i[2];
    end 
    if(N500) begin
      \nz.mem_97_sv2v_reg  <= data_i[1];
    end 
    if(N499) begin
      \nz.mem_96_sv2v_reg  <= data_i[0];
    end 
    if(N498) begin
      \nz.mem_95_sv2v_reg  <= data_i[2];
    end 
    if(N497) begin
      \nz.mem_94_sv2v_reg  <= data_i[1];
    end 
    if(N496) begin
      \nz.mem_93_sv2v_reg  <= data_i[0];
    end 
    if(N495) begin
      \nz.mem_92_sv2v_reg  <= data_i[2];
    end 
    if(N494) begin
      \nz.mem_91_sv2v_reg  <= data_i[1];
    end 
    if(N493) begin
      \nz.mem_90_sv2v_reg  <= data_i[0];
    end 
    if(N492) begin
      \nz.mem_89_sv2v_reg  <= data_i[2];
    end 
    if(N491) begin
      \nz.mem_88_sv2v_reg  <= data_i[1];
    end 
    if(N490) begin
      \nz.mem_87_sv2v_reg  <= data_i[0];
    end 
    if(N489) begin
      \nz.mem_86_sv2v_reg  <= data_i[2];
    end 
    if(N488) begin
      \nz.mem_85_sv2v_reg  <= data_i[1];
    end 
    if(N487) begin
      \nz.mem_84_sv2v_reg  <= data_i[0];
    end 
    if(N486) begin
      \nz.mem_83_sv2v_reg  <= data_i[2];
    end 
    if(N485) begin
      \nz.mem_82_sv2v_reg  <= data_i[1];
    end 
    if(N484) begin
      \nz.mem_81_sv2v_reg  <= data_i[0];
    end 
    if(N483) begin
      \nz.mem_80_sv2v_reg  <= data_i[2];
    end 
    if(N482) begin
      \nz.mem_79_sv2v_reg  <= data_i[1];
    end 
    if(N481) begin
      \nz.mem_78_sv2v_reg  <= data_i[0];
    end 
    if(N480) begin
      \nz.mem_77_sv2v_reg  <= data_i[2];
    end 
    if(N479) begin
      \nz.mem_76_sv2v_reg  <= data_i[1];
    end 
    if(N478) begin
      \nz.mem_75_sv2v_reg  <= data_i[0];
    end 
    if(N477) begin
      \nz.mem_74_sv2v_reg  <= data_i[2];
    end 
    if(N476) begin
      \nz.mem_73_sv2v_reg  <= data_i[1];
    end 
    if(N475) begin
      \nz.mem_72_sv2v_reg  <= data_i[0];
    end 
    if(N474) begin
      \nz.mem_71_sv2v_reg  <= data_i[2];
    end 
    if(N473) begin
      \nz.mem_70_sv2v_reg  <= data_i[1];
    end 
    if(N472) begin
      \nz.mem_69_sv2v_reg  <= data_i[0];
    end 
    if(N471) begin
      \nz.mem_68_sv2v_reg  <= data_i[2];
    end 
    if(N470) begin
      \nz.mem_67_sv2v_reg  <= data_i[1];
    end 
    if(N469) begin
      \nz.mem_66_sv2v_reg  <= data_i[0];
    end 
    if(N468) begin
      \nz.mem_65_sv2v_reg  <= data_i[2];
    end 
    if(N467) begin
      \nz.mem_64_sv2v_reg  <= data_i[1];
    end 
    if(N466) begin
      \nz.mem_63_sv2v_reg  <= data_i[0];
    end 
    if(N465) begin
      \nz.mem_62_sv2v_reg  <= data_i[2];
    end 
    if(N464) begin
      \nz.mem_61_sv2v_reg  <= data_i[1];
    end 
    if(N463) begin
      \nz.mem_60_sv2v_reg  <= data_i[0];
    end 
    if(N462) begin
      \nz.mem_59_sv2v_reg  <= data_i[2];
    end 
    if(N461) begin
      \nz.mem_58_sv2v_reg  <= data_i[1];
    end 
    if(N460) begin
      \nz.mem_57_sv2v_reg  <= data_i[0];
    end 
    if(N459) begin
      \nz.mem_56_sv2v_reg  <= data_i[2];
    end 
    if(N458) begin
      \nz.mem_55_sv2v_reg  <= data_i[1];
    end 
    if(N457) begin
      \nz.mem_54_sv2v_reg  <= data_i[0];
    end 
    if(N456) begin
      \nz.mem_53_sv2v_reg  <= data_i[2];
    end 
    if(N455) begin
      \nz.mem_52_sv2v_reg  <= data_i[1];
    end 
    if(N454) begin
      \nz.mem_51_sv2v_reg  <= data_i[0];
    end 
    if(N453) begin
      \nz.mem_50_sv2v_reg  <= data_i[2];
    end 
    if(N452) begin
      \nz.mem_49_sv2v_reg  <= data_i[1];
    end 
    if(N451) begin
      \nz.mem_48_sv2v_reg  <= data_i[0];
    end 
    if(N450) begin
      \nz.mem_47_sv2v_reg  <= data_i[2];
    end 
    if(N449) begin
      \nz.mem_46_sv2v_reg  <= data_i[1];
    end 
    if(N448) begin
      \nz.mem_45_sv2v_reg  <= data_i[0];
    end 
    if(N447) begin
      \nz.mem_44_sv2v_reg  <= data_i[2];
    end 
    if(N446) begin
      \nz.mem_43_sv2v_reg  <= data_i[1];
    end 
    if(N445) begin
      \nz.mem_42_sv2v_reg  <= data_i[0];
    end 
    if(N444) begin
      \nz.mem_41_sv2v_reg  <= data_i[2];
    end 
    if(N443) begin
      \nz.mem_40_sv2v_reg  <= data_i[1];
    end 
    if(N442) begin
      \nz.mem_39_sv2v_reg  <= data_i[0];
    end 
    if(N441) begin
      \nz.mem_38_sv2v_reg  <= data_i[2];
    end 
    if(N440) begin
      \nz.mem_37_sv2v_reg  <= data_i[1];
    end 
    if(N439) begin
      \nz.mem_36_sv2v_reg  <= data_i[0];
    end 
    if(N438) begin
      \nz.mem_35_sv2v_reg  <= data_i[2];
    end 
    if(N437) begin
      \nz.mem_34_sv2v_reg  <= data_i[1];
    end 
    if(N436) begin
      \nz.mem_33_sv2v_reg  <= data_i[0];
    end 
    if(N435) begin
      \nz.mem_32_sv2v_reg  <= data_i[2];
    end 
    if(N434) begin
      \nz.mem_31_sv2v_reg  <= data_i[1];
    end 
    if(N433) begin
      \nz.mem_30_sv2v_reg  <= data_i[0];
    end 
    if(N432) begin
      \nz.mem_29_sv2v_reg  <= data_i[2];
    end 
    if(N431) begin
      \nz.mem_28_sv2v_reg  <= data_i[1];
    end 
    if(N430) begin
      \nz.mem_27_sv2v_reg  <= data_i[0];
    end 
    if(N429) begin
      \nz.mem_26_sv2v_reg  <= data_i[2];
    end 
    if(N428) begin
      \nz.mem_25_sv2v_reg  <= data_i[1];
    end 
    if(N427) begin
      \nz.mem_24_sv2v_reg  <= data_i[0];
    end 
    if(N426) begin
      \nz.mem_23_sv2v_reg  <= data_i[2];
    end 
    if(N425) begin
      \nz.mem_22_sv2v_reg  <= data_i[1];
    end 
    if(N424) begin
      \nz.mem_21_sv2v_reg  <= data_i[0];
    end 
    if(N423) begin
      \nz.mem_20_sv2v_reg  <= data_i[2];
    end 
    if(N422) begin
      \nz.mem_19_sv2v_reg  <= data_i[1];
    end 
    if(N421) begin
      \nz.mem_18_sv2v_reg  <= data_i[0];
    end 
    if(N420) begin
      \nz.mem_17_sv2v_reg  <= data_i[2];
    end 
    if(N419) begin
      \nz.mem_16_sv2v_reg  <= data_i[1];
    end 
    if(N418) begin
      \nz.mem_15_sv2v_reg  <= data_i[0];
    end 
    if(N417) begin
      \nz.mem_14_sv2v_reg  <= data_i[2];
    end 
    if(N416) begin
      \nz.mem_13_sv2v_reg  <= data_i[1];
    end 
    if(N415) begin
      \nz.mem_12_sv2v_reg  <= data_i[0];
    end 
    if(N414) begin
      \nz.mem_11_sv2v_reg  <= data_i[2];
    end 
    if(N413) begin
      \nz.mem_10_sv2v_reg  <= data_i[1];
    end 
    if(N412) begin
      \nz.mem_9_sv2v_reg  <= data_i[0];
    end 
    if(N411) begin
      \nz.mem_8_sv2v_reg  <= data_i[2];
    end 
    if(N410) begin
      \nz.mem_7_sv2v_reg  <= data_i[1];
    end 
    if(N409) begin
      \nz.mem_6_sv2v_reg  <= data_i[0];
    end 
    if(N408) begin
      \nz.mem_5_sv2v_reg  <= data_i[2];
    end 
    if(N407) begin
      \nz.mem_4_sv2v_reg  <= data_i[1];
    end 
    if(N406) begin
      \nz.mem_3_sv2v_reg  <= data_i[0];
    end 
    if(N405) begin
      \nz.mem_2_sv2v_reg  <= data_i[2];
    end 
    if(N404) begin
      \nz.mem_1_sv2v_reg  <= data_i[1];
    end 
    if(N403) begin
      \nz.mem_0_sv2v_reg  <= data_i[0];
    end 
  end


endmodule



module bsg_mem_1rw_sync_mask_write_bit_width_p3_els_p64_latch_last_read_p1
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [2:0] data_i;
  input [5:0] addr_i;
  input [2:0] w_mask_i;
  output [2:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [2:0] data_o;

  bsg_mem_1rw_sync_mask_write_bit_synth_width_p3_els_p64_latch_last_read_p1
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .addr_i(addr_i),
    .v_i(v_i),
    .w_mask_i(w_mask_i),
    .w_i(w_i),
    .data_o(data_o)
  );


endmodule



module bsg_lru_pseudo_tree_decode_ways_p2
(
  way_id_i,
  data_o,
  mask_o
);

  input [0:0] way_id_i;
  output [0:0] data_o;
  output [0:0] mask_o;
  wire [0:0] data_o,mask_o;
  wire N0;
  assign mask_o[0] = 1'b1;
  assign data_o[0] = 1'b1 & N0;
  assign N0 = ~way_id_i[0];

endmodule



module bsg_lru_pseudo_tree_encode_ways_p2
(
  lru_i,
  way_id_o
);

  input [0:0] lru_i;
  output [0:0] way_id_o;
  wire [0:0] way_id_o;
  assign way_id_o[0] = lru_i[0];

endmodule



module bsg_decode_num_out_p2
(
  i,
  o
);

  input [0:0] i;
  output [1:0] o;
  wire [1:0] o;
  assign o = { 1'b0, 1'b1 } << i[0];

endmodule



module bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2_word_tracking_p1
(
  clk_i,
  reset_i,
  miss_v_i,
  track_miss_i,
  decode_v_i,
  addr_v_i,
  mask_v_i,
  tag_v_i,
  valid_v_i,
  lock_v_i,
  tag_hit_v_i,
  tag_hit_way_id_i,
  tag_hit_found_i,
  sbuf_empty_i,
  tbuf_empty_i,
  dma_cmd_o,
  dma_way_o,
  dma_addr_o,
  dma_done_i,
  track_data_we_o,
  stat_info_i,
  stat_mem_v_o,
  stat_mem_w_o,
  stat_mem_addr_o,
  stat_mem_data_o,
  stat_mem_w_mask_o,
  tag_mem_v_o,
  tag_mem_w_o,
  tag_mem_addr_o,
  tag_mem_data_o,
  tag_mem_w_mask_o,
  track_mem_v_o,
  track_mem_w_o,
  track_mem_addr_o,
  track_mem_w_mask_o,
  track_mem_data_o,
  done_o,
  recover_o,
  chosen_way_o,
  select_snoop_data_r_o,
  ack_i
);

  input [20:0] decode_v_i;
  input [27:0] addr_v_i;
  input [3:0] mask_v_i;
  input [35:0] tag_v_i;
  input [1:0] valid_v_i;
  input [1:0] lock_v_i;
  input [1:0] tag_hit_v_i;
  input [0:0] tag_hit_way_id_i;
  output [3:0] dma_cmd_o;
  output [0:0] dma_way_o;
  output [27:0] dma_addr_o;
  input [2:0] stat_info_i;
  output [5:0] stat_mem_addr_o;
  output [2:0] stat_mem_data_o;
  output [2:0] stat_mem_w_mask_o;
  output [5:0] tag_mem_addr_o;
  output [39:0] tag_mem_data_o;
  output [39:0] tag_mem_w_mask_o;
  output [5:0] track_mem_addr_o;
  output [7:0] track_mem_w_mask_o;
  output [7:0] track_mem_data_o;
  output [0:0] chosen_way_o;
  input clk_i;
  input reset_i;
  input miss_v_i;
  input track_miss_i;
  input tag_hit_found_i;
  input sbuf_empty_i;
  input tbuf_empty_i;
  input dma_done_i;
  input ack_i;
  output track_data_we_o;
  output stat_mem_v_o;
  output stat_mem_w_o;
  output tag_mem_v_o;
  output tag_mem_w_o;
  output track_mem_v_o;
  output track_mem_w_o;
  output done_o;
  output recover_o;
  output select_snoop_data_r_o;
  wire [3:0] dma_cmd_o,miss_state_r,miss_state_n;
  wire [0:0] dma_way_o,chosen_way_o,invalid_way_id,flush_way_r,chosen_way_lru_data,
  chosen_way_lru_mask,modify_mask_lo,modify_data_lo,modified_lru_bits,lru_way_id,
  chosen_way_n;
  wire [27:0] dma_addr_o;
  wire [5:0] stat_mem_addr_o,tag_mem_addr_o,track_mem_addr_o;
  wire [2:0] stat_mem_data_o,stat_mem_w_mask_o;
  wire [39:0] tag_mem_data_o,tag_mem_w_mask_o;
  wire [7:0] track_mem_w_mask_o,track_mem_data_o;
  wire track_data_we_o,stat_mem_v_o,stat_mem_w_o,tag_mem_v_o,tag_mem_w_o,track_mem_v_o,
  track_mem_w_o,done_o,recover_o,select_snoop_data_r_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,
  N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,
  track_mem_data_o_1__3_,_0_net__1_,_0_net__0_,invalid_exist,goto_flush_op,goto_lock_op,
  N27,N28,full_word_op,st_tag_miss_op,N29,N30,select_snoop_data_n,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,
  N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,
  N224,N225,N226,N227;
  wire [1:0] chosen_way_decode,addr_way_v_decode,flush_way_decode;
  reg track_data_we_o_sv2v_reg,miss_state_r_3_sv2v_reg,miss_state_r_2_sv2v_reg,
  miss_state_r_1_sv2v_reg,miss_state_r_0_sv2v_reg,chosen_way_o_0_sv2v_reg,
  flush_way_r_0_sv2v_reg,select_snoop_data_r_o_sv2v_reg;
  assign track_data_we_o = track_data_we_o_sv2v_reg;
  assign miss_state_r[3] = miss_state_r_3_sv2v_reg;
  assign miss_state_r[2] = miss_state_r_2_sv2v_reg;
  assign miss_state_r[1] = miss_state_r_1_sv2v_reg;
  assign miss_state_r[0] = miss_state_r_0_sv2v_reg;
  assign chosen_way_o[0] = chosen_way_o_0_sv2v_reg;
  assign flush_way_r[0] = flush_way_r_0_sv2v_reg;
  assign select_snoop_data_r_o = select_snoop_data_r_o_sv2v_reg;
  assign dma_addr_o[0] = 1'b0;
  assign dma_addr_o[1] = 1'b0;
  assign stat_mem_addr_o[5] = addr_v_i[9];
  assign track_mem_addr_o[5] = stat_mem_addr_o[5];
  assign tag_mem_addr_o[5] = stat_mem_addr_o[5];
  assign stat_mem_addr_o[4] = addr_v_i[8];
  assign track_mem_addr_o[4] = stat_mem_addr_o[4];
  assign tag_mem_addr_o[4] = stat_mem_addr_o[4];
  assign stat_mem_addr_o[3] = addr_v_i[7];
  assign track_mem_addr_o[3] = stat_mem_addr_o[3];
  assign tag_mem_addr_o[3] = stat_mem_addr_o[3];
  assign stat_mem_addr_o[2] = addr_v_i[6];
  assign track_mem_addr_o[2] = stat_mem_addr_o[2];
  assign tag_mem_addr_o[2] = stat_mem_addr_o[2];
  assign stat_mem_addr_o[1] = addr_v_i[5];
  assign track_mem_addr_o[1] = stat_mem_addr_o[1];
  assign tag_mem_addr_o[1] = stat_mem_addr_o[1];
  assign stat_mem_addr_o[0] = addr_v_i[4];
  assign track_mem_addr_o[0] = stat_mem_addr_o[0];
  assign tag_mem_addr_o[0] = stat_mem_addr_o[0];
  assign dma_cmd_o[2] = track_mem_data_o_1__3_;
  assign track_mem_data_o[0] = track_mem_data_o_1__3_;
  assign track_mem_data_o[1] = track_mem_data_o_1__3_;
  assign track_mem_data_o[2] = track_mem_data_o_1__3_;
  assign track_mem_data_o[3] = track_mem_data_o_1__3_;
  assign track_mem_data_o[4] = track_mem_data_o_1__3_;
  assign track_mem_data_o[5] = track_mem_data_o_1__3_;
  assign track_mem_data_o[6] = track_mem_data_o_1__3_;
  assign track_mem_data_o[7] = track_mem_data_o_1__3_;

  bsg_priority_encode_width_p2_lo_to_hi_p1
  invalid_way_pe
  (
    .i({ _0_net__1_, _0_net__0_ }),
    .addr_o(invalid_way_id[0]),
    .v_o(invalid_exist)
  );


  bsg_lru_pseudo_tree_decode_ways_p2
  chosen_way_lru_decode
  (
    .way_id_i(chosen_way_o[0]),
    .data_o(chosen_way_lru_data[0]),
    .mask_o(chosen_way_lru_mask[0])
  );


  bsg_lru_pseudo_tree_backup
  backup_lru
  (
    .disabled_ways_i(lock_v_i),
    .modify_mask_o(modify_mask_lo[0]),
    .modify_data_o(modify_data_lo[0])
  );


  bsg_mux_bitwise
  lru_bit_mux
  (
    .data0_i(stat_info_i[0]),
    .data1_i(modify_data_lo[0]),
    .sel_i(modify_mask_lo[0]),
    .data_o(modified_lru_bits[0])
  );


  bsg_lru_pseudo_tree_encode_ways_p2
  lru_encode
  (
    .lru_i(modified_lru_bits[0]),
    .way_id_o(lru_way_id[0])
  );


  bsg_decode_num_out_p2
  chosen_way_demux
  (
    .i(chosen_way_n[0]),
    .o(chosen_way_decode)
  );


  bsg_decode_num_out_p2
  addr_way_v_demux
  (
    .i(addr_v_i[10]),
    .o(addr_way_v_decode)
  );

  assign N35 = N31 & N32;
  assign N36 = N33 & N34;
  assign N37 = N35 & N36;
  assign N38 = miss_state_r[3] | N32;
  assign N39 = miss_state_r[1] | miss_state_r[0];
  assign N40 = N38 | N39;
  assign N42 = miss_state_r[3] | miss_state_r[2];
  assign N43 = miss_state_r[1] | N34;
  assign N44 = N42 | N43;
  assign N46 = miss_state_r[3] | miss_state_r[2];
  assign N47 = N33 | miss_state_r[0];
  assign N48 = N46 | N47;
  assign N50 = miss_state_r[3] | miss_state_r[2];
  assign N51 = N33 | N34;
  assign N52 = N50 | N51;
  assign N54 = miss_state_r[3] | N32;
  assign N55 = miss_state_r[1] | N34;
  assign N56 = N54 | N55;
  assign N58 = miss_state_r[3] | N32;
  assign N59 = N33 | miss_state_r[0];
  assign N60 = N58 | N59;
  assign N62 = miss_state_r[3] | N32;
  assign N63 = N33 | N34;
  assign N64 = N62 | N63;
  assign N66 = N31 | miss_state_r[2];
  assign N67 = miss_state_r[1] | miss_state_r[0];
  assign N68 = N66 | N67;
  assign N70 = N31 | miss_state_r[2];
  assign N71 = miss_state_r[1] | N34;
  assign N72 = N70 | N71;
  assign N74 = N31 | miss_state_r[2];
  assign N75 = N33 | miss_state_r[0];
  assign N76 = N74 | N75;
  assign N78 = miss_state_r[3] & miss_state_r[1];
  assign N79 = N78 & miss_state_r[0];
  assign N80 = miss_state_r[3] & miss_state_r[2];
  assign N97 = (N96)? stat_info_i[1] : 
               (N0)? stat_info_i[2] : 1'b0;
  assign N0 = N95;
  assign N98 = (N96)? valid_v_i[0] : 
               (N0)? valid_v_i[1] : 1'b0;
  assign N109 = (N108)? stat_info_i[1] : 
                (N1)? stat_info_i[2] : 1'b0;
  assign N1 = N103;
  assign N110 = (N108)? valid_v_i[0] : 
                (N1)? valid_v_i[1] : 1'b0;
  assign N114 = (N113)? tag_v_i[17] : 
                (N2)? tag_v_i[35] : 1'b0;
  assign N2 = dma_way_o[0];
  assign N115 = (N113)? tag_v_i[16] : 
                (N2)? tag_v_i[34] : 1'b0;
  assign N116 = (N113)? tag_v_i[15] : 
                (N2)? tag_v_i[33] : 1'b0;
  assign N117 = (N113)? tag_v_i[14] : 
                (N2)? tag_v_i[32] : 1'b0;
  assign N118 = (N113)? tag_v_i[13] : 
                (N2)? tag_v_i[31] : 1'b0;
  assign N119 = (N113)? tag_v_i[12] : 
                (N2)? tag_v_i[30] : 1'b0;
  assign N120 = (N113)? tag_v_i[11] : 
                (N2)? tag_v_i[29] : 1'b0;
  assign N121 = (N113)? tag_v_i[10] : 
                (N2)? tag_v_i[28] : 1'b0;
  assign N122 = (N113)? tag_v_i[9] : 
                (N2)? tag_v_i[27] : 1'b0;
  assign N123 = (N113)? tag_v_i[8] : 
                (N2)? tag_v_i[26] : 1'b0;
  assign N124 = (N113)? tag_v_i[7] : 
                (N2)? tag_v_i[25] : 1'b0;
  assign N125 = (N113)? tag_v_i[6] : 
                (N2)? tag_v_i[24] : 1'b0;
  assign N126 = (N113)? tag_v_i[5] : 
                (N2)? tag_v_i[23] : 1'b0;
  assign N127 = (N113)? tag_v_i[4] : 
                (N2)? tag_v_i[22] : 1'b0;
  assign N128 = (N113)? tag_v_i[3] : 
                (N2)? tag_v_i[21] : 1'b0;
  assign N129 = (N113)? tag_v_i[2] : 
                (N2)? tag_v_i[20] : 1'b0;
  assign N130 = (N113)? tag_v_i[1] : 
                (N2)? tag_v_i[19] : 1'b0;
  assign N131 = (N113)? tag_v_i[0] : 
                (N2)? tag_v_i[18] : 1'b0;
  assign N133 = (N113)? tag_v_i[17] : 
                (N2)? tag_v_i[35] : 1'b0;
  assign N134 = (N113)? tag_v_i[16] : 
                (N2)? tag_v_i[34] : 1'b0;
  assign N135 = (N113)? tag_v_i[15] : 
                (N2)? tag_v_i[33] : 1'b0;
  assign N136 = (N113)? tag_v_i[14] : 
                (N2)? tag_v_i[32] : 1'b0;
  assign N137 = (N113)? tag_v_i[13] : 
                (N2)? tag_v_i[31] : 1'b0;
  assign N138 = (N113)? tag_v_i[12] : 
                (N2)? tag_v_i[30] : 1'b0;
  assign N139 = (N113)? tag_v_i[11] : 
                (N2)? tag_v_i[29] : 1'b0;
  assign N140 = (N113)? tag_v_i[10] : 
                (N2)? tag_v_i[28] : 1'b0;
  assign N141 = (N113)? tag_v_i[9] : 
                (N2)? tag_v_i[27] : 1'b0;
  assign N142 = (N113)? tag_v_i[8] : 
                (N2)? tag_v_i[26] : 1'b0;
  assign N143 = (N113)? tag_v_i[7] : 
                (N2)? tag_v_i[25] : 1'b0;
  assign N144 = (N113)? tag_v_i[6] : 
                (N2)? tag_v_i[24] : 1'b0;
  assign N145 = (N113)? tag_v_i[5] : 
                (N2)? tag_v_i[23] : 1'b0;
  assign N146 = (N113)? tag_v_i[4] : 
                (N2)? tag_v_i[22] : 1'b0;
  assign N147 = (N113)? tag_v_i[3] : 
                (N2)? tag_v_i[21] : 1'b0;
  assign N148 = (N113)? tag_v_i[2] : 
                (N2)? tag_v_i[20] : 1'b0;
  assign N149 = (N113)? tag_v_i[1] : 
                (N2)? tag_v_i[19] : 1'b0;
  assign N150 = (N113)? tag_v_i[0] : 
                (N2)? tag_v_i[18] : 1'b0;
  assign N166 = (N165)? stat_info_i[1] : 
                (N3)? stat_info_i[2] : 1'b0;
  assign N3 = N164;
  assign N167 = (N165)? valid_v_i[0] : 
                (N3)? valid_v_i[1] : 1'b0;
  assign full_word_op = (N4)? N28 : 
                        (N27)? decode_v_i[20] : 1'b0;
  assign N4 = decode_v_i[17];
  assign dma_way_o[0] = (N5)? flush_way_r[0] : 
                        (N6)? chosen_way_o[0] : 1'b0;
  assign N5 = goto_flush_op;
  assign N6 = N29;
  assign flush_way_decode = (N7)? addr_way_v_decode : 
                            (N30)? tag_hit_v_i : 1'b0;
  assign N7 = decode_v_i[13];
  assign { N89, N88, N87 } = (N5)? { 1'b0, 1'b0, 1'b1 } : 
                             (N174)? { 1'b0, 1'b1, 1'b0 } : 
                             (N177)? { 1'b1, 1'b1, 1'b1 } : 
                             (N86)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign { N92, N91, N90 } = (N8)? { N89, N88, N87 } : 
                             (N83)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = N82;
  assign N95 = (N9)? tag_hit_way_id_i[0] : 
               (N179)? invalid_way_id[0] : 
               (N94)? lru_way_id[0] : 1'b0;
  assign N9 = track_miss_i;
  assign N100 = ~N99;
  assign { N102, N101 } = (N10)? { N100, N99 } : 
                          (N11)? { 1'b1, 1'b0 } : 1'b0;
  assign N10 = dma_done_i;
  assign N11 = N132;
  assign N103 = (N7)? addr_v_i[10] : 
                (N30)? tag_hit_way_id_i[0] : 1'b0;
  assign N112 = ~N111;
  assign N155 = ~N154;
  assign { N159, N158, N157, N156 } = (N10)? { N154, N155, N155, N154 } : 
                                      (N11)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 1'b0;
  assign { N162, N161 } = (N9)? { 1'b0, 1'b0 } : 
                          (N12)? chosen_way_decode : 1'b0;
  assign N12 = N217;
  assign N164 = (N13)? invalid_way_id[0] : 
                (N14)? lru_way_id[0] : 1'b0;
  assign N13 = invalid_exist;
  assign N14 = N163;
  assign N169 = ~N168;
  assign stat_mem_v_o = (N15)? N82 : 
                        (N16)? 1'b0 : 
                        (N17)? 1'b1 : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b0 : 
                        (N20)? N151 : 
                        (N21)? dma_done_i : 
                        (N22)? 1'b0 : 
                        (N23)? 1'b1 : 
                        (N24)? 1'b0 : 
                        (N25)? 1'b0 : 
                        (N26)? 1'b0 : 1'b0;
  assign N15 = N37;
  assign N16 = dma_cmd_o[0];
  assign N17 = N45;
  assign N18 = N49;
  assign N19 = dma_cmd_o[1];
  assign N20 = dma_cmd_o[3];
  assign N21 = track_mem_data_o_1__3_;
  assign N22 = N65;
  assign N23 = N69;
  assign N24 = N73;
  assign N25 = N77;
  assign N26 = N81;
  assign track_mem_v_o = (N15)? N82 : 
                         (N16)? 1'b0 : 
                         (N17)? 1'b0 : 
                         (N18)? 1'b0 : 
                         (N19)? 1'b0 : 
                         (N20)? N153 : 
                         (N21)? dma_done_i : 
                         (N22)? 1'b0 : 
                         (N23)? 1'b1 : 
                         (N24)? 1'b0 : 
                         (N25)? 1'b0 : 
                         (N26)? 1'b0 : 1'b0;
  assign miss_state_n = (N15)? { 1'b0, N92, N91, N90 } : 
                        (N16)? { 1'b0, N102, dma_done_i, N101 } : 
                        (N17)? { N112, 1'b0, N111, 1'b1 } : 
                        (N18)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                        (N19)? { 1'b0, dma_done_i, N132, 1'b1 } : 
                        (N20)? { N159, N158, N157, N156 } : 
                        (N21)? { dma_done_i, N132, N132, dma_done_i } : 
                        (N22)? { N169, 1'b0, N168, N168 } : 
                        (N23)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                        (N24)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                        (N25)? { N170, 1'b0, N170, 1'b0 } : 
                        (N26)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign chosen_way_n[0] = (N15)? chosen_way_o[0] : 
                           (N16)? N95 : 
                           (N17)? chosen_way_o[0] : 
                           (N18)? chosen_way_o[0] : 
                           (N19)? chosen_way_o[0] : 
                           (N20)? chosen_way_o[0] : 
                           (N21)? chosen_way_o[0] : 
                           (N22)? N164 : 
                           (N23)? chosen_way_o[0] : 
                           (N24)? chosen_way_o[0] : 
                           (N25)? chosen_way_o[0] : 
                           (N26)? chosen_way_o[0] : 1'b0;
  assign dma_addr_o[3:2] = (N21)? addr_v_i[3:2] : 
                           (N172)? { 1'b0, 1'b0 } : 1'b0;
  assign dma_addr_o[27:4] = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N16)? { addr_v_i[27:10], stat_mem_addr_o } : 
                            (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, stat_mem_addr_o } : 
                            (N20)? { N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, stat_mem_addr_o } : 
                            (N21)? { addr_v_i[27:10], stat_mem_addr_o } : 
                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N23)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_o = (N15)? 1'b0 : 
                        (N16)? 1'b0 : 
                        (N17)? 1'b1 : 
                        (N18)? 1'b0 : 
                        (N19)? 1'b0 : 
                        (N20)? 1'b1 : 
                        (N21)? 1'b1 : 
                        (N22)? 1'b0 : 
                        (N23)? 1'b1 : 
                        (N24)? 1'b0 : 
                        (N25)? 1'b0 : 
                        (N26)? 1'b0 : 1'b0;
  assign stat_mem_data_o = (N15)? { 1'b0, 1'b0, 1'b0 } : 
                           (N16)? { 1'b0, 1'b0, 1'b0 } : 
                           (N17)? { 1'b0, 1'b0, 1'b0 } : 
                           (N18)? { 1'b0, 1'b0, 1'b0 } : 
                           (N19)? { 1'b0, 1'b0, 1'b0 } : 
                           (N20)? { 1'b1, 1'b1, chosen_way_lru_data[0:0] } : 
                           (N21)? { N160, N160, chosen_way_lru_data[0:0] } : 
                           (N22)? { 1'b0, 1'b0, 1'b0 } : 
                           (N23)? { 1'b1, 1'b1, chosen_way_lru_data[0:0] } : 
                           (N24)? { 1'b0, 1'b0, 1'b0 } : 
                           (N25)? { 1'b0, 1'b0, 1'b0 } : 
                           (N26)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign stat_mem_w_mask_o = (N15)? { 1'b0, 1'b0, 1'b0 } : 
                             (N16)? { 1'b0, 1'b0, 1'b0 } : 
                             (N17)? { flush_way_decode, 1'b0 } : 
                             (N18)? { 1'b0, 1'b0, 1'b0 } : 
                             (N19)? { 1'b0, 1'b0, 1'b0 } : 
                             (N20)? { chosen_way_decode, chosen_way_lru_mask[0:0] } : 
                             (N21)? { N162, N161, chosen_way_lru_mask[0:0] } : 
                             (N22)? { 1'b0, 1'b0, 1'b0 } : 
                             (N23)? { chosen_way_decode, chosen_way_lru_mask[0:0] } : 
                             (N24)? { 1'b0, 1'b0, 1'b0 } : 
                             (N25)? { 1'b0, 1'b0, 1'b0 } : 
                             (N26)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_v_o = (N15)? 1'b0 : 
                       (N16)? 1'b0 : 
                       (N17)? 1'b1 : 
                       (N18)? 1'b1 : 
                       (N19)? 1'b0 : 
                       (N20)? N152 : 
                       (N21)? dma_done_i : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b1 : 
                       (N24)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N26)? 1'b0 : 1'b0;
  assign tag_mem_w_o = (N15)? 1'b0 : 
                       (N16)? 1'b0 : 
                       (N17)? 1'b1 : 
                       (N18)? 1'b1 : 
                       (N19)? 1'b0 : 
                       (N20)? 1'b1 : 
                       (N21)? 1'b1 : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b1 : 
                       (N24)? 1'b0 : 
                       (N25)? 1'b0 : 
                       (N26)? 1'b0 : 1'b0;
  assign tag_mem_w_mask_o = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N17)? { N106, N107, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N104, N105, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N18)? { 1'b0, tag_hit_v_i[1:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, tag_hit_v_i[0:0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N20)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N21)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N23)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                            (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                            (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign tag_mem_data_o = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N18)? { 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, decode_v_i[7:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N20)? { 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10] } : 
                          (N21)? { 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10] } : 
                          (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N23)? { 1'b1, decode_v_i[7:7], addr_v_i[27:10], 1'b1, decode_v_i[7:7], addr_v_i[27:10] } : 
                          (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                          (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign track_mem_w_o = (N15)? 1'b0 : 
                         (N16)? 1'b0 : 
                         (N17)? 1'b0 : 
                         (N18)? 1'b0 : 
                         (N19)? 1'b0 : 
                         (N20)? 1'b1 : 
                         (N21)? 1'b1 : 
                         (N22)? 1'b0 : 
                         (N23)? 1'b1 : 
                         (N24)? 1'b0 : 
                         (N25)? 1'b0 : 
                         (N26)? 1'b0 : 1'b0;
  assign track_mem_w_mask_o = (N15)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N20)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N21)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N23)? { chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode[1:1], chosen_way_decode, chosen_way_decode[0:0], chosen_way_decode[0:0], chosen_way_decode[0:0] } : 
                              (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N25)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                              (N26)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign select_snoop_data_n = (N21)? 1'b1 : 
                               (N25)? 1'b0 : 1'b0;
  assign recover_o = (N15)? 1'b0 : 
                     (N16)? 1'b0 : 
                     (N17)? 1'b0 : 
                     (N18)? 1'b0 : 
                     (N19)? 1'b0 : 
                     (N20)? 1'b0 : 
                     (N21)? 1'b0 : 
                     (N22)? 1'b0 : 
                     (N23)? 1'b0 : 
                     (N24)? 1'b1 : 
                     (N25)? 1'b0 : 
                     (N26)? 1'b0 : 1'b0;
  assign done_o = (N15)? 1'b0 : 
                  (N16)? 1'b0 : 
                  (N17)? 1'b0 : 
                  (N18)? 1'b0 : 
                  (N19)? 1'b0 : 
                  (N20)? 1'b0 : 
                  (N21)? 1'b0 : 
                  (N22)? 1'b0 : 
                  (N23)? 1'b0 : 
                  (N24)? 1'b0 : 
                  (N25)? 1'b1 : 
                  (N26)? 1'b0 : 1'b0;
  assign _0_net__1_ = N205 & N206;
  assign N205 = ~valid_v_i[1];
  assign N206 = ~lock_v_i[1];
  assign _0_net__0_ = N207 & N208;
  assign N207 = ~valid_v_i[0];
  assign N208 = ~lock_v_i[0];
  assign goto_flush_op = N210 | decode_v_i[9];
  assign N210 = N209 | decode_v_i[10];
  assign N209 = decode_v_i[13] | decode_v_i[8];
  assign goto_lock_op = decode_v_i[6] | N211;
  assign N211 = decode_v_i[7] & tag_hit_found_i;
  assign N27 = ~decode_v_i[17];
  assign N28 = N213 & mask_v_i[0];
  assign N213 = N212 & mask_v_i[1];
  assign N212 = mask_v_i[3] & mask_v_i[2];
  assign st_tag_miss_op = N214 & N215;
  assign N214 = decode_v_i[15] & full_word_op;
  assign N215 = ~tag_hit_found_i;
  assign N29 = ~goto_flush_op;
  assign N30 = ~decode_v_i[13];
  assign N31 = ~miss_state_r[3];
  assign N32 = ~miss_state_r[2];
  assign N33 = ~miss_state_r[1];
  assign N34 = ~miss_state_r[0];
  assign N41 = ~N40;
  assign N45 = ~N44;
  assign N49 = ~N48;
  assign N53 = ~N52;
  assign N57 = ~N56;
  assign N61 = ~N60;
  assign N65 = ~N64;
  assign N69 = ~N68;
  assign N73 = ~N72;
  assign N77 = ~N76;
  assign N81 = N79 | N80;
  assign dma_cmd_o[0] = N41;
  assign dma_cmd_o[1] = N53;
  assign dma_cmd_o[3] = N57;
  assign track_mem_data_o_1__3_ = N61;
  assign N82 = N216 & tbuf_empty_i;
  assign N216 = miss_v_i & sbuf_empty_i;
  assign N83 = ~N82;
  assign N84 = goto_lock_op | goto_flush_op;
  assign N85 = st_tag_miss_op | N84;
  assign N86 = ~N85;
  assign N93 = invalid_exist | track_miss_i;
  assign N94 = ~N93;
  assign N96 = ~N95;
  assign N99 = N218 & N98;
  assign N218 = N217 & N97;
  assign N217 = ~track_miss_i;
  assign N104 = N219 & flush_way_decode[0];
  assign N219 = decode_v_i[8] | decode_v_i[9];
  assign N105 = N220 & flush_way_decode[0];
  assign N220 = decode_v_i[8] | decode_v_i[9];
  assign N106 = N221 & flush_way_decode[1];
  assign N221 = decode_v_i[8] | decode_v_i[9];
  assign N107 = N222 & flush_way_decode[1];
  assign N222 = decode_v_i[8] | decode_v_i[9];
  assign N108 = ~N103;
  assign N111 = N224 & N110;
  assign N224 = N223 & N109;
  assign N223 = ~decode_v_i[8];
  assign N113 = ~dma_way_o[0];
  assign N132 = ~dma_done_i;
  assign N151 = dma_done_i & st_tag_miss_op;
  assign N152 = dma_done_i & st_tag_miss_op;
  assign N153 = dma_done_i & st_tag_miss_op;
  assign N154 = N226 | st_tag_miss_op;
  assign N226 = N225 | decode_v_i[10];
  assign N225 = decode_v_i[13] | decode_v_i[9];
  assign N160 = decode_v_i[15] | decode_v_i[4];
  assign N163 = ~invalid_exist;
  assign N165 = ~N164;
  assign N168 = N166 & N167;
  assign N170 = ~ack_i;
  assign N171 = ~track_mem_data_o_1__3_;
  assign N172 = N171;
  assign N173 = ~goto_flush_op;
  assign N174 = goto_lock_op & N173;
  assign N175 = ~goto_lock_op;
  assign N176 = N173 & N175;
  assign N177 = st_tag_miss_op & N176;
  assign N178 = ~track_miss_i;
  assign N179 = invalid_exist & N178;
  assign N180 = track_mem_v_o & N227;
  assign N227 = ~track_mem_w_o;
  assign N181 = N37 | dma_cmd_o[0];
  assign N182 = N181 | N49;
  assign N183 = N182 | dma_cmd_o[1];
  assign N184 = N183 | dma_cmd_o[3];
  assign N185 = N184 | track_mem_data_o_1__3_;
  assign N186 = N185 | N65;
  assign N187 = N186 | N69;
  assign N188 = N187 | N73;
  assign N189 = N188 | N77;
  assign N190 = N189 | N81;
  assign N191 = ~N190;
  assign N192 = N181 | N45;
  assign N193 = N192 | N49;
  assign N194 = N193 | dma_cmd_o[1];
  assign N195 = N194 | dma_cmd_o[3];
  assign N196 = N132 & track_mem_data_o_1__3_;
  assign N197 = N195 | N196;
  assign N198 = N197 | N65;
  assign N199 = N198 | N69;
  assign N200 = N199 | N73;
  assign N201 = N170 & N77;
  assign N202 = N200 | N201;
  assign N203 = N202 | N81;
  assign N204 = ~N203;

  always @(posedge clk_i) begin
    if(reset_i) begin
      track_data_we_o_sv2v_reg <= 1'b0;
      miss_state_r_3_sv2v_reg <= 1'b0;
      miss_state_r_2_sv2v_reg <= 1'b0;
      miss_state_r_1_sv2v_reg <= 1'b0;
      miss_state_r_0_sv2v_reg <= 1'b0;
      chosen_way_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      track_data_we_o_sv2v_reg <= N180;
      miss_state_r_3_sv2v_reg <= miss_state_n[3];
      miss_state_r_2_sv2v_reg <= miss_state_n[2];
      miss_state_r_1_sv2v_reg <= miss_state_n[1];
      miss_state_r_0_sv2v_reg <= miss_state_n[0];
      chosen_way_o_0_sv2v_reg <= chosen_way_n[0];
    end 
    if(reset_i) begin
      flush_way_r_0_sv2v_reg <= 1'b0;
    end else if(N191) begin
      flush_way_r_0_sv2v_reg <= N103;
    end 
    if(reset_i) begin
      select_snoop_data_r_o_sv2v_reg <= 1'b0;
    end else if(N204) begin
      select_snoop_data_r_o_sv2v_reg <= select_snoop_data_n;
    end 
  end


endmodule



module bsg_counter_clear_up_4_0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [2:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire [2:0] count_o;
  wire N0,N1,N4,N5,N6,N8,N9,N10,N11,N12,N13,N14,N15,N2,N3,N7,N30,N16;
  reg count_o_2_sv2v_reg,count_o_1_sv2v_reg,count_o_0_sv2v_reg;
  assign count_o[2] = count_o_2_sv2v_reg;
  assign count_o[1] = count_o_1_sv2v_reg;
  assign count_o[0] = count_o_0_sv2v_reg;
  assign N16 = reset_i | clear_i;
  assign { N8, N6, N5 } = count_o + 1'b1;
  assign N9 = (N0)? 1'b1 : 
              (N7)? 1'b1 : 
              (N3)? 1'b0 : 1'b0;
  assign N0 = clear_i;
  assign N11 = (N1)? 1'b1 : 
               (N30)? 1'b0 : 1'b0;
  assign N1 = up_i;
  assign N10 = (N0)? up_i : 
               (N7)? N5 : 1'b0;
  assign N4 = N15;
  assign N12 = ~reset_i;
  assign N13 = ~clear_i;
  assign N14 = N12 & N13;
  assign N15 = up_i & N14;
  assign N2 = up_i | clear_i;
  assign N3 = ~N2;
  assign N7 = up_i & N13;
  assign N30 = ~up_i;

  always @(posedge clk_i) begin
    if(N16) begin
      count_o_2_sv2v_reg <= 1'b0;
      count_o_1_sv2v_reg <= 1'b0;
    end else if(N11) begin
      count_o_2_sv2v_reg <= N8;
      count_o_1_sv2v_reg <= N6;
    end 
    if(reset_i) begin
      count_o_0_sv2v_reg <= 1'b0;
    end else if(N9) begin
      count_o_0_sv2v_reg <= N10;
    end 
  end


endmodule



module bsg_circular_ptr_slots_p4_max_add_p1
(
  clk,
  reset_i,
  add_i,
  o,
  n_o
);

  input [0:0] add_i;
  output [1:0] o;
  output [1:0] n_o;
  input clk;
  input reset_i;
  wire [1:0] o,n_o,\genblk1.genblk1.ptr_r_p1 ;
  wire N0,N1,N2;
  reg o_1_sv2v_reg,o_0_sv2v_reg;
  assign o[1] = o_1_sv2v_reg;
  assign o[0] = o_0_sv2v_reg;
  assign \genblk1.genblk1.ptr_r_p1  = o + 1'b1;
  assign n_o = (N0)? \genblk1.genblk1.ptr_r_p1  : 
               (N1)? o : 1'b0;
  assign N0 = add_i[0];
  assign N1 = N2;
  assign N2 = ~add_i[0];

  always @(posedge clk) begin
    if(reset_i) begin
      o_1_sv2v_reg <= 1'b0;
      o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      o_1_sv2v_reg <= n_o[1];
      o_0_sv2v_reg <= n_o[0];
    end 
  end


endmodule



module bsg_fifo_tracker_els_p4
(
  clk_i,
  reset_i,
  enq_i,
  deq_i,
  wptr_r_o,
  rptr_r_o,
  rptr_n_o,
  full_o,
  empty_o
);

  output [1:0] wptr_r_o;
  output [1:0] rptr_r_o;
  output [1:0] rptr_n_o;
  input clk_i;
  input reset_i;
  input enq_i;
  input deq_i;
  output full_o;
  output empty_o;
  wire [1:0] wptr_r_o,rptr_r_o,rptr_n_o;
  wire full_o,empty_o,enq_r,deq_r,N0,equal_ptrs,sv2v_dc_1,sv2v_dc_2;
  reg deq_r_sv2v_reg,enq_r_sv2v_reg;
  assign deq_r = deq_r_sv2v_reg;
  assign enq_r = enq_r_sv2v_reg;

  bsg_circular_ptr_slots_p4_max_add_p1
  rptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(deq_i),
    .o(rptr_r_o),
    .n_o(rptr_n_o)
  );


  bsg_circular_ptr_slots_p4_max_add_p1
  wptr
  (
    .clk(clk_i),
    .reset_i(reset_i),
    .add_i(enq_i),
    .o(wptr_r_o),
    .n_o({ sv2v_dc_1, sv2v_dc_2 })
  );

  assign equal_ptrs = rptr_r_o == wptr_r_o;
  assign N0 = enq_i | deq_i;
  assign empty_o = equal_ptrs & deq_r;
  assign full_o = equal_ptrs & enq_r;

  always @(posedge clk_i) begin
    if(reset_i) begin
      deq_r_sv2v_reg <= 1'b1;
      enq_r_sv2v_reg <= 1'b0;
    end else if(N0) begin
      deq_r_sv2v_reg <= deq_i;
      enq_r_sv2v_reg <= enq_i;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;
  wire [127:0] \nz.mem ;
  reg \nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,\nz.mem_125_sv2v_reg ,
  \nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,\nz.mem_121_sv2v_reg ,
  \nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,\nz.mem_118_sv2v_reg ,
  \nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,\nz.mem_114_sv2v_reg ,
  \nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,\nz.mem_110_sv2v_reg ,
  \nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,\nz.mem_107_sv2v_reg ,
  \nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,\nz.mem_103_sv2v_reg ,
  \nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,\nz.mem_99_sv2v_reg ,
  \nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,\nz.mem_96_sv2v_reg ,
  \nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,\nz.mem_92_sv2v_reg ,
  \nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,\nz.mem_88_sv2v_reg ,
  \nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,\nz.mem_84_sv2v_reg ,
  \nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,\nz.mem_80_sv2v_reg ,
  \nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,\nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,
  \nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,\nz.mem_73_sv2v_reg ,
  \nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,\nz.mem_69_sv2v_reg ,
  \nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,\nz.mem_65_sv2v_reg ,
  \nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,
  \nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,
  \nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,
  \nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,
  \nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,
  \nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,
  \nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,
  \nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,
  \nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,
  \nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,
  \nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N8)? \nz.mem [31] : 
                        (N10)? \nz.mem [63] : 
                        (N9)? \nz.mem [95] : 
                        (N11)? \nz.mem [127] : 1'b0;
  assign r_data_o[30] = (N8)? \nz.mem [30] : 
                        (N10)? \nz.mem [62] : 
                        (N9)? \nz.mem [94] : 
                        (N11)? \nz.mem [126] : 1'b0;
  assign r_data_o[29] = (N8)? \nz.mem [29] : 
                        (N10)? \nz.mem [61] : 
                        (N9)? \nz.mem [93] : 
                        (N11)? \nz.mem [125] : 1'b0;
  assign r_data_o[28] = (N8)? \nz.mem [28] : 
                        (N10)? \nz.mem [60] : 
                        (N9)? \nz.mem [92] : 
                        (N11)? \nz.mem [124] : 1'b0;
  assign r_data_o[27] = (N8)? \nz.mem [27] : 
                        (N10)? \nz.mem [59] : 
                        (N9)? \nz.mem [91] : 
                        (N11)? \nz.mem [123] : 1'b0;
  assign r_data_o[26] = (N8)? \nz.mem [26] : 
                        (N10)? \nz.mem [58] : 
                        (N9)? \nz.mem [90] : 
                        (N11)? \nz.mem [122] : 1'b0;
  assign r_data_o[25] = (N8)? \nz.mem [25] : 
                        (N10)? \nz.mem [57] : 
                        (N9)? \nz.mem [89] : 
                        (N11)? \nz.mem [121] : 1'b0;
  assign r_data_o[24] = (N8)? \nz.mem [24] : 
                        (N10)? \nz.mem [56] : 
                        (N9)? \nz.mem [88] : 
                        (N11)? \nz.mem [120] : 1'b0;
  assign r_data_o[23] = (N8)? \nz.mem [23] : 
                        (N10)? \nz.mem [55] : 
                        (N9)? \nz.mem [87] : 
                        (N11)? \nz.mem [119] : 1'b0;
  assign r_data_o[22] = (N8)? \nz.mem [22] : 
                        (N10)? \nz.mem [54] : 
                        (N9)? \nz.mem [86] : 
                        (N11)? \nz.mem [118] : 1'b0;
  assign r_data_o[21] = (N8)? \nz.mem [21] : 
                        (N10)? \nz.mem [53] : 
                        (N9)? \nz.mem [85] : 
                        (N11)? \nz.mem [117] : 1'b0;
  assign r_data_o[20] = (N8)? \nz.mem [20] : 
                        (N10)? \nz.mem [52] : 
                        (N9)? \nz.mem [84] : 
                        (N11)? \nz.mem [116] : 1'b0;
  assign r_data_o[19] = (N8)? \nz.mem [19] : 
                        (N10)? \nz.mem [51] : 
                        (N9)? \nz.mem [83] : 
                        (N11)? \nz.mem [115] : 1'b0;
  assign r_data_o[18] = (N8)? \nz.mem [18] : 
                        (N10)? \nz.mem [50] : 
                        (N9)? \nz.mem [82] : 
                        (N11)? \nz.mem [114] : 1'b0;
  assign r_data_o[17] = (N8)? \nz.mem [17] : 
                        (N10)? \nz.mem [49] : 
                        (N9)? \nz.mem [81] : 
                        (N11)? \nz.mem [113] : 1'b0;
  assign r_data_o[16] = (N8)? \nz.mem [16] : 
                        (N10)? \nz.mem [48] : 
                        (N9)? \nz.mem [80] : 
                        (N11)? \nz.mem [112] : 1'b0;
  assign r_data_o[15] = (N8)? \nz.mem [15] : 
                        (N10)? \nz.mem [47] : 
                        (N9)? \nz.mem [79] : 
                        (N11)? \nz.mem [111] : 1'b0;
  assign r_data_o[14] = (N8)? \nz.mem [14] : 
                        (N10)? \nz.mem [46] : 
                        (N9)? \nz.mem [78] : 
                        (N11)? \nz.mem [110] : 1'b0;
  assign r_data_o[13] = (N8)? \nz.mem [13] : 
                        (N10)? \nz.mem [45] : 
                        (N9)? \nz.mem [77] : 
                        (N11)? \nz.mem [109] : 1'b0;
  assign r_data_o[12] = (N8)? \nz.mem [12] : 
                        (N10)? \nz.mem [44] : 
                        (N9)? \nz.mem [76] : 
                        (N11)? \nz.mem [108] : 1'b0;
  assign r_data_o[11] = (N8)? \nz.mem [11] : 
                        (N10)? \nz.mem [43] : 
                        (N9)? \nz.mem [75] : 
                        (N11)? \nz.mem [107] : 1'b0;
  assign r_data_o[10] = (N8)? \nz.mem [10] : 
                        (N10)? \nz.mem [42] : 
                        (N9)? \nz.mem [74] : 
                        (N11)? \nz.mem [106] : 1'b0;
  assign r_data_o[9] = (N8)? \nz.mem [9] : 
                       (N10)? \nz.mem [41] : 
                       (N9)? \nz.mem [73] : 
                       (N11)? \nz.mem [105] : 1'b0;
  assign r_data_o[8] = (N8)? \nz.mem [8] : 
                       (N10)? \nz.mem [40] : 
                       (N9)? \nz.mem [72] : 
                       (N11)? \nz.mem [104] : 1'b0;
  assign r_data_o[7] = (N8)? \nz.mem [7] : 
                       (N10)? \nz.mem [39] : 
                       (N9)? \nz.mem [71] : 
                       (N11)? \nz.mem [103] : 1'b0;
  assign r_data_o[6] = (N8)? \nz.mem [6] : 
                       (N10)? \nz.mem [38] : 
                       (N9)? \nz.mem [70] : 
                       (N11)? \nz.mem [102] : 1'b0;
  assign r_data_o[5] = (N8)? \nz.mem [5] : 
                       (N10)? \nz.mem [37] : 
                       (N9)? \nz.mem [69] : 
                       (N11)? \nz.mem [101] : 1'b0;
  assign r_data_o[4] = (N8)? \nz.mem [4] : 
                       (N10)? \nz.mem [36] : 
                       (N9)? \nz.mem [68] : 
                       (N11)? \nz.mem [100] : 1'b0;
  assign r_data_o[3] = (N8)? \nz.mem [3] : 
                       (N10)? \nz.mem [35] : 
                       (N9)? \nz.mem [67] : 
                       (N11)? \nz.mem [99] : 1'b0;
  assign r_data_o[2] = (N8)? \nz.mem [2] : 
                       (N10)? \nz.mem [34] : 
                       (N9)? \nz.mem [66] : 
                       (N11)? \nz.mem [98] : 1'b0;
  assign r_data_o[1] = (N8)? \nz.mem [1] : 
                       (N10)? \nz.mem [33] : 
                       (N9)? \nz.mem [65] : 
                       (N11)? \nz.mem [97] : 1'b0;
  assign r_data_o[0] = (N8)? \nz.mem [0] : 
                       (N10)? \nz.mem [32] : 
                       (N9)? \nz.mem [64] : 
                       (N11)? \nz.mem [96] : 1'b0;
  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N20, N19, N18, N17 } = (N4)? { N16, N15, N14, N13 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N20) begin
      \nz.mem_127_sv2v_reg  <= w_data_i[31];
      \nz.mem_126_sv2v_reg  <= w_data_i[30];
      \nz.mem_125_sv2v_reg  <= w_data_i[29];
      \nz.mem_124_sv2v_reg  <= w_data_i[28];
      \nz.mem_123_sv2v_reg  <= w_data_i[27];
      \nz.mem_122_sv2v_reg  <= w_data_i[26];
      \nz.mem_121_sv2v_reg  <= w_data_i[25];
      \nz.mem_120_sv2v_reg  <= w_data_i[24];
      \nz.mem_119_sv2v_reg  <= w_data_i[23];
      \nz.mem_118_sv2v_reg  <= w_data_i[22];
      \nz.mem_117_sv2v_reg  <= w_data_i[21];
      \nz.mem_116_sv2v_reg  <= w_data_i[20];
      \nz.mem_115_sv2v_reg  <= w_data_i[19];
      \nz.mem_114_sv2v_reg  <= w_data_i[18];
      \nz.mem_113_sv2v_reg  <= w_data_i[17];
      \nz.mem_112_sv2v_reg  <= w_data_i[16];
      \nz.mem_111_sv2v_reg  <= w_data_i[15];
      \nz.mem_110_sv2v_reg  <= w_data_i[14];
      \nz.mem_109_sv2v_reg  <= w_data_i[13];
      \nz.mem_108_sv2v_reg  <= w_data_i[12];
      \nz.mem_107_sv2v_reg  <= w_data_i[11];
      \nz.mem_106_sv2v_reg  <= w_data_i[10];
      \nz.mem_105_sv2v_reg  <= w_data_i[9];
      \nz.mem_104_sv2v_reg  <= w_data_i[8];
      \nz.mem_103_sv2v_reg  <= w_data_i[7];
      \nz.mem_102_sv2v_reg  <= w_data_i[6];
      \nz.mem_101_sv2v_reg  <= w_data_i[5];
      \nz.mem_100_sv2v_reg  <= w_data_i[4];
      \nz.mem_99_sv2v_reg  <= w_data_i[3];
      \nz.mem_98_sv2v_reg  <= w_data_i[2];
      \nz.mem_97_sv2v_reg  <= w_data_i[1];
      \nz.mem_96_sv2v_reg  <= w_data_i[0];
    end 
    if(N19) begin
      \nz.mem_95_sv2v_reg  <= w_data_i[31];
      \nz.mem_94_sv2v_reg  <= w_data_i[30];
      \nz.mem_93_sv2v_reg  <= w_data_i[29];
      \nz.mem_92_sv2v_reg  <= w_data_i[28];
      \nz.mem_91_sv2v_reg  <= w_data_i[27];
      \nz.mem_90_sv2v_reg  <= w_data_i[26];
      \nz.mem_89_sv2v_reg  <= w_data_i[25];
      \nz.mem_88_sv2v_reg  <= w_data_i[24];
      \nz.mem_87_sv2v_reg  <= w_data_i[23];
      \nz.mem_86_sv2v_reg  <= w_data_i[22];
      \nz.mem_85_sv2v_reg  <= w_data_i[21];
      \nz.mem_84_sv2v_reg  <= w_data_i[20];
      \nz.mem_83_sv2v_reg  <= w_data_i[19];
      \nz.mem_82_sv2v_reg  <= w_data_i[18];
      \nz.mem_81_sv2v_reg  <= w_data_i[17];
      \nz.mem_80_sv2v_reg  <= w_data_i[16];
      \nz.mem_79_sv2v_reg  <= w_data_i[15];
      \nz.mem_78_sv2v_reg  <= w_data_i[14];
      \nz.mem_77_sv2v_reg  <= w_data_i[13];
      \nz.mem_76_sv2v_reg  <= w_data_i[12];
      \nz.mem_75_sv2v_reg  <= w_data_i[11];
      \nz.mem_74_sv2v_reg  <= w_data_i[10];
      \nz.mem_73_sv2v_reg  <= w_data_i[9];
      \nz.mem_72_sv2v_reg  <= w_data_i[8];
      \nz.mem_71_sv2v_reg  <= w_data_i[7];
      \nz.mem_70_sv2v_reg  <= w_data_i[6];
      \nz.mem_69_sv2v_reg  <= w_data_i[5];
      \nz.mem_68_sv2v_reg  <= w_data_i[4];
      \nz.mem_67_sv2v_reg  <= w_data_i[3];
      \nz.mem_66_sv2v_reg  <= w_data_i[2];
      \nz.mem_65_sv2v_reg  <= w_data_i[1];
      \nz.mem_64_sv2v_reg  <= w_data_i[0];
    end 
    if(N18) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N17) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [31:0] w_data_i;
  input [1:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p4_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enque,full,empty,sv2v_dc_1,sv2v_dc_2;
  wire [1:0] wptr_r,rptr_r;

  bsg_fifo_tracker_els_p4
  ft
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .enq_i(enque),
    .deq_i(yumi_i),
    .wptr_r_o(wptr_r),
    .rptr_r_o(rptr_r),
    .rptr_n_o({ sv2v_dc_1, sv2v_dc_2 }),
    .full_o(full),
    .empty_o(empty)
  );


  bsg_mem_1r1w_width_p32_els_p4_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enque),
    .w_addr_i(wptr_r),
    .w_data_i(data_i),
    .r_v_i(v_o),
    .r_addr_i(rptr_r),
    .r_data_o(data_o)
  );

  assign enque = v_i & ready_o;
  assign ready_o = ~full;
  assign v_o = ~empty;

endmodule



module bsg_fifo_1r1w_small_width_p32_els_p4
(
  clk_i,
  reset_i,
  v_i,
  ready_o,
  data_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o;

  bsg_fifo_1r1w_small_unhardened_width_p32_els_p4_ready_THEN_valid_p0
  \unhardened.un.fifo 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .ready_o(ready_o),
    .data_i(data_i),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );


endmodule



module bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  wire [63:0] \nz.mem ;
  reg \nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,\nz.mem_61_sv2v_reg ,
  \nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,\nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,
  \nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,\nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,
  \nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,\nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,
  \nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,\nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,
  \nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,\nz.mem_42_sv2v_reg ,
  \nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,\nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,
  \nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,\nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,
  \nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,\nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,
  \nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,\nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,
  \nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,\nz.mem_23_sv2v_reg ,
  \nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,\nz.mem_19_sv2v_reg ,
  \nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,\nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,
  \nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,\nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,
  \nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,\nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,
  \nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,\nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,
  \nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,\nz.mem_0_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[31] = (N3)? \nz.mem [31] : 
                        (N0)? \nz.mem [63] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[30] = (N3)? \nz.mem [30] : 
                        (N0)? \nz.mem [62] : 1'b0;
  assign r_data_o[29] = (N3)? \nz.mem [29] : 
                        (N0)? \nz.mem [61] : 1'b0;
  assign r_data_o[28] = (N3)? \nz.mem [28] : 
                        (N0)? \nz.mem [60] : 1'b0;
  assign r_data_o[27] = (N3)? \nz.mem [27] : 
                        (N0)? \nz.mem [59] : 1'b0;
  assign r_data_o[26] = (N3)? \nz.mem [26] : 
                        (N0)? \nz.mem [58] : 1'b0;
  assign r_data_o[25] = (N3)? \nz.mem [25] : 
                        (N0)? \nz.mem [57] : 1'b0;
  assign r_data_o[24] = (N3)? \nz.mem [24] : 
                        (N0)? \nz.mem [56] : 1'b0;
  assign r_data_o[23] = (N3)? \nz.mem [23] : 
                        (N0)? \nz.mem [55] : 1'b0;
  assign r_data_o[22] = (N3)? \nz.mem [22] : 
                        (N0)? \nz.mem [54] : 1'b0;
  assign r_data_o[21] = (N3)? \nz.mem [21] : 
                        (N0)? \nz.mem [53] : 1'b0;
  assign r_data_o[20] = (N3)? \nz.mem [20] : 
                        (N0)? \nz.mem [52] : 1'b0;
  assign r_data_o[19] = (N3)? \nz.mem [19] : 
                        (N0)? \nz.mem [51] : 1'b0;
  assign r_data_o[18] = (N3)? \nz.mem [18] : 
                        (N0)? \nz.mem [50] : 1'b0;
  assign r_data_o[17] = (N3)? \nz.mem [17] : 
                        (N0)? \nz.mem [49] : 1'b0;
  assign r_data_o[16] = (N3)? \nz.mem [16] : 
                        (N0)? \nz.mem [48] : 1'b0;
  assign r_data_o[15] = (N3)? \nz.mem [15] : 
                        (N0)? \nz.mem [47] : 1'b0;
  assign r_data_o[14] = (N3)? \nz.mem [14] : 
                        (N0)? \nz.mem [46] : 1'b0;
  assign r_data_o[13] = (N3)? \nz.mem [13] : 
                        (N0)? \nz.mem [45] : 1'b0;
  assign r_data_o[12] = (N3)? \nz.mem [12] : 
                        (N0)? \nz.mem [44] : 1'b0;
  assign r_data_o[11] = (N3)? \nz.mem [11] : 
                        (N0)? \nz.mem [43] : 1'b0;
  assign r_data_o[10] = (N3)? \nz.mem [10] : 
                        (N0)? \nz.mem [42] : 1'b0;
  assign r_data_o[9] = (N3)? \nz.mem [9] : 
                       (N0)? \nz.mem [41] : 1'b0;
  assign r_data_o[8] = (N3)? \nz.mem [8] : 
                       (N0)? \nz.mem [40] : 1'b0;
  assign r_data_o[7] = (N3)? \nz.mem [7] : 
                       (N0)? \nz.mem [39] : 1'b0;
  assign r_data_o[6] = (N3)? \nz.mem [6] : 
                       (N0)? \nz.mem [38] : 1'b0;
  assign r_data_o[5] = (N3)? \nz.mem [5] : 
                       (N0)? \nz.mem [37] : 1'b0;
  assign r_data_o[4] = (N3)? \nz.mem [4] : 
                       (N0)? \nz.mem [36] : 1'b0;
  assign r_data_o[3] = (N3)? \nz.mem [3] : 
                       (N0)? \nz.mem [35] : 1'b0;
  assign r_data_o[2] = (N3)? \nz.mem [2] : 
                       (N0)? \nz.mem [34] : 1'b0;
  assign r_data_o[1] = (N3)? \nz.mem [1] : 
                       (N0)? \nz.mem [33] : 1'b0;
  assign r_data_o[0] = (N3)? \nz.mem [0] : 
                       (N0)? \nz.mem [32] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      \nz.mem_63_sv2v_reg  <= w_data_i[31];
      \nz.mem_62_sv2v_reg  <= w_data_i[30];
      \nz.mem_61_sv2v_reg  <= w_data_i[29];
      \nz.mem_60_sv2v_reg  <= w_data_i[28];
      \nz.mem_59_sv2v_reg  <= w_data_i[27];
      \nz.mem_58_sv2v_reg  <= w_data_i[26];
      \nz.mem_57_sv2v_reg  <= w_data_i[25];
      \nz.mem_56_sv2v_reg  <= w_data_i[24];
      \nz.mem_55_sv2v_reg  <= w_data_i[23];
      \nz.mem_54_sv2v_reg  <= w_data_i[22];
      \nz.mem_53_sv2v_reg  <= w_data_i[21];
      \nz.mem_52_sv2v_reg  <= w_data_i[20];
      \nz.mem_51_sv2v_reg  <= w_data_i[19];
      \nz.mem_50_sv2v_reg  <= w_data_i[18];
      \nz.mem_49_sv2v_reg  <= w_data_i[17];
      \nz.mem_48_sv2v_reg  <= w_data_i[16];
      \nz.mem_47_sv2v_reg  <= w_data_i[15];
      \nz.mem_46_sv2v_reg  <= w_data_i[14];
      \nz.mem_45_sv2v_reg  <= w_data_i[13];
      \nz.mem_44_sv2v_reg  <= w_data_i[12];
      \nz.mem_43_sv2v_reg  <= w_data_i[11];
      \nz.mem_42_sv2v_reg  <= w_data_i[10];
      \nz.mem_41_sv2v_reg  <= w_data_i[9];
      \nz.mem_40_sv2v_reg  <= w_data_i[8];
      \nz.mem_39_sv2v_reg  <= w_data_i[7];
      \nz.mem_38_sv2v_reg  <= w_data_i[6];
      \nz.mem_37_sv2v_reg  <= w_data_i[5];
      \nz.mem_36_sv2v_reg  <= w_data_i[4];
      \nz.mem_35_sv2v_reg  <= w_data_i[3];
      \nz.mem_34_sv2v_reg  <= w_data_i[2];
      \nz.mem_33_sv2v_reg  <= w_data_i[1];
      \nz.mem_32_sv2v_reg  <= w_data_i[0];
    end 
    if(N7) begin
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [31:0] w_data_i;
  input [0:0] r_addr_i;
  output [31:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [31:0] r_data_o;

  bsg_mem_1r1w_synth_width_p32_els_p2_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p32
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [31:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,enq_i,tail_r,_0_net_,head_r,empty_r,full_r,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,N14;
  reg full_r_sv2v_reg,tail_r_sv2v_reg,head_r_sv2v_reg,empty_r_sv2v_reg;
  assign full_r = full_r_sv2v_reg;
  assign tail_r = tail_r_sv2v_reg;
  assign head_r = head_r_sv2v_reg;
  assign empty_r = empty_r_sv2v_reg;

  bsg_mem_1r1w_width_p32_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign _0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N5;
  assign N5 = ~full_r;
  assign N1 = enq_i;
  assign N0 = ~tail_r;
  assign N2 = ~head_r;
  assign N3 = N7 | N9;
  assign N7 = empty_r & N6;
  assign N6 = ~enq_i;
  assign N9 = N8 & N6;
  assign N8 = N5 & yumi_i;
  assign N4 = N13 | N14;
  assign N13 = N11 & N12;
  assign N11 = N10 & enq_i;
  assign N10 = ~empty_r;
  assign N12 = ~yumi_i;
  assign N14 = full_r & N12;

  always @(posedge clk_i) begin
    if(reset_i) begin
      full_r_sv2v_reg <= 1'b0;
      empty_r_sv2v_reg <= 1'b1;
    end else if(1'b1) begin
      full_r_sv2v_reg <= N4;
      empty_r_sv2v_reg <= N3;
    end 
    if(reset_i) begin
      tail_r_sv2v_reg <= 1'b0;
    end else if(N1) begin
      tail_r_sv2v_reg <= N0;
    end 
    if(reset_i) begin
      head_r_sv2v_reg <= 1'b0;
    end else if(yumi_i) begin
      head_r_sv2v_reg <= N2;
    end 
  end


endmodule



module bsg_expand_bitmask_in_width_p2_expand_p4
(
  i,
  o
);

  input [1:0] i;
  output [7:0] o;
  wire [7:0] o;
  wire o_7_,o_3_;
  assign o_7_ = i[1];
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;
  assign o_3_ = i[0];
  assign o[0] = o_3_;
  assign o[1] = o_3_;
  assign o[2] = o_3_;
  assign o[3] = o_3_;

endmodule



module bsg_mux_width_p4_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [7:0] data_i;
  input [0:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[7] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[6] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[5] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[4] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p1_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [3:0] data_i;
  input [1:0] sel_i;
  output [0:0] data_o;
  wire [0:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[1] : 
                     (N3)? data_i[2] : 
                     (N5)? data_i[3] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_expand_bitmask_in_width_p1_expand_p4
(
  i,
  o
);

  input [0:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire o_3_;
  assign o_3_ = i[0];
  assign o[0] = o_3_;
  assign o[1] = o_3_;
  assign o[2] = o_3_;
  assign o[3] = o_3_;

endmodule



module bsg_mux_width_p32_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [63:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1;
  assign data_o[31] = (N1)? data_i[31] : 
                      (N0)? data_i[63] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[30] = (N1)? data_i[30] : 
                      (N0)? data_i[62] : 1'b0;
  assign data_o[29] = (N1)? data_i[29] : 
                      (N0)? data_i[61] : 1'b0;
  assign data_o[28] = (N1)? data_i[28] : 
                      (N0)? data_i[60] : 1'b0;
  assign data_o[27] = (N1)? data_i[27] : 
                      (N0)? data_i[59] : 1'b0;
  assign data_o[26] = (N1)? data_i[26] : 
                      (N0)? data_i[58] : 1'b0;
  assign data_o[25] = (N1)? data_i[25] : 
                      (N0)? data_i[57] : 1'b0;
  assign data_o[24] = (N1)? data_i[24] : 
                      (N0)? data_i[56] : 1'b0;
  assign data_o[23] = (N1)? data_i[23] : 
                      (N0)? data_i[55] : 1'b0;
  assign data_o[22] = (N1)? data_i[22] : 
                      (N0)? data_i[54] : 1'b0;
  assign data_o[21] = (N1)? data_i[21] : 
                      (N0)? data_i[53] : 1'b0;
  assign data_o[20] = (N1)? data_i[20] : 
                      (N0)? data_i[52] : 1'b0;
  assign data_o[19] = (N1)? data_i[19] : 
                      (N0)? data_i[51] : 1'b0;
  assign data_o[18] = (N1)? data_i[18] : 
                      (N0)? data_i[50] : 1'b0;
  assign data_o[17] = (N1)? data_i[17] : 
                      (N0)? data_i[49] : 1'b0;
  assign data_o[16] = (N1)? data_i[16] : 
                      (N0)? data_i[48] : 1'b0;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[47] : 1'b0;
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[46] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[45] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[44] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[43] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[42] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[41] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[40] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[39] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[38] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[37] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[36] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[35] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[34] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[33] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[32] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_mux_width_p32_els_p1
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  assign data_o[31] = data_i[31];
  assign data_o[30] = data_i[30];
  assign data_o[29] = data_i[29];
  assign data_o[28] = data_i[28];
  assign data_o[27] = data_i[27];
  assign data_o[26] = data_i[26];
  assign data_o[25] = data_i[25];
  assign data_o[24] = data_i[24];
  assign data_o[23] = data_i[23];
  assign data_o[22] = data_i[22];
  assign data_o[21] = data_i[21];
  assign data_o[20] = data_i[20];
  assign data_o[19] = data_i[19];
  assign data_o[18] = data_i[18];
  assign data_o[17] = data_i[17];
  assign data_o[16] = data_i[16];
  assign data_o[15] = data_i[15];
  assign data_o[14] = data_i[14];
  assign data_o[13] = data_i[13];
  assign data_o[12] = data_i[12];
  assign data_o[11] = data_i[11];
  assign data_o[10] = data_i[10];
  assign data_o[9] = data_i[9];
  assign data_o[8] = data_i[8];
  assign data_o[7] = data_i[7];
  assign data_o[6] = data_i[6];
  assign data_o[5] = data_i[5];
  assign data_o[4] = data_i[4];
  assign data_o[3] = data_i[3];
  assign data_o[2] = data_i[2];
  assign data_o[1] = data_i[1];
  assign data_o[0] = data_i[0];

endmodule



module bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2_word_tracking_p1_dma_data_width_p32_debug_p0
(
  clk_i,
  reset_i,
  dma_cmd_i,
  dma_way_i,
  dma_addr_i,
  done_o,
  track_data_we_i,
  snoop_word_o,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  data_mem_v_o,
  data_mem_w_o,
  data_mem_addr_o,
  data_mem_w_mask_o,
  data_mem_data_o,
  data_mem_data_i,
  track_miss_i,
  track_mem_data_i,
  dma_evict_o
);

  input [3:0] dma_cmd_i;
  input [0:0] dma_way_i;
  input [27:0] dma_addr_i;
  output [31:0] snoop_word_o;
  output [32:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  output [7:0] data_mem_addr_o;
  output [7:0] data_mem_w_mask_o;
  output [63:0] data_mem_data_o;
  input [63:0] data_mem_data_i;
  input [7:0] track_mem_data_i;
  input clk_i;
  input reset_i;
  input track_data_we_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  input track_miss_i;
  output done_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output data_mem_v_o;
  output data_mem_w_o;
  output dma_evict_o;
  wire [31:0] snoop_word_o,dma_data_o,out_fifo_data_li,snoop_word_n;
  wire [32:0] dma_pkt_o;
  wire [7:0] data_mem_addr_o,data_mem_w_mask_o,dma_way_mask_expanded,track_mem_data_r;
  wire [63:0] data_mem_data_o;
  wire done_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,data_mem_v_o,data_mem_w_o,
  dma_evict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,dma_pkt_o_31_,dma_pkt_o_30_,
  dma_pkt_o_29_,dma_pkt_o_28_,dma_pkt_o_27_,dma_pkt_o_26_,dma_pkt_o_25_,dma_pkt_o_24_,
  dma_pkt_o_23_,dma_pkt_o_22_,dma_pkt_o_21_,dma_pkt_o_20_,dma_pkt_o_19_,
  dma_pkt_o_18_,dma_pkt_o_17_,dma_pkt_o_16_,dma_pkt_o_15_,dma_pkt_o_14_,data_mem_addr_o_7_,
  data_mem_addr_o_6_,data_mem_addr_o_5_,data_mem_addr_o_4_,data_mem_addr_o_3_,
  data_mem_addr_o_2_,data_mem_data_o_1__31_,data_mem_data_o_1__30_,data_mem_data_o_1__29_,
  data_mem_data_o_1__28_,data_mem_data_o_1__27_,data_mem_data_o_1__26_,
  data_mem_data_o_1__25_,data_mem_data_o_1__24_,data_mem_data_o_1__23_,
  data_mem_data_o_1__22_,data_mem_data_o_1__21_,data_mem_data_o_1__20_,data_mem_data_o_1__19_,
  data_mem_data_o_1__18_,data_mem_data_o_1__17_,data_mem_data_o_1__16_,
  data_mem_data_o_1__15_,data_mem_data_o_1__14_,data_mem_data_o_1__13_,data_mem_data_o_1__12_,
  data_mem_data_o_1__11_,data_mem_data_o_1__10_,data_mem_data_o_1__9_,
  data_mem_data_o_1__8_,data_mem_data_o_1__7_,data_mem_data_o_1__6_,data_mem_data_o_1__5_,
  data_mem_data_o_1__4_,data_mem_data_o_1__3_,data_mem_data_o_1__2_,data_mem_data_o_1__1_,
  data_mem_data_o_1__0_,counter_clear,counter_up,in_fifo_v_lo,in_fifo_yumi_li,
  out_fifo_v_li,out_fifo_ready_lo,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,
  N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,
  N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,
  N66,N67,N68,N69,N70,N71,snoop_word_we,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89;
  wire [2:2] counter_r;
  wire [1:0] dma_way_mask,dma_state_r,dma_state_n;
  wire [3:0] track_data_way_picked,track_bits_offset_picked_expanded,
  data_mem_w_mask_way_picked;
  wire [0:0] track_bits_offset_picked;
  reg track_mem_data_r_7_sv2v_reg,track_mem_data_r_6_sv2v_reg,
  track_mem_data_r_5_sv2v_reg,track_mem_data_r_4_sv2v_reg,track_mem_data_r_3_sv2v_reg,
  track_mem_data_r_2_sv2v_reg,track_mem_data_r_1_sv2v_reg,track_mem_data_r_0_sv2v_reg,
  dma_state_r_1_sv2v_reg,dma_state_r_0_sv2v_reg,snoop_word_o_31_sv2v_reg,snoop_word_o_30_sv2v_reg,
  snoop_word_o_29_sv2v_reg,snoop_word_o_28_sv2v_reg,snoop_word_o_27_sv2v_reg,
  snoop_word_o_26_sv2v_reg,snoop_word_o_25_sv2v_reg,snoop_word_o_24_sv2v_reg,
  snoop_word_o_23_sv2v_reg,snoop_word_o_22_sv2v_reg,snoop_word_o_21_sv2v_reg,
  snoop_word_o_20_sv2v_reg,snoop_word_o_19_sv2v_reg,snoop_word_o_18_sv2v_reg,
  snoop_word_o_17_sv2v_reg,snoop_word_o_16_sv2v_reg,snoop_word_o_15_sv2v_reg,snoop_word_o_14_sv2v_reg,
  snoop_word_o_13_sv2v_reg,snoop_word_o_12_sv2v_reg,snoop_word_o_11_sv2v_reg,
  snoop_word_o_10_sv2v_reg,snoop_word_o_9_sv2v_reg,snoop_word_o_8_sv2v_reg,
  snoop_word_o_7_sv2v_reg,snoop_word_o_6_sv2v_reg,snoop_word_o_5_sv2v_reg,
  snoop_word_o_4_sv2v_reg,snoop_word_o_3_sv2v_reg,snoop_word_o_2_sv2v_reg,snoop_word_o_1_sv2v_reg,
  snoop_word_o_0_sv2v_reg;
  assign track_mem_data_r[7] = track_mem_data_r_7_sv2v_reg;
  assign track_mem_data_r[6] = track_mem_data_r_6_sv2v_reg;
  assign track_mem_data_r[5] = track_mem_data_r_5_sv2v_reg;
  assign track_mem_data_r[4] = track_mem_data_r_4_sv2v_reg;
  assign track_mem_data_r[3] = track_mem_data_r_3_sv2v_reg;
  assign track_mem_data_r[2] = track_mem_data_r_2_sv2v_reg;
  assign track_mem_data_r[1] = track_mem_data_r_1_sv2v_reg;
  assign track_mem_data_r[0] = track_mem_data_r_0_sv2v_reg;
  assign dma_state_r[1] = dma_state_r_1_sv2v_reg;
  assign dma_state_r[0] = dma_state_r_0_sv2v_reg;
  assign snoop_word_o[31] = snoop_word_o_31_sv2v_reg;
  assign snoop_word_o[30] = snoop_word_o_30_sv2v_reg;
  assign snoop_word_o[29] = snoop_word_o_29_sv2v_reg;
  assign snoop_word_o[28] = snoop_word_o_28_sv2v_reg;
  assign snoop_word_o[27] = snoop_word_o_27_sv2v_reg;
  assign snoop_word_o[26] = snoop_word_o_26_sv2v_reg;
  assign snoop_word_o[25] = snoop_word_o_25_sv2v_reg;
  assign snoop_word_o[24] = snoop_word_o_24_sv2v_reg;
  assign snoop_word_o[23] = snoop_word_o_23_sv2v_reg;
  assign snoop_word_o[22] = snoop_word_o_22_sv2v_reg;
  assign snoop_word_o[21] = snoop_word_o_21_sv2v_reg;
  assign snoop_word_o[20] = snoop_word_o_20_sv2v_reg;
  assign snoop_word_o[19] = snoop_word_o_19_sv2v_reg;
  assign snoop_word_o[18] = snoop_word_o_18_sv2v_reg;
  assign snoop_word_o[17] = snoop_word_o_17_sv2v_reg;
  assign snoop_word_o[16] = snoop_word_o_16_sv2v_reg;
  assign snoop_word_o[15] = snoop_word_o_15_sv2v_reg;
  assign snoop_word_o[14] = snoop_word_o_14_sv2v_reg;
  assign snoop_word_o[13] = snoop_word_o_13_sv2v_reg;
  assign snoop_word_o[12] = snoop_word_o_12_sv2v_reg;
  assign snoop_word_o[11] = snoop_word_o_11_sv2v_reg;
  assign snoop_word_o[10] = snoop_word_o_10_sv2v_reg;
  assign snoop_word_o[9] = snoop_word_o_9_sv2v_reg;
  assign snoop_word_o[8] = snoop_word_o_8_sv2v_reg;
  assign snoop_word_o[7] = snoop_word_o_7_sv2v_reg;
  assign snoop_word_o[6] = snoop_word_o_6_sv2v_reg;
  assign snoop_word_o[5] = snoop_word_o_5_sv2v_reg;
  assign snoop_word_o[4] = snoop_word_o_4_sv2v_reg;
  assign snoop_word_o[3] = snoop_word_o_3_sv2v_reg;
  assign snoop_word_o[2] = snoop_word_o_2_sv2v_reg;
  assign snoop_word_o[1] = snoop_word_o_1_sv2v_reg;
  assign snoop_word_o[0] = snoop_word_o_0_sv2v_reg;
  assign dma_pkt_o[4] = 1'b0;
  assign dma_pkt_o[5] = 1'b0;
  assign dma_pkt_o[6] = 1'b0;
  assign dma_pkt_o[7] = 1'b0;
  assign dma_pkt_o_31_ = dma_addr_i[27];
  assign dma_pkt_o[31] = dma_pkt_o_31_;
  assign dma_pkt_o_30_ = dma_addr_i[26];
  assign dma_pkt_o[30] = dma_pkt_o_30_;
  assign dma_pkt_o_29_ = dma_addr_i[25];
  assign dma_pkt_o[29] = dma_pkt_o_29_;
  assign dma_pkt_o_28_ = dma_addr_i[24];
  assign dma_pkt_o[28] = dma_pkt_o_28_;
  assign dma_pkt_o_27_ = dma_addr_i[23];
  assign dma_pkt_o[27] = dma_pkt_o_27_;
  assign dma_pkt_o_26_ = dma_addr_i[22];
  assign dma_pkt_o[26] = dma_pkt_o_26_;
  assign dma_pkt_o_25_ = dma_addr_i[21];
  assign dma_pkt_o[25] = dma_pkt_o_25_;
  assign dma_pkt_o_24_ = dma_addr_i[20];
  assign dma_pkt_o[24] = dma_pkt_o_24_;
  assign dma_pkt_o_23_ = dma_addr_i[19];
  assign dma_pkt_o[23] = dma_pkt_o_23_;
  assign dma_pkt_o_22_ = dma_addr_i[18];
  assign dma_pkt_o[22] = dma_pkt_o_22_;
  assign dma_pkt_o_21_ = dma_addr_i[17];
  assign dma_pkt_o[21] = dma_pkt_o_21_;
  assign dma_pkt_o_20_ = dma_addr_i[16];
  assign dma_pkt_o[20] = dma_pkt_o_20_;
  assign dma_pkt_o_19_ = dma_addr_i[15];
  assign dma_pkt_o[19] = dma_pkt_o_19_;
  assign dma_pkt_o_18_ = dma_addr_i[14];
  assign dma_pkt_o[18] = dma_pkt_o_18_;
  assign dma_pkt_o_17_ = dma_addr_i[13];
  assign dma_pkt_o[17] = dma_pkt_o_17_;
  assign dma_pkt_o_16_ = dma_addr_i[12];
  assign dma_pkt_o[16] = dma_pkt_o_16_;
  assign dma_pkt_o_15_ = dma_addr_i[11];
  assign dma_pkt_o[15] = dma_pkt_o_15_;
  assign dma_pkt_o_14_ = dma_addr_i[10];
  assign dma_pkt_o[14] = dma_pkt_o_14_;
  assign data_mem_addr_o_7_ = dma_addr_i[9];
  assign dma_pkt_o[13] = data_mem_addr_o_7_;
  assign data_mem_addr_o[7] = data_mem_addr_o_7_;
  assign data_mem_addr_o_6_ = dma_addr_i[8];
  assign dma_pkt_o[12] = data_mem_addr_o_6_;
  assign data_mem_addr_o[6] = data_mem_addr_o_6_;
  assign data_mem_addr_o_5_ = dma_addr_i[7];
  assign dma_pkt_o[11] = data_mem_addr_o_5_;
  assign data_mem_addr_o[5] = data_mem_addr_o_5_;
  assign data_mem_addr_o_4_ = dma_addr_i[6];
  assign dma_pkt_o[10] = data_mem_addr_o_4_;
  assign data_mem_addr_o[4] = data_mem_addr_o_4_;
  assign data_mem_addr_o_3_ = dma_addr_i[5];
  assign dma_pkt_o[9] = data_mem_addr_o_3_;
  assign data_mem_addr_o[3] = data_mem_addr_o_3_;
  assign data_mem_addr_o_2_ = dma_addr_i[4];
  assign dma_pkt_o[8] = data_mem_addr_o_2_;
  assign data_mem_addr_o[2] = data_mem_addr_o_2_;
  assign data_mem_data_o[31] = data_mem_data_o_1__31_;
  assign data_mem_data_o[63] = data_mem_data_o_1__31_;
  assign data_mem_data_o[30] = data_mem_data_o_1__30_;
  assign data_mem_data_o[62] = data_mem_data_o_1__30_;
  assign data_mem_data_o[29] = data_mem_data_o_1__29_;
  assign data_mem_data_o[61] = data_mem_data_o_1__29_;
  assign data_mem_data_o[28] = data_mem_data_o_1__28_;
  assign data_mem_data_o[60] = data_mem_data_o_1__28_;
  assign data_mem_data_o[27] = data_mem_data_o_1__27_;
  assign data_mem_data_o[59] = data_mem_data_o_1__27_;
  assign data_mem_data_o[26] = data_mem_data_o_1__26_;
  assign data_mem_data_o[58] = data_mem_data_o_1__26_;
  assign data_mem_data_o[25] = data_mem_data_o_1__25_;
  assign data_mem_data_o[57] = data_mem_data_o_1__25_;
  assign data_mem_data_o[24] = data_mem_data_o_1__24_;
  assign data_mem_data_o[56] = data_mem_data_o_1__24_;
  assign data_mem_data_o[23] = data_mem_data_o_1__23_;
  assign data_mem_data_o[55] = data_mem_data_o_1__23_;
  assign data_mem_data_o[22] = data_mem_data_o_1__22_;
  assign data_mem_data_o[54] = data_mem_data_o_1__22_;
  assign data_mem_data_o[21] = data_mem_data_o_1__21_;
  assign data_mem_data_o[53] = data_mem_data_o_1__21_;
  assign data_mem_data_o[20] = data_mem_data_o_1__20_;
  assign data_mem_data_o[52] = data_mem_data_o_1__20_;
  assign data_mem_data_o[19] = data_mem_data_o_1__19_;
  assign data_mem_data_o[51] = data_mem_data_o_1__19_;
  assign data_mem_data_o[18] = data_mem_data_o_1__18_;
  assign data_mem_data_o[50] = data_mem_data_o_1__18_;
  assign data_mem_data_o[17] = data_mem_data_o_1__17_;
  assign data_mem_data_o[49] = data_mem_data_o_1__17_;
  assign data_mem_data_o[16] = data_mem_data_o_1__16_;
  assign data_mem_data_o[48] = data_mem_data_o_1__16_;
  assign data_mem_data_o[15] = data_mem_data_o_1__15_;
  assign data_mem_data_o[47] = data_mem_data_o_1__15_;
  assign data_mem_data_o[14] = data_mem_data_o_1__14_;
  assign data_mem_data_o[46] = data_mem_data_o_1__14_;
  assign data_mem_data_o[13] = data_mem_data_o_1__13_;
  assign data_mem_data_o[45] = data_mem_data_o_1__13_;
  assign data_mem_data_o[12] = data_mem_data_o_1__12_;
  assign data_mem_data_o[44] = data_mem_data_o_1__12_;
  assign data_mem_data_o[11] = data_mem_data_o_1__11_;
  assign data_mem_data_o[43] = data_mem_data_o_1__11_;
  assign data_mem_data_o[10] = data_mem_data_o_1__10_;
  assign data_mem_data_o[42] = data_mem_data_o_1__10_;
  assign data_mem_data_o[9] = data_mem_data_o_1__9_;
  assign data_mem_data_o[41] = data_mem_data_o_1__9_;
  assign data_mem_data_o[8] = data_mem_data_o_1__8_;
  assign data_mem_data_o[40] = data_mem_data_o_1__8_;
  assign data_mem_data_o[7] = data_mem_data_o_1__7_;
  assign data_mem_data_o[39] = data_mem_data_o_1__7_;
  assign data_mem_data_o[6] = data_mem_data_o_1__6_;
  assign data_mem_data_o[38] = data_mem_data_o_1__6_;
  assign data_mem_data_o[5] = data_mem_data_o_1__5_;
  assign data_mem_data_o[37] = data_mem_data_o_1__5_;
  assign data_mem_data_o[4] = data_mem_data_o_1__4_;
  assign data_mem_data_o[36] = data_mem_data_o_1__4_;
  assign data_mem_data_o[3] = data_mem_data_o_1__3_;
  assign data_mem_data_o[35] = data_mem_data_o_1__3_;
  assign data_mem_data_o[2] = data_mem_data_o_1__2_;
  assign data_mem_data_o[34] = data_mem_data_o_1__2_;
  assign data_mem_data_o[1] = data_mem_data_o_1__1_;
  assign data_mem_data_o[33] = data_mem_data_o_1__1_;
  assign data_mem_data_o[0] = data_mem_data_o_1__0_;
  assign data_mem_data_o[32] = data_mem_data_o_1__0_;

  bsg_counter_clear_up_4_0
  dma_counter
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(counter_clear),
    .up_i(counter_up),
    .count_o({ counter_r[2:2], data_mem_addr_o[1:0] })
  );


  bsg_fifo_1r1w_small_width_p32_els_p4
  in_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(dma_data_v_i),
    .ready_o(dma_data_ready_o),
    .data_i(dma_data_i),
    .v_o(in_fifo_v_lo),
    .data_o({ data_mem_data_o_1__31_, data_mem_data_o_1__30_, data_mem_data_o_1__29_, data_mem_data_o_1__28_, data_mem_data_o_1__27_, data_mem_data_o_1__26_, data_mem_data_o_1__25_, data_mem_data_o_1__24_, data_mem_data_o_1__23_, data_mem_data_o_1__22_, data_mem_data_o_1__21_, data_mem_data_o_1__20_, data_mem_data_o_1__19_, data_mem_data_o_1__18_, data_mem_data_o_1__17_, data_mem_data_o_1__16_, data_mem_data_o_1__15_, data_mem_data_o_1__14_, data_mem_data_o_1__13_, data_mem_data_o_1__12_, data_mem_data_o_1__11_, data_mem_data_o_1__10_, data_mem_data_o_1__9_, data_mem_data_o_1__8_, data_mem_data_o_1__7_, data_mem_data_o_1__6_, data_mem_data_o_1__5_, data_mem_data_o_1__4_, data_mem_data_o_1__3_, data_mem_data_o_1__2_, data_mem_data_o_1__1_, data_mem_data_o_1__0_ }),
    .yumi_i(in_fifo_yumi_li)
  );


  bsg_two_fifo_width_p32
  out_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(out_fifo_ready_lo),
    .data_i(out_fifo_data_li),
    .v_i(out_fifo_v_li),
    .v_o(dma_data_v_o),
    .data_o(dma_data_o),
    .yumi_i(dma_data_yumi_i)
  );


  bsg_decode_num_out_p2
  dma_way_demux
  (
    .i(dma_way_i[0]),
    .o(dma_way_mask)
  );


  bsg_expand_bitmask_in_width_p2_expand_p4
  expand0
  (
    .i(dma_way_mask),
    .o(dma_way_mask_expanded)
  );


  bsg_mux_width_p4_els_p2
  track_way_mux
  (
    .data_i(track_mem_data_r),
    .sel_i(dma_way_i[0]),
    .data_o(track_data_way_picked)
  );


  bsg_mux_width_p1_els_p4
  track_offset_mux
  (
    .data_i(track_data_way_picked),
    .sel_i(data_mem_addr_o[1:0]),
    .data_o(track_bits_offset_picked[0])
  );


  bsg_expand_bitmask_in_width_p1_expand_p4
  expand1
  (
    .i(track_bits_offset_picked[0]),
    .o(track_bits_offset_picked_expanded)
  );


  bsg_mux_width_p32_els_p2
  write_data_mux
  (
    .data_i(data_mem_data_i),
    .sel_i(dma_way_i[0]),
    .data_o(out_fifo_data_li)
  );

  assign N18 = N17 & N85;
  assign N19 = dma_state_r[1] | N85;
  assign N21 = N17 | dma_state_r[0];
  assign N23 = dma_state_r[1] & dma_state_r[0];
  assign N24 = dma_cmd_i[1] | N41;
  assign N25 = N27 | N24;
  assign N27 = dma_cmd_i[3] | dma_cmd_i[2];
  assign N28 = N40 | dma_cmd_i[0];
  assign N29 = N27 | N28;
  assign N31 = dma_cmd_i[3] | N39;
  assign N32 = N31 | N35;
  assign N34 = N38 | dma_cmd_i[2];
  assign N35 = dma_cmd_i[1] | dma_cmd_i[0];
  assign N36 = N34 | N35;
  assign N42 = N38 & N39;
  assign N43 = N40 & N41;
  assign N44 = N42 & N43;
  assign N71 = data_mem_addr_o[1:0] == dma_addr_i[3:2];

  bsg_mux_width_p32_els_p1
  snoop_mux0
  (
    .data_i({ data_mem_data_o_1__31_, data_mem_data_o_1__30_, data_mem_data_o_1__29_, data_mem_data_o_1__28_, data_mem_data_o_1__27_, data_mem_data_o_1__26_, data_mem_data_o_1__25_, data_mem_data_o_1__24_, data_mem_data_o_1__23_, data_mem_data_o_1__22_, data_mem_data_o_1__21_, data_mem_data_o_1__20_, data_mem_data_o_1__19_, data_mem_data_o_1__18_, data_mem_data_o_1__17_, data_mem_data_o_1__16_, data_mem_data_o_1__15_, data_mem_data_o_1__14_, data_mem_data_o_1__13_, data_mem_data_o_1__12_, data_mem_data_o_1__11_, data_mem_data_o_1__10_, data_mem_data_o_1__9_, data_mem_data_o_1__8_, data_mem_data_o_1__7_, data_mem_data_o_1__6_, data_mem_data_o_1__5_, data_mem_data_o_1__4_, data_mem_data_o_1__3_, data_mem_data_o_1__2_, data_mem_data_o_1__1_, data_mem_data_o_1__0_ }),
    .sel_i(dma_addr_i[2]),
    .data_o(snoop_word_n)
  );

  assign N76 = ~counter_r[2];
  assign N77 = data_mem_addr_o[1] | N76;
  assign N78 = data_mem_addr_o[0] | N77;
  assign N79 = ~N78;
  assign N80 = ~data_mem_addr_o[1];
  assign N81 = ~data_mem_addr_o[0];
  assign N82 = N80 | counter_r[2];
  assign N83 = N81 | N82;
  assign N84 = ~N83;
  assign N85 = ~dma_state_r[0];
  assign N86 = N85 | dma_state_r[1];
  assign N87 = ~N86;
  assign data_mem_w_mask_way_picked = (N0)? { N13, N14, N15, N16 } : 
                                      (N12)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign N0 = track_miss_i;
  assign N50 = (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N1 = N26;
  assign N2 = N30;
  assign N3 = N33;
  assign N4 = N37;
  assign N5 = N44;
  assign { N55, N54, N53, N52, N51 } = (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N2)? { 1'b1, track_data_way_picked } : 
                                       (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                       (N49)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N56 = (N1)? dma_pkt_yumi_i : 
               (N2)? dma_pkt_yumi_i : 
               (N3)? 1'b0 : 
               (N4)? 1'b0 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N57 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b1 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N58 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? 1'b1 : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N59 = (N1)? 1'b0 : 
               (N2)? 1'b0 : 
               (N3)? 1'b0 : 
               (N4)? track_bits_offset_picked[0] : 
               (N5)? 1'b0 : 
               (N49)? 1'b0 : 1'b0;
  assign N61 = ~N60;
  assign N66 = ~N65;
  assign counter_clear = (N6)? N57 : 
                         (N7)? N63 : 
                         (N8)? N68 : 
                         (N9)? 1'b0 : 1'b0;
  assign N6 = N18;
  assign N7 = N20;
  assign N8 = N22;
  assign N9 = N23;
  assign counter_up = (N6)? N58 : 
                      (N7)? N62 : 
                      (N8)? N67 : 
                      (N9)? 1'b0 : 1'b0;
  assign data_mem_v_o = (N6)? N59 : 
                        (N7)? in_fifo_v_lo : 
                        (N8)? N69 : 
                        (N9)? 1'b0 : 1'b0;
  assign dma_pkt_v_o = (N6)? N50 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b0 : 
                       (N9)? 1'b0 : 1'b0;
  assign { dma_pkt_o[32:32], dma_pkt_o[3:0] } = (N6)? { N55, N54, N53, N52, N51 } : 
                                                (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N8)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign done_o = (N6)? N56 : 
                  (N7)? N64 : 
                  (N8)? N70 : 
                  (N9)? 1'b0 : 1'b0;
  assign dma_state_n = (N6)? { N37, N33 } : 
                       (N7)? { 1'b0, N61 } : 
                       (N8)? { N66, 1'b0 } : 
                       (N9)? { 1'b0, 1'b0 } : 1'b0;
  assign data_mem_w_o = (N6)? 1'b0 : 
                        (N7)? in_fifo_v_lo : 
                        (N8)? 1'b0 : 
                        (N9)? 1'b0 : 1'b0;
  assign in_fifo_yumi_li = (N6)? 1'b0 : 
                           (N7)? in_fifo_v_lo : 
                           (N8)? 1'b0 : 
                           (N9)? 1'b0 : 1'b0;
  assign out_fifo_v_li = (N6)? 1'b0 : 
                         (N7)? 1'b0 : 
                         (N8)? 1'b1 : 
                         (N9)? 1'b0 : 1'b0;
  assign dma_evict_o = (N6)? 1'b0 : 
                       (N7)? 1'b0 : 
                       (N8)? 1'b1 : 
                       (N9)? 1'b0 : 1'b0;
  assign N74 = (N10)? 1'b0 : 
               (N11)? snoop_word_we : 1'b0;
  assign N10 = N73;
  assign N11 = N72;
  assign N75 = (N10)? 1'b0 : 
               (N11)? track_data_we_i : 1'b0;
  assign N12 = ~track_miss_i;
  assign N13 = ~track_bits_offset_picked_expanded[3];
  assign N14 = ~track_bits_offset_picked_expanded[2];
  assign N15 = ~track_bits_offset_picked_expanded[1];
  assign N16 = ~track_bits_offset_picked_expanded[0];
  assign data_mem_w_mask_o[7] = dma_way_mask_expanded[7] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[6] = dma_way_mask_expanded[6] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[5] = dma_way_mask_expanded[5] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[4] = dma_way_mask_expanded[4] & data_mem_w_mask_way_picked[0];
  assign data_mem_w_mask_o[3] = dma_way_mask_expanded[3] & data_mem_w_mask_way_picked[3];
  assign data_mem_w_mask_o[2] = dma_way_mask_expanded[2] & data_mem_w_mask_way_picked[2];
  assign data_mem_w_mask_o[1] = dma_way_mask_expanded[1] & data_mem_w_mask_way_picked[1];
  assign data_mem_w_mask_o[0] = dma_way_mask_expanded[0] & data_mem_w_mask_way_picked[0];
  assign N17 = ~dma_state_r[1];
  assign N20 = ~N19;
  assign N22 = ~N21;
  assign N26 = ~N25;
  assign N30 = ~N29;
  assign N33 = ~N32;
  assign N37 = ~N36;
  assign N38 = ~dma_cmd_i[3];
  assign N39 = ~dma_cmd_i[2];
  assign N40 = ~dma_cmd_i[1];
  assign N41 = ~dma_cmd_i[0];
  assign N45 = N30 | N26;
  assign N46 = N33 | N45;
  assign N47 = N37 | N46;
  assign N48 = N44 | N47;
  assign N49 = ~N48;
  assign N60 = N84 & in_fifo_v_lo;
  assign N62 = in_fifo_v_lo & N83;
  assign N63 = in_fifo_v_lo & N84;
  assign N64 = N84 & in_fifo_v_lo;
  assign N65 = N79 & out_fifo_ready_lo;
  assign N67 = out_fifo_ready_lo & N78;
  assign N68 = out_fifo_ready_lo & N79;
  assign N69 = N88 & track_bits_offset_picked[0];
  assign N88 = out_fifo_ready_lo & N78;
  assign N70 = N79 & out_fifo_ready_lo;
  assign snoop_word_we = N89 & N71;
  assign N89 = N87 & in_fifo_v_lo;
  assign N72 = ~reset_i;
  assign N73 = reset_i;

  always @(posedge clk_i) begin
    if(N75) begin
      track_mem_data_r_7_sv2v_reg <= track_mem_data_i[7];
      track_mem_data_r_6_sv2v_reg <= track_mem_data_i[6];
      track_mem_data_r_5_sv2v_reg <= track_mem_data_i[5];
      track_mem_data_r_4_sv2v_reg <= track_mem_data_i[4];
      track_mem_data_r_3_sv2v_reg <= track_mem_data_i[3];
      track_mem_data_r_2_sv2v_reg <= track_mem_data_i[2];
      track_mem_data_r_1_sv2v_reg <= track_mem_data_i[1];
      track_mem_data_r_0_sv2v_reg <= track_mem_data_i[0];
    end 
    if(reset_i) begin
      dma_state_r_1_sv2v_reg <= 1'b0;
      dma_state_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      dma_state_r_1_sv2v_reg <= dma_state_n[1];
      dma_state_r_0_sv2v_reg <= dma_state_n[0];
    end 
    if(N74) begin
      snoop_word_o_31_sv2v_reg <= snoop_word_n[31];
      snoop_word_o_30_sv2v_reg <= snoop_word_n[30];
      snoop_word_o_29_sv2v_reg <= snoop_word_n[29];
      snoop_word_o_28_sv2v_reg <= snoop_word_n[28];
      snoop_word_o_27_sv2v_reg <= snoop_word_n[27];
      snoop_word_o_26_sv2v_reg <= snoop_word_n[26];
      snoop_word_o_25_sv2v_reg <= snoop_word_n[25];
      snoop_word_o_24_sv2v_reg <= snoop_word_n[24];
      snoop_word_o_23_sv2v_reg <= snoop_word_n[23];
      snoop_word_o_22_sv2v_reg <= snoop_word_n[22];
      snoop_word_o_21_sv2v_reg <= snoop_word_n[21];
      snoop_word_o_20_sv2v_reg <= snoop_word_n[20];
      snoop_word_o_19_sv2v_reg <= snoop_word_n[19];
      snoop_word_o_18_sv2v_reg <= snoop_word_n[18];
      snoop_word_o_17_sv2v_reg <= snoop_word_n[17];
      snoop_word_o_16_sv2v_reg <= snoop_word_n[16];
      snoop_word_o_15_sv2v_reg <= snoop_word_n[15];
      snoop_word_o_14_sv2v_reg <= snoop_word_n[14];
      snoop_word_o_13_sv2v_reg <= snoop_word_n[13];
      snoop_word_o_12_sv2v_reg <= snoop_word_n[12];
      snoop_word_o_11_sv2v_reg <= snoop_word_n[11];
      snoop_word_o_10_sv2v_reg <= snoop_word_n[10];
      snoop_word_o_9_sv2v_reg <= snoop_word_n[9];
      snoop_word_o_8_sv2v_reg <= snoop_word_n[8];
      snoop_word_o_7_sv2v_reg <= snoop_word_n[7];
      snoop_word_o_6_sv2v_reg <= snoop_word_n[6];
      snoop_word_o_5_sv2v_reg <= snoop_word_n[5];
      snoop_word_o_4_sv2v_reg <= snoop_word_n[4];
      snoop_word_o_3_sv2v_reg <= snoop_word_n[3];
      snoop_word_o_2_sv2v_reg <= snoop_word_n[2];
      snoop_word_o_1_sv2v_reg <= snoop_word_n[1];
      snoop_word_o_0_sv2v_reg <= snoop_word_n[0];
    end 
  end


endmodule



module bsg_cache_buffer_queue_width_p65
(
  clk_i,
  reset_i,
  v_i,
  data_i,
  v_o,
  data_o,
  yumi_i,
  el0_valid_o,
  el1_valid_o,
  el0_snoop_o,
  el1_snoop_o,
  empty_o,
  full_o
);

  input [64:0] data_i;
  output [64:0] data_o;
  output [64:0] el0_snoop_o;
  output [64:0] el1_snoop_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output v_o;
  output el0_valid_o;
  output el1_valid_o;
  output empty_o;
  output full_o;
  wire [64:0] data_o,el0_snoop_o,el1_snoop_o;
  wire v_o,el0_valid_o,el1_valid_o,empty_o,full_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,
  N11,N12,N13,N14,N15,el0_enable,el1_enable,mux0_sel,mux1_sel,N16,N17,N18,N19,N20,
  N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,
  N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,
  N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,
  N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91;
  wire [1:0] num_els_r;
  reg num_els_r_1_sv2v_reg,num_els_r_0_sv2v_reg,el0_snoop_o_64_sv2v_reg,
  el0_snoop_o_63_sv2v_reg,el0_snoop_o_62_sv2v_reg,el0_snoop_o_61_sv2v_reg,
  el0_snoop_o_60_sv2v_reg,el0_snoop_o_59_sv2v_reg,el0_snoop_o_58_sv2v_reg,el0_snoop_o_57_sv2v_reg,
  el0_snoop_o_56_sv2v_reg,el0_snoop_o_55_sv2v_reg,el0_snoop_o_54_sv2v_reg,
  el0_snoop_o_53_sv2v_reg,el0_snoop_o_52_sv2v_reg,el0_snoop_o_51_sv2v_reg,
  el0_snoop_o_50_sv2v_reg,el0_snoop_o_49_sv2v_reg,el0_snoop_o_48_sv2v_reg,el0_snoop_o_47_sv2v_reg,
  el0_snoop_o_46_sv2v_reg,el0_snoop_o_45_sv2v_reg,el0_snoop_o_44_sv2v_reg,
  el0_snoop_o_43_sv2v_reg,el0_snoop_o_42_sv2v_reg,el0_snoop_o_41_sv2v_reg,
  el0_snoop_o_40_sv2v_reg,el0_snoop_o_39_sv2v_reg,el0_snoop_o_38_sv2v_reg,el0_snoop_o_37_sv2v_reg,
  el0_snoop_o_36_sv2v_reg,el0_snoop_o_35_sv2v_reg,el0_snoop_o_34_sv2v_reg,
  el0_snoop_o_33_sv2v_reg,el0_snoop_o_32_sv2v_reg,el0_snoop_o_31_sv2v_reg,
  el0_snoop_o_30_sv2v_reg,el0_snoop_o_29_sv2v_reg,el0_snoop_o_28_sv2v_reg,el0_snoop_o_27_sv2v_reg,
  el0_snoop_o_26_sv2v_reg,el0_snoop_o_25_sv2v_reg,el0_snoop_o_24_sv2v_reg,
  el0_snoop_o_23_sv2v_reg,el0_snoop_o_22_sv2v_reg,el0_snoop_o_21_sv2v_reg,
  el0_snoop_o_20_sv2v_reg,el0_snoop_o_19_sv2v_reg,el0_snoop_o_18_sv2v_reg,el0_snoop_o_17_sv2v_reg,
  el0_snoop_o_16_sv2v_reg,el0_snoop_o_15_sv2v_reg,el0_snoop_o_14_sv2v_reg,
  el0_snoop_o_13_sv2v_reg,el0_snoop_o_12_sv2v_reg,el0_snoop_o_11_sv2v_reg,
  el0_snoop_o_10_sv2v_reg,el0_snoop_o_9_sv2v_reg,el0_snoop_o_8_sv2v_reg,el0_snoop_o_7_sv2v_reg,
  el0_snoop_o_6_sv2v_reg,el0_snoop_o_5_sv2v_reg,el0_snoop_o_4_sv2v_reg,
  el0_snoop_o_3_sv2v_reg,el0_snoop_o_2_sv2v_reg,el0_snoop_o_1_sv2v_reg,el0_snoop_o_0_sv2v_reg,
  el1_snoop_o_64_sv2v_reg,el1_snoop_o_63_sv2v_reg,el1_snoop_o_62_sv2v_reg,
  el1_snoop_o_61_sv2v_reg,el1_snoop_o_60_sv2v_reg,el1_snoop_o_59_sv2v_reg,el1_snoop_o_58_sv2v_reg,
  el1_snoop_o_57_sv2v_reg,el1_snoop_o_56_sv2v_reg,el1_snoop_o_55_sv2v_reg,
  el1_snoop_o_54_sv2v_reg,el1_snoop_o_53_sv2v_reg,el1_snoop_o_52_sv2v_reg,
  el1_snoop_o_51_sv2v_reg,el1_snoop_o_50_sv2v_reg,el1_snoop_o_49_sv2v_reg,el1_snoop_o_48_sv2v_reg,
  el1_snoop_o_47_sv2v_reg,el1_snoop_o_46_sv2v_reg,el1_snoop_o_45_sv2v_reg,
  el1_snoop_o_44_sv2v_reg,el1_snoop_o_43_sv2v_reg,el1_snoop_o_42_sv2v_reg,
  el1_snoop_o_41_sv2v_reg,el1_snoop_o_40_sv2v_reg,el1_snoop_o_39_sv2v_reg,el1_snoop_o_38_sv2v_reg,
  el1_snoop_o_37_sv2v_reg,el1_snoop_o_36_sv2v_reg,el1_snoop_o_35_sv2v_reg,
  el1_snoop_o_34_sv2v_reg,el1_snoop_o_33_sv2v_reg,el1_snoop_o_32_sv2v_reg,
  el1_snoop_o_31_sv2v_reg,el1_snoop_o_30_sv2v_reg,el1_snoop_o_29_sv2v_reg,el1_snoop_o_28_sv2v_reg,
  el1_snoop_o_27_sv2v_reg,el1_snoop_o_26_sv2v_reg,el1_snoop_o_25_sv2v_reg,
  el1_snoop_o_24_sv2v_reg,el1_snoop_o_23_sv2v_reg,el1_snoop_o_22_sv2v_reg,
  el1_snoop_o_21_sv2v_reg,el1_snoop_o_20_sv2v_reg,el1_snoop_o_19_sv2v_reg,el1_snoop_o_18_sv2v_reg,
  el1_snoop_o_17_sv2v_reg,el1_snoop_o_16_sv2v_reg,el1_snoop_o_15_sv2v_reg,
  el1_snoop_o_14_sv2v_reg,el1_snoop_o_13_sv2v_reg,el1_snoop_o_12_sv2v_reg,
  el1_snoop_o_11_sv2v_reg,el1_snoop_o_10_sv2v_reg,el1_snoop_o_9_sv2v_reg,el1_snoop_o_8_sv2v_reg,
  el1_snoop_o_7_sv2v_reg,el1_snoop_o_6_sv2v_reg,el1_snoop_o_5_sv2v_reg,
  el1_snoop_o_4_sv2v_reg,el1_snoop_o_3_sv2v_reg,el1_snoop_o_2_sv2v_reg,el1_snoop_o_1_sv2v_reg,
  el1_snoop_o_0_sv2v_reg;
  assign num_els_r[1] = num_els_r_1_sv2v_reg;
  assign num_els_r[0] = num_els_r_0_sv2v_reg;
  assign el0_snoop_o[64] = el0_snoop_o_64_sv2v_reg;
  assign el0_snoop_o[63] = el0_snoop_o_63_sv2v_reg;
  assign el0_snoop_o[62] = el0_snoop_o_62_sv2v_reg;
  assign el0_snoop_o[61] = el0_snoop_o_61_sv2v_reg;
  assign el0_snoop_o[60] = el0_snoop_o_60_sv2v_reg;
  assign el0_snoop_o[59] = el0_snoop_o_59_sv2v_reg;
  assign el0_snoop_o[58] = el0_snoop_o_58_sv2v_reg;
  assign el0_snoop_o[57] = el0_snoop_o_57_sv2v_reg;
  assign el0_snoop_o[56] = el0_snoop_o_56_sv2v_reg;
  assign el0_snoop_o[55] = el0_snoop_o_55_sv2v_reg;
  assign el0_snoop_o[54] = el0_snoop_o_54_sv2v_reg;
  assign el0_snoop_o[53] = el0_snoop_o_53_sv2v_reg;
  assign el0_snoop_o[52] = el0_snoop_o_52_sv2v_reg;
  assign el0_snoop_o[51] = el0_snoop_o_51_sv2v_reg;
  assign el0_snoop_o[50] = el0_snoop_o_50_sv2v_reg;
  assign el0_snoop_o[49] = el0_snoop_o_49_sv2v_reg;
  assign el0_snoop_o[48] = el0_snoop_o_48_sv2v_reg;
  assign el0_snoop_o[47] = el0_snoop_o_47_sv2v_reg;
  assign el0_snoop_o[46] = el0_snoop_o_46_sv2v_reg;
  assign el0_snoop_o[45] = el0_snoop_o_45_sv2v_reg;
  assign el0_snoop_o[44] = el0_snoop_o_44_sv2v_reg;
  assign el0_snoop_o[43] = el0_snoop_o_43_sv2v_reg;
  assign el0_snoop_o[42] = el0_snoop_o_42_sv2v_reg;
  assign el0_snoop_o[41] = el0_snoop_o_41_sv2v_reg;
  assign el0_snoop_o[40] = el0_snoop_o_40_sv2v_reg;
  assign el0_snoop_o[39] = el0_snoop_o_39_sv2v_reg;
  assign el0_snoop_o[38] = el0_snoop_o_38_sv2v_reg;
  assign el0_snoop_o[37] = el0_snoop_o_37_sv2v_reg;
  assign el0_snoop_o[36] = el0_snoop_o_36_sv2v_reg;
  assign el0_snoop_o[35] = el0_snoop_o_35_sv2v_reg;
  assign el0_snoop_o[34] = el0_snoop_o_34_sv2v_reg;
  assign el0_snoop_o[33] = el0_snoop_o_33_sv2v_reg;
  assign el0_snoop_o[32] = el0_snoop_o_32_sv2v_reg;
  assign el0_snoop_o[31] = el0_snoop_o_31_sv2v_reg;
  assign el0_snoop_o[30] = el0_snoop_o_30_sv2v_reg;
  assign el0_snoop_o[29] = el0_snoop_o_29_sv2v_reg;
  assign el0_snoop_o[28] = el0_snoop_o_28_sv2v_reg;
  assign el0_snoop_o[27] = el0_snoop_o_27_sv2v_reg;
  assign el0_snoop_o[26] = el0_snoop_o_26_sv2v_reg;
  assign el0_snoop_o[25] = el0_snoop_o_25_sv2v_reg;
  assign el0_snoop_o[24] = el0_snoop_o_24_sv2v_reg;
  assign el0_snoop_o[23] = el0_snoop_o_23_sv2v_reg;
  assign el0_snoop_o[22] = el0_snoop_o_22_sv2v_reg;
  assign el0_snoop_o[21] = el0_snoop_o_21_sv2v_reg;
  assign el0_snoop_o[20] = el0_snoop_o_20_sv2v_reg;
  assign el0_snoop_o[19] = el0_snoop_o_19_sv2v_reg;
  assign el0_snoop_o[18] = el0_snoop_o_18_sv2v_reg;
  assign el0_snoop_o[17] = el0_snoop_o_17_sv2v_reg;
  assign el0_snoop_o[16] = el0_snoop_o_16_sv2v_reg;
  assign el0_snoop_o[15] = el0_snoop_o_15_sv2v_reg;
  assign el0_snoop_o[14] = el0_snoop_o_14_sv2v_reg;
  assign el0_snoop_o[13] = el0_snoop_o_13_sv2v_reg;
  assign el0_snoop_o[12] = el0_snoop_o_12_sv2v_reg;
  assign el0_snoop_o[11] = el0_snoop_o_11_sv2v_reg;
  assign el0_snoop_o[10] = el0_snoop_o_10_sv2v_reg;
  assign el0_snoop_o[9] = el0_snoop_o_9_sv2v_reg;
  assign el0_snoop_o[8] = el0_snoop_o_8_sv2v_reg;
  assign el0_snoop_o[7] = el0_snoop_o_7_sv2v_reg;
  assign el0_snoop_o[6] = el0_snoop_o_6_sv2v_reg;
  assign el0_snoop_o[5] = el0_snoop_o_5_sv2v_reg;
  assign el0_snoop_o[4] = el0_snoop_o_4_sv2v_reg;
  assign el0_snoop_o[3] = el0_snoop_o_3_sv2v_reg;
  assign el0_snoop_o[2] = el0_snoop_o_2_sv2v_reg;
  assign el0_snoop_o[1] = el0_snoop_o_1_sv2v_reg;
  assign el0_snoop_o[0] = el0_snoop_o_0_sv2v_reg;
  assign el1_snoop_o[64] = el1_snoop_o_64_sv2v_reg;
  assign el1_snoop_o[63] = el1_snoop_o_63_sv2v_reg;
  assign el1_snoop_o[62] = el1_snoop_o_62_sv2v_reg;
  assign el1_snoop_o[61] = el1_snoop_o_61_sv2v_reg;
  assign el1_snoop_o[60] = el1_snoop_o_60_sv2v_reg;
  assign el1_snoop_o[59] = el1_snoop_o_59_sv2v_reg;
  assign el1_snoop_o[58] = el1_snoop_o_58_sv2v_reg;
  assign el1_snoop_o[57] = el1_snoop_o_57_sv2v_reg;
  assign el1_snoop_o[56] = el1_snoop_o_56_sv2v_reg;
  assign el1_snoop_o[55] = el1_snoop_o_55_sv2v_reg;
  assign el1_snoop_o[54] = el1_snoop_o_54_sv2v_reg;
  assign el1_snoop_o[53] = el1_snoop_o_53_sv2v_reg;
  assign el1_snoop_o[52] = el1_snoop_o_52_sv2v_reg;
  assign el1_snoop_o[51] = el1_snoop_o_51_sv2v_reg;
  assign el1_snoop_o[50] = el1_snoop_o_50_sv2v_reg;
  assign el1_snoop_o[49] = el1_snoop_o_49_sv2v_reg;
  assign el1_snoop_o[48] = el1_snoop_o_48_sv2v_reg;
  assign el1_snoop_o[47] = el1_snoop_o_47_sv2v_reg;
  assign el1_snoop_o[46] = el1_snoop_o_46_sv2v_reg;
  assign el1_snoop_o[45] = el1_snoop_o_45_sv2v_reg;
  assign el1_snoop_o[44] = el1_snoop_o_44_sv2v_reg;
  assign el1_snoop_o[43] = el1_snoop_o_43_sv2v_reg;
  assign el1_snoop_o[42] = el1_snoop_o_42_sv2v_reg;
  assign el1_snoop_o[41] = el1_snoop_o_41_sv2v_reg;
  assign el1_snoop_o[40] = el1_snoop_o_40_sv2v_reg;
  assign el1_snoop_o[39] = el1_snoop_o_39_sv2v_reg;
  assign el1_snoop_o[38] = el1_snoop_o_38_sv2v_reg;
  assign el1_snoop_o[37] = el1_snoop_o_37_sv2v_reg;
  assign el1_snoop_o[36] = el1_snoop_o_36_sv2v_reg;
  assign el1_snoop_o[35] = el1_snoop_o_35_sv2v_reg;
  assign el1_snoop_o[34] = el1_snoop_o_34_sv2v_reg;
  assign el1_snoop_o[33] = el1_snoop_o_33_sv2v_reg;
  assign el1_snoop_o[32] = el1_snoop_o_32_sv2v_reg;
  assign el1_snoop_o[31] = el1_snoop_o_31_sv2v_reg;
  assign el1_snoop_o[30] = el1_snoop_o_30_sv2v_reg;
  assign el1_snoop_o[29] = el1_snoop_o_29_sv2v_reg;
  assign el1_snoop_o[28] = el1_snoop_o_28_sv2v_reg;
  assign el1_snoop_o[27] = el1_snoop_o_27_sv2v_reg;
  assign el1_snoop_o[26] = el1_snoop_o_26_sv2v_reg;
  assign el1_snoop_o[25] = el1_snoop_o_25_sv2v_reg;
  assign el1_snoop_o[24] = el1_snoop_o_24_sv2v_reg;
  assign el1_snoop_o[23] = el1_snoop_o_23_sv2v_reg;
  assign el1_snoop_o[22] = el1_snoop_o_22_sv2v_reg;
  assign el1_snoop_o[21] = el1_snoop_o_21_sv2v_reg;
  assign el1_snoop_o[20] = el1_snoop_o_20_sv2v_reg;
  assign el1_snoop_o[19] = el1_snoop_o_19_sv2v_reg;
  assign el1_snoop_o[18] = el1_snoop_o_18_sv2v_reg;
  assign el1_snoop_o[17] = el1_snoop_o_17_sv2v_reg;
  assign el1_snoop_o[16] = el1_snoop_o_16_sv2v_reg;
  assign el1_snoop_o[15] = el1_snoop_o_15_sv2v_reg;
  assign el1_snoop_o[14] = el1_snoop_o_14_sv2v_reg;
  assign el1_snoop_o[13] = el1_snoop_o_13_sv2v_reg;
  assign el1_snoop_o[12] = el1_snoop_o_12_sv2v_reg;
  assign el1_snoop_o[11] = el1_snoop_o_11_sv2v_reg;
  assign el1_snoop_o[10] = el1_snoop_o_10_sv2v_reg;
  assign el1_snoop_o[9] = el1_snoop_o_9_sv2v_reg;
  assign el1_snoop_o[8] = el1_snoop_o_8_sv2v_reg;
  assign el1_snoop_o[7] = el1_snoop_o_7_sv2v_reg;
  assign el1_snoop_o[6] = el1_snoop_o_6_sv2v_reg;
  assign el1_snoop_o[5] = el1_snoop_o_5_sv2v_reg;
  assign el1_snoop_o[4] = el1_snoop_o_4_sv2v_reg;
  assign el1_snoop_o[3] = el1_snoop_o_3_sv2v_reg;
  assign el1_snoop_o[2] = el1_snoop_o_2_sv2v_reg;
  assign el1_snoop_o[1] = el1_snoop_o_1_sv2v_reg;
  assign el1_snoop_o[0] = el1_snoop_o_0_sv2v_reg;
  assign N10 = N8 & N9;
  assign N11 = num_els_r[1] | N9;
  assign N13 = N8 | num_els_r[0];
  assign N15 = num_els_r[1] & num_els_r[0];
  assign { N20, N19 } = num_els_r + v_i;
  assign { N23, N22 } = { N20, N19 } - N21;
  assign v_o = (N0)? v_i : 
               (N1)? 1'b1 : 
               (N2)? 1'b1 : 
               (N3)? 1'b0 : 1'b0;
  assign N0 = N10;
  assign N1 = N12;
  assign N2 = N14;
  assign N3 = N15;
  assign empty_o = (N0)? 1'b1 : 
                   (N1)? 1'b0 : 
                   (N2)? 1'b0 : 
                   (N3)? 1'b0 : 1'b0;
  assign full_o = (N0)? 1'b0 : 
                  (N1)? 1'b0 : 
                  (N2)? 1'b1 : 
                  (N3)? 1'b0 : 1'b0;
  assign el0_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b0 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el1_valid_o = (N0)? 1'b0 : 
                       (N1)? 1'b1 : 
                       (N2)? 1'b1 : 
                       (N3)? 1'b0 : 1'b0;
  assign el0_enable = (N0)? 1'b0 : 
                      (N1)? N16 : 
                      (N2)? N17 : 
                      (N3)? 1'b0 : 1'b0;
  assign el1_enable = (N0)? N16 : 
                      (N1)? N17 : 
                      (N2)? yumi_i : 
                      (N3)? 1'b0 : 1'b0;
  assign mux0_sel = (N0)? 1'b0 : 
                    (N1)? 1'b0 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign mux1_sel = (N0)? 1'b0 : 
                    (N1)? 1'b1 : 
                    (N2)? 1'b1 : 
                    (N3)? 1'b0 : 1'b0;
  assign { N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25 } = (N4)? el0_snoop_o : 
                                                                                                                                                                                                                                                                                                                                                   (N5)? data_i : 1'b0;
  assign N4 = mux0_sel;
  assign N5 = N24;
  assign data_o = (N6)? el1_snoop_o : 
                  (N7)? data_i : 1'b0;
  assign N6 = mux1_sel;
  assign N7 = N90;
  assign N8 = ~num_els_r[1];
  assign N9 = ~num_els_r[0];
  assign N12 = ~N11;
  assign N14 = ~N13;
  assign N16 = v_i & N91;
  assign N91 = ~yumi_i;
  assign N17 = v_i & yumi_i;
  assign N18 = ~reset_i;
  assign N21 = v_o & yumi_i;
  assign N24 = ~mux0_sel;
  assign N90 = ~mux1_sel;

  always @(posedge clk_i) begin
    if(reset_i) begin
      num_els_r_1_sv2v_reg <= 1'b0;
      num_els_r_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      num_els_r_1_sv2v_reg <= N23;
      num_els_r_0_sv2v_reg <= N22;
    end 
    if(el0_enable) begin
      el0_snoop_o_64_sv2v_reg <= data_i[64];
      el0_snoop_o_63_sv2v_reg <= data_i[63];
      el0_snoop_o_62_sv2v_reg <= data_i[62];
      el0_snoop_o_61_sv2v_reg <= data_i[61];
      el0_snoop_o_60_sv2v_reg <= data_i[60];
      el0_snoop_o_59_sv2v_reg <= data_i[59];
      el0_snoop_o_58_sv2v_reg <= data_i[58];
      el0_snoop_o_57_sv2v_reg <= data_i[57];
      el0_snoop_o_56_sv2v_reg <= data_i[56];
      el0_snoop_o_55_sv2v_reg <= data_i[55];
      el0_snoop_o_54_sv2v_reg <= data_i[54];
      el0_snoop_o_53_sv2v_reg <= data_i[53];
      el0_snoop_o_52_sv2v_reg <= data_i[52];
      el0_snoop_o_51_sv2v_reg <= data_i[51];
      el0_snoop_o_50_sv2v_reg <= data_i[50];
      el0_snoop_o_49_sv2v_reg <= data_i[49];
      el0_snoop_o_48_sv2v_reg <= data_i[48];
      el0_snoop_o_47_sv2v_reg <= data_i[47];
      el0_snoop_o_46_sv2v_reg <= data_i[46];
      el0_snoop_o_45_sv2v_reg <= data_i[45];
      el0_snoop_o_44_sv2v_reg <= data_i[44];
      el0_snoop_o_43_sv2v_reg <= data_i[43];
      el0_snoop_o_42_sv2v_reg <= data_i[42];
      el0_snoop_o_41_sv2v_reg <= data_i[41];
      el0_snoop_o_40_sv2v_reg <= data_i[40];
      el0_snoop_o_39_sv2v_reg <= data_i[39];
      el0_snoop_o_38_sv2v_reg <= data_i[38];
      el0_snoop_o_37_sv2v_reg <= data_i[37];
      el0_snoop_o_36_sv2v_reg <= data_i[36];
      el0_snoop_o_35_sv2v_reg <= data_i[35];
      el0_snoop_o_34_sv2v_reg <= data_i[34];
      el0_snoop_o_33_sv2v_reg <= data_i[33];
      el0_snoop_o_32_sv2v_reg <= data_i[32];
      el0_snoop_o_31_sv2v_reg <= data_i[31];
      el0_snoop_o_30_sv2v_reg <= data_i[30];
      el0_snoop_o_29_sv2v_reg <= data_i[29];
      el0_snoop_o_28_sv2v_reg <= data_i[28];
      el0_snoop_o_27_sv2v_reg <= data_i[27];
      el0_snoop_o_26_sv2v_reg <= data_i[26];
      el0_snoop_o_25_sv2v_reg <= data_i[25];
      el0_snoop_o_24_sv2v_reg <= data_i[24];
      el0_snoop_o_23_sv2v_reg <= data_i[23];
      el0_snoop_o_22_sv2v_reg <= data_i[22];
      el0_snoop_o_21_sv2v_reg <= data_i[21];
      el0_snoop_o_20_sv2v_reg <= data_i[20];
      el0_snoop_o_19_sv2v_reg <= data_i[19];
      el0_snoop_o_18_sv2v_reg <= data_i[18];
      el0_snoop_o_17_sv2v_reg <= data_i[17];
      el0_snoop_o_16_sv2v_reg <= data_i[16];
      el0_snoop_o_15_sv2v_reg <= data_i[15];
      el0_snoop_o_14_sv2v_reg <= data_i[14];
      el0_snoop_o_13_sv2v_reg <= data_i[13];
      el0_snoop_o_12_sv2v_reg <= data_i[12];
      el0_snoop_o_11_sv2v_reg <= data_i[11];
      el0_snoop_o_10_sv2v_reg <= data_i[10];
      el0_snoop_o_9_sv2v_reg <= data_i[9];
      el0_snoop_o_8_sv2v_reg <= data_i[8];
      el0_snoop_o_7_sv2v_reg <= data_i[7];
      el0_snoop_o_6_sv2v_reg <= data_i[6];
      el0_snoop_o_5_sv2v_reg <= data_i[5];
      el0_snoop_o_4_sv2v_reg <= data_i[4];
      el0_snoop_o_3_sv2v_reg <= data_i[3];
      el0_snoop_o_2_sv2v_reg <= data_i[2];
      el0_snoop_o_1_sv2v_reg <= data_i[1];
      el0_snoop_o_0_sv2v_reg <= data_i[0];
    end 
    if(el1_enable) begin
      el1_snoop_o_64_sv2v_reg <= N89;
      el1_snoop_o_63_sv2v_reg <= N88;
      el1_snoop_o_62_sv2v_reg <= N87;
      el1_snoop_o_61_sv2v_reg <= N86;
      el1_snoop_o_60_sv2v_reg <= N85;
      el1_snoop_o_59_sv2v_reg <= N84;
      el1_snoop_o_58_sv2v_reg <= N83;
      el1_snoop_o_57_sv2v_reg <= N82;
      el1_snoop_o_56_sv2v_reg <= N81;
      el1_snoop_o_55_sv2v_reg <= N80;
      el1_snoop_o_54_sv2v_reg <= N79;
      el1_snoop_o_53_sv2v_reg <= N78;
      el1_snoop_o_52_sv2v_reg <= N77;
      el1_snoop_o_51_sv2v_reg <= N76;
      el1_snoop_o_50_sv2v_reg <= N75;
      el1_snoop_o_49_sv2v_reg <= N74;
      el1_snoop_o_48_sv2v_reg <= N73;
      el1_snoop_o_47_sv2v_reg <= N72;
      el1_snoop_o_46_sv2v_reg <= N71;
      el1_snoop_o_45_sv2v_reg <= N70;
      el1_snoop_o_44_sv2v_reg <= N69;
      el1_snoop_o_43_sv2v_reg <= N68;
      el1_snoop_o_42_sv2v_reg <= N67;
      el1_snoop_o_41_sv2v_reg <= N66;
      el1_snoop_o_40_sv2v_reg <= N65;
      el1_snoop_o_39_sv2v_reg <= N64;
      el1_snoop_o_38_sv2v_reg <= N63;
      el1_snoop_o_37_sv2v_reg <= N62;
      el1_snoop_o_36_sv2v_reg <= N61;
      el1_snoop_o_35_sv2v_reg <= N60;
      el1_snoop_o_34_sv2v_reg <= N59;
      el1_snoop_o_33_sv2v_reg <= N58;
      el1_snoop_o_32_sv2v_reg <= N57;
      el1_snoop_o_31_sv2v_reg <= N56;
      el1_snoop_o_30_sv2v_reg <= N55;
      el1_snoop_o_29_sv2v_reg <= N54;
      el1_snoop_o_28_sv2v_reg <= N53;
      el1_snoop_o_27_sv2v_reg <= N52;
      el1_snoop_o_26_sv2v_reg <= N51;
      el1_snoop_o_25_sv2v_reg <= N50;
      el1_snoop_o_24_sv2v_reg <= N49;
      el1_snoop_o_23_sv2v_reg <= N48;
      el1_snoop_o_22_sv2v_reg <= N47;
      el1_snoop_o_21_sv2v_reg <= N46;
      el1_snoop_o_20_sv2v_reg <= N45;
      el1_snoop_o_19_sv2v_reg <= N44;
      el1_snoop_o_18_sv2v_reg <= N43;
      el1_snoop_o_17_sv2v_reg <= N42;
      el1_snoop_o_16_sv2v_reg <= N41;
      el1_snoop_o_15_sv2v_reg <= N40;
      el1_snoop_o_14_sv2v_reg <= N39;
      el1_snoop_o_13_sv2v_reg <= N38;
      el1_snoop_o_12_sv2v_reg <= N37;
      el1_snoop_o_11_sv2v_reg <= N36;
      el1_snoop_o_10_sv2v_reg <= N35;
      el1_snoop_o_9_sv2v_reg <= N34;
      el1_snoop_o_8_sv2v_reg <= N33;
      el1_snoop_o_7_sv2v_reg <= N32;
      el1_snoop_o_6_sv2v_reg <= N31;
      el1_snoop_o_5_sv2v_reg <= N30;
      el1_snoop_o_4_sv2v_reg <= N29;
      el1_snoop_o_3_sv2v_reg <= N28;
      el1_snoop_o_2_sv2v_reg <= N27;
      el1_snoop_o_1_sv2v_reg <= N26;
      el1_snoop_o_0_sv2v_reg <= N25;
    end 
  end


endmodule



module bsg_mux_segmented_segments_p4_segment_width_p8
(
  data0_i,
  data1_i,
  sel_i,
  data_o
);

  input [31:0] data0_i;
  input [31:0] data1_i;
  input [3:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7;
  assign data_o[7:0] = (N0)? data1_i[7:0] : 
                       (N4)? data0_i[7:0] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[15:8] = (N1)? data1_i[15:8] : 
                        (N5)? data0_i[15:8] : 1'b0;
  assign N1 = sel_i[1];
  assign data_o[23:16] = (N2)? data1_i[23:16] : 
                         (N6)? data0_i[23:16] : 1'b0;
  assign N2 = sel_i[2];
  assign data_o[31:24] = (N3)? data1_i[31:24] : 
                         (N7)? data0_i[31:24] : 1'b0;
  assign N3 = sel_i[3];
  assign N4 = ~sel_i[0];
  assign N5 = ~sel_i[1];
  assign N6 = ~sel_i[2];
  assign N7 = ~sel_i[3];

endmodule



module bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p2
(
  clk_i,
  reset_i,
  sbuf_entry_i,
  v_i,
  sbuf_entry_o,
  v_o,
  yumi_i,
  empty_o,
  full_o,
  bypass_addr_i,
  bypass_v_i,
  bypass_data_o,
  bypass_mask_o
);

  input [64:0] sbuf_entry_i;
  output [64:0] sbuf_entry_o;
  input [27:0] bypass_addr_i;
  output [31:0] bypass_data_o;
  output [3:0] bypass_mask_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input bypass_v_i;
  output v_o;
  output empty_o;
  output full_o;
  wire [64:0] sbuf_entry_o,el0,el1;
  wire [31:0] bypass_data_o,el0or1_data,bypass_data_n;
  wire [3:0] bypass_mask_o,bypass_mask_n;
  wire v_o,empty_o,full_o,N0,el0_valid,el1_valid,tag_hit0_n,tag_hit1_n,tag_hit2_n,
  _2_net__3_,_2_net__2_,_2_net__1_,_2_net__0_,_4_net__3_,_4_net__2_,_4_net__1_,
  _4_net__0_,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  wire [3:3] tag_hit0x4,tag_hit1x4,tag_hit2x4;
  reg bypass_data_o_31_sv2v_reg,bypass_data_o_30_sv2v_reg,bypass_data_o_29_sv2v_reg,
  bypass_data_o_28_sv2v_reg,bypass_data_o_27_sv2v_reg,bypass_data_o_26_sv2v_reg,
  bypass_data_o_25_sv2v_reg,bypass_data_o_24_sv2v_reg,bypass_data_o_23_sv2v_reg,
  bypass_data_o_22_sv2v_reg,bypass_data_o_21_sv2v_reg,bypass_data_o_20_sv2v_reg,
  bypass_data_o_19_sv2v_reg,bypass_data_o_18_sv2v_reg,bypass_data_o_17_sv2v_reg,
  bypass_data_o_16_sv2v_reg,bypass_data_o_15_sv2v_reg,bypass_data_o_14_sv2v_reg,
  bypass_data_o_13_sv2v_reg,bypass_data_o_12_sv2v_reg,bypass_data_o_11_sv2v_reg,
  bypass_data_o_10_sv2v_reg,bypass_data_o_9_sv2v_reg,bypass_data_o_8_sv2v_reg,
  bypass_data_o_7_sv2v_reg,bypass_data_o_6_sv2v_reg,bypass_data_o_5_sv2v_reg,
  bypass_data_o_4_sv2v_reg,bypass_data_o_3_sv2v_reg,bypass_data_o_2_sv2v_reg,bypass_data_o_1_sv2v_reg,
  bypass_data_o_0_sv2v_reg,bypass_mask_o_3_sv2v_reg,bypass_mask_o_2_sv2v_reg,
  bypass_mask_o_1_sv2v_reg,bypass_mask_o_0_sv2v_reg;
  assign bypass_data_o[31] = bypass_data_o_31_sv2v_reg;
  assign bypass_data_o[30] = bypass_data_o_30_sv2v_reg;
  assign bypass_data_o[29] = bypass_data_o_29_sv2v_reg;
  assign bypass_data_o[28] = bypass_data_o_28_sv2v_reg;
  assign bypass_data_o[27] = bypass_data_o_27_sv2v_reg;
  assign bypass_data_o[26] = bypass_data_o_26_sv2v_reg;
  assign bypass_data_o[25] = bypass_data_o_25_sv2v_reg;
  assign bypass_data_o[24] = bypass_data_o_24_sv2v_reg;
  assign bypass_data_o[23] = bypass_data_o_23_sv2v_reg;
  assign bypass_data_o[22] = bypass_data_o_22_sv2v_reg;
  assign bypass_data_o[21] = bypass_data_o_21_sv2v_reg;
  assign bypass_data_o[20] = bypass_data_o_20_sv2v_reg;
  assign bypass_data_o[19] = bypass_data_o_19_sv2v_reg;
  assign bypass_data_o[18] = bypass_data_o_18_sv2v_reg;
  assign bypass_data_o[17] = bypass_data_o_17_sv2v_reg;
  assign bypass_data_o[16] = bypass_data_o_16_sv2v_reg;
  assign bypass_data_o[15] = bypass_data_o_15_sv2v_reg;
  assign bypass_data_o[14] = bypass_data_o_14_sv2v_reg;
  assign bypass_data_o[13] = bypass_data_o_13_sv2v_reg;
  assign bypass_data_o[12] = bypass_data_o_12_sv2v_reg;
  assign bypass_data_o[11] = bypass_data_o_11_sv2v_reg;
  assign bypass_data_o[10] = bypass_data_o_10_sv2v_reg;
  assign bypass_data_o[9] = bypass_data_o_9_sv2v_reg;
  assign bypass_data_o[8] = bypass_data_o_8_sv2v_reg;
  assign bypass_data_o[7] = bypass_data_o_7_sv2v_reg;
  assign bypass_data_o[6] = bypass_data_o_6_sv2v_reg;
  assign bypass_data_o[5] = bypass_data_o_5_sv2v_reg;
  assign bypass_data_o[4] = bypass_data_o_4_sv2v_reg;
  assign bypass_data_o[3] = bypass_data_o_3_sv2v_reg;
  assign bypass_data_o[2] = bypass_data_o_2_sv2v_reg;
  assign bypass_data_o[1] = bypass_data_o_1_sv2v_reg;
  assign bypass_data_o[0] = bypass_data_o_0_sv2v_reg;
  assign bypass_mask_o[3] = bypass_mask_o_3_sv2v_reg;
  assign bypass_mask_o[2] = bypass_mask_o_2_sv2v_reg;
  assign bypass_mask_o[1] = bypass_mask_o_1_sv2v_reg;
  assign bypass_mask_o[0] = bypass_mask_o_0_sv2v_reg;

  bsg_cache_buffer_queue_width_p65
  q0
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .data_i(sbuf_entry_i),
    .v_o(v_o),
    .data_o(sbuf_entry_o),
    .yumi_i(yumi_i),
    .el0_valid_o(el0_valid),
    .el1_valid_o(el1_valid),
    .el0_snoop_o(el0),
    .el1_snoop_o(el1),
    .empty_o(empty_o),
    .full_o(full_o)
  );

  assign tag_hit0_n = bypass_addr_i[27:2] == el0[64:39];
  assign tag_hit1_n = bypass_addr_i[27:2] == el1[64:39];
  assign tag_hit2_n = bypass_addr_i[27:2] == sbuf_entry_i[64:39];

  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge0
  (
    .data0_i(el1[36:5]),
    .data1_i(el0[36:5]),
    .sel_i({ _2_net__3_, _2_net__2_, _2_net__1_, _2_net__0_ }),
    .data_o(el0or1_data)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  mux_segmented_merge1
  (
    .data0_i(el0or1_data),
    .data1_i(sbuf_entry_i[36:5]),
    .sel_i({ _4_net__3_, _4_net__2_, _4_net__1_, _4_net__0_ }),
    .data_o(bypass_data_n)
  );

  assign N2 = (N0)? 1'b1 : 
              (N1)? 1'b0 : 1'b0;
  assign N0 = bypass_v_i;
  assign tag_hit0x4[3] = tag_hit0_n & el0_valid;
  assign tag_hit1x4[3] = tag_hit1_n & el1_valid;
  assign tag_hit2x4[3] = tag_hit2_n & v_i;
  assign bypass_mask_n[3] = N5 | N6;
  assign N5 = N3 | N4;
  assign N3 = tag_hit0x4[3] & el0[4];
  assign N4 = tag_hit1x4[3] & el1[4];
  assign N6 = tag_hit2x4[3] & sbuf_entry_i[4];
  assign bypass_mask_n[2] = N9 | N10;
  assign N9 = N7 | N8;
  assign N7 = tag_hit0x4[3] & el0[3];
  assign N8 = tag_hit1x4[3] & el1[3];
  assign N10 = tag_hit2x4[3] & sbuf_entry_i[3];
  assign bypass_mask_n[1] = N13 | N14;
  assign N13 = N11 | N12;
  assign N11 = tag_hit0x4[3] & el0[2];
  assign N12 = tag_hit1x4[3] & el1[2];
  assign N14 = tag_hit2x4[3] & sbuf_entry_i[2];
  assign bypass_mask_n[0] = N17 | N18;
  assign N17 = N15 | N16;
  assign N15 = tag_hit0x4[3] & el0[1];
  assign N16 = tag_hit1x4[3] & el1[1];
  assign N18 = tag_hit2x4[3] & sbuf_entry_i[1];
  assign _2_net__3_ = tag_hit0x4[3] & el0[4];
  assign _2_net__2_ = tag_hit0x4[3] & el0[3];
  assign _2_net__1_ = tag_hit0x4[3] & el0[2];
  assign _2_net__0_ = tag_hit0x4[3] & el0[1];
  assign _4_net__3_ = tag_hit2x4[3] & sbuf_entry_i[4];
  assign _4_net__2_ = tag_hit2x4[3] & sbuf_entry_i[3];
  assign _4_net__1_ = tag_hit2x4[3] & sbuf_entry_i[2];
  assign _4_net__0_ = tag_hit2x4[3] & sbuf_entry_i[1];
  assign N1 = ~bypass_v_i;

  always @(posedge clk_i) begin
    if(reset_i) begin
      bypass_data_o_31_sv2v_reg <= 1'b0;
      bypass_data_o_30_sv2v_reg <= 1'b0;
      bypass_data_o_29_sv2v_reg <= 1'b0;
      bypass_data_o_28_sv2v_reg <= 1'b0;
      bypass_data_o_27_sv2v_reg <= 1'b0;
      bypass_data_o_26_sv2v_reg <= 1'b0;
      bypass_data_o_25_sv2v_reg <= 1'b0;
      bypass_data_o_24_sv2v_reg <= 1'b0;
      bypass_data_o_23_sv2v_reg <= 1'b0;
      bypass_data_o_22_sv2v_reg <= 1'b0;
      bypass_data_o_21_sv2v_reg <= 1'b0;
      bypass_data_o_20_sv2v_reg <= 1'b0;
      bypass_data_o_19_sv2v_reg <= 1'b0;
      bypass_data_o_18_sv2v_reg <= 1'b0;
      bypass_data_o_17_sv2v_reg <= 1'b0;
      bypass_data_o_16_sv2v_reg <= 1'b0;
      bypass_data_o_15_sv2v_reg <= 1'b0;
      bypass_data_o_14_sv2v_reg <= 1'b0;
      bypass_data_o_13_sv2v_reg <= 1'b0;
      bypass_data_o_12_sv2v_reg <= 1'b0;
      bypass_data_o_11_sv2v_reg <= 1'b0;
      bypass_data_o_10_sv2v_reg <= 1'b0;
      bypass_data_o_9_sv2v_reg <= 1'b0;
      bypass_data_o_8_sv2v_reg <= 1'b0;
      bypass_data_o_7_sv2v_reg <= 1'b0;
      bypass_data_o_6_sv2v_reg <= 1'b0;
      bypass_data_o_5_sv2v_reg <= 1'b0;
      bypass_data_o_4_sv2v_reg <= 1'b0;
      bypass_data_o_3_sv2v_reg <= 1'b0;
      bypass_data_o_2_sv2v_reg <= 1'b0;
      bypass_data_o_1_sv2v_reg <= 1'b0;
      bypass_data_o_0_sv2v_reg <= 1'b0;
      bypass_mask_o_3_sv2v_reg <= 1'b0;
      bypass_mask_o_2_sv2v_reg <= 1'b0;
      bypass_mask_o_1_sv2v_reg <= 1'b0;
      bypass_mask_o_0_sv2v_reg <= 1'b0;
    end else if(N2) begin
      bypass_data_o_31_sv2v_reg <= bypass_data_n[31];
      bypass_data_o_30_sv2v_reg <= bypass_data_n[30];
      bypass_data_o_29_sv2v_reg <= bypass_data_n[29];
      bypass_data_o_28_sv2v_reg <= bypass_data_n[28];
      bypass_data_o_27_sv2v_reg <= bypass_data_n[27];
      bypass_data_o_26_sv2v_reg <= bypass_data_n[26];
      bypass_data_o_25_sv2v_reg <= bypass_data_n[25];
      bypass_data_o_24_sv2v_reg <= bypass_data_n[24];
      bypass_data_o_23_sv2v_reg <= bypass_data_n[23];
      bypass_data_o_22_sv2v_reg <= bypass_data_n[22];
      bypass_data_o_21_sv2v_reg <= bypass_data_n[21];
      bypass_data_o_20_sv2v_reg <= bypass_data_n[20];
      bypass_data_o_19_sv2v_reg <= bypass_data_n[19];
      bypass_data_o_18_sv2v_reg <= bypass_data_n[18];
      bypass_data_o_17_sv2v_reg <= bypass_data_n[17];
      bypass_data_o_16_sv2v_reg <= bypass_data_n[16];
      bypass_data_o_15_sv2v_reg <= bypass_data_n[15];
      bypass_data_o_14_sv2v_reg <= bypass_data_n[14];
      bypass_data_o_13_sv2v_reg <= bypass_data_n[13];
      bypass_data_o_12_sv2v_reg <= bypass_data_n[12];
      bypass_data_o_11_sv2v_reg <= bypass_data_n[11];
      bypass_data_o_10_sv2v_reg <= bypass_data_n[10];
      bypass_data_o_9_sv2v_reg <= bypass_data_n[9];
      bypass_data_o_8_sv2v_reg <= bypass_data_n[8];
      bypass_data_o_7_sv2v_reg <= bypass_data_n[7];
      bypass_data_o_6_sv2v_reg <= bypass_data_n[6];
      bypass_data_o_5_sv2v_reg <= bypass_data_n[5];
      bypass_data_o_4_sv2v_reg <= bypass_data_n[4];
      bypass_data_o_3_sv2v_reg <= bypass_data_n[3];
      bypass_data_o_2_sv2v_reg <= bypass_data_n[2];
      bypass_data_o_1_sv2v_reg <= bypass_data_n[1];
      bypass_data_o_0_sv2v_reg <= bypass_data_n[0];
      bypass_mask_o_3_sv2v_reg <= bypass_mask_n[3];
      bypass_mask_o_2_sv2v_reg <= bypass_mask_n[2];
      bypass_mask_o_1_sv2v_reg <= bypass_mask_n[1];
      bypass_mask_o_0_sv2v_reg <= bypass_mask_n[0];
    end 
  end


endmodule



module bsg_decode_num_out_p1
(
  i,
  o
);

  input [0:0] i;
  output [0:0] o;
  wire [0:0] o;
  assign o[0] = 1'b1;

endmodule



module bsg_mux_width_p32_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [95:0] data_i;
  input [1:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[31] = (N2)? data_i[31] : 
                      (N3)? data_i[63] : 
                      (N4)? data_i[95] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[30] = (N2)? data_i[30] : 
                      (N3)? data_i[62] : 
                      (N4)? data_i[94] : 1'b0;
  assign data_o[29] = (N2)? data_i[29] : 
                      (N3)? data_i[61] : 
                      (N4)? data_i[93] : 1'b0;
  assign data_o[28] = (N2)? data_i[28] : 
                      (N3)? data_i[60] : 
                      (N4)? data_i[92] : 1'b0;
  assign data_o[27] = (N2)? data_i[27] : 
                      (N3)? data_i[59] : 
                      (N4)? data_i[91] : 1'b0;
  assign data_o[26] = (N2)? data_i[26] : 
                      (N3)? data_i[58] : 
                      (N4)? data_i[90] : 1'b0;
  assign data_o[25] = (N2)? data_i[25] : 
                      (N3)? data_i[57] : 
                      (N4)? data_i[89] : 1'b0;
  assign data_o[24] = (N2)? data_i[24] : 
                      (N3)? data_i[56] : 
                      (N4)? data_i[88] : 1'b0;
  assign data_o[23] = (N2)? data_i[23] : 
                      (N3)? data_i[55] : 
                      (N4)? data_i[87] : 1'b0;
  assign data_o[22] = (N2)? data_i[22] : 
                      (N3)? data_i[54] : 
                      (N4)? data_i[86] : 1'b0;
  assign data_o[21] = (N2)? data_i[21] : 
                      (N3)? data_i[53] : 
                      (N4)? data_i[85] : 1'b0;
  assign data_o[20] = (N2)? data_i[20] : 
                      (N3)? data_i[52] : 
                      (N4)? data_i[84] : 1'b0;
  assign data_o[19] = (N2)? data_i[19] : 
                      (N3)? data_i[51] : 
                      (N4)? data_i[83] : 1'b0;
  assign data_o[18] = (N2)? data_i[18] : 
                      (N3)? data_i[50] : 
                      (N4)? data_i[82] : 1'b0;
  assign data_o[17] = (N2)? data_i[17] : 
                      (N3)? data_i[49] : 
                      (N4)? data_i[81] : 1'b0;
  assign data_o[16] = (N2)? data_i[16] : 
                      (N3)? data_i[48] : 
                      (N4)? data_i[80] : 1'b0;
  assign data_o[15] = (N2)? data_i[15] : 
                      (N3)? data_i[47] : 
                      (N4)? data_i[79] : 1'b0;
  assign data_o[14] = (N2)? data_i[14] : 
                      (N3)? data_i[46] : 
                      (N4)? data_i[78] : 1'b0;
  assign data_o[13] = (N2)? data_i[13] : 
                      (N3)? data_i[45] : 
                      (N4)? data_i[77] : 1'b0;
  assign data_o[12] = (N2)? data_i[12] : 
                      (N3)? data_i[44] : 
                      (N4)? data_i[76] : 1'b0;
  assign data_o[11] = (N2)? data_i[11] : 
                      (N3)? data_i[43] : 
                      (N4)? data_i[75] : 1'b0;
  assign data_o[10] = (N2)? data_i[10] : 
                      (N3)? data_i[42] : 
                      (N4)? data_i[74] : 1'b0;
  assign data_o[9] = (N2)? data_i[9] : 
                     (N3)? data_i[41] : 
                     (N4)? data_i[73] : 1'b0;
  assign data_o[8] = (N2)? data_i[8] : 
                     (N3)? data_i[40] : 
                     (N4)? data_i[72] : 1'b0;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N3)? data_i[39] : 
                     (N4)? data_i[71] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N3)? data_i[38] : 
                     (N4)? data_i[70] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N3)? data_i[37] : 
                     (N4)? data_i[69] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N3)? data_i[36] : 
                     (N4)? data_i[68] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[35] : 
                     (N4)? data_i[67] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[34] : 
                     (N4)? data_i[66] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[33] : 
                     (N4)? data_i[65] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[32] : 
                     (N4)? data_i[64] : 1'b0;

endmodule



module bsg_mux_width_p4_els_p3
(
  data_i,
  sel_i,
  data_o
);

  input [11:0] data_i;
  input [1:0] sel_i;
  output [3:0] data_o;
  wire [3:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign N5 = N0 & N1;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign data_o[3] = (N2)? data_i[3] : 
                     (N3)? data_i[7] : 
                     (N4)? data_i[11] : 1'b0;
  assign N2 = N5;
  assign N3 = sel_i[0];
  assign N4 = sel_i[1];
  assign data_o[2] = (N2)? data_i[2] : 
                     (N3)? data_i[6] : 
                     (N4)? data_i[10] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N3)? data_i[5] : 
                     (N4)? data_i[9] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N3)? data_i[4] : 
                     (N4)? data_i[8] : 1'b0;

endmodule



module bsg_decode_num_out_p4
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_expand_bitmask_in_width_p4_expand_p1
(
  i,
  o
);

  input [3:0] i;
  output [3:0] o;
  wire [3:0] o;
  assign o[3] = i[3];
  assign o[2] = i[2];
  assign o[1] = i[1];
  assign o[0] = i[0];

endmodule



module bsg_expand_bitmask_in_width_p2_expand_p2
(
  i,
  o
);

  input [1:0] i;
  output [3:0] o;
  wire [3:0] o;
  wire o_3_,o_1_;
  assign o_3_ = i[1];
  assign o[2] = o_3_;
  assign o[3] = o_3_;
  assign o_1_ = i[0];
  assign o[0] = o_1_;
  assign o[1] = o_1_;

endmodule



module bsg_expand_bitmask_in_width_p4_expand_p8
(
  i,
  o
);

  input [3:0] i;
  output [31:0] o;
  wire [31:0] o;
  wire o_31_,o_23_,o_15_,o_7_;
  assign o_31_ = i[3];
  assign o[24] = o_31_;
  assign o[25] = o_31_;
  assign o[26] = o_31_;
  assign o[27] = o_31_;
  assign o[28] = o_31_;
  assign o[29] = o_31_;
  assign o[30] = o_31_;
  assign o[31] = o_31_;
  assign o_23_ = i[2];
  assign o[16] = o_23_;
  assign o[17] = o_23_;
  assign o[18] = o_23_;
  assign o[19] = o_23_;
  assign o[20] = o_23_;
  assign o[21] = o_23_;
  assign o[22] = o_23_;
  assign o[23] = o_23_;
  assign o_15_ = i[1];
  assign o[8] = o_15_;
  assign o[9] = o_15_;
  assign o[10] = o_15_;
  assign o[11] = o_15_;
  assign o[12] = o_15_;
  assign o[13] = o_15_;
  assign o[14] = o_15_;
  assign o[15] = o_15_;
  assign o_7_ = i[0];
  assign o[0] = o_7_;
  assign o[1] = o_7_;
  assign o[2] = o_7_;
  assign o[3] = o_7_;
  assign o[4] = o_7_;
  assign o[5] = o_7_;
  assign o[6] = o_7_;
  assign o[7] = o_7_;

endmodule



module bsg_mux_width_p8_els_p4
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [1:0] sel_i;
  output [7:0] data_o;
  wire [7:0] data_o;
  wire N0,N1,N2,N3,N4,N5;
  assign data_o[7] = (N2)? data_i[7] : 
                     (N4)? data_i[15] : 
                     (N3)? data_i[23] : 
                     (N5)? data_i[31] : 1'b0;
  assign data_o[6] = (N2)? data_i[6] : 
                     (N4)? data_i[14] : 
                     (N3)? data_i[22] : 
                     (N5)? data_i[30] : 1'b0;
  assign data_o[5] = (N2)? data_i[5] : 
                     (N4)? data_i[13] : 
                     (N3)? data_i[21] : 
                     (N5)? data_i[29] : 1'b0;
  assign data_o[4] = (N2)? data_i[4] : 
                     (N4)? data_i[12] : 
                     (N3)? data_i[20] : 
                     (N5)? data_i[28] : 1'b0;
  assign data_o[3] = (N2)? data_i[3] : 
                     (N4)? data_i[11] : 
                     (N3)? data_i[19] : 
                     (N5)? data_i[27] : 1'b0;
  assign data_o[2] = (N2)? data_i[2] : 
                     (N4)? data_i[10] : 
                     (N3)? data_i[18] : 
                     (N5)? data_i[26] : 1'b0;
  assign data_o[1] = (N2)? data_i[1] : 
                     (N4)? data_i[9] : 
                     (N3)? data_i[17] : 
                     (N5)? data_i[25] : 1'b0;
  assign data_o[0] = (N2)? data_i[0] : 
                     (N4)? data_i[8] : 
                     (N3)? data_i[16] : 
                     (N5)? data_i[24] : 1'b0;
  assign N0 = ~sel_i[0];
  assign N1 = ~sel_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & sel_i[1];
  assign N4 = sel_i[0] & N1;
  assign N5 = sel_i[0] & sel_i[1];

endmodule



module bsg_mux_width_p16_els_p2
(
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [0:0] sel_i;
  output [15:0] data_o;
  wire [15:0] data_o;
  wire N0,N1;
  assign data_o[15] = (N1)? data_i[15] : 
                      (N0)? data_i[31] : 1'b0;
  assign N0 = sel_i[0];
  assign data_o[14] = (N1)? data_i[14] : 
                      (N0)? data_i[30] : 1'b0;
  assign data_o[13] = (N1)? data_i[13] : 
                      (N0)? data_i[29] : 1'b0;
  assign data_o[12] = (N1)? data_i[12] : 
                      (N0)? data_i[28] : 1'b0;
  assign data_o[11] = (N1)? data_i[11] : 
                      (N0)? data_i[27] : 1'b0;
  assign data_o[10] = (N1)? data_i[10] : 
                      (N0)? data_i[26] : 1'b0;
  assign data_o[9] = (N1)? data_i[9] : 
                     (N0)? data_i[25] : 1'b0;
  assign data_o[8] = (N1)? data_i[8] : 
                     (N0)? data_i[24] : 1'b0;
  assign data_o[7] = (N1)? data_i[7] : 
                     (N0)? data_i[23] : 1'b0;
  assign data_o[6] = (N1)? data_i[6] : 
                     (N0)? data_i[22] : 1'b0;
  assign data_o[5] = (N1)? data_i[5] : 
                     (N0)? data_i[21] : 1'b0;
  assign data_o[4] = (N1)? data_i[4] : 
                     (N0)? data_i[20] : 1'b0;
  assign data_o[3] = (N1)? data_i[3] : 
                     (N0)? data_i[19] : 1'b0;
  assign data_o[2] = (N1)? data_i[2] : 
                     (N0)? data_i[18] : 1'b0;
  assign data_o[1] = (N1)? data_i[1] : 
                     (N0)? data_i[17] : 1'b0;
  assign data_o[0] = (N1)? data_i[0] : 
                     (N0)? data_i[16] : 1'b0;
  assign N1 = ~sel_i[0];

endmodule



module bsg_cache
(
  clk_i,
  reset_i,
  cache_pkt_i,
  v_i,
  yumi_o,
  data_o,
  v_o,
  yumi_i,
  dma_pkt_o,
  dma_pkt_v_o,
  dma_pkt_yumi_i,
  dma_data_i,
  dma_data_v_i,
  dma_data_ready_o,
  dma_data_o,
  dma_data_v_o,
  dma_data_yumi_i,
  v_we_o
);

  input [69:0] cache_pkt_i;
  output [31:0] data_o;
  output [32:0] dma_pkt_o;
  input [31:0] dma_data_i;
  output [31:0] dma_data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  input dma_pkt_yumi_i;
  input dma_data_v_i;
  input dma_data_yumi_i;
  output yumi_o;
  output v_o;
  output dma_pkt_v_o;
  output dma_data_ready_o;
  output dma_data_v_o;
  output v_we_o;
  wire [31:0] data_o,dma_data_o,data_tl_r,data_v_r,snoop_word_lo,bypass_data_lo,sbuf_data_in,
  atomic_mem_data,atomic_alu_result,\sbuf_in_sel_2_.slice_data ,ld_data_way_picked,
  ld_data_offset_picked,bypass_data_masked,snoop_or_ld_data,expanded_mask_v,
  ld_data_masked,ld_data_final_lo;
  wire [32:0] dma_pkt_o;
  wire yumi_o,v_o,dma_pkt_v_o,dma_data_ready_o,dma_data_v_o,v_we_o,N0,N1,N3,N4,N5,N6,
  N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,tl_we,
  sbuf_hazard,N65,N66,v_tl_r,N67,N68,N69,N70,N71,tag_mem_v_li,tag_mem_w_li,data_mem_v_li,
  data_mem_w_li,track_mem_v_li,track_mem_w_li,N72,N73,N74,v_v_r,N75,N76,N77,N78,
  N79,N80,N81,N82,tag_hit_found,N83,N84,N85,N86,partial_st,N87,N88,N89,N90,
  partial_st_tl,N91,N92,N93,N94,N95,partial_st_v,ld_st_amo_tag_miss,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,bypass_track_lo,track_miss,N108,N109,tagfl_hit,
  aflinv_hit,N110,N111,N112,N113,N114,N115,alock_miss,N116,N117,N118,N119,N120,
  aunlock_hit,miss_v,retval_op_v,stat_mem_v_li,stat_mem_w_li,sbuf_empty_lo,
  tbuf_empty_lo,dma_done_li,miss_track_data_we_lo,miss_stat_mem_v_lo,miss_stat_mem_w_lo,
  miss_tag_mem_v_lo,miss_tag_mem_w_lo,miss_track_mem_v_lo,miss_track_mem_w_lo,
  recover_lo,miss_done_lo,_1_net_,select_snoop_data_r_lo,dma_data_mem_v_lo,
  dma_data_mem_w_lo,dma_evict_lo,sbuf_entry_li_data__31_,sbuf_entry_li_data__30_,
  sbuf_entry_li_data__29_,sbuf_entry_li_data__28_,sbuf_entry_li_data__27_,sbuf_entry_li_data__26_,
  sbuf_entry_li_data__25_,sbuf_entry_li_data__24_,sbuf_entry_li_data__23_,
  sbuf_entry_li_data__22_,sbuf_entry_li_data__21_,sbuf_entry_li_data__20_,
  sbuf_entry_li_data__19_,sbuf_entry_li_data__18_,sbuf_entry_li_data__17_,sbuf_entry_li_data__16_,
  sbuf_entry_li_data__15_,sbuf_entry_li_data__14_,sbuf_entry_li_data__13_,
  sbuf_entry_li_data__12_,sbuf_entry_li_data__11_,sbuf_entry_li_data__10_,
  sbuf_entry_li_data__9_,sbuf_entry_li_data__8_,sbuf_entry_li_data__7_,sbuf_entry_li_data__6_,
  sbuf_entry_li_data__5_,sbuf_entry_li_data__4_,sbuf_entry_li_data__3_,
  sbuf_entry_li_data__2_,sbuf_entry_li_data__1_,sbuf_entry_li_data__0_,sbuf_entry_li_mask__3_,
  sbuf_entry_li_mask__2_,sbuf_entry_li_mask__1_,sbuf_entry_li_mask__0_,
  sbuf_entry_li_way_id__0_,sbuf_v_li,sbuf_v_lo,sbuf_yumi_li,sbuf_full_lo,sbuf_bypass_v_li,N121,
  N122,N123,N124,N125,N126,N127,N128,N129,N130,ld_data_final_li_1__31_,
  ld_data_final_li_1__30_,ld_data_final_li_1__29_,ld_data_final_li_1__28_,
  ld_data_final_li_1__27_,ld_data_final_li_1__26_,ld_data_final_li_1__25_,ld_data_final_li_1__24_,
  ld_data_final_li_1__23_,ld_data_final_li_1__22_,ld_data_final_li_1__21_,
  ld_data_final_li_1__20_,ld_data_final_li_1__19_,ld_data_final_li_1__18_,
  ld_data_final_li_1__17_,ld_data_final_li_1__16_,ld_data_final_li_0__31_,ld_data_final_li_0__30_,
  ld_data_final_li_0__29_,ld_data_final_li_0__28_,ld_data_final_li_0__27_,
  ld_data_final_li_0__26_,ld_data_final_li_0__25_,ld_data_final_li_0__24_,
  ld_data_final_li_0__23_,ld_data_final_li_0__22_,ld_data_final_li_0__21_,ld_data_final_li_0__20_,
  ld_data_final_li_0__19_,ld_data_final_li_0__18_,ld_data_final_li_0__17_,
  ld_data_final_li_0__16_,ld_data_final_li_0__15_,ld_data_final_li_0__14_,
  ld_data_final_li_0__13_,ld_data_final_li_0__12_,ld_data_final_li_0__11_,ld_data_final_li_0__10_,
  ld_data_final_li_0__9_,ld_data_final_li_0__8_,N131,N132,N133,N134,N135,N136,N137,
  N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,
  N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,
  N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,
  N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,
  N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,tbuf_v_li,tbuf_v_lo,tbuf_yumi_li,
  tbuf_full_lo,tbuf_bypass_v_li,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,tl_ready,N545,N546,tagst_write_en,N547,N548,N549,N550,N551,N552,
  N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
  N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,
  N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N2,
  N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,
  N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,
  N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,
  N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,
  N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,
  N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,
  N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,
  N712,N713,N714,N715,N716,N717,N718,N719,N720,N721;
  wire [20:0] decode,decode_tl_r,decode_v_r;
  wire [3:0] mask_tl_r,mask_v_r,dma_cmd_lo,bypass_mask_lo,sbuf_expand_mask,sbuf_mask_in,
  \sbuf_in_sel_0_.decode_lo ,tbuf_word_offset_decode;
  wire [27:0] addr_tl_r,addr_v_r,dma_addr_lo,tbuf_addr_lo;
  wire [5:0] tag_mem_addr_li,track_mem_addr_li,stat_mem_addr_li,miss_stat_mem_addr_lo,
  miss_tag_mem_addr_lo,miss_track_mem_addr_lo;
  wire [39:0] tag_mem_data_li,tag_mem_w_mask_li,tag_mem_data_lo,miss_tag_mem_data_lo,
  miss_tag_mem_w_mask_lo;
  wire [7:0] data_mem_addr_li,data_mem_w_mask_li,track_mem_data_li,track_mem_w_mask_li,
  track_mem_data_lo,track_data_v_r,miss_track_mem_w_mask_lo,miss_track_mem_data_lo,
  dma_data_mem_addr_lo,dma_data_mem_w_mask_lo,sbuf_data_mem_w_mask,
  tbuf_track_mem_w_mask,\ld_data_sel_0_.byte_sel ;
  wire [63:0] data_mem_data_li,data_mem_data_lo,ld_data_v_r,dma_data_mem_data_lo;
  wire [1:0] valid_v_r,lock_v_r,tag_hit_v,sbuf_way_decode,\sbuf_in_sel_1_.decode_lo ,
  tbuf_way_decode,addr_way_decode;
  wire [35:0] tag_v_r;
  wire [0:0] tag_hit_way_id,dma_way_lo,chosen_way_lo,sbuf_burst_offset_decode,
  \sbuf_in_sel_2_.decode_lo ,tbuf_way_li,tbuf_way_lo,plru_decode_data_lo,plru_decode_mask_lo;
  wire [2:0] stat_mem_data_li,stat_mem_w_mask_li,stat_mem_data_lo,miss_stat_mem_data_lo,
  miss_stat_mem_w_mask_lo;
  wire [64:0] sbuf_entry_lo;
  wire [11:0] sbuf_mask_in_mux_li;
  wire [15:0] \ld_data_sel_1_.byte_sel ;
  reg data_tl_r_31_sv2v_reg,data_tl_r_30_sv2v_reg,data_tl_r_29_sv2v_reg,
  data_tl_r_28_sv2v_reg,data_tl_r_27_sv2v_reg,data_tl_r_26_sv2v_reg,data_tl_r_25_sv2v_reg,
  data_tl_r_24_sv2v_reg,data_tl_r_23_sv2v_reg,data_tl_r_22_sv2v_reg,
  data_tl_r_21_sv2v_reg,data_tl_r_20_sv2v_reg,data_tl_r_19_sv2v_reg,data_tl_r_18_sv2v_reg,
  data_tl_r_17_sv2v_reg,data_tl_r_16_sv2v_reg,data_tl_r_15_sv2v_reg,data_tl_r_14_sv2v_reg,
  data_tl_r_13_sv2v_reg,data_tl_r_12_sv2v_reg,data_tl_r_11_sv2v_reg,
  data_tl_r_10_sv2v_reg,data_tl_r_9_sv2v_reg,data_tl_r_8_sv2v_reg,data_tl_r_7_sv2v_reg,
  data_tl_r_6_sv2v_reg,data_tl_r_5_sv2v_reg,data_tl_r_4_sv2v_reg,data_tl_r_3_sv2v_reg,
  data_tl_r_2_sv2v_reg,data_tl_r_1_sv2v_reg,data_tl_r_0_sv2v_reg,v_tl_r_sv2v_reg,
  decode_tl_r_20_sv2v_reg,decode_tl_r_19_sv2v_reg,decode_tl_r_18_sv2v_reg,
  decode_tl_r_17_sv2v_reg,decode_tl_r_16_sv2v_reg,decode_tl_r_15_sv2v_reg,decode_tl_r_14_sv2v_reg,
  decode_tl_r_13_sv2v_reg,decode_tl_r_12_sv2v_reg,decode_tl_r_11_sv2v_reg,
  decode_tl_r_10_sv2v_reg,decode_tl_r_9_sv2v_reg,decode_tl_r_8_sv2v_reg,
  decode_tl_r_7_sv2v_reg,decode_tl_r_6_sv2v_reg,decode_tl_r_5_sv2v_reg,decode_tl_r_4_sv2v_reg,
  decode_tl_r_3_sv2v_reg,decode_tl_r_2_sv2v_reg,decode_tl_r_1_sv2v_reg,
  decode_tl_r_0_sv2v_reg,mask_tl_r_3_sv2v_reg,mask_tl_r_2_sv2v_reg,mask_tl_r_1_sv2v_reg,
  mask_tl_r_0_sv2v_reg,addr_tl_r_27_sv2v_reg,addr_tl_r_26_sv2v_reg,addr_tl_r_25_sv2v_reg,
  addr_tl_r_24_sv2v_reg,addr_tl_r_23_sv2v_reg,addr_tl_r_22_sv2v_reg,
  addr_tl_r_21_sv2v_reg,addr_tl_r_20_sv2v_reg,addr_tl_r_19_sv2v_reg,addr_tl_r_18_sv2v_reg,
  addr_tl_r_17_sv2v_reg,addr_tl_r_16_sv2v_reg,addr_tl_r_15_sv2v_reg,addr_tl_r_14_sv2v_reg,
  addr_tl_r_13_sv2v_reg,addr_tl_r_12_sv2v_reg,addr_tl_r_11_sv2v_reg,
  addr_tl_r_10_sv2v_reg,addr_tl_r_9_sv2v_reg,addr_tl_r_8_sv2v_reg,addr_tl_r_7_sv2v_reg,
  addr_tl_r_6_sv2v_reg,addr_tl_r_5_sv2v_reg,addr_tl_r_4_sv2v_reg,addr_tl_r_3_sv2v_reg,
  addr_tl_r_2_sv2v_reg,addr_tl_r_1_sv2v_reg,addr_tl_r_0_sv2v_reg,ld_data_v_r_63_sv2v_reg,
  ld_data_v_r_62_sv2v_reg,ld_data_v_r_61_sv2v_reg,ld_data_v_r_60_sv2v_reg,
  ld_data_v_r_59_sv2v_reg,ld_data_v_r_58_sv2v_reg,ld_data_v_r_57_sv2v_reg,
  ld_data_v_r_56_sv2v_reg,ld_data_v_r_55_sv2v_reg,ld_data_v_r_54_sv2v_reg,ld_data_v_r_53_sv2v_reg,
  ld_data_v_r_52_sv2v_reg,ld_data_v_r_51_sv2v_reg,ld_data_v_r_50_sv2v_reg,
  ld_data_v_r_49_sv2v_reg,ld_data_v_r_48_sv2v_reg,ld_data_v_r_47_sv2v_reg,
  ld_data_v_r_46_sv2v_reg,ld_data_v_r_45_sv2v_reg,ld_data_v_r_44_sv2v_reg,ld_data_v_r_43_sv2v_reg,
  ld_data_v_r_42_sv2v_reg,ld_data_v_r_41_sv2v_reg,ld_data_v_r_40_sv2v_reg,
  ld_data_v_r_39_sv2v_reg,ld_data_v_r_38_sv2v_reg,ld_data_v_r_37_sv2v_reg,
  ld_data_v_r_36_sv2v_reg,ld_data_v_r_35_sv2v_reg,ld_data_v_r_34_sv2v_reg,ld_data_v_r_33_sv2v_reg,
  ld_data_v_r_32_sv2v_reg,ld_data_v_r_31_sv2v_reg,ld_data_v_r_30_sv2v_reg,
  ld_data_v_r_29_sv2v_reg,ld_data_v_r_28_sv2v_reg,ld_data_v_r_27_sv2v_reg,
  ld_data_v_r_26_sv2v_reg,ld_data_v_r_25_sv2v_reg,ld_data_v_r_24_sv2v_reg,ld_data_v_r_23_sv2v_reg,
  ld_data_v_r_22_sv2v_reg,ld_data_v_r_21_sv2v_reg,ld_data_v_r_20_sv2v_reg,
  ld_data_v_r_19_sv2v_reg,ld_data_v_r_18_sv2v_reg,ld_data_v_r_17_sv2v_reg,
  ld_data_v_r_16_sv2v_reg,ld_data_v_r_15_sv2v_reg,ld_data_v_r_14_sv2v_reg,ld_data_v_r_13_sv2v_reg,
  ld_data_v_r_12_sv2v_reg,ld_data_v_r_11_sv2v_reg,ld_data_v_r_10_sv2v_reg,
  ld_data_v_r_9_sv2v_reg,ld_data_v_r_8_sv2v_reg,ld_data_v_r_7_sv2v_reg,
  ld_data_v_r_6_sv2v_reg,ld_data_v_r_5_sv2v_reg,ld_data_v_r_4_sv2v_reg,ld_data_v_r_3_sv2v_reg,
  ld_data_v_r_2_sv2v_reg,ld_data_v_r_1_sv2v_reg,ld_data_v_r_0_sv2v_reg,v_v_r_sv2v_reg,
  track_data_v_r_7_sv2v_reg,track_data_v_r_6_sv2v_reg,track_data_v_r_5_sv2v_reg,
  track_data_v_r_4_sv2v_reg,track_data_v_r_3_sv2v_reg,track_data_v_r_2_sv2v_reg,
  track_data_v_r_1_sv2v_reg,track_data_v_r_0_sv2v_reg,mask_v_r_3_sv2v_reg,
  mask_v_r_2_sv2v_reg,mask_v_r_1_sv2v_reg,mask_v_r_0_sv2v_reg,decode_v_r_20_sv2v_reg,
  decode_v_r_19_sv2v_reg,decode_v_r_18_sv2v_reg,decode_v_r_17_sv2v_reg,decode_v_r_16_sv2v_reg,
  decode_v_r_15_sv2v_reg,decode_v_r_14_sv2v_reg,decode_v_r_13_sv2v_reg,
  decode_v_r_12_sv2v_reg,decode_v_r_11_sv2v_reg,decode_v_r_10_sv2v_reg,decode_v_r_9_sv2v_reg,
  decode_v_r_8_sv2v_reg,decode_v_r_7_sv2v_reg,decode_v_r_6_sv2v_reg,
  decode_v_r_5_sv2v_reg,decode_v_r_4_sv2v_reg,decode_v_r_3_sv2v_reg,decode_v_r_2_sv2v_reg,
  decode_v_r_1_sv2v_reg,decode_v_r_0_sv2v_reg,addr_v_r_27_sv2v_reg,addr_v_r_26_sv2v_reg,
  addr_v_r_25_sv2v_reg,addr_v_r_24_sv2v_reg,addr_v_r_23_sv2v_reg,
  addr_v_r_22_sv2v_reg,addr_v_r_21_sv2v_reg,addr_v_r_20_sv2v_reg,addr_v_r_19_sv2v_reg,
  addr_v_r_18_sv2v_reg,addr_v_r_17_sv2v_reg,addr_v_r_16_sv2v_reg,addr_v_r_15_sv2v_reg,
  addr_v_r_14_sv2v_reg,addr_v_r_13_sv2v_reg,addr_v_r_12_sv2v_reg,addr_v_r_11_sv2v_reg,
  addr_v_r_10_sv2v_reg,addr_v_r_9_sv2v_reg,addr_v_r_8_sv2v_reg,addr_v_r_7_sv2v_reg,
  addr_v_r_6_sv2v_reg,addr_v_r_5_sv2v_reg,addr_v_r_4_sv2v_reg,addr_v_r_3_sv2v_reg,
  addr_v_r_2_sv2v_reg,addr_v_r_1_sv2v_reg,addr_v_r_0_sv2v_reg,data_v_r_31_sv2v_reg,
  data_v_r_30_sv2v_reg,data_v_r_29_sv2v_reg,data_v_r_28_sv2v_reg,data_v_r_27_sv2v_reg,
  data_v_r_26_sv2v_reg,data_v_r_25_sv2v_reg,data_v_r_24_sv2v_reg,
  data_v_r_23_sv2v_reg,data_v_r_22_sv2v_reg,data_v_r_21_sv2v_reg,data_v_r_20_sv2v_reg,
  data_v_r_19_sv2v_reg,data_v_r_18_sv2v_reg,data_v_r_17_sv2v_reg,data_v_r_16_sv2v_reg,
  data_v_r_15_sv2v_reg,data_v_r_14_sv2v_reg,data_v_r_13_sv2v_reg,data_v_r_12_sv2v_reg,
  data_v_r_11_sv2v_reg,data_v_r_10_sv2v_reg,data_v_r_9_sv2v_reg,data_v_r_8_sv2v_reg,
  data_v_r_7_sv2v_reg,data_v_r_6_sv2v_reg,data_v_r_5_sv2v_reg,data_v_r_4_sv2v_reg,
  data_v_r_3_sv2v_reg,data_v_r_2_sv2v_reg,data_v_r_1_sv2v_reg,data_v_r_0_sv2v_reg,
  valid_v_r_1_sv2v_reg,valid_v_r_0_sv2v_reg,lock_v_r_1_sv2v_reg,lock_v_r_0_sv2v_reg,
  tag_v_r_35_sv2v_reg,tag_v_r_34_sv2v_reg,tag_v_r_33_sv2v_reg,tag_v_r_32_sv2v_reg,
  tag_v_r_31_sv2v_reg,tag_v_r_30_sv2v_reg,tag_v_r_29_sv2v_reg,tag_v_r_28_sv2v_reg,
  tag_v_r_27_sv2v_reg,tag_v_r_26_sv2v_reg,tag_v_r_25_sv2v_reg,tag_v_r_24_sv2v_reg,
  tag_v_r_23_sv2v_reg,tag_v_r_22_sv2v_reg,tag_v_r_21_sv2v_reg,tag_v_r_20_sv2v_reg,
  tag_v_r_19_sv2v_reg,tag_v_r_18_sv2v_reg,tag_v_r_17_sv2v_reg,tag_v_r_16_sv2v_reg,
  tag_v_r_15_sv2v_reg,tag_v_r_14_sv2v_reg,tag_v_r_13_sv2v_reg,tag_v_r_12_sv2v_reg,
  tag_v_r_11_sv2v_reg,tag_v_r_10_sv2v_reg,tag_v_r_9_sv2v_reg,tag_v_r_8_sv2v_reg,
  tag_v_r_7_sv2v_reg,tag_v_r_6_sv2v_reg,tag_v_r_5_sv2v_reg,tag_v_r_4_sv2v_reg,
  tag_v_r_3_sv2v_reg,tag_v_r_2_sv2v_reg,tag_v_r_1_sv2v_reg,tag_v_r_0_sv2v_reg;
  assign data_tl_r[31] = data_tl_r_31_sv2v_reg;
  assign data_tl_r[30] = data_tl_r_30_sv2v_reg;
  assign data_tl_r[29] = data_tl_r_29_sv2v_reg;
  assign data_tl_r[28] = data_tl_r_28_sv2v_reg;
  assign data_tl_r[27] = data_tl_r_27_sv2v_reg;
  assign data_tl_r[26] = data_tl_r_26_sv2v_reg;
  assign data_tl_r[25] = data_tl_r_25_sv2v_reg;
  assign data_tl_r[24] = data_tl_r_24_sv2v_reg;
  assign data_tl_r[23] = data_tl_r_23_sv2v_reg;
  assign data_tl_r[22] = data_tl_r_22_sv2v_reg;
  assign data_tl_r[21] = data_tl_r_21_sv2v_reg;
  assign data_tl_r[20] = data_tl_r_20_sv2v_reg;
  assign data_tl_r[19] = data_tl_r_19_sv2v_reg;
  assign data_tl_r[18] = data_tl_r_18_sv2v_reg;
  assign data_tl_r[17] = data_tl_r_17_sv2v_reg;
  assign data_tl_r[16] = data_tl_r_16_sv2v_reg;
  assign data_tl_r[15] = data_tl_r_15_sv2v_reg;
  assign data_tl_r[14] = data_tl_r_14_sv2v_reg;
  assign data_tl_r[13] = data_tl_r_13_sv2v_reg;
  assign data_tl_r[12] = data_tl_r_12_sv2v_reg;
  assign data_tl_r[11] = data_tl_r_11_sv2v_reg;
  assign data_tl_r[10] = data_tl_r_10_sv2v_reg;
  assign data_tl_r[9] = data_tl_r_9_sv2v_reg;
  assign data_tl_r[8] = data_tl_r_8_sv2v_reg;
  assign data_tl_r[7] = data_tl_r_7_sv2v_reg;
  assign data_tl_r[6] = data_tl_r_6_sv2v_reg;
  assign data_tl_r[5] = data_tl_r_5_sv2v_reg;
  assign data_tl_r[4] = data_tl_r_4_sv2v_reg;
  assign data_tl_r[3] = data_tl_r_3_sv2v_reg;
  assign data_tl_r[2] = data_tl_r_2_sv2v_reg;
  assign data_tl_r[1] = data_tl_r_1_sv2v_reg;
  assign data_tl_r[0] = data_tl_r_0_sv2v_reg;
  assign v_tl_r = v_tl_r_sv2v_reg;
  assign decode_tl_r[20] = decode_tl_r_20_sv2v_reg;
  assign decode_tl_r[19] = decode_tl_r_19_sv2v_reg;
  assign decode_tl_r[18] = decode_tl_r_18_sv2v_reg;
  assign decode_tl_r[17] = decode_tl_r_17_sv2v_reg;
  assign decode_tl_r[16] = decode_tl_r_16_sv2v_reg;
  assign decode_tl_r[15] = decode_tl_r_15_sv2v_reg;
  assign decode_tl_r[14] = decode_tl_r_14_sv2v_reg;
  assign decode_tl_r[13] = decode_tl_r_13_sv2v_reg;
  assign decode_tl_r[12] = decode_tl_r_12_sv2v_reg;
  assign decode_tl_r[11] = decode_tl_r_11_sv2v_reg;
  assign decode_tl_r[10] = decode_tl_r_10_sv2v_reg;
  assign decode_tl_r[9] = decode_tl_r_9_sv2v_reg;
  assign decode_tl_r[8] = decode_tl_r_8_sv2v_reg;
  assign decode_tl_r[7] = decode_tl_r_7_sv2v_reg;
  assign decode_tl_r[6] = decode_tl_r_6_sv2v_reg;
  assign decode_tl_r[5] = decode_tl_r_5_sv2v_reg;
  assign decode_tl_r[4] = decode_tl_r_4_sv2v_reg;
  assign decode_tl_r[3] = decode_tl_r_3_sv2v_reg;
  assign decode_tl_r[2] = decode_tl_r_2_sv2v_reg;
  assign decode_tl_r[1] = decode_tl_r_1_sv2v_reg;
  assign decode_tl_r[0] = decode_tl_r_0_sv2v_reg;
  assign mask_tl_r[3] = mask_tl_r_3_sv2v_reg;
  assign mask_tl_r[2] = mask_tl_r_2_sv2v_reg;
  assign mask_tl_r[1] = mask_tl_r_1_sv2v_reg;
  assign mask_tl_r[0] = mask_tl_r_0_sv2v_reg;
  assign addr_tl_r[27] = addr_tl_r_27_sv2v_reg;
  assign addr_tl_r[26] = addr_tl_r_26_sv2v_reg;
  assign addr_tl_r[25] = addr_tl_r_25_sv2v_reg;
  assign addr_tl_r[24] = addr_tl_r_24_sv2v_reg;
  assign addr_tl_r[23] = addr_tl_r_23_sv2v_reg;
  assign addr_tl_r[22] = addr_tl_r_22_sv2v_reg;
  assign addr_tl_r[21] = addr_tl_r_21_sv2v_reg;
  assign addr_tl_r[20] = addr_tl_r_20_sv2v_reg;
  assign addr_tl_r[19] = addr_tl_r_19_sv2v_reg;
  assign addr_tl_r[18] = addr_tl_r_18_sv2v_reg;
  assign addr_tl_r[17] = addr_tl_r_17_sv2v_reg;
  assign addr_tl_r[16] = addr_tl_r_16_sv2v_reg;
  assign addr_tl_r[15] = addr_tl_r_15_sv2v_reg;
  assign addr_tl_r[14] = addr_tl_r_14_sv2v_reg;
  assign addr_tl_r[13] = addr_tl_r_13_sv2v_reg;
  assign addr_tl_r[12] = addr_tl_r_12_sv2v_reg;
  assign addr_tl_r[11] = addr_tl_r_11_sv2v_reg;
  assign addr_tl_r[10] = addr_tl_r_10_sv2v_reg;
  assign addr_tl_r[9] = addr_tl_r_9_sv2v_reg;
  assign addr_tl_r[8] = addr_tl_r_8_sv2v_reg;
  assign addr_tl_r[7] = addr_tl_r_7_sv2v_reg;
  assign addr_tl_r[6] = addr_tl_r_6_sv2v_reg;
  assign addr_tl_r[5] = addr_tl_r_5_sv2v_reg;
  assign addr_tl_r[4] = addr_tl_r_4_sv2v_reg;
  assign addr_tl_r[3] = addr_tl_r_3_sv2v_reg;
  assign addr_tl_r[2] = addr_tl_r_2_sv2v_reg;
  assign addr_tl_r[1] = addr_tl_r_1_sv2v_reg;
  assign addr_tl_r[0] = addr_tl_r_0_sv2v_reg;
  assign ld_data_v_r[63] = ld_data_v_r_63_sv2v_reg;
  assign ld_data_v_r[62] = ld_data_v_r_62_sv2v_reg;
  assign ld_data_v_r[61] = ld_data_v_r_61_sv2v_reg;
  assign ld_data_v_r[60] = ld_data_v_r_60_sv2v_reg;
  assign ld_data_v_r[59] = ld_data_v_r_59_sv2v_reg;
  assign ld_data_v_r[58] = ld_data_v_r_58_sv2v_reg;
  assign ld_data_v_r[57] = ld_data_v_r_57_sv2v_reg;
  assign ld_data_v_r[56] = ld_data_v_r_56_sv2v_reg;
  assign ld_data_v_r[55] = ld_data_v_r_55_sv2v_reg;
  assign ld_data_v_r[54] = ld_data_v_r_54_sv2v_reg;
  assign ld_data_v_r[53] = ld_data_v_r_53_sv2v_reg;
  assign ld_data_v_r[52] = ld_data_v_r_52_sv2v_reg;
  assign ld_data_v_r[51] = ld_data_v_r_51_sv2v_reg;
  assign ld_data_v_r[50] = ld_data_v_r_50_sv2v_reg;
  assign ld_data_v_r[49] = ld_data_v_r_49_sv2v_reg;
  assign ld_data_v_r[48] = ld_data_v_r_48_sv2v_reg;
  assign ld_data_v_r[47] = ld_data_v_r_47_sv2v_reg;
  assign ld_data_v_r[46] = ld_data_v_r_46_sv2v_reg;
  assign ld_data_v_r[45] = ld_data_v_r_45_sv2v_reg;
  assign ld_data_v_r[44] = ld_data_v_r_44_sv2v_reg;
  assign ld_data_v_r[43] = ld_data_v_r_43_sv2v_reg;
  assign ld_data_v_r[42] = ld_data_v_r_42_sv2v_reg;
  assign ld_data_v_r[41] = ld_data_v_r_41_sv2v_reg;
  assign ld_data_v_r[40] = ld_data_v_r_40_sv2v_reg;
  assign ld_data_v_r[39] = ld_data_v_r_39_sv2v_reg;
  assign ld_data_v_r[38] = ld_data_v_r_38_sv2v_reg;
  assign ld_data_v_r[37] = ld_data_v_r_37_sv2v_reg;
  assign ld_data_v_r[36] = ld_data_v_r_36_sv2v_reg;
  assign ld_data_v_r[35] = ld_data_v_r_35_sv2v_reg;
  assign ld_data_v_r[34] = ld_data_v_r_34_sv2v_reg;
  assign ld_data_v_r[33] = ld_data_v_r_33_sv2v_reg;
  assign ld_data_v_r[32] = ld_data_v_r_32_sv2v_reg;
  assign ld_data_v_r[31] = ld_data_v_r_31_sv2v_reg;
  assign ld_data_v_r[30] = ld_data_v_r_30_sv2v_reg;
  assign ld_data_v_r[29] = ld_data_v_r_29_sv2v_reg;
  assign ld_data_v_r[28] = ld_data_v_r_28_sv2v_reg;
  assign ld_data_v_r[27] = ld_data_v_r_27_sv2v_reg;
  assign ld_data_v_r[26] = ld_data_v_r_26_sv2v_reg;
  assign ld_data_v_r[25] = ld_data_v_r_25_sv2v_reg;
  assign ld_data_v_r[24] = ld_data_v_r_24_sv2v_reg;
  assign ld_data_v_r[23] = ld_data_v_r_23_sv2v_reg;
  assign ld_data_v_r[22] = ld_data_v_r_22_sv2v_reg;
  assign ld_data_v_r[21] = ld_data_v_r_21_sv2v_reg;
  assign ld_data_v_r[20] = ld_data_v_r_20_sv2v_reg;
  assign ld_data_v_r[19] = ld_data_v_r_19_sv2v_reg;
  assign ld_data_v_r[18] = ld_data_v_r_18_sv2v_reg;
  assign ld_data_v_r[17] = ld_data_v_r_17_sv2v_reg;
  assign ld_data_v_r[16] = ld_data_v_r_16_sv2v_reg;
  assign ld_data_v_r[15] = ld_data_v_r_15_sv2v_reg;
  assign ld_data_v_r[14] = ld_data_v_r_14_sv2v_reg;
  assign ld_data_v_r[13] = ld_data_v_r_13_sv2v_reg;
  assign ld_data_v_r[12] = ld_data_v_r_12_sv2v_reg;
  assign ld_data_v_r[11] = ld_data_v_r_11_sv2v_reg;
  assign ld_data_v_r[10] = ld_data_v_r_10_sv2v_reg;
  assign ld_data_v_r[9] = ld_data_v_r_9_sv2v_reg;
  assign ld_data_v_r[8] = ld_data_v_r_8_sv2v_reg;
  assign ld_data_v_r[7] = ld_data_v_r_7_sv2v_reg;
  assign ld_data_v_r[6] = ld_data_v_r_6_sv2v_reg;
  assign ld_data_v_r[5] = ld_data_v_r_5_sv2v_reg;
  assign ld_data_v_r[4] = ld_data_v_r_4_sv2v_reg;
  assign ld_data_v_r[3] = ld_data_v_r_3_sv2v_reg;
  assign ld_data_v_r[2] = ld_data_v_r_2_sv2v_reg;
  assign ld_data_v_r[1] = ld_data_v_r_1_sv2v_reg;
  assign ld_data_v_r[0] = ld_data_v_r_0_sv2v_reg;
  assign v_v_r = v_v_r_sv2v_reg;
  assign track_data_v_r[7] = track_data_v_r_7_sv2v_reg;
  assign track_data_v_r[6] = track_data_v_r_6_sv2v_reg;
  assign track_data_v_r[5] = track_data_v_r_5_sv2v_reg;
  assign track_data_v_r[4] = track_data_v_r_4_sv2v_reg;
  assign track_data_v_r[3] = track_data_v_r_3_sv2v_reg;
  assign track_data_v_r[2] = track_data_v_r_2_sv2v_reg;
  assign track_data_v_r[1] = track_data_v_r_1_sv2v_reg;
  assign track_data_v_r[0] = track_data_v_r_0_sv2v_reg;
  assign mask_v_r[3] = mask_v_r_3_sv2v_reg;
  assign mask_v_r[2] = mask_v_r_2_sv2v_reg;
  assign mask_v_r[1] = mask_v_r_1_sv2v_reg;
  assign mask_v_r[0] = mask_v_r_0_sv2v_reg;
  assign decode_v_r[20] = decode_v_r_20_sv2v_reg;
  assign decode_v_r[19] = decode_v_r_19_sv2v_reg;
  assign decode_v_r[18] = decode_v_r_18_sv2v_reg;
  assign decode_v_r[17] = decode_v_r_17_sv2v_reg;
  assign decode_v_r[16] = decode_v_r_16_sv2v_reg;
  assign decode_v_r[15] = decode_v_r_15_sv2v_reg;
  assign decode_v_r[14] = decode_v_r_14_sv2v_reg;
  assign decode_v_r[13] = decode_v_r_13_sv2v_reg;
  assign decode_v_r[12] = decode_v_r_12_sv2v_reg;
  assign decode_v_r[11] = decode_v_r_11_sv2v_reg;
  assign decode_v_r[10] = decode_v_r_10_sv2v_reg;
  assign decode_v_r[9] = decode_v_r_9_sv2v_reg;
  assign decode_v_r[8] = decode_v_r_8_sv2v_reg;
  assign decode_v_r[7] = decode_v_r_7_sv2v_reg;
  assign decode_v_r[6] = decode_v_r_6_sv2v_reg;
  assign decode_v_r[5] = decode_v_r_5_sv2v_reg;
  assign decode_v_r[4] = decode_v_r_4_sv2v_reg;
  assign decode_v_r[3] = decode_v_r_3_sv2v_reg;
  assign decode_v_r[2] = decode_v_r_2_sv2v_reg;
  assign decode_v_r[1] = decode_v_r_1_sv2v_reg;
  assign decode_v_r[0] = decode_v_r_0_sv2v_reg;
  assign addr_v_r[27] = addr_v_r_27_sv2v_reg;
  assign addr_v_r[26] = addr_v_r_26_sv2v_reg;
  assign addr_v_r[25] = addr_v_r_25_sv2v_reg;
  assign addr_v_r[24] = addr_v_r_24_sv2v_reg;
  assign addr_v_r[23] = addr_v_r_23_sv2v_reg;
  assign addr_v_r[22] = addr_v_r_22_sv2v_reg;
  assign addr_v_r[21] = addr_v_r_21_sv2v_reg;
  assign addr_v_r[20] = addr_v_r_20_sv2v_reg;
  assign addr_v_r[19] = addr_v_r_19_sv2v_reg;
  assign addr_v_r[18] = addr_v_r_18_sv2v_reg;
  assign addr_v_r[17] = addr_v_r_17_sv2v_reg;
  assign addr_v_r[16] = addr_v_r_16_sv2v_reg;
  assign addr_v_r[15] = addr_v_r_15_sv2v_reg;
  assign addr_v_r[14] = addr_v_r_14_sv2v_reg;
  assign addr_v_r[13] = addr_v_r_13_sv2v_reg;
  assign addr_v_r[12] = addr_v_r_12_sv2v_reg;
  assign addr_v_r[11] = addr_v_r_11_sv2v_reg;
  assign addr_v_r[10] = addr_v_r_10_sv2v_reg;
  assign addr_v_r[9] = addr_v_r_9_sv2v_reg;
  assign addr_v_r[8] = addr_v_r_8_sv2v_reg;
  assign addr_v_r[7] = addr_v_r_7_sv2v_reg;
  assign addr_v_r[6] = addr_v_r_6_sv2v_reg;
  assign addr_v_r[5] = addr_v_r_5_sv2v_reg;
  assign addr_v_r[4] = addr_v_r_4_sv2v_reg;
  assign addr_v_r[3] = addr_v_r_3_sv2v_reg;
  assign addr_v_r[2] = addr_v_r_2_sv2v_reg;
  assign addr_v_r[1] = addr_v_r_1_sv2v_reg;
  assign addr_v_r[0] = addr_v_r_0_sv2v_reg;
  assign data_v_r[31] = data_v_r_31_sv2v_reg;
  assign data_v_r[30] = data_v_r_30_sv2v_reg;
  assign data_v_r[29] = data_v_r_29_sv2v_reg;
  assign data_v_r[28] = data_v_r_28_sv2v_reg;
  assign data_v_r[27] = data_v_r_27_sv2v_reg;
  assign data_v_r[26] = data_v_r_26_sv2v_reg;
  assign data_v_r[25] = data_v_r_25_sv2v_reg;
  assign data_v_r[24] = data_v_r_24_sv2v_reg;
  assign data_v_r[23] = data_v_r_23_sv2v_reg;
  assign data_v_r[22] = data_v_r_22_sv2v_reg;
  assign data_v_r[21] = data_v_r_21_sv2v_reg;
  assign data_v_r[20] = data_v_r_20_sv2v_reg;
  assign data_v_r[19] = data_v_r_19_sv2v_reg;
  assign data_v_r[18] = data_v_r_18_sv2v_reg;
  assign data_v_r[17] = data_v_r_17_sv2v_reg;
  assign data_v_r[16] = data_v_r_16_sv2v_reg;
  assign data_v_r[15] = data_v_r_15_sv2v_reg;
  assign data_v_r[14] = data_v_r_14_sv2v_reg;
  assign data_v_r[13] = data_v_r_13_sv2v_reg;
  assign data_v_r[12] = data_v_r_12_sv2v_reg;
  assign data_v_r[11] = data_v_r_11_sv2v_reg;
  assign data_v_r[10] = data_v_r_10_sv2v_reg;
  assign data_v_r[9] = data_v_r_9_sv2v_reg;
  assign data_v_r[8] = data_v_r_8_sv2v_reg;
  assign data_v_r[7] = data_v_r_7_sv2v_reg;
  assign data_v_r[6] = data_v_r_6_sv2v_reg;
  assign data_v_r[5] = data_v_r_5_sv2v_reg;
  assign data_v_r[4] = data_v_r_4_sv2v_reg;
  assign data_v_r[3] = data_v_r_3_sv2v_reg;
  assign data_v_r[2] = data_v_r_2_sv2v_reg;
  assign data_v_r[1] = data_v_r_1_sv2v_reg;
  assign data_v_r[0] = data_v_r_0_sv2v_reg;
  assign valid_v_r[1] = valid_v_r_1_sv2v_reg;
  assign valid_v_r[0] = valid_v_r_0_sv2v_reg;
  assign lock_v_r[1] = lock_v_r_1_sv2v_reg;
  assign lock_v_r[0] = lock_v_r_0_sv2v_reg;
  assign tag_v_r[35] = tag_v_r_35_sv2v_reg;
  assign tag_v_r[34] = tag_v_r_34_sv2v_reg;
  assign tag_v_r[33] = tag_v_r_33_sv2v_reg;
  assign tag_v_r[32] = tag_v_r_32_sv2v_reg;
  assign tag_v_r[31] = tag_v_r_31_sv2v_reg;
  assign tag_v_r[30] = tag_v_r_30_sv2v_reg;
  assign tag_v_r[29] = tag_v_r_29_sv2v_reg;
  assign tag_v_r[28] = tag_v_r_28_sv2v_reg;
  assign tag_v_r[27] = tag_v_r_27_sv2v_reg;
  assign tag_v_r[26] = tag_v_r_26_sv2v_reg;
  assign tag_v_r[25] = tag_v_r_25_sv2v_reg;
  assign tag_v_r[24] = tag_v_r_24_sv2v_reg;
  assign tag_v_r[23] = tag_v_r_23_sv2v_reg;
  assign tag_v_r[22] = tag_v_r_22_sv2v_reg;
  assign tag_v_r[21] = tag_v_r_21_sv2v_reg;
  assign tag_v_r[20] = tag_v_r_20_sv2v_reg;
  assign tag_v_r[19] = tag_v_r_19_sv2v_reg;
  assign tag_v_r[18] = tag_v_r_18_sv2v_reg;
  assign tag_v_r[17] = tag_v_r_17_sv2v_reg;
  assign tag_v_r[16] = tag_v_r_16_sv2v_reg;
  assign tag_v_r[15] = tag_v_r_15_sv2v_reg;
  assign tag_v_r[14] = tag_v_r_14_sv2v_reg;
  assign tag_v_r[13] = tag_v_r_13_sv2v_reg;
  assign tag_v_r[12] = tag_v_r_12_sv2v_reg;
  assign tag_v_r[11] = tag_v_r_11_sv2v_reg;
  assign tag_v_r[10] = tag_v_r_10_sv2v_reg;
  assign tag_v_r[9] = tag_v_r_9_sv2v_reg;
  assign tag_v_r[8] = tag_v_r_8_sv2v_reg;
  assign tag_v_r[7] = tag_v_r_7_sv2v_reg;
  assign tag_v_r[6] = tag_v_r_6_sv2v_reg;
  assign tag_v_r[5] = tag_v_r_5_sv2v_reg;
  assign tag_v_r[4] = tag_v_r_4_sv2v_reg;
  assign tag_v_r[3] = tag_v_r_3_sv2v_reg;
  assign tag_v_r[2] = tag_v_r_2_sv2v_reg;
  assign tag_v_r[1] = tag_v_r_1_sv2v_reg;
  assign tag_v_r[0] = tag_v_r_0_sv2v_reg;

  bsg_cache_decode
  decode0
  (
    .opcode_i(cache_pkt_i[69:64]),
    .decode_o(decode)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p40_els_p64_latch_last_read_p1
  tag_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(tag_mem_data_li),
    .addr_i(tag_mem_addr_li),
    .v_i(tag_mem_v_li),
    .w_mask_i(tag_mem_w_mask_li),
    .w_i(tag_mem_w_li),
    .data_o(tag_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_byte_els_p256_data_width_p64_latch_last_read_p1
  data_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(data_mem_v_li),
    .w_i(data_mem_w_li),
    .addr_i(data_mem_addr_li),
    .data_i(data_mem_data_li),
    .write_mask_i(data_mem_w_mask_li),
    .data_o(data_mem_data_lo)
  );


  bsg_mem_1rw_sync_mask_write_bit_width_p8_els_p64_latch_last_read_p1
  \track_mem_gen.track_mem 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(track_mem_data_li),
    .addr_i(track_mem_addr_li),
    .v_i(track_mem_v_li),
    .w_mask_i(track_mem_w_mask_li),
    .w_i(track_mem_w_li),
    .data_o(track_mem_data_lo)
  );

  assign N81 = addr_v_r[27:10] == tag_v_r[17:0];
  assign N82 = addr_v_r[27:10] == tag_v_r[35:18];

  bsg_priority_encode_width_p2_lo_to_hi_p1
  tag_hit_pe
  (
    .i(tag_hit_v),
    .addr_o(tag_hit_way_id[0]),
    .v_o(tag_hit_found)
  );

  assign N97 = (N96)? track_data_v_r[3] : 
               (N0)? track_data_v_r[7] : 1'b0;
  assign N0 = tag_hit_way_id[0];
  assign N98 = (N96)? track_data_v_r[2] : 
               (N0)? track_data_v_r[6] : 1'b0;
  assign N99 = (N96)? track_data_v_r[1] : 
               (N0)? track_data_v_r[5] : 1'b0;
  assign N100 = (N96)? track_data_v_r[0] : 
                (N0)? track_data_v_r[4] : 1'b0;
  assign N107 = (N103)? N100 : 
                (N105)? N99 : 
                (N104)? N98 : 
                (N106)? N97 : 1'b0;
  assign N109 = (N108)? valid_v_r[0] : 
                (N1)? valid_v_r[1] : 1'b0;
  assign N1 = addr_v_r[10];
  assign N113 = (N112)? lock_v_r[0] : 
                (N0)? lock_v_r[1] : 1'b0;
  assign N119 = (N118)? lock_v_r[0] : 
                (N0)? lock_v_r[1] : 1'b0;

  bsg_mem_1rw_sync_mask_write_bit_width_p3_els_p64_latch_last_read_p1
  stat_mem
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(stat_mem_data_li),
    .addr_i(stat_mem_addr_li),
    .v_i(stat_mem_v_li),
    .w_mask_i(stat_mem_w_mask_li),
    .w_i(stat_mem_w_li),
    .data_o(stat_mem_data_lo)
  );


  bsg_cache_miss_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2_word_tracking_p1
  miss
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .miss_v_i(miss_v),
    .track_miss_i(track_miss),
    .decode_v_i(decode_v_r),
    .addr_v_i(addr_v_r),
    .mask_v_i(mask_v_r),
    .tag_v_i(tag_v_r),
    .valid_v_i(valid_v_r),
    .lock_v_i(lock_v_r),
    .tag_hit_v_i(tag_hit_v),
    .tag_hit_way_id_i(tag_hit_way_id[0]),
    .tag_hit_found_i(tag_hit_found),
    .sbuf_empty_i(sbuf_empty_lo),
    .tbuf_empty_i(tbuf_empty_lo),
    .dma_cmd_o(dma_cmd_lo),
    .dma_way_o(dma_way_lo[0]),
    .dma_addr_o(dma_addr_lo),
    .dma_done_i(dma_done_li),
    .track_data_we_o(miss_track_data_we_lo),
    .stat_info_i(stat_mem_data_lo),
    .stat_mem_v_o(miss_stat_mem_v_lo),
    .stat_mem_w_o(miss_stat_mem_w_lo),
    .stat_mem_addr_o(miss_stat_mem_addr_lo),
    .stat_mem_data_o(miss_stat_mem_data_lo),
    .stat_mem_w_mask_o(miss_stat_mem_w_mask_lo),
    .tag_mem_v_o(miss_tag_mem_v_lo),
    .tag_mem_w_o(miss_tag_mem_w_lo),
    .tag_mem_addr_o(miss_tag_mem_addr_lo),
    .tag_mem_data_o(miss_tag_mem_data_lo),
    .tag_mem_w_mask_o(miss_tag_mem_w_mask_lo),
    .track_mem_v_o(miss_track_mem_v_lo),
    .track_mem_w_o(miss_track_mem_w_lo),
    .track_mem_addr_o(miss_track_mem_addr_lo),
    .track_mem_w_mask_o(miss_track_mem_w_mask_lo),
    .track_mem_data_o(miss_track_mem_data_lo),
    .done_o(miss_done_lo),
    .recover_o(recover_lo),
    .chosen_way_o(chosen_way_lo[0]),
    .select_snoop_data_r_o(select_snoop_data_r_lo),
    .ack_i(_1_net_)
  );


  bsg_cache_dma_addr_width_p28_data_width_p32_block_size_in_words_p4_sets_p64_ways_p2_word_tracking_p1_dma_data_width_p32_debug_p0
  dma
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .dma_cmd_i(dma_cmd_lo),
    .dma_way_i(dma_way_lo[0]),
    .dma_addr_i(dma_addr_lo),
    .done_o(dma_done_li),
    .track_data_we_i(miss_track_data_we_lo),
    .snoop_word_o(snoop_word_lo),
    .dma_pkt_o(dma_pkt_o),
    .dma_pkt_v_o(dma_pkt_v_o),
    .dma_pkt_yumi_i(dma_pkt_yumi_i),
    .dma_data_i(dma_data_i),
    .dma_data_v_i(dma_data_v_i),
    .dma_data_ready_o(dma_data_ready_o),
    .dma_data_o(dma_data_o),
    .dma_data_v_o(dma_data_v_o),
    .dma_data_yumi_i(dma_data_yumi_i),
    .data_mem_v_o(dma_data_mem_v_lo),
    .data_mem_w_o(dma_data_mem_w_lo),
    .data_mem_addr_o(dma_data_mem_addr_lo),
    .data_mem_w_mask_o(dma_data_mem_w_mask_lo),
    .data_mem_data_o(dma_data_mem_data_lo),
    .data_mem_data_i(data_mem_data_lo),
    .track_miss_i(track_miss),
    .track_mem_data_i(track_mem_data_lo),
    .dma_evict_o(dma_evict_lo)
  );


  bsg_cache_sbuf_data_width_p32_addr_width_p28_ways_p2
  sbuf
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .sbuf_entry_i({ addr_v_r, sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_, sbuf_entry_li_way_id__0_ }),
    .v_i(sbuf_v_li),
    .sbuf_entry_o(sbuf_entry_lo),
    .v_o(sbuf_v_lo),
    .yumi_i(sbuf_yumi_li),
    .empty_o(sbuf_empty_lo),
    .full_o(sbuf_full_lo),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(sbuf_bypass_v_li),
    .bypass_data_o(bypass_data_lo),
    .bypass_mask_o(bypass_mask_lo)
  );


  bsg_decode_num_out_p2
  sbuf_way_demux
  (
    .i(sbuf_entry_lo[0]),
    .o(sbuf_way_decode)
  );


  bsg_decode_num_out_p1
  sbuf_bo_demux
  (
    .i(sbuf_entry_lo[39]),
    .o(sbuf_burst_offset_decode[0])
  );


  bsg_expand_bitmask_in_width_p1_expand_p4
  expand0
  (
    .i(sbuf_burst_offset_decode[0]),
    .o(sbuf_expand_mask)
  );


  bsg_mux_width_p32_els_p3
  sbuf_data_in_mux
  (
    .data_i({ \sbuf_in_sel_2_.slice_data , data_v_r[15:0], data_v_r[15:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0], data_v_r[7:0] }),
    .sel_i(decode_v_r[20:19]),
    .data_o(sbuf_data_in)
  );


  bsg_mux_width_p4_els_p3
  sbuf_mask_in_mux
  (
    .data_i(sbuf_mask_in_mux_li),
    .sel_i(decode_v_r[20:19]),
    .data_o(sbuf_mask_in)
  );

  assign N133 = N132 | decode_v_r[3];
  assign N134 = decode_v_r[2] | decode_v_r[1];
  assign N135 = N133 | N134;
  assign N136 = N135 | decode_v_r[0];
  assign N140 = N132 | decode_v_r[3];
  assign N141 = decode_v_r[2] | N138;
  assign N142 = N140 | N141;
  assign N143 = N142 | N139;
  assign N146 = N132 | decode_v_r[3];
  assign N147 = N145 | decode_v_r[1];
  assign N148 = N146 | N147;
  assign N149 = N148 | decode_v_r[0];
  assign N152 = N132 | decode_v_r[3];
  assign N153 = decode_v_r[2] | N151;
  assign N154 = N152 | N153;
  assign N155 = N154 | decode_v_r[0];
  assign N158 = N132 | decode_v_r[3];
  assign N159 = decode_v_r[2] | decode_v_r[1];
  assign N160 = N158 | N159;
  assign N161 = N160 | N157;
  assign N165 = N132 | decode_v_r[3];
  assign N166 = N163 | decode_v_r[1];
  assign N167 = N165 | N166;
  assign N168 = N167 | N164;
  assign N172 = N132 | decode_v_r[3];
  assign N173 = N170 | N171;
  assign N174 = N172 | N173;
  assign N175 = N174 | decode_v_r[0];
  assign N180 = N132 | decode_v_r[3];
  assign N181 = N177 | N178;
  assign N182 = N180 | N181;
  assign N183 = N182 | N179;
  assign N186 = N132 | N185;
  assign N187 = decode_v_r[2] | decode_v_r[1];
  assign N188 = N186 | N187;
  assign N189 = N188 | decode_v_r[0];
  assign N191 = N131 & decode_v_r[3];
  assign N192 = N191 & decode_v_r[0];
  assign N193 = N131 & decode_v_r[3];
  assign N194 = N193 & decode_v_r[1];
  assign N195 = N131 & decode_v_r[3];
  assign N196 = N195 & decode_v_r[2];
  assign N326 = $signed(data_v_r) < $signed(atomic_mem_data);
  assign N360 = $signed(data_v_r) > $signed(atomic_mem_data);
  assign N394 = data_v_r < atomic_mem_data;
  assign N428 = data_v_r > atomic_mem_data;

  bsg_decode_num_out_p4
  \sbuf_in_sel_0_.dec 
  (
    .i(addr_v_r[1:0]),
    .o(\sbuf_in_sel_0_.decode_lo )
  );


  bsg_expand_bitmask_in_width_p4_expand_p1
  \sbuf_in_sel_0_.exp 
  (
    .i(\sbuf_in_sel_0_.decode_lo ),
    .o(sbuf_mask_in_mux_li[3:0])
  );


  bsg_decode_num_out_p2
  \sbuf_in_sel_1_.dec 
  (
    .i(addr_v_r[1]),
    .o(\sbuf_in_sel_1_.decode_lo )
  );


  bsg_expand_bitmask_in_width_p2_expand_p2
  \sbuf_in_sel_1_.exp 
  (
    .i(\sbuf_in_sel_1_.decode_lo ),
    .o(sbuf_mask_in_mux_li[7:4])
  );


  bsg_decode_num_out_p1
  \sbuf_in_sel_2_.dec 
  (
    .i(addr_v_r[2]),
    .o(\sbuf_in_sel_2_.decode_lo [0])
  );


  bsg_expand_bitmask_in_width_p1_expand_p4
  \sbuf_in_sel_2_.exp 
  (
    .i(\sbuf_in_sel_2_.decode_lo [0]),
    .o(sbuf_mask_in_mux_li[11:8])
  );


  bsg_cache_tbuf
  \tbuf_gen.tbuf 
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .addr_i(addr_v_r),
    .way_i(tbuf_way_li[0]),
    .v_i(tbuf_v_li),
    .addr_o(tbuf_addr_lo),
    .way_o(tbuf_way_lo[0]),
    .v_o(tbuf_v_lo),
    .yumi_i(tbuf_yumi_li),
    .empty_o(tbuf_empty_lo),
    .full_o(tbuf_full_lo),
    .bypass_addr_i(addr_tl_r),
    .bypass_v_i(tbuf_bypass_v_li),
    .bypass_track_o(bypass_track_lo)
  );


  bsg_decode_num_out_p2
  tbuf_way_demux
  (
    .i(tbuf_way_lo[0]),
    .o(tbuf_way_decode)
  );


  bsg_decode_num_out_p4
  tbuf_wo_demux
  (
    .i(tbuf_addr_lo[3:2]),
    .o(tbuf_word_offset_decode)
  );


  bsg_mux_width_p32_els_p2
  ld_data_mux
  (
    .data_i(ld_data_v_r),
    .sel_i(tag_hit_way_id[0]),
    .data_o(ld_data_way_picked)
  );


  bsg_mux_width_p32_els_p1
  mux00
  (
    .data_i(ld_data_way_picked),
    .sel_i(addr_v_r[2]),
    .data_o(ld_data_offset_picked)
  );


  bsg_mux_segmented_segments_p4_segment_width_p8
  bypass_mux_segmented
  (
    .data0_i(ld_data_offset_picked),
    .data1_i(bypass_data_lo),
    .sel_i(bypass_mask_lo),
    .data_o(bypass_data_masked)
  );


  bsg_expand_bitmask_in_width_p4_expand_p8
  mask_v_expand
  (
    .i(mask_v_r),
    .o(expanded_mask_v)
  );


  bsg_mux_width_p8_els_p4
  \ld_data_sel_0_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1:0]),
    .data_o(\ld_data_sel_0_.byte_sel )
  );


  bsg_mux_width_p16_els_p2
  \ld_data_sel_1_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[1]),
    .data_o(\ld_data_sel_1_.byte_sel )
  );


  bsg_mux_width_p32_els_p1
  \ld_data_sel_2_.byte_mux 
  (
    .data_i(snoop_or_ld_data),
    .sel_i(addr_v_r[2]),
    .data_o(atomic_mem_data)
  );


  bsg_mux_width_p32_els_p3
  ld_data_size_mux
  (
    .data_i({ atomic_mem_data, ld_data_final_li_1__31_, ld_data_final_li_1__30_, ld_data_final_li_1__29_, ld_data_final_li_1__28_, ld_data_final_li_1__27_, ld_data_final_li_1__26_, ld_data_final_li_1__25_, ld_data_final_li_1__24_, ld_data_final_li_1__23_, ld_data_final_li_1__22_, ld_data_final_li_1__21_, ld_data_final_li_1__20_, ld_data_final_li_1__19_, ld_data_final_li_1__18_, ld_data_final_li_1__17_, ld_data_final_li_1__16_, \ld_data_sel_1_.byte_sel , ld_data_final_li_0__31_, ld_data_final_li_0__30_, ld_data_final_li_0__29_, ld_data_final_li_0__28_, ld_data_final_li_0__27_, ld_data_final_li_0__26_, ld_data_final_li_0__25_, ld_data_final_li_0__24_, ld_data_final_li_0__23_, ld_data_final_li_0__22_, ld_data_final_li_0__21_, ld_data_final_li_0__20_, ld_data_final_li_0__19_, ld_data_final_li_0__18_, ld_data_final_li_0__17_, ld_data_final_li_0__16_, ld_data_final_li_0__15_, ld_data_final_li_0__14_, ld_data_final_li_0__13_, ld_data_final_li_0__12_, ld_data_final_li_0__11_, ld_data_final_li_0__10_, ld_data_final_li_0__9_, ld_data_final_li_0__8_, \ld_data_sel_0_.byte_sel  }),
    .sel_i(decode_v_r[20:19]),
    .data_o(ld_data_final_lo)
  );

  assign N477 = (N476)? lock_v_r[0] : 
                (N1)? lock_v_r[1] : 1'b0;
  assign N479 = (N478)? valid_v_r[0] : 
                (N1)? valid_v_r[1] : 1'b0;
  assign N481 = (N480)? tag_v_r[17] : 
                (N1)? tag_v_r[35] : 1'b0;
  assign N482 = (N480)? tag_v_r[16] : 
                (N1)? tag_v_r[34] : 1'b0;
  assign N483 = (N480)? tag_v_r[15] : 
                (N1)? tag_v_r[33] : 1'b0;
  assign N484 = (N480)? tag_v_r[14] : 
                (N1)? tag_v_r[32] : 1'b0;
  assign N485 = (N480)? tag_v_r[13] : 
                (N1)? tag_v_r[31] : 1'b0;
  assign N486 = (N480)? tag_v_r[12] : 
                (N1)? tag_v_r[30] : 1'b0;
  assign N487 = (N480)? tag_v_r[11] : 
                (N1)? tag_v_r[29] : 1'b0;
  assign N488 = (N480)? tag_v_r[10] : 
                (N1)? tag_v_r[28] : 1'b0;
  assign N489 = (N480)? tag_v_r[9] : 
                (N1)? tag_v_r[27] : 1'b0;
  assign N490 = (N480)? tag_v_r[8] : 
                (N1)? tag_v_r[26] : 1'b0;
  assign N491 = (N480)? tag_v_r[7] : 
                (N1)? tag_v_r[25] : 1'b0;
  assign N492 = (N480)? tag_v_r[6] : 
                (N1)? tag_v_r[24] : 1'b0;
  assign N493 = (N480)? tag_v_r[5] : 
                (N1)? tag_v_r[23] : 1'b0;
  assign N494 = (N480)? tag_v_r[4] : 
                (N1)? tag_v_r[22] : 1'b0;
  assign N495 = (N480)? tag_v_r[3] : 
                (N1)? tag_v_r[21] : 1'b0;
  assign N496 = (N480)? tag_v_r[2] : 
                (N1)? tag_v_r[20] : 1'b0;
  assign N497 = (N480)? tag_v_r[1] : 
                (N1)? tag_v_r[19] : 1'b0;
  assign N498 = (N480)? tag_v_r[0] : 
                (N1)? tag_v_r[18] : 1'b0;

  bsg_decode_num_out_p2
  addr_way_demux
  (
    .i(cache_pkt_i[46]),
    .o(addr_way_decode)
  );


  bsg_lru_pseudo_tree_decode_ways_p2
  plru_decode
  (
    .way_id_i(tag_hit_way_id[0]),
    .data_o(plru_decode_data_lo[0]),
    .mask_o(plru_decode_mask_lo[0])
  );

  assign { N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294 } = data_v_r + atomic_mem_data;
  assign N67 = (N3)? 1'b1 : 
               (N71)? 1'b1 : 
               (N66)? 1'b0 : 1'b0;
  assign N3 = tl_we;
  assign N68 = (N3)? v_i : 
               (N71)? 1'b0 : 1'b0;
  assign N69 = (N3)? v_i : 
               (N71)? 1'b0 : 
               (N66)? 1'b0 : 1'b0;
  assign N75 = (N4)? 1'b1 : 
               (N2)? 1'b0 : 1'b0;
  assign N4 = v_we_o;
  assign N76 = (N4)? v_tl_r : 
               (N2)? 1'b0 : 1'b0;
  assign N77 = (N4)? v_tl_r : 
               (N2)? 1'b0 : 1'b0;
  assign N78 = (N5)? 1'b0 : 
               (N80)? v_tl_r : 
               (N74)? 1'b0 : 1'b0;
  assign N5 = N72;
  assign N86 = (N6)? N84 : 
               (N83)? N85 : 1'b0;
  assign N6 = decode[17];
  assign N90 = (N7)? N88 : 
               (N87)? N89 : 1'b0;
  assign N7 = decode_tl_r[17];
  assign N95 = (N8)? N93 : 
               (N92)? N94 : 1'b0;
  assign N8 = N91;
  assign N115 = (N9)? N114 : 
                (N10)? 1'b1 : 1'b0;
  assign N9 = N111;
  assign N10 = N110;
  assign N120 = (N11)? N119 : 
                (N12)? 1'b0 : 1'b0;
  assign N11 = N117;
  assign N12 = N116;
  assign sbuf_data_mem_w_mask[3:0] = (N13)? { N122, N123, N124, N125 } : 
                                     (N121)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = sbuf_way_decode[0];
  assign sbuf_data_mem_w_mask[7:4] = (N14)? { N127, N128, N129, N130 } : 
                                     (N126)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = sbuf_way_decode[1];
  assign { N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328 } = (N15)? data_v_r : 
                                                                                                                                                                                                              (N327)? atomic_mem_data : 1'b0;
  assign N15 = N326;
  assign { N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362 } = (N16)? data_v_r : 
                                                                                                                                                                                                              (N361)? atomic_mem_data : 1'b0;
  assign N16 = N360;
  assign { N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396 } = (N17)? data_v_r : 
                                                                                                                                                                                                              (N395)? atomic_mem_data : 1'b0;
  assign N17 = N394;
  assign { N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430 } = (N18)? data_v_r : 
                                                                                                                                                                                                              (N429)? atomic_mem_data : 1'b0;
  assign N18 = N428;
  assign atomic_alu_result = (N19)? data_v_r : 
                             (N20)? { N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229 } : 
                             (N21)? { N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261 } : 
                             (N22)? { N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293 } : 
                             (N23)? { N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294 } : 
                             (N24)? { N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328 } : 
                             (N25)? { N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362 } : 
                             (N26)? { N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396 } : 
                             (N27)? { N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430 } : 
                             (N28)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                             (N29)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N19 = N137;
  assign N20 = N144;
  assign N21 = N150;
  assign N22 = N156;
  assign N23 = N162;
  assign N24 = N169;
  assign N25 = N176;
  assign N26 = N184;
  assign N27 = N190;
  assign N28 = N132;
  assign N29 = N197;
  assign \sbuf_in_sel_2_.slice_data  = (N30)? atomic_alu_result : 
                                       (N463)? data_v_r : 1'b0;
  assign N30 = N462;
  assign { sbuf_entry_li_data__31_, sbuf_entry_li_data__30_, sbuf_entry_li_data__29_, sbuf_entry_li_data__28_, sbuf_entry_li_data__27_, sbuf_entry_li_data__26_, sbuf_entry_li_data__25_, sbuf_entry_li_data__24_, sbuf_entry_li_data__23_, sbuf_entry_li_data__22_, sbuf_entry_li_data__21_, sbuf_entry_li_data__20_, sbuf_entry_li_data__19_, sbuf_entry_li_data__18_, sbuf_entry_li_data__17_, sbuf_entry_li_data__16_, sbuf_entry_li_data__15_, sbuf_entry_li_data__14_, sbuf_entry_li_data__13_, sbuf_entry_li_data__12_, sbuf_entry_li_data__11_, sbuf_entry_li_data__10_, sbuf_entry_li_data__9_, sbuf_entry_li_data__8_, sbuf_entry_li_data__7_, sbuf_entry_li_data__6_, sbuf_entry_li_data__5_, sbuf_entry_li_data__4_, sbuf_entry_li_data__3_, sbuf_entry_li_data__2_, sbuf_entry_li_data__1_, sbuf_entry_li_data__0_, sbuf_entry_li_mask__3_, sbuf_entry_li_mask__2_, sbuf_entry_li_mask__1_, sbuf_entry_li_mask__0_ } = (N31)? { data_v_r, mask_v_r } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N465)? { sbuf_data_in, sbuf_mask_in } : 1'b0;
  assign N31 = N464;
  assign tbuf_track_mem_w_mask[3:0] = (N32)? tbuf_word_offset_decode : 
                                      (N466)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = tbuf_way_decode[0];
  assign tbuf_track_mem_w_mask[7:4] = (N33)? tbuf_word_offset_decode : 
                                      (N467)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N33 = tbuf_way_decode[1];
  assign snoop_or_ld_data = (N34)? snoop_word_lo : 
                            (N35)? bypass_data_masked : 1'b0;
  assign N34 = select_snoop_data_r_lo;
  assign N35 = N468;
  assign { N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499 } = (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N477, N479 } : 
                                                                                                                                                                                                              (N532)? { 1'b0, 1'b0, 1'b0, 1'b0, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, addr_v_r[9:4], 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                              (N535)? ld_data_masked : 
                                                                                                                                                                                                              (N475)? ld_data_final_lo : 1'b0;
  assign N36 = N470;
  assign data_o = (N37)? { N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499 } : 
                  (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N37 = retval_op_v;
  assign N38 = N469;
  assign N538 = (N39)? miss_done_lo : 
                (N40)? 1'b1 : 1'b0;
  assign N39 = N537;
  assign N40 = N536;
  assign v_we_o = (N41)? N540 : 
                  (N42)? 1'b1 : 1'b0;
  assign N41 = v_v_r;
  assign N42 = N539;
  assign N544 = (N43)? N543 : 
                (N44)? 1'b1 : 1'b0;
  assign N43 = N542;
  assign N44 = N541;
  assign N546 = (N45)? v_we_o : 
                (N46)? 1'b1 : 1'b0;
  assign N45 = v_tl_r;
  assign N46 = N545;
  assign tag_mem_w_li = (N47)? N549 : 
                        (N48)? tagst_write_en : 1'b0;
  assign N47 = N548;
  assign N48 = N547;
  assign { N559, N558, N557, N556, N555, N554 } = (N49)? addr_tl_r[9:4] : 
                                                  (N561)? miss_tag_mem_addr_lo : 
                                                  (N553)? cache_pkt_i[45:40] : 1'b0;
  assign N49 = recover_lo;
  assign tag_mem_addr_li = (N50)? { N559, N558, N557, N556, N555, N554 } : 
                           (N51)? cache_pkt_i[45:40] : 1'b0;
  assign N50 = N551;
  assign N51 = N550;
  assign tag_mem_data_li = (N50)? miss_tag_mem_data_lo : 
                           (N51)? { cache_pkt_i[35:34], cache_pkt_i[21:4], cache_pkt_i[35:34], cache_pkt_i[21:4] } : 1'b0;
  assign tag_mem_w_mask_li = (N50)? miss_tag_mem_w_mask_lo : 
                             (N51)? { addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode[1:1], addr_way_decode, addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0], addr_way_decode[0:0] } : 1'b0;
  assign data_mem_data_li = (N52)? dma_data_mem_data_lo : 
                            (N53)? { sbuf_entry_lo[36:5], sbuf_entry_lo[36:5] } : 1'b0;
  assign N52 = dma_data_mem_w_lo;
  assign N53 = N562;
  assign data_mem_addr_li = (N49)? addr_tl_r[9:2] : 
                            (N567)? dma_data_mem_addr_lo : 
                            (N570)? cache_pkt_i[45:38] : 
                            (N566)? sbuf_entry_lo[46:39] : 1'b0;
  assign data_mem_w_mask_li = (N52)? dma_data_mem_w_mask_lo : 
                              (N53)? sbuf_data_mem_w_mask : 1'b0;
  assign track_mem_w_li = (N54)? miss_track_mem_w_lo : 
                          (N55)? N571 : 1'b0;
  assign N54 = miss_track_mem_v_lo;
  assign N55 = N641;
  assign track_mem_data_li = (N54)? miss_track_mem_data_lo : 
                             (N55)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 1'b0;
  assign track_mem_w_mask_li = (N54)? miss_track_mem_w_mask_lo : 
                               (N55)? tbuf_track_mem_w_mask : 1'b0;
  assign track_mem_addr_li = (N49)? addr_tl_r[9:4] : 
                             (N576)? miss_track_mem_addr_lo : 
                             (N579)? cache_pkt_i[45:40] : 
                             (N575)? tbuf_addr_lo[9:4] : 1'b0;
  assign { N592, N591, N590 } = (N56)? { 1'b0, 1'b0, 1'b0 } : 
                                (N585)? { N586, N587, plru_decode_data_lo[0:0] } : 1'b0;
  assign N56 = N584;
  assign { N595, N594, N593 } = (N56)? { 1'b1, 1'b1, 1'b1 } : 
                                (N585)? { N588, N589, plru_decode_mask_lo[0:0] } : 1'b0;
  assign stat_mem_v_li = (N57)? miss_stat_mem_v_lo : 
                         (N58)? N582 : 1'b0;
  assign N57 = N581;
  assign N58 = N580;
  assign stat_mem_w_li = (N57)? miss_stat_mem_w_lo : 
                         (N58)? N583 : 1'b0;
  assign stat_mem_addr_li = (N57)? miss_stat_mem_addr_lo : 
                            (N58)? addr_v_r[9:4] : 1'b0;
  assign stat_mem_data_li = (N57)? miss_stat_mem_data_lo : 
                            (N58)? { N592, N591, N590 } : 1'b0;
  assign stat_mem_w_mask_li = (N57)? miss_stat_mem_w_mask_lo : 
                              (N58)? { N595, N594, N593 } : 1'b0;
  assign sbuf_entry_li_way_id__0_ = (N59)? chosen_way_lo[0] : 
                                    (N60)? tag_hit_way_id[0] : 1'b0;
  assign N59 = N597;
  assign N60 = N596;
  assign tbuf_way_li[0] = (N61)? chosen_way_lo[0] : 
                          (N62)? tag_hit_way_id[0] : 1'b0;
  assign N61 = N599;
  assign N62 = N598;
  assign N600 = ~decode_v_r[0];
  assign N601 = N63 & N600;
  assign N63 = ~decode_v_r[1];
  assign N131 = N64 & N601;
  assign N64 = ~decode_v_r[3];
  assign N65 = sbuf_hazard | tl_we;
  assign N66 = ~N65;
  assign N70 = ~tl_we;
  assign N71 = sbuf_hazard & N70;
  assign N72 = reset_i;
  assign N73 = v_we_o | N72;
  assign N74 = ~N73;
  assign N79 = ~N72;
  assign N80 = v_we_o & N79;
  assign tag_hit_v[0] = N81 & valid_v_r[0];
  assign tag_hit_v[1] = N82 & valid_v_r[1];
  assign N83 = ~decode[17];
  assign N84 = ~N604;
  assign N604 = N603 & cache_pkt_i[0];
  assign N603 = N602 & cache_pkt_i[1];
  assign N602 = cache_pkt_i[3] & cache_pkt_i[2];
  assign N85 = ~decode[20];
  assign partial_st = decode[15] & N86;
  assign N87 = ~decode_tl_r[17];
  assign N88 = ~N607;
  assign N607 = N606 & mask_tl_r[0];
  assign N606 = N605 & mask_tl_r[1];
  assign N605 = mask_tl_r[3] & mask_tl_r[2];
  assign N89 = ~decode_tl_r[20];
  assign partial_st_tl = decode_tl_r[15] & N90;
  assign N91 = decode_v_r[17];
  assign N92 = ~N91;
  assign N93 = ~N610;
  assign N610 = N609 & mask_v_r[0];
  assign N609 = N608 & mask_v_r[1];
  assign N608 = mask_v_r[3] & mask_v_r[2];
  assign N94 = ~decode_v_r[20];
  assign partial_st_v = decode_v_r[15] & N95;
  assign ld_st_amo_tag_miss = N612 & N613;
  assign N612 = N611 | decode_v_r[4];
  assign N611 = decode_v_r[16] | decode_v_r[15];
  assign N613 = ~tag_hit_found;
  assign N96 = ~tag_hit_way_id[0];
  assign N101 = ~addr_v_r[2];
  assign N102 = ~addr_v_r[3];
  assign N103 = N101 & N102;
  assign N104 = N101 & addr_v_r[3];
  assign N105 = addr_v_r[2] & N102;
  assign N106 = addr_v_r[2] & addr_v_r[3];
  assign track_miss = N616 & N618;
  assign N616 = N615 & tag_hit_found;
  assign N615 = N614 | partial_st_v;
  assign N614 = decode_v_r[16] | decode_v_r[4];
  assign N618 = ~N617;
  assign N617 = N107 | bypass_track_lo;
  assign N108 = ~addr_v_r[10];
  assign tagfl_hit = decode_v_r[13] & N109;
  assign aflinv_hit = N620 & tag_hit_found;
  assign N620 = N619 | decode_v_r[8];
  assign N619 = decode_v_r[10] | decode_v_r[9];
  assign N110 = ~tag_hit_found;
  assign N111 = tag_hit_found;
  assign N112 = ~tag_hit_way_id[0];
  assign N114 = ~N113;
  assign alock_miss = decode_v_r[7] & N115;
  assign N116 = ~tag_hit_found;
  assign N117 = tag_hit_found;
  assign N118 = ~tag_hit_way_id[0];
  assign aunlock_hit = decode_v_r[6] & N120;
  assign miss_v = N622 & N627;
  assign N622 = N621 & v_v_r;
  assign N621 = ~decode_v_r[14];
  assign N627 = N626 | aunlock_hit;
  assign N626 = N625 | alock_miss;
  assign N625 = N624 | aflinv_hit;
  assign N624 = N623 | tagfl_hit;
  assign N623 = ld_st_amo_tag_miss | track_miss;
  assign retval_op_v = N629 | decode_v_r[4];
  assign N629 = N628 | decode_v_r[11];
  assign N628 = decode_v_r[16] | decode_v_r[12];
  assign _1_net_ = v_o & yumi_i;
  assign N121 = ~sbuf_way_decode[0];
  assign N122 = sbuf_expand_mask[3] & sbuf_entry_lo[4];
  assign N123 = sbuf_expand_mask[2] & sbuf_entry_lo[3];
  assign N124 = sbuf_expand_mask[1] & sbuf_entry_lo[2];
  assign N125 = sbuf_expand_mask[0] & sbuf_entry_lo[1];
  assign N126 = ~sbuf_way_decode[1];
  assign N127 = sbuf_expand_mask[3] & sbuf_entry_lo[4];
  assign N128 = sbuf_expand_mask[2] & sbuf_entry_lo[3];
  assign N129 = sbuf_expand_mask[1] & sbuf_entry_lo[2];
  assign N130 = sbuf_expand_mask[0] & sbuf_entry_lo[1];
  assign N132 = ~N131;
  assign N137 = ~N136;
  assign N138 = ~decode_v_r[1];
  assign N139 = ~decode_v_r[0];
  assign N144 = ~N143;
  assign N145 = ~decode_v_r[2];
  assign N150 = ~N149;
  assign N151 = ~decode_v_r[1];
  assign N156 = ~N155;
  assign N157 = ~decode_v_r[0];
  assign N162 = ~N161;
  assign N163 = ~decode_v_r[2];
  assign N164 = ~decode_v_r[0];
  assign N169 = ~N168;
  assign N170 = ~decode_v_r[2];
  assign N171 = ~decode_v_r[1];
  assign N176 = ~N175;
  assign N177 = ~decode_v_r[2];
  assign N178 = ~decode_v_r[1];
  assign N179 = ~decode_v_r[0];
  assign N184 = ~N183;
  assign N185 = ~decode_v_r[3];
  assign N190 = ~N189;
  assign N197 = N192 | N630;
  assign N630 = N194 | N196;
  assign N198 = data_v_r[31] & atomic_mem_data[31];
  assign N199 = data_v_r[30] & atomic_mem_data[30];
  assign N200 = data_v_r[29] & atomic_mem_data[29];
  assign N201 = data_v_r[28] & atomic_mem_data[28];
  assign N202 = data_v_r[27] & atomic_mem_data[27];
  assign N203 = data_v_r[26] & atomic_mem_data[26];
  assign N204 = data_v_r[25] & atomic_mem_data[25];
  assign N205 = data_v_r[24] & atomic_mem_data[24];
  assign N206 = data_v_r[23] & atomic_mem_data[23];
  assign N207 = data_v_r[22] & atomic_mem_data[22];
  assign N208 = data_v_r[21] & atomic_mem_data[21];
  assign N209 = data_v_r[20] & atomic_mem_data[20];
  assign N210 = data_v_r[19] & atomic_mem_data[19];
  assign N211 = data_v_r[18] & atomic_mem_data[18];
  assign N212 = data_v_r[17] & atomic_mem_data[17];
  assign N213 = data_v_r[16] & atomic_mem_data[16];
  assign N214 = data_v_r[15] & atomic_mem_data[15];
  assign N215 = data_v_r[14] & atomic_mem_data[14];
  assign N216 = data_v_r[13] & atomic_mem_data[13];
  assign N217 = data_v_r[12] & atomic_mem_data[12];
  assign N218 = data_v_r[11] & atomic_mem_data[11];
  assign N219 = data_v_r[10] & atomic_mem_data[10];
  assign N220 = data_v_r[9] & atomic_mem_data[9];
  assign N221 = data_v_r[8] & atomic_mem_data[8];
  assign N222 = data_v_r[7] & atomic_mem_data[7];
  assign N223 = data_v_r[6] & atomic_mem_data[6];
  assign N224 = data_v_r[5] & atomic_mem_data[5];
  assign N225 = data_v_r[4] & atomic_mem_data[4];
  assign N226 = data_v_r[3] & atomic_mem_data[3];
  assign N227 = data_v_r[2] & atomic_mem_data[2];
  assign N228 = data_v_r[1] & atomic_mem_data[1];
  assign N229 = data_v_r[0] & atomic_mem_data[0];
  assign N230 = data_v_r[31] | atomic_mem_data[31];
  assign N231 = data_v_r[30] | atomic_mem_data[30];
  assign N232 = data_v_r[29] | atomic_mem_data[29];
  assign N233 = data_v_r[28] | atomic_mem_data[28];
  assign N234 = data_v_r[27] | atomic_mem_data[27];
  assign N235 = data_v_r[26] | atomic_mem_data[26];
  assign N236 = data_v_r[25] | atomic_mem_data[25];
  assign N237 = data_v_r[24] | atomic_mem_data[24];
  assign N238 = data_v_r[23] | atomic_mem_data[23];
  assign N239 = data_v_r[22] | atomic_mem_data[22];
  assign N240 = data_v_r[21] | atomic_mem_data[21];
  assign N241 = data_v_r[20] | atomic_mem_data[20];
  assign N242 = data_v_r[19] | atomic_mem_data[19];
  assign N243 = data_v_r[18] | atomic_mem_data[18];
  assign N244 = data_v_r[17] | atomic_mem_data[17];
  assign N245 = data_v_r[16] | atomic_mem_data[16];
  assign N246 = data_v_r[15] | atomic_mem_data[15];
  assign N247 = data_v_r[14] | atomic_mem_data[14];
  assign N248 = data_v_r[13] | atomic_mem_data[13];
  assign N249 = data_v_r[12] | atomic_mem_data[12];
  assign N250 = data_v_r[11] | atomic_mem_data[11];
  assign N251 = data_v_r[10] | atomic_mem_data[10];
  assign N252 = data_v_r[9] | atomic_mem_data[9];
  assign N253 = data_v_r[8] | atomic_mem_data[8];
  assign N254 = data_v_r[7] | atomic_mem_data[7];
  assign N255 = data_v_r[6] | atomic_mem_data[6];
  assign N256 = data_v_r[5] | atomic_mem_data[5];
  assign N257 = data_v_r[4] | atomic_mem_data[4];
  assign N258 = data_v_r[3] | atomic_mem_data[3];
  assign N259 = data_v_r[2] | atomic_mem_data[2];
  assign N260 = data_v_r[1] | atomic_mem_data[1];
  assign N261 = data_v_r[0] | atomic_mem_data[0];
  assign N262 = data_v_r[31] ^ atomic_mem_data[31];
  assign N263 = data_v_r[30] ^ atomic_mem_data[30];
  assign N264 = data_v_r[29] ^ atomic_mem_data[29];
  assign N265 = data_v_r[28] ^ atomic_mem_data[28];
  assign N266 = data_v_r[27] ^ atomic_mem_data[27];
  assign N267 = data_v_r[26] ^ atomic_mem_data[26];
  assign N268 = data_v_r[25] ^ atomic_mem_data[25];
  assign N269 = data_v_r[24] ^ atomic_mem_data[24];
  assign N270 = data_v_r[23] ^ atomic_mem_data[23];
  assign N271 = data_v_r[22] ^ atomic_mem_data[22];
  assign N272 = data_v_r[21] ^ atomic_mem_data[21];
  assign N273 = data_v_r[20] ^ atomic_mem_data[20];
  assign N274 = data_v_r[19] ^ atomic_mem_data[19];
  assign N275 = data_v_r[18] ^ atomic_mem_data[18];
  assign N276 = data_v_r[17] ^ atomic_mem_data[17];
  assign N277 = data_v_r[16] ^ atomic_mem_data[16];
  assign N278 = data_v_r[15] ^ atomic_mem_data[15];
  assign N279 = data_v_r[14] ^ atomic_mem_data[14];
  assign N280 = data_v_r[13] ^ atomic_mem_data[13];
  assign N281 = data_v_r[12] ^ atomic_mem_data[12];
  assign N282 = data_v_r[11] ^ atomic_mem_data[11];
  assign N283 = data_v_r[10] ^ atomic_mem_data[10];
  assign N284 = data_v_r[9] ^ atomic_mem_data[9];
  assign N285 = data_v_r[8] ^ atomic_mem_data[8];
  assign N286 = data_v_r[7] ^ atomic_mem_data[7];
  assign N287 = data_v_r[6] ^ atomic_mem_data[6];
  assign N288 = data_v_r[5] ^ atomic_mem_data[5];
  assign N289 = data_v_r[4] ^ atomic_mem_data[4];
  assign N290 = data_v_r[3] ^ atomic_mem_data[3];
  assign N291 = data_v_r[2] ^ atomic_mem_data[2];
  assign N292 = data_v_r[1] ^ atomic_mem_data[1];
  assign N293 = data_v_r[0] ^ atomic_mem_data[0];
  assign N327 = ~N326;
  assign N361 = ~N360;
  assign N395 = ~N394;
  assign N429 = ~N428;
  assign N462 = decode_v_r[4];
  assign N463 = ~N462;
  assign N464 = decode_v_r[17];
  assign N465 = ~N464;
  assign N466 = ~tbuf_way_decode[0];
  assign N467 = ~tbuf_way_decode[1];
  assign N468 = ~select_snoop_data_r_lo;
  assign ld_data_masked[31] = snoop_or_ld_data[31] & expanded_mask_v[31];
  assign ld_data_masked[30] = snoop_or_ld_data[30] & expanded_mask_v[30];
  assign ld_data_masked[29] = snoop_or_ld_data[29] & expanded_mask_v[29];
  assign ld_data_masked[28] = snoop_or_ld_data[28] & expanded_mask_v[28];
  assign ld_data_masked[27] = snoop_or_ld_data[27] & expanded_mask_v[27];
  assign ld_data_masked[26] = snoop_or_ld_data[26] & expanded_mask_v[26];
  assign ld_data_masked[25] = snoop_or_ld_data[25] & expanded_mask_v[25];
  assign ld_data_masked[24] = snoop_or_ld_data[24] & expanded_mask_v[24];
  assign ld_data_masked[23] = snoop_or_ld_data[23] & expanded_mask_v[23];
  assign ld_data_masked[22] = snoop_or_ld_data[22] & expanded_mask_v[22];
  assign ld_data_masked[21] = snoop_or_ld_data[21] & expanded_mask_v[21];
  assign ld_data_masked[20] = snoop_or_ld_data[20] & expanded_mask_v[20];
  assign ld_data_masked[19] = snoop_or_ld_data[19] & expanded_mask_v[19];
  assign ld_data_masked[18] = snoop_or_ld_data[18] & expanded_mask_v[18];
  assign ld_data_masked[17] = snoop_or_ld_data[17] & expanded_mask_v[17];
  assign ld_data_masked[16] = snoop_or_ld_data[16] & expanded_mask_v[16];
  assign ld_data_masked[15] = snoop_or_ld_data[15] & expanded_mask_v[15];
  assign ld_data_masked[14] = snoop_or_ld_data[14] & expanded_mask_v[14];
  assign ld_data_masked[13] = snoop_or_ld_data[13] & expanded_mask_v[13];
  assign ld_data_masked[12] = snoop_or_ld_data[12] & expanded_mask_v[12];
  assign ld_data_masked[11] = snoop_or_ld_data[11] & expanded_mask_v[11];
  assign ld_data_masked[10] = snoop_or_ld_data[10] & expanded_mask_v[10];
  assign ld_data_masked[9] = snoop_or_ld_data[9] & expanded_mask_v[9];
  assign ld_data_masked[8] = snoop_or_ld_data[8] & expanded_mask_v[8];
  assign ld_data_masked[7] = snoop_or_ld_data[7] & expanded_mask_v[7];
  assign ld_data_masked[6] = snoop_or_ld_data[6] & expanded_mask_v[6];
  assign ld_data_masked[5] = snoop_or_ld_data[5] & expanded_mask_v[5];
  assign ld_data_masked[4] = snoop_or_ld_data[4] & expanded_mask_v[4];
  assign ld_data_masked[3] = snoop_or_ld_data[3] & expanded_mask_v[3];
  assign ld_data_masked[2] = snoop_or_ld_data[2] & expanded_mask_v[2];
  assign ld_data_masked[1] = snoop_or_ld_data[1] & expanded_mask_v[1];
  assign ld_data_masked[0] = snoop_or_ld_data[0] & expanded_mask_v[0];
  assign ld_data_final_li_0__31_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__30_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__29_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__28_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__27_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__26_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__25_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__24_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__23_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__22_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__21_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__20_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__19_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__18_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__17_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__16_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__15_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__14_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__13_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__12_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__11_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__10_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__9_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_0__8_ = decode_v_r[18] & \ld_data_sel_0_.byte_sel [7];
  assign ld_data_final_li_1__31_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__30_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__29_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__28_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__27_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__26_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__25_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__24_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__23_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__22_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__21_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__20_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__19_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__18_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__17_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign ld_data_final_li_1__16_ = decode_v_r[18] & \ld_data_sel_1_.byte_sel [15];
  assign N469 = ~retval_op_v;
  assign N470 = decode_v_r[12];
  assign N471 = decode_v_r[11];
  assign N472 = decode_v_r[17];
  assign N473 = N471 | N470;
  assign N474 = N472 | N473;
  assign N475 = ~N474;
  assign N476 = ~addr_v_r[10];
  assign N478 = ~addr_v_r[10];
  assign N480 = ~addr_v_r[10];
  assign N531 = ~N470;
  assign N532 = N471 & N531;
  assign N533 = ~N471;
  assign N534 = N531 & N533;
  assign N535 = N472 & N534;
  assign N536 = ~miss_v;
  assign N537 = miss_v;
  assign v_o = v_v_r & N538;
  assign N539 = ~v_v_r;
  assign N540 = v_o & yumi_i;
  assign sbuf_hazard = N634 & N636;
  assign N634 = sbuf_full_lo & N633;
  assign N633 = N631 & N632;
  assign N631 = v_o & yumi_i;
  assign N632 = decode_v_r[15] | decode_v_r[4];
  assign N636 = v_i & N635;
  assign N635 = decode[16] | decode[4];
  assign N541 = ~miss_v;
  assign N542 = miss_v;
  assign N543 = N646 & N647;
  assign N646 = N644 & N645;
  assign N644 = N642 & N643;
  assign N642 = N640 & N641;
  assign N640 = N638 & N639;
  assign N638 = ~N637;
  assign N637 = decode[14] & v_i;
  assign N639 = ~miss_tag_mem_v_lo;
  assign N641 = ~miss_track_mem_v_lo;
  assign N643 = ~dma_data_mem_v_lo;
  assign N645 = ~recover_lo;
  assign N647 = ~dma_evict_lo;
  assign tl_ready = N544 & N648;
  assign N648 = ~sbuf_hazard;
  assign N545 = ~v_tl_r;
  assign tl_we = tl_ready & N546;
  assign yumi_o = v_i & tl_we;
  assign tagst_write_en = decode[14] & yumi_o;
  assign tag_mem_v_li = N653 | N654;
  assign N653 = N652 | miss_tag_mem_v_lo;
  assign N652 = N649 | N651;
  assign N649 = decode[5] & yumi_o;
  assign N651 = N650 & v_tl_r;
  assign N650 = recover_lo & decode_tl_r[5];
  assign N654 = decode[14] & yumi_o;
  assign N547 = ~miss_v;
  assign N548 = miss_v;
  assign N549 = miss_tag_mem_v_lo & miss_tag_mem_w_lo;
  assign N550 = ~miss_v;
  assign N551 = miss_v;
  assign N552 = miss_tag_mem_v_lo | recover_lo;
  assign N553 = ~N552;
  assign N560 = ~recover_lo;
  assign N561 = miss_tag_mem_v_lo & N560;
  assign data_mem_v_li = N661 | N662;
  assign N661 = N660 | dma_data_mem_v_lo;
  assign N660 = N656 | N659;
  assign N656 = yumi_o & N655;
  assign N655 = decode[16] | decode[4];
  assign N659 = N657 & N658;
  assign N657 = v_tl_r & recover_lo;
  assign N658 = decode_tl_r[16] | decode_tl_r[4];
  assign N662 = sbuf_v_lo & sbuf_yumi_li;
  assign data_mem_w_li = dma_data_mem_w_lo | N663;
  assign N663 = sbuf_v_lo & sbuf_yumi_li;
  assign N562 = ~dma_data_mem_w_lo;
  assign N563 = N664 & yumi_o;
  assign N664 = decode[16] | decode[4];
  assign N564 = dma_data_mem_v_lo | recover_lo;
  assign N565 = N563 | N564;
  assign N566 = ~N565;
  assign N567 = dma_data_mem_v_lo & N560;
  assign N568 = ~dma_data_mem_v_lo;
  assign N569 = N560 & N568;
  assign N570 = N563 & N569;
  assign track_mem_v_li = N673 | N674;
  assign N673 = N672 | miss_track_mem_v_lo;
  assign N672 = N667 | N671;
  assign N667 = yumi_o & N666;
  assign N666 = N665 | partial_st;
  assign N665 = decode[16] | decode[4];
  assign N671 = N668 & N670;
  assign N668 = v_tl_r & recover_lo;
  assign N670 = N669 | partial_st_tl;
  assign N669 = decode_tl_r[16] | decode_tl_r[4];
  assign N674 = tbuf_v_lo & tbuf_yumi_li;
  assign N571 = tbuf_v_lo & tbuf_yumi_li;
  assign N572 = N676 & yumi_o;
  assign N676 = N675 | partial_st;
  assign N675 = decode[16] | decode[4];
  assign N573 = miss_track_mem_v_lo | recover_lo;
  assign N574 = N572 | N573;
  assign N575 = ~N574;
  assign N576 = miss_track_mem_v_lo & N560;
  assign N577 = ~miss_track_mem_v_lo;
  assign N578 = N560 & N577;
  assign N579 = N572 & N578;
  assign N580 = ~miss_v;
  assign N581 = miss_v;
  assign N582 = N680 & yumi_i;
  assign N680 = N679 & v_o;
  assign N679 = N678 | decode_v_r[4];
  assign N678 = N677 | decode_v_r[14];
  assign N677 = decode_v_r[15] | decode_v_r[16];
  assign N583 = N684 & yumi_i;
  assign N684 = N683 & v_o;
  assign N683 = N682 | decode_v_r[4];
  assign N682 = N681 | decode_v_r[14];
  assign N681 = decode_v_r[15] | decode_v_r[16];
  assign N584 = decode_v_r[14];
  assign N585 = ~N584;
  assign N586 = decode_v_r[15] | decode_v_r[4];
  assign N587 = decode_v_r[15] | decode_v_r[4];
  assign N588 = N685 & tag_hit_v[1];
  assign N685 = decode_v_r[15] | decode_v_r[4];
  assign N589 = N686 & tag_hit_v[0];
  assign N686 = decode_v_r[15] | decode_v_r[4];
  assign sbuf_v_li = N688 & yumi_i;
  assign N688 = N687 & v_o;
  assign N687 = decode_v_r[15] | decode_v_r[4];
  assign N596 = ~miss_v;
  assign N597 = miss_v;
  assign sbuf_yumi_li = N693 & N700;
  assign N693 = N692 & N643;
  assign N692 = sbuf_v_lo & N691;
  assign N691 = ~N690;
  assign N690 = N689 & yumi_o;
  assign N689 = decode[16] | decode[4];
  assign N700 = ~N699;
  assign N699 = N697 & N698;
  assign N697 = N695 & N696;
  assign N695 = v_tl_r & N694;
  assign N694 = decode_tl_r[16] | decode_tl_r[4];
  assign N696 = ~v_we_o;
  assign N698 = ~miss_v;
  assign sbuf_bypass_v_li = N702 & v_we_o;
  assign N702 = N701 & v_tl_r;
  assign N701 = decode_tl_r[16] | decode_tl_r[4];
  assign tbuf_v_li = N705 & yumi_i;
  assign N705 = N704 & v_o;
  assign N704 = decode_v_r[15] & N703;
  assign N703 = ~partial_st_v;
  assign N598 = ~miss_v;
  assign N599 = miss_v;
  assign tbuf_yumi_li = N711 & N718;
  assign N711 = N710 & N641;
  assign N710 = tbuf_v_lo & N709;
  assign N709 = ~N708;
  assign N708 = N707 & yumi_o;
  assign N707 = N706 | partial_st;
  assign N706 = decode[16] | decode[4];
  assign N718 = ~N717;
  assign N717 = N715 & N716;
  assign N715 = N714 & N696;
  assign N714 = v_tl_r & N713;
  assign N713 = N712 | partial_st_tl;
  assign N712 = decode_tl_r[16] | decode_tl_r[4];
  assign N716 = ~miss_v;
  assign tbuf_bypass_v_li = N721 & v_we_o;
  assign N721 = N720 & v_tl_r;
  assign N720 = N719 | partial_st_tl;
  assign N719 = decode_tl_r[16] | decode_tl_r[4];
  assign N2 = ~v_we_o;

  always @(posedge clk_i) begin
    if(reset_i) begin
      data_tl_r_31_sv2v_reg <= 1'b0;
      data_tl_r_30_sv2v_reg <= 1'b0;
      data_tl_r_29_sv2v_reg <= 1'b0;
      data_tl_r_28_sv2v_reg <= 1'b0;
      data_tl_r_27_sv2v_reg <= 1'b0;
      data_tl_r_26_sv2v_reg <= 1'b0;
      data_tl_r_25_sv2v_reg <= 1'b0;
      data_tl_r_24_sv2v_reg <= 1'b0;
      data_tl_r_23_sv2v_reg <= 1'b0;
      data_tl_r_22_sv2v_reg <= 1'b0;
      data_tl_r_21_sv2v_reg <= 1'b0;
      data_tl_r_20_sv2v_reg <= 1'b0;
      data_tl_r_19_sv2v_reg <= 1'b0;
      data_tl_r_18_sv2v_reg <= 1'b0;
      data_tl_r_17_sv2v_reg <= 1'b0;
      data_tl_r_16_sv2v_reg <= 1'b0;
      data_tl_r_15_sv2v_reg <= 1'b0;
      data_tl_r_14_sv2v_reg <= 1'b0;
      data_tl_r_13_sv2v_reg <= 1'b0;
      data_tl_r_12_sv2v_reg <= 1'b0;
      data_tl_r_11_sv2v_reg <= 1'b0;
      data_tl_r_10_sv2v_reg <= 1'b0;
      data_tl_r_9_sv2v_reg <= 1'b0;
      data_tl_r_8_sv2v_reg <= 1'b0;
      data_tl_r_7_sv2v_reg <= 1'b0;
      data_tl_r_6_sv2v_reg <= 1'b0;
      data_tl_r_5_sv2v_reg <= 1'b0;
      data_tl_r_4_sv2v_reg <= 1'b0;
      data_tl_r_3_sv2v_reg <= 1'b0;
      data_tl_r_2_sv2v_reg <= 1'b0;
      data_tl_r_1_sv2v_reg <= 1'b0;
      data_tl_r_0_sv2v_reg <= 1'b0;
      decode_tl_r_20_sv2v_reg <= 1'b0;
      decode_tl_r_19_sv2v_reg <= 1'b0;
      decode_tl_r_18_sv2v_reg <= 1'b0;
      decode_tl_r_17_sv2v_reg <= 1'b0;
      decode_tl_r_16_sv2v_reg <= 1'b0;
      decode_tl_r_15_sv2v_reg <= 1'b0;
      decode_tl_r_14_sv2v_reg <= 1'b0;
      decode_tl_r_13_sv2v_reg <= 1'b0;
      decode_tl_r_12_sv2v_reg <= 1'b0;
      decode_tl_r_11_sv2v_reg <= 1'b0;
      decode_tl_r_10_sv2v_reg <= 1'b0;
      decode_tl_r_9_sv2v_reg <= 1'b0;
      decode_tl_r_8_sv2v_reg <= 1'b0;
      decode_tl_r_7_sv2v_reg <= 1'b0;
      decode_tl_r_6_sv2v_reg <= 1'b0;
      decode_tl_r_5_sv2v_reg <= 1'b0;
      decode_tl_r_4_sv2v_reg <= 1'b0;
      decode_tl_r_3_sv2v_reg <= 1'b0;
      decode_tl_r_2_sv2v_reg <= 1'b0;
      decode_tl_r_1_sv2v_reg <= 1'b0;
      decode_tl_r_0_sv2v_reg <= 1'b0;
      mask_tl_r_3_sv2v_reg <= 1'b0;
      mask_tl_r_2_sv2v_reg <= 1'b0;
      mask_tl_r_1_sv2v_reg <= 1'b0;
      mask_tl_r_0_sv2v_reg <= 1'b0;
      addr_tl_r_27_sv2v_reg <= 1'b0;
      addr_tl_r_26_sv2v_reg <= 1'b0;
      addr_tl_r_25_sv2v_reg <= 1'b0;
      addr_tl_r_24_sv2v_reg <= 1'b0;
      addr_tl_r_23_sv2v_reg <= 1'b0;
      addr_tl_r_22_sv2v_reg <= 1'b0;
      addr_tl_r_21_sv2v_reg <= 1'b0;
      addr_tl_r_20_sv2v_reg <= 1'b0;
      addr_tl_r_19_sv2v_reg <= 1'b0;
      addr_tl_r_18_sv2v_reg <= 1'b0;
      addr_tl_r_17_sv2v_reg <= 1'b0;
      addr_tl_r_16_sv2v_reg <= 1'b0;
      addr_tl_r_15_sv2v_reg <= 1'b0;
      addr_tl_r_14_sv2v_reg <= 1'b0;
      addr_tl_r_13_sv2v_reg <= 1'b0;
      addr_tl_r_12_sv2v_reg <= 1'b0;
      addr_tl_r_11_sv2v_reg <= 1'b0;
      addr_tl_r_10_sv2v_reg <= 1'b0;
      addr_tl_r_9_sv2v_reg <= 1'b0;
      addr_tl_r_8_sv2v_reg <= 1'b0;
      addr_tl_r_7_sv2v_reg <= 1'b0;
      addr_tl_r_6_sv2v_reg <= 1'b0;
      addr_tl_r_5_sv2v_reg <= 1'b0;
      addr_tl_r_4_sv2v_reg <= 1'b0;
      addr_tl_r_3_sv2v_reg <= 1'b0;
      addr_tl_r_2_sv2v_reg <= 1'b0;
      addr_tl_r_1_sv2v_reg <= 1'b0;
      addr_tl_r_0_sv2v_reg <= 1'b0;
    end else if(N69) begin
      data_tl_r_31_sv2v_reg <= cache_pkt_i[35];
      data_tl_r_30_sv2v_reg <= cache_pkt_i[34];
      data_tl_r_29_sv2v_reg <= cache_pkt_i[33];
      data_tl_r_28_sv2v_reg <= cache_pkt_i[32];
      data_tl_r_27_sv2v_reg <= cache_pkt_i[31];
      data_tl_r_26_sv2v_reg <= cache_pkt_i[30];
      data_tl_r_25_sv2v_reg <= cache_pkt_i[29];
      data_tl_r_24_sv2v_reg <= cache_pkt_i[28];
      data_tl_r_23_sv2v_reg <= cache_pkt_i[27];
      data_tl_r_22_sv2v_reg <= cache_pkt_i[26];
      data_tl_r_21_sv2v_reg <= cache_pkt_i[25];
      data_tl_r_20_sv2v_reg <= cache_pkt_i[24];
      data_tl_r_19_sv2v_reg <= cache_pkt_i[23];
      data_tl_r_18_sv2v_reg <= cache_pkt_i[22];
      data_tl_r_17_sv2v_reg <= cache_pkt_i[21];
      data_tl_r_16_sv2v_reg <= cache_pkt_i[20];
      data_tl_r_15_sv2v_reg <= cache_pkt_i[19];
      data_tl_r_14_sv2v_reg <= cache_pkt_i[18];
      data_tl_r_13_sv2v_reg <= cache_pkt_i[17];
      data_tl_r_12_sv2v_reg <= cache_pkt_i[16];
      data_tl_r_11_sv2v_reg <= cache_pkt_i[15];
      data_tl_r_10_sv2v_reg <= cache_pkt_i[14];
      data_tl_r_9_sv2v_reg <= cache_pkt_i[13];
      data_tl_r_8_sv2v_reg <= cache_pkt_i[12];
      data_tl_r_7_sv2v_reg <= cache_pkt_i[11];
      data_tl_r_6_sv2v_reg <= cache_pkt_i[10];
      data_tl_r_5_sv2v_reg <= cache_pkt_i[9];
      data_tl_r_4_sv2v_reg <= cache_pkt_i[8];
      data_tl_r_3_sv2v_reg <= cache_pkt_i[7];
      data_tl_r_2_sv2v_reg <= cache_pkt_i[6];
      data_tl_r_1_sv2v_reg <= cache_pkt_i[5];
      data_tl_r_0_sv2v_reg <= cache_pkt_i[4];
      decode_tl_r_20_sv2v_reg <= decode[20];
      decode_tl_r_19_sv2v_reg <= decode[19];
      decode_tl_r_18_sv2v_reg <= decode[18];
      decode_tl_r_17_sv2v_reg <= decode[17];
      decode_tl_r_16_sv2v_reg <= decode[16];
      decode_tl_r_15_sv2v_reg <= decode[15];
      decode_tl_r_14_sv2v_reg <= decode[14];
      decode_tl_r_13_sv2v_reg <= decode[13];
      decode_tl_r_12_sv2v_reg <= decode[12];
      decode_tl_r_11_sv2v_reg <= decode[11];
      decode_tl_r_10_sv2v_reg <= decode[10];
      decode_tl_r_9_sv2v_reg <= decode[9];
      decode_tl_r_8_sv2v_reg <= decode[8];
      decode_tl_r_7_sv2v_reg <= decode[7];
      decode_tl_r_6_sv2v_reg <= decode[6];
      decode_tl_r_5_sv2v_reg <= decode[5];
      decode_tl_r_4_sv2v_reg <= decode[4];
      decode_tl_r_3_sv2v_reg <= decode[3];
      decode_tl_r_2_sv2v_reg <= decode[2];
      decode_tl_r_1_sv2v_reg <= decode[1];
      decode_tl_r_0_sv2v_reg <= decode[0];
      mask_tl_r_3_sv2v_reg <= cache_pkt_i[3];
      mask_tl_r_2_sv2v_reg <= cache_pkt_i[2];
      mask_tl_r_1_sv2v_reg <= cache_pkt_i[1];
      mask_tl_r_0_sv2v_reg <= cache_pkt_i[0];
      addr_tl_r_27_sv2v_reg <= cache_pkt_i[63];
      addr_tl_r_26_sv2v_reg <= cache_pkt_i[62];
      addr_tl_r_25_sv2v_reg <= cache_pkt_i[61];
      addr_tl_r_24_sv2v_reg <= cache_pkt_i[60];
      addr_tl_r_23_sv2v_reg <= cache_pkt_i[59];
      addr_tl_r_22_sv2v_reg <= cache_pkt_i[58];
      addr_tl_r_21_sv2v_reg <= cache_pkt_i[57];
      addr_tl_r_20_sv2v_reg <= cache_pkt_i[56];
      addr_tl_r_19_sv2v_reg <= cache_pkt_i[55];
      addr_tl_r_18_sv2v_reg <= cache_pkt_i[54];
      addr_tl_r_17_sv2v_reg <= cache_pkt_i[53];
      addr_tl_r_16_sv2v_reg <= cache_pkt_i[52];
      addr_tl_r_15_sv2v_reg <= cache_pkt_i[51];
      addr_tl_r_14_sv2v_reg <= cache_pkt_i[50];
      addr_tl_r_13_sv2v_reg <= cache_pkt_i[49];
      addr_tl_r_12_sv2v_reg <= cache_pkt_i[48];
      addr_tl_r_11_sv2v_reg <= cache_pkt_i[47];
      addr_tl_r_10_sv2v_reg <= cache_pkt_i[46];
      addr_tl_r_9_sv2v_reg <= cache_pkt_i[45];
      addr_tl_r_8_sv2v_reg <= cache_pkt_i[44];
      addr_tl_r_7_sv2v_reg <= cache_pkt_i[43];
      addr_tl_r_6_sv2v_reg <= cache_pkt_i[42];
      addr_tl_r_5_sv2v_reg <= cache_pkt_i[41];
      addr_tl_r_4_sv2v_reg <= cache_pkt_i[40];
      addr_tl_r_3_sv2v_reg <= cache_pkt_i[39];
      addr_tl_r_2_sv2v_reg <= cache_pkt_i[38];
      addr_tl_r_1_sv2v_reg <= cache_pkt_i[37];
      addr_tl_r_0_sv2v_reg <= cache_pkt_i[36];
    end 
    if(reset_i) begin
      v_tl_r_sv2v_reg <= 1'b0;
    end else if(N67) begin
      v_tl_r_sv2v_reg <= N68;
    end 
    if(N78) begin
      ld_data_v_r_63_sv2v_reg <= data_mem_data_lo[63];
      ld_data_v_r_62_sv2v_reg <= data_mem_data_lo[62];
      ld_data_v_r_61_sv2v_reg <= data_mem_data_lo[61];
      ld_data_v_r_60_sv2v_reg <= data_mem_data_lo[60];
      ld_data_v_r_59_sv2v_reg <= data_mem_data_lo[59];
      ld_data_v_r_58_sv2v_reg <= data_mem_data_lo[58];
      ld_data_v_r_57_sv2v_reg <= data_mem_data_lo[57];
      ld_data_v_r_56_sv2v_reg <= data_mem_data_lo[56];
      ld_data_v_r_55_sv2v_reg <= data_mem_data_lo[55];
      ld_data_v_r_54_sv2v_reg <= data_mem_data_lo[54];
      ld_data_v_r_53_sv2v_reg <= data_mem_data_lo[53];
      ld_data_v_r_52_sv2v_reg <= data_mem_data_lo[52];
      ld_data_v_r_51_sv2v_reg <= data_mem_data_lo[51];
      ld_data_v_r_50_sv2v_reg <= data_mem_data_lo[50];
      ld_data_v_r_49_sv2v_reg <= data_mem_data_lo[49];
      ld_data_v_r_48_sv2v_reg <= data_mem_data_lo[48];
      ld_data_v_r_47_sv2v_reg <= data_mem_data_lo[47];
      ld_data_v_r_46_sv2v_reg <= data_mem_data_lo[46];
      ld_data_v_r_45_sv2v_reg <= data_mem_data_lo[45];
      ld_data_v_r_44_sv2v_reg <= data_mem_data_lo[44];
      ld_data_v_r_43_sv2v_reg <= data_mem_data_lo[43];
      ld_data_v_r_42_sv2v_reg <= data_mem_data_lo[42];
      ld_data_v_r_41_sv2v_reg <= data_mem_data_lo[41];
      ld_data_v_r_40_sv2v_reg <= data_mem_data_lo[40];
      ld_data_v_r_39_sv2v_reg <= data_mem_data_lo[39];
      ld_data_v_r_38_sv2v_reg <= data_mem_data_lo[38];
      ld_data_v_r_37_sv2v_reg <= data_mem_data_lo[37];
      ld_data_v_r_36_sv2v_reg <= data_mem_data_lo[36];
      ld_data_v_r_35_sv2v_reg <= data_mem_data_lo[35];
      ld_data_v_r_34_sv2v_reg <= data_mem_data_lo[34];
      ld_data_v_r_33_sv2v_reg <= data_mem_data_lo[33];
      ld_data_v_r_32_sv2v_reg <= data_mem_data_lo[32];
      ld_data_v_r_31_sv2v_reg <= data_mem_data_lo[31];
      ld_data_v_r_30_sv2v_reg <= data_mem_data_lo[30];
      ld_data_v_r_29_sv2v_reg <= data_mem_data_lo[29];
      ld_data_v_r_28_sv2v_reg <= data_mem_data_lo[28];
      ld_data_v_r_27_sv2v_reg <= data_mem_data_lo[27];
      ld_data_v_r_26_sv2v_reg <= data_mem_data_lo[26];
      ld_data_v_r_25_sv2v_reg <= data_mem_data_lo[25];
      ld_data_v_r_24_sv2v_reg <= data_mem_data_lo[24];
      ld_data_v_r_23_sv2v_reg <= data_mem_data_lo[23];
      ld_data_v_r_22_sv2v_reg <= data_mem_data_lo[22];
      ld_data_v_r_21_sv2v_reg <= data_mem_data_lo[21];
      ld_data_v_r_20_sv2v_reg <= data_mem_data_lo[20];
      ld_data_v_r_19_sv2v_reg <= data_mem_data_lo[19];
      ld_data_v_r_18_sv2v_reg <= data_mem_data_lo[18];
      ld_data_v_r_17_sv2v_reg <= data_mem_data_lo[17];
      ld_data_v_r_16_sv2v_reg <= data_mem_data_lo[16];
      ld_data_v_r_15_sv2v_reg <= data_mem_data_lo[15];
      ld_data_v_r_14_sv2v_reg <= data_mem_data_lo[14];
      ld_data_v_r_13_sv2v_reg <= data_mem_data_lo[13];
      ld_data_v_r_12_sv2v_reg <= data_mem_data_lo[12];
      ld_data_v_r_11_sv2v_reg <= data_mem_data_lo[11];
      ld_data_v_r_10_sv2v_reg <= data_mem_data_lo[10];
      ld_data_v_r_9_sv2v_reg <= data_mem_data_lo[9];
      ld_data_v_r_8_sv2v_reg <= data_mem_data_lo[8];
      ld_data_v_r_7_sv2v_reg <= data_mem_data_lo[7];
      ld_data_v_r_6_sv2v_reg <= data_mem_data_lo[6];
      ld_data_v_r_5_sv2v_reg <= data_mem_data_lo[5];
      ld_data_v_r_4_sv2v_reg <= data_mem_data_lo[4];
      ld_data_v_r_3_sv2v_reg <= data_mem_data_lo[3];
      ld_data_v_r_2_sv2v_reg <= data_mem_data_lo[2];
      ld_data_v_r_1_sv2v_reg <= data_mem_data_lo[1];
      ld_data_v_r_0_sv2v_reg <= data_mem_data_lo[0];
    end 
    if(reset_i) begin
      v_v_r_sv2v_reg <= 1'b0;
    end else if(N75) begin
      v_v_r_sv2v_reg <= v_tl_r;
    end 
    if(reset_i) begin
      track_data_v_r_7_sv2v_reg <= 1'b0;
      track_data_v_r_6_sv2v_reg <= 1'b0;
      track_data_v_r_5_sv2v_reg <= 1'b0;
      track_data_v_r_4_sv2v_reg <= 1'b0;
      track_data_v_r_3_sv2v_reg <= 1'b0;
      track_data_v_r_2_sv2v_reg <= 1'b0;
      track_data_v_r_1_sv2v_reg <= 1'b0;
      track_data_v_r_0_sv2v_reg <= 1'b0;
      mask_v_r_0_sv2v_reg <= 1'b0;
      lock_v_r_1_sv2v_reg <= 1'b0;
      lock_v_r_0_sv2v_reg <= 1'b0;
      tag_v_r_35_sv2v_reg <= 1'b0;
      tag_v_r_34_sv2v_reg <= 1'b0;
      tag_v_r_33_sv2v_reg <= 1'b0;
      tag_v_r_32_sv2v_reg <= 1'b0;
      tag_v_r_31_sv2v_reg <= 1'b0;
      tag_v_r_30_sv2v_reg <= 1'b0;
      tag_v_r_29_sv2v_reg <= 1'b0;
      tag_v_r_28_sv2v_reg <= 1'b0;
      tag_v_r_27_sv2v_reg <= 1'b0;
      tag_v_r_26_sv2v_reg <= 1'b0;
      tag_v_r_25_sv2v_reg <= 1'b0;
      tag_v_r_24_sv2v_reg <= 1'b0;
      tag_v_r_23_sv2v_reg <= 1'b0;
      tag_v_r_22_sv2v_reg <= 1'b0;
      tag_v_r_21_sv2v_reg <= 1'b0;
      tag_v_r_20_sv2v_reg <= 1'b0;
      tag_v_r_19_sv2v_reg <= 1'b0;
      tag_v_r_18_sv2v_reg <= 1'b0;
      tag_v_r_17_sv2v_reg <= 1'b0;
      tag_v_r_16_sv2v_reg <= 1'b0;
      tag_v_r_15_sv2v_reg <= 1'b0;
      tag_v_r_14_sv2v_reg <= 1'b0;
      tag_v_r_13_sv2v_reg <= 1'b0;
      tag_v_r_12_sv2v_reg <= 1'b0;
      tag_v_r_11_sv2v_reg <= 1'b0;
    end else if(N76) begin
      track_data_v_r_7_sv2v_reg <= track_mem_data_lo[7];
      track_data_v_r_6_sv2v_reg <= track_mem_data_lo[6];
      track_data_v_r_5_sv2v_reg <= track_mem_data_lo[5];
      track_data_v_r_4_sv2v_reg <= track_mem_data_lo[4];
      track_data_v_r_3_sv2v_reg <= track_mem_data_lo[3];
      track_data_v_r_2_sv2v_reg <= track_mem_data_lo[2];
      track_data_v_r_1_sv2v_reg <= track_mem_data_lo[1];
      track_data_v_r_0_sv2v_reg <= track_mem_data_lo[0];
      mask_v_r_0_sv2v_reg <= mask_tl_r[0];
      lock_v_r_1_sv2v_reg <= tag_mem_data_lo[38];
      lock_v_r_0_sv2v_reg <= tag_mem_data_lo[18];
      tag_v_r_35_sv2v_reg <= tag_mem_data_lo[37];
      tag_v_r_34_sv2v_reg <= tag_mem_data_lo[36];
      tag_v_r_33_sv2v_reg <= tag_mem_data_lo[35];
      tag_v_r_32_sv2v_reg <= tag_mem_data_lo[34];
      tag_v_r_31_sv2v_reg <= tag_mem_data_lo[33];
      tag_v_r_30_sv2v_reg <= tag_mem_data_lo[32];
      tag_v_r_29_sv2v_reg <= tag_mem_data_lo[31];
      tag_v_r_28_sv2v_reg <= tag_mem_data_lo[30];
      tag_v_r_27_sv2v_reg <= tag_mem_data_lo[29];
      tag_v_r_26_sv2v_reg <= tag_mem_data_lo[28];
      tag_v_r_25_sv2v_reg <= tag_mem_data_lo[27];
      tag_v_r_24_sv2v_reg <= tag_mem_data_lo[26];
      tag_v_r_23_sv2v_reg <= tag_mem_data_lo[25];
      tag_v_r_22_sv2v_reg <= tag_mem_data_lo[24];
      tag_v_r_21_sv2v_reg <= tag_mem_data_lo[23];
      tag_v_r_20_sv2v_reg <= tag_mem_data_lo[22];
      tag_v_r_19_sv2v_reg <= tag_mem_data_lo[21];
      tag_v_r_18_sv2v_reg <= tag_mem_data_lo[20];
      tag_v_r_17_sv2v_reg <= tag_mem_data_lo[17];
      tag_v_r_16_sv2v_reg <= tag_mem_data_lo[16];
      tag_v_r_15_sv2v_reg <= tag_mem_data_lo[15];
      tag_v_r_14_sv2v_reg <= tag_mem_data_lo[14];
      tag_v_r_13_sv2v_reg <= tag_mem_data_lo[13];
      tag_v_r_12_sv2v_reg <= tag_mem_data_lo[12];
      tag_v_r_11_sv2v_reg <= tag_mem_data_lo[11];
    end 
    if(reset_i) begin
      mask_v_r_3_sv2v_reg <= 1'b0;
      mask_v_r_2_sv2v_reg <= 1'b0;
      mask_v_r_1_sv2v_reg <= 1'b0;
      decode_v_r_20_sv2v_reg <= 1'b0;
      decode_v_r_19_sv2v_reg <= 1'b0;
      decode_v_r_18_sv2v_reg <= 1'b0;
      decode_v_r_17_sv2v_reg <= 1'b0;
      decode_v_r_16_sv2v_reg <= 1'b0;
      decode_v_r_15_sv2v_reg <= 1'b0;
      decode_v_r_14_sv2v_reg <= 1'b0;
      decode_v_r_13_sv2v_reg <= 1'b0;
      decode_v_r_12_sv2v_reg <= 1'b0;
      decode_v_r_11_sv2v_reg <= 1'b0;
      decode_v_r_10_sv2v_reg <= 1'b0;
      decode_v_r_9_sv2v_reg <= 1'b0;
      decode_v_r_8_sv2v_reg <= 1'b0;
      decode_v_r_7_sv2v_reg <= 1'b0;
      decode_v_r_6_sv2v_reg <= 1'b0;
      decode_v_r_5_sv2v_reg <= 1'b0;
      decode_v_r_4_sv2v_reg <= 1'b0;
      decode_v_r_3_sv2v_reg <= 1'b0;
      decode_v_r_2_sv2v_reg <= 1'b0;
      decode_v_r_1_sv2v_reg <= 1'b0;
      decode_v_r_0_sv2v_reg <= 1'b0;
      addr_v_r_27_sv2v_reg <= 1'b0;
      addr_v_r_26_sv2v_reg <= 1'b0;
      addr_v_r_25_sv2v_reg <= 1'b0;
      addr_v_r_24_sv2v_reg <= 1'b0;
      addr_v_r_23_sv2v_reg <= 1'b0;
      addr_v_r_22_sv2v_reg <= 1'b0;
      addr_v_r_21_sv2v_reg <= 1'b0;
      addr_v_r_20_sv2v_reg <= 1'b0;
      addr_v_r_19_sv2v_reg <= 1'b0;
      addr_v_r_18_sv2v_reg <= 1'b0;
      addr_v_r_17_sv2v_reg <= 1'b0;
      addr_v_r_16_sv2v_reg <= 1'b0;
      addr_v_r_15_sv2v_reg <= 1'b0;
      addr_v_r_14_sv2v_reg <= 1'b0;
      addr_v_r_13_sv2v_reg <= 1'b0;
      addr_v_r_12_sv2v_reg <= 1'b0;
      addr_v_r_11_sv2v_reg <= 1'b0;
      addr_v_r_10_sv2v_reg <= 1'b0;
      addr_v_r_9_sv2v_reg <= 1'b0;
      addr_v_r_8_sv2v_reg <= 1'b0;
      addr_v_r_7_sv2v_reg <= 1'b0;
      addr_v_r_6_sv2v_reg <= 1'b0;
      addr_v_r_5_sv2v_reg <= 1'b0;
      addr_v_r_4_sv2v_reg <= 1'b0;
      addr_v_r_3_sv2v_reg <= 1'b0;
      addr_v_r_2_sv2v_reg <= 1'b0;
      addr_v_r_1_sv2v_reg <= 1'b0;
      addr_v_r_0_sv2v_reg <= 1'b0;
      data_v_r_31_sv2v_reg <= 1'b0;
      data_v_r_30_sv2v_reg <= 1'b0;
      data_v_r_29_sv2v_reg <= 1'b0;
      data_v_r_28_sv2v_reg <= 1'b0;
      data_v_r_27_sv2v_reg <= 1'b0;
      data_v_r_26_sv2v_reg <= 1'b0;
      data_v_r_25_sv2v_reg <= 1'b0;
      data_v_r_24_sv2v_reg <= 1'b0;
      data_v_r_23_sv2v_reg <= 1'b0;
      data_v_r_22_sv2v_reg <= 1'b0;
      data_v_r_21_sv2v_reg <= 1'b0;
      data_v_r_20_sv2v_reg <= 1'b0;
      data_v_r_19_sv2v_reg <= 1'b0;
      data_v_r_18_sv2v_reg <= 1'b0;
      data_v_r_17_sv2v_reg <= 1'b0;
      data_v_r_16_sv2v_reg <= 1'b0;
      data_v_r_15_sv2v_reg <= 1'b0;
      data_v_r_14_sv2v_reg <= 1'b0;
      data_v_r_13_sv2v_reg <= 1'b0;
      data_v_r_12_sv2v_reg <= 1'b0;
      data_v_r_11_sv2v_reg <= 1'b0;
      data_v_r_10_sv2v_reg <= 1'b0;
      data_v_r_9_sv2v_reg <= 1'b0;
      data_v_r_8_sv2v_reg <= 1'b0;
      data_v_r_7_sv2v_reg <= 1'b0;
      data_v_r_6_sv2v_reg <= 1'b0;
      data_v_r_5_sv2v_reg <= 1'b0;
      data_v_r_4_sv2v_reg <= 1'b0;
      data_v_r_3_sv2v_reg <= 1'b0;
      data_v_r_2_sv2v_reg <= 1'b0;
      data_v_r_1_sv2v_reg <= 1'b0;
      data_v_r_0_sv2v_reg <= 1'b0;
      valid_v_r_1_sv2v_reg <= 1'b0;
      valid_v_r_0_sv2v_reg <= 1'b0;
      tag_v_r_10_sv2v_reg <= 1'b0;
      tag_v_r_9_sv2v_reg <= 1'b0;
      tag_v_r_8_sv2v_reg <= 1'b0;
      tag_v_r_7_sv2v_reg <= 1'b0;
      tag_v_r_6_sv2v_reg <= 1'b0;
      tag_v_r_5_sv2v_reg <= 1'b0;
      tag_v_r_4_sv2v_reg <= 1'b0;
      tag_v_r_3_sv2v_reg <= 1'b0;
      tag_v_r_2_sv2v_reg <= 1'b0;
      tag_v_r_1_sv2v_reg <= 1'b0;
      tag_v_r_0_sv2v_reg <= 1'b0;
    end else if(N77) begin
      mask_v_r_3_sv2v_reg <= mask_tl_r[3];
      mask_v_r_2_sv2v_reg <= mask_tl_r[2];
      mask_v_r_1_sv2v_reg <= mask_tl_r[1];
      decode_v_r_20_sv2v_reg <= decode_tl_r[20];
      decode_v_r_19_sv2v_reg <= decode_tl_r[19];
      decode_v_r_18_sv2v_reg <= decode_tl_r[18];
      decode_v_r_17_sv2v_reg <= decode_tl_r[17];
      decode_v_r_16_sv2v_reg <= decode_tl_r[16];
      decode_v_r_15_sv2v_reg <= decode_tl_r[15];
      decode_v_r_14_sv2v_reg <= decode_tl_r[14];
      decode_v_r_13_sv2v_reg <= decode_tl_r[13];
      decode_v_r_12_sv2v_reg <= decode_tl_r[12];
      decode_v_r_11_sv2v_reg <= decode_tl_r[11];
      decode_v_r_10_sv2v_reg <= decode_tl_r[10];
      decode_v_r_9_sv2v_reg <= decode_tl_r[9];
      decode_v_r_8_sv2v_reg <= decode_tl_r[8];
      decode_v_r_7_sv2v_reg <= decode_tl_r[7];
      decode_v_r_6_sv2v_reg <= decode_tl_r[6];
      decode_v_r_5_sv2v_reg <= decode_tl_r[5];
      decode_v_r_4_sv2v_reg <= decode_tl_r[4];
      decode_v_r_3_sv2v_reg <= decode_tl_r[3];
      decode_v_r_2_sv2v_reg <= decode_tl_r[2];
      decode_v_r_1_sv2v_reg <= decode_tl_r[1];
      decode_v_r_0_sv2v_reg <= decode_tl_r[0];
      addr_v_r_27_sv2v_reg <= addr_tl_r[27];
      addr_v_r_26_sv2v_reg <= addr_tl_r[26];
      addr_v_r_25_sv2v_reg <= addr_tl_r[25];
      addr_v_r_24_sv2v_reg <= addr_tl_r[24];
      addr_v_r_23_sv2v_reg <= addr_tl_r[23];
      addr_v_r_22_sv2v_reg <= addr_tl_r[22];
      addr_v_r_21_sv2v_reg <= addr_tl_r[21];
      addr_v_r_20_sv2v_reg <= addr_tl_r[20];
      addr_v_r_19_sv2v_reg <= addr_tl_r[19];
      addr_v_r_18_sv2v_reg <= addr_tl_r[18];
      addr_v_r_17_sv2v_reg <= addr_tl_r[17];
      addr_v_r_16_sv2v_reg <= addr_tl_r[16];
      addr_v_r_15_sv2v_reg <= addr_tl_r[15];
      addr_v_r_14_sv2v_reg <= addr_tl_r[14];
      addr_v_r_13_sv2v_reg <= addr_tl_r[13];
      addr_v_r_12_sv2v_reg <= addr_tl_r[12];
      addr_v_r_11_sv2v_reg <= addr_tl_r[11];
      addr_v_r_10_sv2v_reg <= addr_tl_r[10];
      addr_v_r_9_sv2v_reg <= addr_tl_r[9];
      addr_v_r_8_sv2v_reg <= addr_tl_r[8];
      addr_v_r_7_sv2v_reg <= addr_tl_r[7];
      addr_v_r_6_sv2v_reg <= addr_tl_r[6];
      addr_v_r_5_sv2v_reg <= addr_tl_r[5];
      addr_v_r_4_sv2v_reg <= addr_tl_r[4];
      addr_v_r_3_sv2v_reg <= addr_tl_r[3];
      addr_v_r_2_sv2v_reg <= addr_tl_r[2];
      addr_v_r_1_sv2v_reg <= addr_tl_r[1];
      addr_v_r_0_sv2v_reg <= addr_tl_r[0];
      data_v_r_31_sv2v_reg <= data_tl_r[31];
      data_v_r_30_sv2v_reg <= data_tl_r[30];
      data_v_r_29_sv2v_reg <= data_tl_r[29];
      data_v_r_28_sv2v_reg <= data_tl_r[28];
      data_v_r_27_sv2v_reg <= data_tl_r[27];
      data_v_r_26_sv2v_reg <= data_tl_r[26];
      data_v_r_25_sv2v_reg <= data_tl_r[25];
      data_v_r_24_sv2v_reg <= data_tl_r[24];
      data_v_r_23_sv2v_reg <= data_tl_r[23];
      data_v_r_22_sv2v_reg <= data_tl_r[22];
      data_v_r_21_sv2v_reg <= data_tl_r[21];
      data_v_r_20_sv2v_reg <= data_tl_r[20];
      data_v_r_19_sv2v_reg <= data_tl_r[19];
      data_v_r_18_sv2v_reg <= data_tl_r[18];
      data_v_r_17_sv2v_reg <= data_tl_r[17];
      data_v_r_16_sv2v_reg <= data_tl_r[16];
      data_v_r_15_sv2v_reg <= data_tl_r[15];
      data_v_r_14_sv2v_reg <= data_tl_r[14];
      data_v_r_13_sv2v_reg <= data_tl_r[13];
      data_v_r_12_sv2v_reg <= data_tl_r[12];
      data_v_r_11_sv2v_reg <= data_tl_r[11];
      data_v_r_10_sv2v_reg <= data_tl_r[10];
      data_v_r_9_sv2v_reg <= data_tl_r[9];
      data_v_r_8_sv2v_reg <= data_tl_r[8];
      data_v_r_7_sv2v_reg <= data_tl_r[7];
      data_v_r_6_sv2v_reg <= data_tl_r[6];
      data_v_r_5_sv2v_reg <= data_tl_r[5];
      data_v_r_4_sv2v_reg <= data_tl_r[4];
      data_v_r_3_sv2v_reg <= data_tl_r[3];
      data_v_r_2_sv2v_reg <= data_tl_r[2];
      data_v_r_1_sv2v_reg <= data_tl_r[1];
      data_v_r_0_sv2v_reg <= data_tl_r[0];
      valid_v_r_1_sv2v_reg <= tag_mem_data_lo[39];
      valid_v_r_0_sv2v_reg <= tag_mem_data_lo[19];
      tag_v_r_10_sv2v_reg <= tag_mem_data_lo[10];
      tag_v_r_9_sv2v_reg <= tag_mem_data_lo[9];
      tag_v_r_8_sv2v_reg <= tag_mem_data_lo[8];
      tag_v_r_7_sv2v_reg <= tag_mem_data_lo[7];
      tag_v_r_6_sv2v_reg <= tag_mem_data_lo[6];
      tag_v_r_5_sv2v_reg <= tag_mem_data_lo[5];
      tag_v_r_4_sv2v_reg <= tag_mem_data_lo[4];
      tag_v_r_3_sv2v_reg <= tag_mem_data_lo[3];
      tag_v_r_2_sv2v_reg <= tag_mem_data_lo[2];
      tag_v_r_1_sv2v_reg <= tag_mem_data_lo[1];
      tag_v_r_0_sv2v_reg <= tag_mem_data_lo[0];
    end 
  end


endmodule

