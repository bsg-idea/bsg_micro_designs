

module top
(
  L_clk_i,
  L_reset_i,
  L_en_o,
  L_v_o,
  L_data_o,
  L_ready_i,
  L_v_i,
  L_data_i,
  L_yumi_o,
  R_clk_i,
  R_reset_i,
  R_en_i,
  R_v_i,
  R_data_i,
  R_ready_o,
  R_v_o,
  R_data_o,
  R_yumi_i
);

  output [49:0] L_data_o;
  input [49:0] L_data_i;
  input [49:0] R_data_i;
  output [49:0] R_data_o;
  input L_clk_i;
  input L_reset_i;
  input L_ready_i;
  input L_v_i;
  input R_clk_i;
  input R_reset_i;
  input R_en_i;
  input R_v_i;
  input R_yumi_i;
  output L_en_o;
  output L_v_o;
  output L_yumi_o;
  output R_ready_o;
  output R_v_o;

  bsg_fsb_node_async_buffer
  wrapper
  (
    .L_data_o(L_data_o),
    .L_data_i(L_data_i),
    .R_data_i(R_data_i),
    .R_data_o(R_data_o),
    .L_clk_i(L_clk_i),
    .L_reset_i(L_reset_i),
    .L_ready_i(L_ready_i),
    .L_v_i(L_v_i),
    .R_clk_i(R_clk_i),
    .R_reset_i(R_reset_i),
    .R_en_i(R_en_i),
    .R_v_i(R_v_i),
    .R_yumi_i(R_yumi_i),
    .L_en_o(L_en_o),
    .L_v_o(L_v_o),
    .L_yumi_o(L_yumi_o),
    .R_ready_o(R_ready_o),
    .R_v_o(R_v_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p50_els_p64_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [49:0] w_data_i;
  input [5:0] r_addr_i;
  output [49:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [49:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294;
  wire [3199:0] \nz.mem ;
  reg \nz.mem_3199_sv2v_reg ,\nz.mem_3198_sv2v_reg ,\nz.mem_3197_sv2v_reg ,
  \nz.mem_3196_sv2v_reg ,\nz.mem_3195_sv2v_reg ,\nz.mem_3194_sv2v_reg ,
  \nz.mem_3193_sv2v_reg ,\nz.mem_3192_sv2v_reg ,\nz.mem_3191_sv2v_reg ,\nz.mem_3190_sv2v_reg ,
  \nz.mem_3189_sv2v_reg ,\nz.mem_3188_sv2v_reg ,\nz.mem_3187_sv2v_reg ,
  \nz.mem_3186_sv2v_reg ,\nz.mem_3185_sv2v_reg ,\nz.mem_3184_sv2v_reg ,\nz.mem_3183_sv2v_reg ,
  \nz.mem_3182_sv2v_reg ,\nz.mem_3181_sv2v_reg ,\nz.mem_3180_sv2v_reg ,
  \nz.mem_3179_sv2v_reg ,\nz.mem_3178_sv2v_reg ,\nz.mem_3177_sv2v_reg ,\nz.mem_3176_sv2v_reg ,
  \nz.mem_3175_sv2v_reg ,\nz.mem_3174_sv2v_reg ,\nz.mem_3173_sv2v_reg ,
  \nz.mem_3172_sv2v_reg ,\nz.mem_3171_sv2v_reg ,\nz.mem_3170_sv2v_reg ,\nz.mem_3169_sv2v_reg ,
  \nz.mem_3168_sv2v_reg ,\nz.mem_3167_sv2v_reg ,\nz.mem_3166_sv2v_reg ,
  \nz.mem_3165_sv2v_reg ,\nz.mem_3164_sv2v_reg ,\nz.mem_3163_sv2v_reg ,\nz.mem_3162_sv2v_reg ,
  \nz.mem_3161_sv2v_reg ,\nz.mem_3160_sv2v_reg ,\nz.mem_3159_sv2v_reg ,
  \nz.mem_3158_sv2v_reg ,\nz.mem_3157_sv2v_reg ,\nz.mem_3156_sv2v_reg ,\nz.mem_3155_sv2v_reg ,
  \nz.mem_3154_sv2v_reg ,\nz.mem_3153_sv2v_reg ,\nz.mem_3152_sv2v_reg ,
  \nz.mem_3151_sv2v_reg ,\nz.mem_3150_sv2v_reg ,\nz.mem_3149_sv2v_reg ,\nz.mem_3148_sv2v_reg ,
  \nz.mem_3147_sv2v_reg ,\nz.mem_3146_sv2v_reg ,\nz.mem_3145_sv2v_reg ,
  \nz.mem_3144_sv2v_reg ,\nz.mem_3143_sv2v_reg ,\nz.mem_3142_sv2v_reg ,\nz.mem_3141_sv2v_reg ,
  \nz.mem_3140_sv2v_reg ,\nz.mem_3139_sv2v_reg ,\nz.mem_3138_sv2v_reg ,
  \nz.mem_3137_sv2v_reg ,\nz.mem_3136_sv2v_reg ,\nz.mem_3135_sv2v_reg ,\nz.mem_3134_sv2v_reg ,
  \nz.mem_3133_sv2v_reg ,\nz.mem_3132_sv2v_reg ,\nz.mem_3131_sv2v_reg ,
  \nz.mem_3130_sv2v_reg ,\nz.mem_3129_sv2v_reg ,\nz.mem_3128_sv2v_reg ,\nz.mem_3127_sv2v_reg ,
  \nz.mem_3126_sv2v_reg ,\nz.mem_3125_sv2v_reg ,\nz.mem_3124_sv2v_reg ,
  \nz.mem_3123_sv2v_reg ,\nz.mem_3122_sv2v_reg ,\nz.mem_3121_sv2v_reg ,\nz.mem_3120_sv2v_reg ,
  \nz.mem_3119_sv2v_reg ,\nz.mem_3118_sv2v_reg ,\nz.mem_3117_sv2v_reg ,
  \nz.mem_3116_sv2v_reg ,\nz.mem_3115_sv2v_reg ,\nz.mem_3114_sv2v_reg ,
  \nz.mem_3113_sv2v_reg ,\nz.mem_3112_sv2v_reg ,\nz.mem_3111_sv2v_reg ,\nz.mem_3110_sv2v_reg ,
  \nz.mem_3109_sv2v_reg ,\nz.mem_3108_sv2v_reg ,\nz.mem_3107_sv2v_reg ,
  \nz.mem_3106_sv2v_reg ,\nz.mem_3105_sv2v_reg ,\nz.mem_3104_sv2v_reg ,\nz.mem_3103_sv2v_reg ,
  \nz.mem_3102_sv2v_reg ,\nz.mem_3101_sv2v_reg ,\nz.mem_3100_sv2v_reg ,
  \nz.mem_3099_sv2v_reg ,\nz.mem_3098_sv2v_reg ,\nz.mem_3097_sv2v_reg ,\nz.mem_3096_sv2v_reg ,
  \nz.mem_3095_sv2v_reg ,\nz.mem_3094_sv2v_reg ,\nz.mem_3093_sv2v_reg ,
  \nz.mem_3092_sv2v_reg ,\nz.mem_3091_sv2v_reg ,\nz.mem_3090_sv2v_reg ,\nz.mem_3089_sv2v_reg ,
  \nz.mem_3088_sv2v_reg ,\nz.mem_3087_sv2v_reg ,\nz.mem_3086_sv2v_reg ,
  \nz.mem_3085_sv2v_reg ,\nz.mem_3084_sv2v_reg ,\nz.mem_3083_sv2v_reg ,\nz.mem_3082_sv2v_reg ,
  \nz.mem_3081_sv2v_reg ,\nz.mem_3080_sv2v_reg ,\nz.mem_3079_sv2v_reg ,
  \nz.mem_3078_sv2v_reg ,\nz.mem_3077_sv2v_reg ,\nz.mem_3076_sv2v_reg ,\nz.mem_3075_sv2v_reg ,
  \nz.mem_3074_sv2v_reg ,\nz.mem_3073_sv2v_reg ,\nz.mem_3072_sv2v_reg ,
  \nz.mem_3071_sv2v_reg ,\nz.mem_3070_sv2v_reg ,\nz.mem_3069_sv2v_reg ,\nz.mem_3068_sv2v_reg ,
  \nz.mem_3067_sv2v_reg ,\nz.mem_3066_sv2v_reg ,\nz.mem_3065_sv2v_reg ,
  \nz.mem_3064_sv2v_reg ,\nz.mem_3063_sv2v_reg ,\nz.mem_3062_sv2v_reg ,\nz.mem_3061_sv2v_reg ,
  \nz.mem_3060_sv2v_reg ,\nz.mem_3059_sv2v_reg ,\nz.mem_3058_sv2v_reg ,
  \nz.mem_3057_sv2v_reg ,\nz.mem_3056_sv2v_reg ,\nz.mem_3055_sv2v_reg ,\nz.mem_3054_sv2v_reg ,
  \nz.mem_3053_sv2v_reg ,\nz.mem_3052_sv2v_reg ,\nz.mem_3051_sv2v_reg ,
  \nz.mem_3050_sv2v_reg ,\nz.mem_3049_sv2v_reg ,\nz.mem_3048_sv2v_reg ,\nz.mem_3047_sv2v_reg ,
  \nz.mem_3046_sv2v_reg ,\nz.mem_3045_sv2v_reg ,\nz.mem_3044_sv2v_reg ,
  \nz.mem_3043_sv2v_reg ,\nz.mem_3042_sv2v_reg ,\nz.mem_3041_sv2v_reg ,\nz.mem_3040_sv2v_reg ,
  \nz.mem_3039_sv2v_reg ,\nz.mem_3038_sv2v_reg ,\nz.mem_3037_sv2v_reg ,
  \nz.mem_3036_sv2v_reg ,\nz.mem_3035_sv2v_reg ,\nz.mem_3034_sv2v_reg ,
  \nz.mem_3033_sv2v_reg ,\nz.mem_3032_sv2v_reg ,\nz.mem_3031_sv2v_reg ,\nz.mem_3030_sv2v_reg ,
  \nz.mem_3029_sv2v_reg ,\nz.mem_3028_sv2v_reg ,\nz.mem_3027_sv2v_reg ,
  \nz.mem_3026_sv2v_reg ,\nz.mem_3025_sv2v_reg ,\nz.mem_3024_sv2v_reg ,\nz.mem_3023_sv2v_reg ,
  \nz.mem_3022_sv2v_reg ,\nz.mem_3021_sv2v_reg ,\nz.mem_3020_sv2v_reg ,
  \nz.mem_3019_sv2v_reg ,\nz.mem_3018_sv2v_reg ,\nz.mem_3017_sv2v_reg ,\nz.mem_3016_sv2v_reg ,
  \nz.mem_3015_sv2v_reg ,\nz.mem_3014_sv2v_reg ,\nz.mem_3013_sv2v_reg ,
  \nz.mem_3012_sv2v_reg ,\nz.mem_3011_sv2v_reg ,\nz.mem_3010_sv2v_reg ,\nz.mem_3009_sv2v_reg ,
  \nz.mem_3008_sv2v_reg ,\nz.mem_3007_sv2v_reg ,\nz.mem_3006_sv2v_reg ,
  \nz.mem_3005_sv2v_reg ,\nz.mem_3004_sv2v_reg ,\nz.mem_3003_sv2v_reg ,\nz.mem_3002_sv2v_reg ,
  \nz.mem_3001_sv2v_reg ,\nz.mem_3000_sv2v_reg ,\nz.mem_2999_sv2v_reg ,
  \nz.mem_2998_sv2v_reg ,\nz.mem_2997_sv2v_reg ,\nz.mem_2996_sv2v_reg ,\nz.mem_2995_sv2v_reg ,
  \nz.mem_2994_sv2v_reg ,\nz.mem_2993_sv2v_reg ,\nz.mem_2992_sv2v_reg ,
  \nz.mem_2991_sv2v_reg ,\nz.mem_2990_sv2v_reg ,\nz.mem_2989_sv2v_reg ,\nz.mem_2988_sv2v_reg ,
  \nz.mem_2987_sv2v_reg ,\nz.mem_2986_sv2v_reg ,\nz.mem_2985_sv2v_reg ,
  \nz.mem_2984_sv2v_reg ,\nz.mem_2983_sv2v_reg ,\nz.mem_2982_sv2v_reg ,\nz.mem_2981_sv2v_reg ,
  \nz.mem_2980_sv2v_reg ,\nz.mem_2979_sv2v_reg ,\nz.mem_2978_sv2v_reg ,
  \nz.mem_2977_sv2v_reg ,\nz.mem_2976_sv2v_reg ,\nz.mem_2975_sv2v_reg ,\nz.mem_2974_sv2v_reg ,
  \nz.mem_2973_sv2v_reg ,\nz.mem_2972_sv2v_reg ,\nz.mem_2971_sv2v_reg ,
  \nz.mem_2970_sv2v_reg ,\nz.mem_2969_sv2v_reg ,\nz.mem_2968_sv2v_reg ,\nz.mem_2967_sv2v_reg ,
  \nz.mem_2966_sv2v_reg ,\nz.mem_2965_sv2v_reg ,\nz.mem_2964_sv2v_reg ,
  \nz.mem_2963_sv2v_reg ,\nz.mem_2962_sv2v_reg ,\nz.mem_2961_sv2v_reg ,\nz.mem_2960_sv2v_reg ,
  \nz.mem_2959_sv2v_reg ,\nz.mem_2958_sv2v_reg ,\nz.mem_2957_sv2v_reg ,
  \nz.mem_2956_sv2v_reg ,\nz.mem_2955_sv2v_reg ,\nz.mem_2954_sv2v_reg ,
  \nz.mem_2953_sv2v_reg ,\nz.mem_2952_sv2v_reg ,\nz.mem_2951_sv2v_reg ,\nz.mem_2950_sv2v_reg ,
  \nz.mem_2949_sv2v_reg ,\nz.mem_2948_sv2v_reg ,\nz.mem_2947_sv2v_reg ,
  \nz.mem_2946_sv2v_reg ,\nz.mem_2945_sv2v_reg ,\nz.mem_2944_sv2v_reg ,\nz.mem_2943_sv2v_reg ,
  \nz.mem_2942_sv2v_reg ,\nz.mem_2941_sv2v_reg ,\nz.mem_2940_sv2v_reg ,
  \nz.mem_2939_sv2v_reg ,\nz.mem_2938_sv2v_reg ,\nz.mem_2937_sv2v_reg ,\nz.mem_2936_sv2v_reg ,
  \nz.mem_2935_sv2v_reg ,\nz.mem_2934_sv2v_reg ,\nz.mem_2933_sv2v_reg ,
  \nz.mem_2932_sv2v_reg ,\nz.mem_2931_sv2v_reg ,\nz.mem_2930_sv2v_reg ,\nz.mem_2929_sv2v_reg ,
  \nz.mem_2928_sv2v_reg ,\nz.mem_2927_sv2v_reg ,\nz.mem_2926_sv2v_reg ,
  \nz.mem_2925_sv2v_reg ,\nz.mem_2924_sv2v_reg ,\nz.mem_2923_sv2v_reg ,\nz.mem_2922_sv2v_reg ,
  \nz.mem_2921_sv2v_reg ,\nz.mem_2920_sv2v_reg ,\nz.mem_2919_sv2v_reg ,
  \nz.mem_2918_sv2v_reg ,\nz.mem_2917_sv2v_reg ,\nz.mem_2916_sv2v_reg ,\nz.mem_2915_sv2v_reg ,
  \nz.mem_2914_sv2v_reg ,\nz.mem_2913_sv2v_reg ,\nz.mem_2912_sv2v_reg ,
  \nz.mem_2911_sv2v_reg ,\nz.mem_2910_sv2v_reg ,\nz.mem_2909_sv2v_reg ,\nz.mem_2908_sv2v_reg ,
  \nz.mem_2907_sv2v_reg ,\nz.mem_2906_sv2v_reg ,\nz.mem_2905_sv2v_reg ,
  \nz.mem_2904_sv2v_reg ,\nz.mem_2903_sv2v_reg ,\nz.mem_2902_sv2v_reg ,\nz.mem_2901_sv2v_reg ,
  \nz.mem_2900_sv2v_reg ,\nz.mem_2899_sv2v_reg ,\nz.mem_2898_sv2v_reg ,
  \nz.mem_2897_sv2v_reg ,\nz.mem_2896_sv2v_reg ,\nz.mem_2895_sv2v_reg ,\nz.mem_2894_sv2v_reg ,
  \nz.mem_2893_sv2v_reg ,\nz.mem_2892_sv2v_reg ,\nz.mem_2891_sv2v_reg ,
  \nz.mem_2890_sv2v_reg ,\nz.mem_2889_sv2v_reg ,\nz.mem_2888_sv2v_reg ,\nz.mem_2887_sv2v_reg ,
  \nz.mem_2886_sv2v_reg ,\nz.mem_2885_sv2v_reg ,\nz.mem_2884_sv2v_reg ,
  \nz.mem_2883_sv2v_reg ,\nz.mem_2882_sv2v_reg ,\nz.mem_2881_sv2v_reg ,\nz.mem_2880_sv2v_reg ,
  \nz.mem_2879_sv2v_reg ,\nz.mem_2878_sv2v_reg ,\nz.mem_2877_sv2v_reg ,
  \nz.mem_2876_sv2v_reg ,\nz.mem_2875_sv2v_reg ,\nz.mem_2874_sv2v_reg ,
  \nz.mem_2873_sv2v_reg ,\nz.mem_2872_sv2v_reg ,\nz.mem_2871_sv2v_reg ,\nz.mem_2870_sv2v_reg ,
  \nz.mem_2869_sv2v_reg ,\nz.mem_2868_sv2v_reg ,\nz.mem_2867_sv2v_reg ,
  \nz.mem_2866_sv2v_reg ,\nz.mem_2865_sv2v_reg ,\nz.mem_2864_sv2v_reg ,\nz.mem_2863_sv2v_reg ,
  \nz.mem_2862_sv2v_reg ,\nz.mem_2861_sv2v_reg ,\nz.mem_2860_sv2v_reg ,
  \nz.mem_2859_sv2v_reg ,\nz.mem_2858_sv2v_reg ,\nz.mem_2857_sv2v_reg ,\nz.mem_2856_sv2v_reg ,
  \nz.mem_2855_sv2v_reg ,\nz.mem_2854_sv2v_reg ,\nz.mem_2853_sv2v_reg ,
  \nz.mem_2852_sv2v_reg ,\nz.mem_2851_sv2v_reg ,\nz.mem_2850_sv2v_reg ,\nz.mem_2849_sv2v_reg ,
  \nz.mem_2848_sv2v_reg ,\nz.mem_2847_sv2v_reg ,\nz.mem_2846_sv2v_reg ,
  \nz.mem_2845_sv2v_reg ,\nz.mem_2844_sv2v_reg ,\nz.mem_2843_sv2v_reg ,\nz.mem_2842_sv2v_reg ,
  \nz.mem_2841_sv2v_reg ,\nz.mem_2840_sv2v_reg ,\nz.mem_2839_sv2v_reg ,
  \nz.mem_2838_sv2v_reg ,\nz.mem_2837_sv2v_reg ,\nz.mem_2836_sv2v_reg ,\nz.mem_2835_sv2v_reg ,
  \nz.mem_2834_sv2v_reg ,\nz.mem_2833_sv2v_reg ,\nz.mem_2832_sv2v_reg ,
  \nz.mem_2831_sv2v_reg ,\nz.mem_2830_sv2v_reg ,\nz.mem_2829_sv2v_reg ,\nz.mem_2828_sv2v_reg ,
  \nz.mem_2827_sv2v_reg ,\nz.mem_2826_sv2v_reg ,\nz.mem_2825_sv2v_reg ,
  \nz.mem_2824_sv2v_reg ,\nz.mem_2823_sv2v_reg ,\nz.mem_2822_sv2v_reg ,\nz.mem_2821_sv2v_reg ,
  \nz.mem_2820_sv2v_reg ,\nz.mem_2819_sv2v_reg ,\nz.mem_2818_sv2v_reg ,
  \nz.mem_2817_sv2v_reg ,\nz.mem_2816_sv2v_reg ,\nz.mem_2815_sv2v_reg ,\nz.mem_2814_sv2v_reg ,
  \nz.mem_2813_sv2v_reg ,\nz.mem_2812_sv2v_reg ,\nz.mem_2811_sv2v_reg ,
  \nz.mem_2810_sv2v_reg ,\nz.mem_2809_sv2v_reg ,\nz.mem_2808_sv2v_reg ,\nz.mem_2807_sv2v_reg ,
  \nz.mem_2806_sv2v_reg ,\nz.mem_2805_sv2v_reg ,\nz.mem_2804_sv2v_reg ,
  \nz.mem_2803_sv2v_reg ,\nz.mem_2802_sv2v_reg ,\nz.mem_2801_sv2v_reg ,\nz.mem_2800_sv2v_reg ,
  \nz.mem_2799_sv2v_reg ,\nz.mem_2798_sv2v_reg ,\nz.mem_2797_sv2v_reg ,
  \nz.mem_2796_sv2v_reg ,\nz.mem_2795_sv2v_reg ,\nz.mem_2794_sv2v_reg ,
  \nz.mem_2793_sv2v_reg ,\nz.mem_2792_sv2v_reg ,\nz.mem_2791_sv2v_reg ,\nz.mem_2790_sv2v_reg ,
  \nz.mem_2789_sv2v_reg ,\nz.mem_2788_sv2v_reg ,\nz.mem_2787_sv2v_reg ,
  \nz.mem_2786_sv2v_reg ,\nz.mem_2785_sv2v_reg ,\nz.mem_2784_sv2v_reg ,\nz.mem_2783_sv2v_reg ,
  \nz.mem_2782_sv2v_reg ,\nz.mem_2781_sv2v_reg ,\nz.mem_2780_sv2v_reg ,
  \nz.mem_2779_sv2v_reg ,\nz.mem_2778_sv2v_reg ,\nz.mem_2777_sv2v_reg ,\nz.mem_2776_sv2v_reg ,
  \nz.mem_2775_sv2v_reg ,\nz.mem_2774_sv2v_reg ,\nz.mem_2773_sv2v_reg ,
  \nz.mem_2772_sv2v_reg ,\nz.mem_2771_sv2v_reg ,\nz.mem_2770_sv2v_reg ,\nz.mem_2769_sv2v_reg ,
  \nz.mem_2768_sv2v_reg ,\nz.mem_2767_sv2v_reg ,\nz.mem_2766_sv2v_reg ,
  \nz.mem_2765_sv2v_reg ,\nz.mem_2764_sv2v_reg ,\nz.mem_2763_sv2v_reg ,\nz.mem_2762_sv2v_reg ,
  \nz.mem_2761_sv2v_reg ,\nz.mem_2760_sv2v_reg ,\nz.mem_2759_sv2v_reg ,
  \nz.mem_2758_sv2v_reg ,\nz.mem_2757_sv2v_reg ,\nz.mem_2756_sv2v_reg ,\nz.mem_2755_sv2v_reg ,
  \nz.mem_2754_sv2v_reg ,\nz.mem_2753_sv2v_reg ,\nz.mem_2752_sv2v_reg ,
  \nz.mem_2751_sv2v_reg ,\nz.mem_2750_sv2v_reg ,\nz.mem_2749_sv2v_reg ,\nz.mem_2748_sv2v_reg ,
  \nz.mem_2747_sv2v_reg ,\nz.mem_2746_sv2v_reg ,\nz.mem_2745_sv2v_reg ,
  \nz.mem_2744_sv2v_reg ,\nz.mem_2743_sv2v_reg ,\nz.mem_2742_sv2v_reg ,\nz.mem_2741_sv2v_reg ,
  \nz.mem_2740_sv2v_reg ,\nz.mem_2739_sv2v_reg ,\nz.mem_2738_sv2v_reg ,
  \nz.mem_2737_sv2v_reg ,\nz.mem_2736_sv2v_reg ,\nz.mem_2735_sv2v_reg ,\nz.mem_2734_sv2v_reg ,
  \nz.mem_2733_sv2v_reg ,\nz.mem_2732_sv2v_reg ,\nz.mem_2731_sv2v_reg ,
  \nz.mem_2730_sv2v_reg ,\nz.mem_2729_sv2v_reg ,\nz.mem_2728_sv2v_reg ,\nz.mem_2727_sv2v_reg ,
  \nz.mem_2726_sv2v_reg ,\nz.mem_2725_sv2v_reg ,\nz.mem_2724_sv2v_reg ,
  \nz.mem_2723_sv2v_reg ,\nz.mem_2722_sv2v_reg ,\nz.mem_2721_sv2v_reg ,\nz.mem_2720_sv2v_reg ,
  \nz.mem_2719_sv2v_reg ,\nz.mem_2718_sv2v_reg ,\nz.mem_2717_sv2v_reg ,
  \nz.mem_2716_sv2v_reg ,\nz.mem_2715_sv2v_reg ,\nz.mem_2714_sv2v_reg ,
  \nz.mem_2713_sv2v_reg ,\nz.mem_2712_sv2v_reg ,\nz.mem_2711_sv2v_reg ,\nz.mem_2710_sv2v_reg ,
  \nz.mem_2709_sv2v_reg ,\nz.mem_2708_sv2v_reg ,\nz.mem_2707_sv2v_reg ,
  \nz.mem_2706_sv2v_reg ,\nz.mem_2705_sv2v_reg ,\nz.mem_2704_sv2v_reg ,\nz.mem_2703_sv2v_reg ,
  \nz.mem_2702_sv2v_reg ,\nz.mem_2701_sv2v_reg ,\nz.mem_2700_sv2v_reg ,
  \nz.mem_2699_sv2v_reg ,\nz.mem_2698_sv2v_reg ,\nz.mem_2697_sv2v_reg ,\nz.mem_2696_sv2v_reg ,
  \nz.mem_2695_sv2v_reg ,\nz.mem_2694_sv2v_reg ,\nz.mem_2693_sv2v_reg ,
  \nz.mem_2692_sv2v_reg ,\nz.mem_2691_sv2v_reg ,\nz.mem_2690_sv2v_reg ,\nz.mem_2689_sv2v_reg ,
  \nz.mem_2688_sv2v_reg ,\nz.mem_2687_sv2v_reg ,\nz.mem_2686_sv2v_reg ,
  \nz.mem_2685_sv2v_reg ,\nz.mem_2684_sv2v_reg ,\nz.mem_2683_sv2v_reg ,\nz.mem_2682_sv2v_reg ,
  \nz.mem_2681_sv2v_reg ,\nz.mem_2680_sv2v_reg ,\nz.mem_2679_sv2v_reg ,
  \nz.mem_2678_sv2v_reg ,\nz.mem_2677_sv2v_reg ,\nz.mem_2676_sv2v_reg ,\nz.mem_2675_sv2v_reg ,
  \nz.mem_2674_sv2v_reg ,\nz.mem_2673_sv2v_reg ,\nz.mem_2672_sv2v_reg ,
  \nz.mem_2671_sv2v_reg ,\nz.mem_2670_sv2v_reg ,\nz.mem_2669_sv2v_reg ,\nz.mem_2668_sv2v_reg ,
  \nz.mem_2667_sv2v_reg ,\nz.mem_2666_sv2v_reg ,\nz.mem_2665_sv2v_reg ,
  \nz.mem_2664_sv2v_reg ,\nz.mem_2663_sv2v_reg ,\nz.mem_2662_sv2v_reg ,\nz.mem_2661_sv2v_reg ,
  \nz.mem_2660_sv2v_reg ,\nz.mem_2659_sv2v_reg ,\nz.mem_2658_sv2v_reg ,
  \nz.mem_2657_sv2v_reg ,\nz.mem_2656_sv2v_reg ,\nz.mem_2655_sv2v_reg ,\nz.mem_2654_sv2v_reg ,
  \nz.mem_2653_sv2v_reg ,\nz.mem_2652_sv2v_reg ,\nz.mem_2651_sv2v_reg ,
  \nz.mem_2650_sv2v_reg ,\nz.mem_2649_sv2v_reg ,\nz.mem_2648_sv2v_reg ,\nz.mem_2647_sv2v_reg ,
  \nz.mem_2646_sv2v_reg ,\nz.mem_2645_sv2v_reg ,\nz.mem_2644_sv2v_reg ,
  \nz.mem_2643_sv2v_reg ,\nz.mem_2642_sv2v_reg ,\nz.mem_2641_sv2v_reg ,\nz.mem_2640_sv2v_reg ,
  \nz.mem_2639_sv2v_reg ,\nz.mem_2638_sv2v_reg ,\nz.mem_2637_sv2v_reg ,
  \nz.mem_2636_sv2v_reg ,\nz.mem_2635_sv2v_reg ,\nz.mem_2634_sv2v_reg ,
  \nz.mem_2633_sv2v_reg ,\nz.mem_2632_sv2v_reg ,\nz.mem_2631_sv2v_reg ,\nz.mem_2630_sv2v_reg ,
  \nz.mem_2629_sv2v_reg ,\nz.mem_2628_sv2v_reg ,\nz.mem_2627_sv2v_reg ,
  \nz.mem_2626_sv2v_reg ,\nz.mem_2625_sv2v_reg ,\nz.mem_2624_sv2v_reg ,\nz.mem_2623_sv2v_reg ,
  \nz.mem_2622_sv2v_reg ,\nz.mem_2621_sv2v_reg ,\nz.mem_2620_sv2v_reg ,
  \nz.mem_2619_sv2v_reg ,\nz.mem_2618_sv2v_reg ,\nz.mem_2617_sv2v_reg ,\nz.mem_2616_sv2v_reg ,
  \nz.mem_2615_sv2v_reg ,\nz.mem_2614_sv2v_reg ,\nz.mem_2613_sv2v_reg ,
  \nz.mem_2612_sv2v_reg ,\nz.mem_2611_sv2v_reg ,\nz.mem_2610_sv2v_reg ,\nz.mem_2609_sv2v_reg ,
  \nz.mem_2608_sv2v_reg ,\nz.mem_2607_sv2v_reg ,\nz.mem_2606_sv2v_reg ,
  \nz.mem_2605_sv2v_reg ,\nz.mem_2604_sv2v_reg ,\nz.mem_2603_sv2v_reg ,\nz.mem_2602_sv2v_reg ,
  \nz.mem_2601_sv2v_reg ,\nz.mem_2600_sv2v_reg ,\nz.mem_2599_sv2v_reg ,
  \nz.mem_2598_sv2v_reg ,\nz.mem_2597_sv2v_reg ,\nz.mem_2596_sv2v_reg ,\nz.mem_2595_sv2v_reg ,
  \nz.mem_2594_sv2v_reg ,\nz.mem_2593_sv2v_reg ,\nz.mem_2592_sv2v_reg ,
  \nz.mem_2591_sv2v_reg ,\nz.mem_2590_sv2v_reg ,\nz.mem_2589_sv2v_reg ,\nz.mem_2588_sv2v_reg ,
  \nz.mem_2587_sv2v_reg ,\nz.mem_2586_sv2v_reg ,\nz.mem_2585_sv2v_reg ,
  \nz.mem_2584_sv2v_reg ,\nz.mem_2583_sv2v_reg ,\nz.mem_2582_sv2v_reg ,\nz.mem_2581_sv2v_reg ,
  \nz.mem_2580_sv2v_reg ,\nz.mem_2579_sv2v_reg ,\nz.mem_2578_sv2v_reg ,
  \nz.mem_2577_sv2v_reg ,\nz.mem_2576_sv2v_reg ,\nz.mem_2575_sv2v_reg ,\nz.mem_2574_sv2v_reg ,
  \nz.mem_2573_sv2v_reg ,\nz.mem_2572_sv2v_reg ,\nz.mem_2571_sv2v_reg ,
  \nz.mem_2570_sv2v_reg ,\nz.mem_2569_sv2v_reg ,\nz.mem_2568_sv2v_reg ,\nz.mem_2567_sv2v_reg ,
  \nz.mem_2566_sv2v_reg ,\nz.mem_2565_sv2v_reg ,\nz.mem_2564_sv2v_reg ,
  \nz.mem_2563_sv2v_reg ,\nz.mem_2562_sv2v_reg ,\nz.mem_2561_sv2v_reg ,\nz.mem_2560_sv2v_reg ,
  \nz.mem_2559_sv2v_reg ,\nz.mem_2558_sv2v_reg ,\nz.mem_2557_sv2v_reg ,
  \nz.mem_2556_sv2v_reg ,\nz.mem_2555_sv2v_reg ,\nz.mem_2554_sv2v_reg ,
  \nz.mem_2553_sv2v_reg ,\nz.mem_2552_sv2v_reg ,\nz.mem_2551_sv2v_reg ,\nz.mem_2550_sv2v_reg ,
  \nz.mem_2549_sv2v_reg ,\nz.mem_2548_sv2v_reg ,\nz.mem_2547_sv2v_reg ,
  \nz.mem_2546_sv2v_reg ,\nz.mem_2545_sv2v_reg ,\nz.mem_2544_sv2v_reg ,\nz.mem_2543_sv2v_reg ,
  \nz.mem_2542_sv2v_reg ,\nz.mem_2541_sv2v_reg ,\nz.mem_2540_sv2v_reg ,
  \nz.mem_2539_sv2v_reg ,\nz.mem_2538_sv2v_reg ,\nz.mem_2537_sv2v_reg ,\nz.mem_2536_sv2v_reg ,
  \nz.mem_2535_sv2v_reg ,\nz.mem_2534_sv2v_reg ,\nz.mem_2533_sv2v_reg ,
  \nz.mem_2532_sv2v_reg ,\nz.mem_2531_sv2v_reg ,\nz.mem_2530_sv2v_reg ,\nz.mem_2529_sv2v_reg ,
  \nz.mem_2528_sv2v_reg ,\nz.mem_2527_sv2v_reg ,\nz.mem_2526_sv2v_reg ,
  \nz.mem_2525_sv2v_reg ,\nz.mem_2524_sv2v_reg ,\nz.mem_2523_sv2v_reg ,\nz.mem_2522_sv2v_reg ,
  \nz.mem_2521_sv2v_reg ,\nz.mem_2520_sv2v_reg ,\nz.mem_2519_sv2v_reg ,
  \nz.mem_2518_sv2v_reg ,\nz.mem_2517_sv2v_reg ,\nz.mem_2516_sv2v_reg ,\nz.mem_2515_sv2v_reg ,
  \nz.mem_2514_sv2v_reg ,\nz.mem_2513_sv2v_reg ,\nz.mem_2512_sv2v_reg ,
  \nz.mem_2511_sv2v_reg ,\nz.mem_2510_sv2v_reg ,\nz.mem_2509_sv2v_reg ,\nz.mem_2508_sv2v_reg ,
  \nz.mem_2507_sv2v_reg ,\nz.mem_2506_sv2v_reg ,\nz.mem_2505_sv2v_reg ,
  \nz.mem_2504_sv2v_reg ,\nz.mem_2503_sv2v_reg ,\nz.mem_2502_sv2v_reg ,\nz.mem_2501_sv2v_reg ,
  \nz.mem_2500_sv2v_reg ,\nz.mem_2499_sv2v_reg ,\nz.mem_2498_sv2v_reg ,
  \nz.mem_2497_sv2v_reg ,\nz.mem_2496_sv2v_reg ,\nz.mem_2495_sv2v_reg ,\nz.mem_2494_sv2v_reg ,
  \nz.mem_2493_sv2v_reg ,\nz.mem_2492_sv2v_reg ,\nz.mem_2491_sv2v_reg ,
  \nz.mem_2490_sv2v_reg ,\nz.mem_2489_sv2v_reg ,\nz.mem_2488_sv2v_reg ,\nz.mem_2487_sv2v_reg ,
  \nz.mem_2486_sv2v_reg ,\nz.mem_2485_sv2v_reg ,\nz.mem_2484_sv2v_reg ,
  \nz.mem_2483_sv2v_reg ,\nz.mem_2482_sv2v_reg ,\nz.mem_2481_sv2v_reg ,\nz.mem_2480_sv2v_reg ,
  \nz.mem_2479_sv2v_reg ,\nz.mem_2478_sv2v_reg ,\nz.mem_2477_sv2v_reg ,
  \nz.mem_2476_sv2v_reg ,\nz.mem_2475_sv2v_reg ,\nz.mem_2474_sv2v_reg ,
  \nz.mem_2473_sv2v_reg ,\nz.mem_2472_sv2v_reg ,\nz.mem_2471_sv2v_reg ,\nz.mem_2470_sv2v_reg ,
  \nz.mem_2469_sv2v_reg ,\nz.mem_2468_sv2v_reg ,\nz.mem_2467_sv2v_reg ,
  \nz.mem_2466_sv2v_reg ,\nz.mem_2465_sv2v_reg ,\nz.mem_2464_sv2v_reg ,\nz.mem_2463_sv2v_reg ,
  \nz.mem_2462_sv2v_reg ,\nz.mem_2461_sv2v_reg ,\nz.mem_2460_sv2v_reg ,
  \nz.mem_2459_sv2v_reg ,\nz.mem_2458_sv2v_reg ,\nz.mem_2457_sv2v_reg ,\nz.mem_2456_sv2v_reg ,
  \nz.mem_2455_sv2v_reg ,\nz.mem_2454_sv2v_reg ,\nz.mem_2453_sv2v_reg ,
  \nz.mem_2452_sv2v_reg ,\nz.mem_2451_sv2v_reg ,\nz.mem_2450_sv2v_reg ,\nz.mem_2449_sv2v_reg ,
  \nz.mem_2448_sv2v_reg ,\nz.mem_2447_sv2v_reg ,\nz.mem_2446_sv2v_reg ,
  \nz.mem_2445_sv2v_reg ,\nz.mem_2444_sv2v_reg ,\nz.mem_2443_sv2v_reg ,\nz.mem_2442_sv2v_reg ,
  \nz.mem_2441_sv2v_reg ,\nz.mem_2440_sv2v_reg ,\nz.mem_2439_sv2v_reg ,
  \nz.mem_2438_sv2v_reg ,\nz.mem_2437_sv2v_reg ,\nz.mem_2436_sv2v_reg ,\nz.mem_2435_sv2v_reg ,
  \nz.mem_2434_sv2v_reg ,\nz.mem_2433_sv2v_reg ,\nz.mem_2432_sv2v_reg ,
  \nz.mem_2431_sv2v_reg ,\nz.mem_2430_sv2v_reg ,\nz.mem_2429_sv2v_reg ,\nz.mem_2428_sv2v_reg ,
  \nz.mem_2427_sv2v_reg ,\nz.mem_2426_sv2v_reg ,\nz.mem_2425_sv2v_reg ,
  \nz.mem_2424_sv2v_reg ,\nz.mem_2423_sv2v_reg ,\nz.mem_2422_sv2v_reg ,\nz.mem_2421_sv2v_reg ,
  \nz.mem_2420_sv2v_reg ,\nz.mem_2419_sv2v_reg ,\nz.mem_2418_sv2v_reg ,
  \nz.mem_2417_sv2v_reg ,\nz.mem_2416_sv2v_reg ,\nz.mem_2415_sv2v_reg ,\nz.mem_2414_sv2v_reg ,
  \nz.mem_2413_sv2v_reg ,\nz.mem_2412_sv2v_reg ,\nz.mem_2411_sv2v_reg ,
  \nz.mem_2410_sv2v_reg ,\nz.mem_2409_sv2v_reg ,\nz.mem_2408_sv2v_reg ,\nz.mem_2407_sv2v_reg ,
  \nz.mem_2406_sv2v_reg ,\nz.mem_2405_sv2v_reg ,\nz.mem_2404_sv2v_reg ,
  \nz.mem_2403_sv2v_reg ,\nz.mem_2402_sv2v_reg ,\nz.mem_2401_sv2v_reg ,\nz.mem_2400_sv2v_reg ,
  \nz.mem_2399_sv2v_reg ,\nz.mem_2398_sv2v_reg ,\nz.mem_2397_sv2v_reg ,
  \nz.mem_2396_sv2v_reg ,\nz.mem_2395_sv2v_reg ,\nz.mem_2394_sv2v_reg ,
  \nz.mem_2393_sv2v_reg ,\nz.mem_2392_sv2v_reg ,\nz.mem_2391_sv2v_reg ,\nz.mem_2390_sv2v_reg ,
  \nz.mem_2389_sv2v_reg ,\nz.mem_2388_sv2v_reg ,\nz.mem_2387_sv2v_reg ,
  \nz.mem_2386_sv2v_reg ,\nz.mem_2385_sv2v_reg ,\nz.mem_2384_sv2v_reg ,\nz.mem_2383_sv2v_reg ,
  \nz.mem_2382_sv2v_reg ,\nz.mem_2381_sv2v_reg ,\nz.mem_2380_sv2v_reg ,
  \nz.mem_2379_sv2v_reg ,\nz.mem_2378_sv2v_reg ,\nz.mem_2377_sv2v_reg ,\nz.mem_2376_sv2v_reg ,
  \nz.mem_2375_sv2v_reg ,\nz.mem_2374_sv2v_reg ,\nz.mem_2373_sv2v_reg ,
  \nz.mem_2372_sv2v_reg ,\nz.mem_2371_sv2v_reg ,\nz.mem_2370_sv2v_reg ,\nz.mem_2369_sv2v_reg ,
  \nz.mem_2368_sv2v_reg ,\nz.mem_2367_sv2v_reg ,\nz.mem_2366_sv2v_reg ,
  \nz.mem_2365_sv2v_reg ,\nz.mem_2364_sv2v_reg ,\nz.mem_2363_sv2v_reg ,\nz.mem_2362_sv2v_reg ,
  \nz.mem_2361_sv2v_reg ,\nz.mem_2360_sv2v_reg ,\nz.mem_2359_sv2v_reg ,
  \nz.mem_2358_sv2v_reg ,\nz.mem_2357_sv2v_reg ,\nz.mem_2356_sv2v_reg ,\nz.mem_2355_sv2v_reg ,
  \nz.mem_2354_sv2v_reg ,\nz.mem_2353_sv2v_reg ,\nz.mem_2352_sv2v_reg ,
  \nz.mem_2351_sv2v_reg ,\nz.mem_2350_sv2v_reg ,\nz.mem_2349_sv2v_reg ,\nz.mem_2348_sv2v_reg ,
  \nz.mem_2347_sv2v_reg ,\nz.mem_2346_sv2v_reg ,\nz.mem_2345_sv2v_reg ,
  \nz.mem_2344_sv2v_reg ,\nz.mem_2343_sv2v_reg ,\nz.mem_2342_sv2v_reg ,\nz.mem_2341_sv2v_reg ,
  \nz.mem_2340_sv2v_reg ,\nz.mem_2339_sv2v_reg ,\nz.mem_2338_sv2v_reg ,
  \nz.mem_2337_sv2v_reg ,\nz.mem_2336_sv2v_reg ,\nz.mem_2335_sv2v_reg ,\nz.mem_2334_sv2v_reg ,
  \nz.mem_2333_sv2v_reg ,\nz.mem_2332_sv2v_reg ,\nz.mem_2331_sv2v_reg ,
  \nz.mem_2330_sv2v_reg ,\nz.mem_2329_sv2v_reg ,\nz.mem_2328_sv2v_reg ,\nz.mem_2327_sv2v_reg ,
  \nz.mem_2326_sv2v_reg ,\nz.mem_2325_sv2v_reg ,\nz.mem_2324_sv2v_reg ,
  \nz.mem_2323_sv2v_reg ,\nz.mem_2322_sv2v_reg ,\nz.mem_2321_sv2v_reg ,\nz.mem_2320_sv2v_reg ,
  \nz.mem_2319_sv2v_reg ,\nz.mem_2318_sv2v_reg ,\nz.mem_2317_sv2v_reg ,
  \nz.mem_2316_sv2v_reg ,\nz.mem_2315_sv2v_reg ,\nz.mem_2314_sv2v_reg ,
  \nz.mem_2313_sv2v_reg ,\nz.mem_2312_sv2v_reg ,\nz.mem_2311_sv2v_reg ,\nz.mem_2310_sv2v_reg ,
  \nz.mem_2309_sv2v_reg ,\nz.mem_2308_sv2v_reg ,\nz.mem_2307_sv2v_reg ,
  \nz.mem_2306_sv2v_reg ,\nz.mem_2305_sv2v_reg ,\nz.mem_2304_sv2v_reg ,\nz.mem_2303_sv2v_reg ,
  \nz.mem_2302_sv2v_reg ,\nz.mem_2301_sv2v_reg ,\nz.mem_2300_sv2v_reg ,
  \nz.mem_2299_sv2v_reg ,\nz.mem_2298_sv2v_reg ,\nz.mem_2297_sv2v_reg ,\nz.mem_2296_sv2v_reg ,
  \nz.mem_2295_sv2v_reg ,\nz.mem_2294_sv2v_reg ,\nz.mem_2293_sv2v_reg ,
  \nz.mem_2292_sv2v_reg ,\nz.mem_2291_sv2v_reg ,\nz.mem_2290_sv2v_reg ,\nz.mem_2289_sv2v_reg ,
  \nz.mem_2288_sv2v_reg ,\nz.mem_2287_sv2v_reg ,\nz.mem_2286_sv2v_reg ,
  \nz.mem_2285_sv2v_reg ,\nz.mem_2284_sv2v_reg ,\nz.mem_2283_sv2v_reg ,\nz.mem_2282_sv2v_reg ,
  \nz.mem_2281_sv2v_reg ,\nz.mem_2280_sv2v_reg ,\nz.mem_2279_sv2v_reg ,
  \nz.mem_2278_sv2v_reg ,\nz.mem_2277_sv2v_reg ,\nz.mem_2276_sv2v_reg ,\nz.mem_2275_sv2v_reg ,
  \nz.mem_2274_sv2v_reg ,\nz.mem_2273_sv2v_reg ,\nz.mem_2272_sv2v_reg ,
  \nz.mem_2271_sv2v_reg ,\nz.mem_2270_sv2v_reg ,\nz.mem_2269_sv2v_reg ,\nz.mem_2268_sv2v_reg ,
  \nz.mem_2267_sv2v_reg ,\nz.mem_2266_sv2v_reg ,\nz.mem_2265_sv2v_reg ,
  \nz.mem_2264_sv2v_reg ,\nz.mem_2263_sv2v_reg ,\nz.mem_2262_sv2v_reg ,\nz.mem_2261_sv2v_reg ,
  \nz.mem_2260_sv2v_reg ,\nz.mem_2259_sv2v_reg ,\nz.mem_2258_sv2v_reg ,
  \nz.mem_2257_sv2v_reg ,\nz.mem_2256_sv2v_reg ,\nz.mem_2255_sv2v_reg ,\nz.mem_2254_sv2v_reg ,
  \nz.mem_2253_sv2v_reg ,\nz.mem_2252_sv2v_reg ,\nz.mem_2251_sv2v_reg ,
  \nz.mem_2250_sv2v_reg ,\nz.mem_2249_sv2v_reg ,\nz.mem_2248_sv2v_reg ,\nz.mem_2247_sv2v_reg ,
  \nz.mem_2246_sv2v_reg ,\nz.mem_2245_sv2v_reg ,\nz.mem_2244_sv2v_reg ,
  \nz.mem_2243_sv2v_reg ,\nz.mem_2242_sv2v_reg ,\nz.mem_2241_sv2v_reg ,\nz.mem_2240_sv2v_reg ,
  \nz.mem_2239_sv2v_reg ,\nz.mem_2238_sv2v_reg ,\nz.mem_2237_sv2v_reg ,
  \nz.mem_2236_sv2v_reg ,\nz.mem_2235_sv2v_reg ,\nz.mem_2234_sv2v_reg ,
  \nz.mem_2233_sv2v_reg ,\nz.mem_2232_sv2v_reg ,\nz.mem_2231_sv2v_reg ,\nz.mem_2230_sv2v_reg ,
  \nz.mem_2229_sv2v_reg ,\nz.mem_2228_sv2v_reg ,\nz.mem_2227_sv2v_reg ,
  \nz.mem_2226_sv2v_reg ,\nz.mem_2225_sv2v_reg ,\nz.mem_2224_sv2v_reg ,\nz.mem_2223_sv2v_reg ,
  \nz.mem_2222_sv2v_reg ,\nz.mem_2221_sv2v_reg ,\nz.mem_2220_sv2v_reg ,
  \nz.mem_2219_sv2v_reg ,\nz.mem_2218_sv2v_reg ,\nz.mem_2217_sv2v_reg ,\nz.mem_2216_sv2v_reg ,
  \nz.mem_2215_sv2v_reg ,\nz.mem_2214_sv2v_reg ,\nz.mem_2213_sv2v_reg ,
  \nz.mem_2212_sv2v_reg ,\nz.mem_2211_sv2v_reg ,\nz.mem_2210_sv2v_reg ,\nz.mem_2209_sv2v_reg ,
  \nz.mem_2208_sv2v_reg ,\nz.mem_2207_sv2v_reg ,\nz.mem_2206_sv2v_reg ,
  \nz.mem_2205_sv2v_reg ,\nz.mem_2204_sv2v_reg ,\nz.mem_2203_sv2v_reg ,\nz.mem_2202_sv2v_reg ,
  \nz.mem_2201_sv2v_reg ,\nz.mem_2200_sv2v_reg ,\nz.mem_2199_sv2v_reg ,
  \nz.mem_2198_sv2v_reg ,\nz.mem_2197_sv2v_reg ,\nz.mem_2196_sv2v_reg ,\nz.mem_2195_sv2v_reg ,
  \nz.mem_2194_sv2v_reg ,\nz.mem_2193_sv2v_reg ,\nz.mem_2192_sv2v_reg ,
  \nz.mem_2191_sv2v_reg ,\nz.mem_2190_sv2v_reg ,\nz.mem_2189_sv2v_reg ,\nz.mem_2188_sv2v_reg ,
  \nz.mem_2187_sv2v_reg ,\nz.mem_2186_sv2v_reg ,\nz.mem_2185_sv2v_reg ,
  \nz.mem_2184_sv2v_reg ,\nz.mem_2183_sv2v_reg ,\nz.mem_2182_sv2v_reg ,\nz.mem_2181_sv2v_reg ,
  \nz.mem_2180_sv2v_reg ,\nz.mem_2179_sv2v_reg ,\nz.mem_2178_sv2v_reg ,
  \nz.mem_2177_sv2v_reg ,\nz.mem_2176_sv2v_reg ,\nz.mem_2175_sv2v_reg ,\nz.mem_2174_sv2v_reg ,
  \nz.mem_2173_sv2v_reg ,\nz.mem_2172_sv2v_reg ,\nz.mem_2171_sv2v_reg ,
  \nz.mem_2170_sv2v_reg ,\nz.mem_2169_sv2v_reg ,\nz.mem_2168_sv2v_reg ,\nz.mem_2167_sv2v_reg ,
  \nz.mem_2166_sv2v_reg ,\nz.mem_2165_sv2v_reg ,\nz.mem_2164_sv2v_reg ,
  \nz.mem_2163_sv2v_reg ,\nz.mem_2162_sv2v_reg ,\nz.mem_2161_sv2v_reg ,\nz.mem_2160_sv2v_reg ,
  \nz.mem_2159_sv2v_reg ,\nz.mem_2158_sv2v_reg ,\nz.mem_2157_sv2v_reg ,
  \nz.mem_2156_sv2v_reg ,\nz.mem_2155_sv2v_reg ,\nz.mem_2154_sv2v_reg ,
  \nz.mem_2153_sv2v_reg ,\nz.mem_2152_sv2v_reg ,\nz.mem_2151_sv2v_reg ,\nz.mem_2150_sv2v_reg ,
  \nz.mem_2149_sv2v_reg ,\nz.mem_2148_sv2v_reg ,\nz.mem_2147_sv2v_reg ,
  \nz.mem_2146_sv2v_reg ,\nz.mem_2145_sv2v_reg ,\nz.mem_2144_sv2v_reg ,\nz.mem_2143_sv2v_reg ,
  \nz.mem_2142_sv2v_reg ,\nz.mem_2141_sv2v_reg ,\nz.mem_2140_sv2v_reg ,
  \nz.mem_2139_sv2v_reg ,\nz.mem_2138_sv2v_reg ,\nz.mem_2137_sv2v_reg ,\nz.mem_2136_sv2v_reg ,
  \nz.mem_2135_sv2v_reg ,\nz.mem_2134_sv2v_reg ,\nz.mem_2133_sv2v_reg ,
  \nz.mem_2132_sv2v_reg ,\nz.mem_2131_sv2v_reg ,\nz.mem_2130_sv2v_reg ,\nz.mem_2129_sv2v_reg ,
  \nz.mem_2128_sv2v_reg ,\nz.mem_2127_sv2v_reg ,\nz.mem_2126_sv2v_reg ,
  \nz.mem_2125_sv2v_reg ,\nz.mem_2124_sv2v_reg ,\nz.mem_2123_sv2v_reg ,\nz.mem_2122_sv2v_reg ,
  \nz.mem_2121_sv2v_reg ,\nz.mem_2120_sv2v_reg ,\nz.mem_2119_sv2v_reg ,
  \nz.mem_2118_sv2v_reg ,\nz.mem_2117_sv2v_reg ,\nz.mem_2116_sv2v_reg ,\nz.mem_2115_sv2v_reg ,
  \nz.mem_2114_sv2v_reg ,\nz.mem_2113_sv2v_reg ,\nz.mem_2112_sv2v_reg ,
  \nz.mem_2111_sv2v_reg ,\nz.mem_2110_sv2v_reg ,\nz.mem_2109_sv2v_reg ,\nz.mem_2108_sv2v_reg ,
  \nz.mem_2107_sv2v_reg ,\nz.mem_2106_sv2v_reg ,\nz.mem_2105_sv2v_reg ,
  \nz.mem_2104_sv2v_reg ,\nz.mem_2103_sv2v_reg ,\nz.mem_2102_sv2v_reg ,\nz.mem_2101_sv2v_reg ,
  \nz.mem_2100_sv2v_reg ,\nz.mem_2099_sv2v_reg ,\nz.mem_2098_sv2v_reg ,
  \nz.mem_2097_sv2v_reg ,\nz.mem_2096_sv2v_reg ,\nz.mem_2095_sv2v_reg ,\nz.mem_2094_sv2v_reg ,
  \nz.mem_2093_sv2v_reg ,\nz.mem_2092_sv2v_reg ,\nz.mem_2091_sv2v_reg ,
  \nz.mem_2090_sv2v_reg ,\nz.mem_2089_sv2v_reg ,\nz.mem_2088_sv2v_reg ,\nz.mem_2087_sv2v_reg ,
  \nz.mem_2086_sv2v_reg ,\nz.mem_2085_sv2v_reg ,\nz.mem_2084_sv2v_reg ,
  \nz.mem_2083_sv2v_reg ,\nz.mem_2082_sv2v_reg ,\nz.mem_2081_sv2v_reg ,\nz.mem_2080_sv2v_reg ,
  \nz.mem_2079_sv2v_reg ,\nz.mem_2078_sv2v_reg ,\nz.mem_2077_sv2v_reg ,
  \nz.mem_2076_sv2v_reg ,\nz.mem_2075_sv2v_reg ,\nz.mem_2074_sv2v_reg ,
  \nz.mem_2073_sv2v_reg ,\nz.mem_2072_sv2v_reg ,\nz.mem_2071_sv2v_reg ,\nz.mem_2070_sv2v_reg ,
  \nz.mem_2069_sv2v_reg ,\nz.mem_2068_sv2v_reg ,\nz.mem_2067_sv2v_reg ,
  \nz.mem_2066_sv2v_reg ,\nz.mem_2065_sv2v_reg ,\nz.mem_2064_sv2v_reg ,\nz.mem_2063_sv2v_reg ,
  \nz.mem_2062_sv2v_reg ,\nz.mem_2061_sv2v_reg ,\nz.mem_2060_sv2v_reg ,
  \nz.mem_2059_sv2v_reg ,\nz.mem_2058_sv2v_reg ,\nz.mem_2057_sv2v_reg ,\nz.mem_2056_sv2v_reg ,
  \nz.mem_2055_sv2v_reg ,\nz.mem_2054_sv2v_reg ,\nz.mem_2053_sv2v_reg ,
  \nz.mem_2052_sv2v_reg ,\nz.mem_2051_sv2v_reg ,\nz.mem_2050_sv2v_reg ,\nz.mem_2049_sv2v_reg ,
  \nz.mem_2048_sv2v_reg ,\nz.mem_2047_sv2v_reg ,\nz.mem_2046_sv2v_reg ,
  \nz.mem_2045_sv2v_reg ,\nz.mem_2044_sv2v_reg ,\nz.mem_2043_sv2v_reg ,\nz.mem_2042_sv2v_reg ,
  \nz.mem_2041_sv2v_reg ,\nz.mem_2040_sv2v_reg ,\nz.mem_2039_sv2v_reg ,
  \nz.mem_2038_sv2v_reg ,\nz.mem_2037_sv2v_reg ,\nz.mem_2036_sv2v_reg ,\nz.mem_2035_sv2v_reg ,
  \nz.mem_2034_sv2v_reg ,\nz.mem_2033_sv2v_reg ,\nz.mem_2032_sv2v_reg ,
  \nz.mem_2031_sv2v_reg ,\nz.mem_2030_sv2v_reg ,\nz.mem_2029_sv2v_reg ,\nz.mem_2028_sv2v_reg ,
  \nz.mem_2027_sv2v_reg ,\nz.mem_2026_sv2v_reg ,\nz.mem_2025_sv2v_reg ,
  \nz.mem_2024_sv2v_reg ,\nz.mem_2023_sv2v_reg ,\nz.mem_2022_sv2v_reg ,\nz.mem_2021_sv2v_reg ,
  \nz.mem_2020_sv2v_reg ,\nz.mem_2019_sv2v_reg ,\nz.mem_2018_sv2v_reg ,
  \nz.mem_2017_sv2v_reg ,\nz.mem_2016_sv2v_reg ,\nz.mem_2015_sv2v_reg ,\nz.mem_2014_sv2v_reg ,
  \nz.mem_2013_sv2v_reg ,\nz.mem_2012_sv2v_reg ,\nz.mem_2011_sv2v_reg ,
  \nz.mem_2010_sv2v_reg ,\nz.mem_2009_sv2v_reg ,\nz.mem_2008_sv2v_reg ,\nz.mem_2007_sv2v_reg ,
  \nz.mem_2006_sv2v_reg ,\nz.mem_2005_sv2v_reg ,\nz.mem_2004_sv2v_reg ,
  \nz.mem_2003_sv2v_reg ,\nz.mem_2002_sv2v_reg ,\nz.mem_2001_sv2v_reg ,\nz.mem_2000_sv2v_reg ,
  \nz.mem_1999_sv2v_reg ,\nz.mem_1998_sv2v_reg ,\nz.mem_1997_sv2v_reg ,
  \nz.mem_1996_sv2v_reg ,\nz.mem_1995_sv2v_reg ,\nz.mem_1994_sv2v_reg ,
  \nz.mem_1993_sv2v_reg ,\nz.mem_1992_sv2v_reg ,\nz.mem_1991_sv2v_reg ,\nz.mem_1990_sv2v_reg ,
  \nz.mem_1989_sv2v_reg ,\nz.mem_1988_sv2v_reg ,\nz.mem_1987_sv2v_reg ,
  \nz.mem_1986_sv2v_reg ,\nz.mem_1985_sv2v_reg ,\nz.mem_1984_sv2v_reg ,\nz.mem_1983_sv2v_reg ,
  \nz.mem_1982_sv2v_reg ,\nz.mem_1981_sv2v_reg ,\nz.mem_1980_sv2v_reg ,
  \nz.mem_1979_sv2v_reg ,\nz.mem_1978_sv2v_reg ,\nz.mem_1977_sv2v_reg ,\nz.mem_1976_sv2v_reg ,
  \nz.mem_1975_sv2v_reg ,\nz.mem_1974_sv2v_reg ,\nz.mem_1973_sv2v_reg ,
  \nz.mem_1972_sv2v_reg ,\nz.mem_1971_sv2v_reg ,\nz.mem_1970_sv2v_reg ,\nz.mem_1969_sv2v_reg ,
  \nz.mem_1968_sv2v_reg ,\nz.mem_1967_sv2v_reg ,\nz.mem_1966_sv2v_reg ,
  \nz.mem_1965_sv2v_reg ,\nz.mem_1964_sv2v_reg ,\nz.mem_1963_sv2v_reg ,\nz.mem_1962_sv2v_reg ,
  \nz.mem_1961_sv2v_reg ,\nz.mem_1960_sv2v_reg ,\nz.mem_1959_sv2v_reg ,
  \nz.mem_1958_sv2v_reg ,\nz.mem_1957_sv2v_reg ,\nz.mem_1956_sv2v_reg ,\nz.mem_1955_sv2v_reg ,
  \nz.mem_1954_sv2v_reg ,\nz.mem_1953_sv2v_reg ,\nz.mem_1952_sv2v_reg ,
  \nz.mem_1951_sv2v_reg ,\nz.mem_1950_sv2v_reg ,\nz.mem_1949_sv2v_reg ,\nz.mem_1948_sv2v_reg ,
  \nz.mem_1947_sv2v_reg ,\nz.mem_1946_sv2v_reg ,\nz.mem_1945_sv2v_reg ,
  \nz.mem_1944_sv2v_reg ,\nz.mem_1943_sv2v_reg ,\nz.mem_1942_sv2v_reg ,\nz.mem_1941_sv2v_reg ,
  \nz.mem_1940_sv2v_reg ,\nz.mem_1939_sv2v_reg ,\nz.mem_1938_sv2v_reg ,
  \nz.mem_1937_sv2v_reg ,\nz.mem_1936_sv2v_reg ,\nz.mem_1935_sv2v_reg ,\nz.mem_1934_sv2v_reg ,
  \nz.mem_1933_sv2v_reg ,\nz.mem_1932_sv2v_reg ,\nz.mem_1931_sv2v_reg ,
  \nz.mem_1930_sv2v_reg ,\nz.mem_1929_sv2v_reg ,\nz.mem_1928_sv2v_reg ,\nz.mem_1927_sv2v_reg ,
  \nz.mem_1926_sv2v_reg ,\nz.mem_1925_sv2v_reg ,\nz.mem_1924_sv2v_reg ,
  \nz.mem_1923_sv2v_reg ,\nz.mem_1922_sv2v_reg ,\nz.mem_1921_sv2v_reg ,\nz.mem_1920_sv2v_reg ,
  \nz.mem_1919_sv2v_reg ,\nz.mem_1918_sv2v_reg ,\nz.mem_1917_sv2v_reg ,
  \nz.mem_1916_sv2v_reg ,\nz.mem_1915_sv2v_reg ,\nz.mem_1914_sv2v_reg ,
  \nz.mem_1913_sv2v_reg ,\nz.mem_1912_sv2v_reg ,\nz.mem_1911_sv2v_reg ,\nz.mem_1910_sv2v_reg ,
  \nz.mem_1909_sv2v_reg ,\nz.mem_1908_sv2v_reg ,\nz.mem_1907_sv2v_reg ,
  \nz.mem_1906_sv2v_reg ,\nz.mem_1905_sv2v_reg ,\nz.mem_1904_sv2v_reg ,\nz.mem_1903_sv2v_reg ,
  \nz.mem_1902_sv2v_reg ,\nz.mem_1901_sv2v_reg ,\nz.mem_1900_sv2v_reg ,
  \nz.mem_1899_sv2v_reg ,\nz.mem_1898_sv2v_reg ,\nz.mem_1897_sv2v_reg ,\nz.mem_1896_sv2v_reg ,
  \nz.mem_1895_sv2v_reg ,\nz.mem_1894_sv2v_reg ,\nz.mem_1893_sv2v_reg ,
  \nz.mem_1892_sv2v_reg ,\nz.mem_1891_sv2v_reg ,\nz.mem_1890_sv2v_reg ,\nz.mem_1889_sv2v_reg ,
  \nz.mem_1888_sv2v_reg ,\nz.mem_1887_sv2v_reg ,\nz.mem_1886_sv2v_reg ,
  \nz.mem_1885_sv2v_reg ,\nz.mem_1884_sv2v_reg ,\nz.mem_1883_sv2v_reg ,\nz.mem_1882_sv2v_reg ,
  \nz.mem_1881_sv2v_reg ,\nz.mem_1880_sv2v_reg ,\nz.mem_1879_sv2v_reg ,
  \nz.mem_1878_sv2v_reg ,\nz.mem_1877_sv2v_reg ,\nz.mem_1876_sv2v_reg ,\nz.mem_1875_sv2v_reg ,
  \nz.mem_1874_sv2v_reg ,\nz.mem_1873_sv2v_reg ,\nz.mem_1872_sv2v_reg ,
  \nz.mem_1871_sv2v_reg ,\nz.mem_1870_sv2v_reg ,\nz.mem_1869_sv2v_reg ,\nz.mem_1868_sv2v_reg ,
  \nz.mem_1867_sv2v_reg ,\nz.mem_1866_sv2v_reg ,\nz.mem_1865_sv2v_reg ,
  \nz.mem_1864_sv2v_reg ,\nz.mem_1863_sv2v_reg ,\nz.mem_1862_sv2v_reg ,\nz.mem_1861_sv2v_reg ,
  \nz.mem_1860_sv2v_reg ,\nz.mem_1859_sv2v_reg ,\nz.mem_1858_sv2v_reg ,
  \nz.mem_1857_sv2v_reg ,\nz.mem_1856_sv2v_reg ,\nz.mem_1855_sv2v_reg ,\nz.mem_1854_sv2v_reg ,
  \nz.mem_1853_sv2v_reg ,\nz.mem_1852_sv2v_reg ,\nz.mem_1851_sv2v_reg ,
  \nz.mem_1850_sv2v_reg ,\nz.mem_1849_sv2v_reg ,\nz.mem_1848_sv2v_reg ,\nz.mem_1847_sv2v_reg ,
  \nz.mem_1846_sv2v_reg ,\nz.mem_1845_sv2v_reg ,\nz.mem_1844_sv2v_reg ,
  \nz.mem_1843_sv2v_reg ,\nz.mem_1842_sv2v_reg ,\nz.mem_1841_sv2v_reg ,\nz.mem_1840_sv2v_reg ,
  \nz.mem_1839_sv2v_reg ,\nz.mem_1838_sv2v_reg ,\nz.mem_1837_sv2v_reg ,
  \nz.mem_1836_sv2v_reg ,\nz.mem_1835_sv2v_reg ,\nz.mem_1834_sv2v_reg ,
  \nz.mem_1833_sv2v_reg ,\nz.mem_1832_sv2v_reg ,\nz.mem_1831_sv2v_reg ,\nz.mem_1830_sv2v_reg ,
  \nz.mem_1829_sv2v_reg ,\nz.mem_1828_sv2v_reg ,\nz.mem_1827_sv2v_reg ,
  \nz.mem_1826_sv2v_reg ,\nz.mem_1825_sv2v_reg ,\nz.mem_1824_sv2v_reg ,\nz.mem_1823_sv2v_reg ,
  \nz.mem_1822_sv2v_reg ,\nz.mem_1821_sv2v_reg ,\nz.mem_1820_sv2v_reg ,
  \nz.mem_1819_sv2v_reg ,\nz.mem_1818_sv2v_reg ,\nz.mem_1817_sv2v_reg ,\nz.mem_1816_sv2v_reg ,
  \nz.mem_1815_sv2v_reg ,\nz.mem_1814_sv2v_reg ,\nz.mem_1813_sv2v_reg ,
  \nz.mem_1812_sv2v_reg ,\nz.mem_1811_sv2v_reg ,\nz.mem_1810_sv2v_reg ,\nz.mem_1809_sv2v_reg ,
  \nz.mem_1808_sv2v_reg ,\nz.mem_1807_sv2v_reg ,\nz.mem_1806_sv2v_reg ,
  \nz.mem_1805_sv2v_reg ,\nz.mem_1804_sv2v_reg ,\nz.mem_1803_sv2v_reg ,\nz.mem_1802_sv2v_reg ,
  \nz.mem_1801_sv2v_reg ,\nz.mem_1800_sv2v_reg ,\nz.mem_1799_sv2v_reg ,
  \nz.mem_1798_sv2v_reg ,\nz.mem_1797_sv2v_reg ,\nz.mem_1796_sv2v_reg ,\nz.mem_1795_sv2v_reg ,
  \nz.mem_1794_sv2v_reg ,\nz.mem_1793_sv2v_reg ,\nz.mem_1792_sv2v_reg ,
  \nz.mem_1791_sv2v_reg ,\nz.mem_1790_sv2v_reg ,\nz.mem_1789_sv2v_reg ,\nz.mem_1788_sv2v_reg ,
  \nz.mem_1787_sv2v_reg ,\nz.mem_1786_sv2v_reg ,\nz.mem_1785_sv2v_reg ,
  \nz.mem_1784_sv2v_reg ,\nz.mem_1783_sv2v_reg ,\nz.mem_1782_sv2v_reg ,\nz.mem_1781_sv2v_reg ,
  \nz.mem_1780_sv2v_reg ,\nz.mem_1779_sv2v_reg ,\nz.mem_1778_sv2v_reg ,
  \nz.mem_1777_sv2v_reg ,\nz.mem_1776_sv2v_reg ,\nz.mem_1775_sv2v_reg ,\nz.mem_1774_sv2v_reg ,
  \nz.mem_1773_sv2v_reg ,\nz.mem_1772_sv2v_reg ,\nz.mem_1771_sv2v_reg ,
  \nz.mem_1770_sv2v_reg ,\nz.mem_1769_sv2v_reg ,\nz.mem_1768_sv2v_reg ,\nz.mem_1767_sv2v_reg ,
  \nz.mem_1766_sv2v_reg ,\nz.mem_1765_sv2v_reg ,\nz.mem_1764_sv2v_reg ,
  \nz.mem_1763_sv2v_reg ,\nz.mem_1762_sv2v_reg ,\nz.mem_1761_sv2v_reg ,\nz.mem_1760_sv2v_reg ,
  \nz.mem_1759_sv2v_reg ,\nz.mem_1758_sv2v_reg ,\nz.mem_1757_sv2v_reg ,
  \nz.mem_1756_sv2v_reg ,\nz.mem_1755_sv2v_reg ,\nz.mem_1754_sv2v_reg ,
  \nz.mem_1753_sv2v_reg ,\nz.mem_1752_sv2v_reg ,\nz.mem_1751_sv2v_reg ,\nz.mem_1750_sv2v_reg ,
  \nz.mem_1749_sv2v_reg ,\nz.mem_1748_sv2v_reg ,\nz.mem_1747_sv2v_reg ,
  \nz.mem_1746_sv2v_reg ,\nz.mem_1745_sv2v_reg ,\nz.mem_1744_sv2v_reg ,\nz.mem_1743_sv2v_reg ,
  \nz.mem_1742_sv2v_reg ,\nz.mem_1741_sv2v_reg ,\nz.mem_1740_sv2v_reg ,
  \nz.mem_1739_sv2v_reg ,\nz.mem_1738_sv2v_reg ,\nz.mem_1737_sv2v_reg ,\nz.mem_1736_sv2v_reg ,
  \nz.mem_1735_sv2v_reg ,\nz.mem_1734_sv2v_reg ,\nz.mem_1733_sv2v_reg ,
  \nz.mem_1732_sv2v_reg ,\nz.mem_1731_sv2v_reg ,\nz.mem_1730_sv2v_reg ,\nz.mem_1729_sv2v_reg ,
  \nz.mem_1728_sv2v_reg ,\nz.mem_1727_sv2v_reg ,\nz.mem_1726_sv2v_reg ,
  \nz.mem_1725_sv2v_reg ,\nz.mem_1724_sv2v_reg ,\nz.mem_1723_sv2v_reg ,\nz.mem_1722_sv2v_reg ,
  \nz.mem_1721_sv2v_reg ,\nz.mem_1720_sv2v_reg ,\nz.mem_1719_sv2v_reg ,
  \nz.mem_1718_sv2v_reg ,\nz.mem_1717_sv2v_reg ,\nz.mem_1716_sv2v_reg ,\nz.mem_1715_sv2v_reg ,
  \nz.mem_1714_sv2v_reg ,\nz.mem_1713_sv2v_reg ,\nz.mem_1712_sv2v_reg ,
  \nz.mem_1711_sv2v_reg ,\nz.mem_1710_sv2v_reg ,\nz.mem_1709_sv2v_reg ,\nz.mem_1708_sv2v_reg ,
  \nz.mem_1707_sv2v_reg ,\nz.mem_1706_sv2v_reg ,\nz.mem_1705_sv2v_reg ,
  \nz.mem_1704_sv2v_reg ,\nz.mem_1703_sv2v_reg ,\nz.mem_1702_sv2v_reg ,\nz.mem_1701_sv2v_reg ,
  \nz.mem_1700_sv2v_reg ,\nz.mem_1699_sv2v_reg ,\nz.mem_1698_sv2v_reg ,
  \nz.mem_1697_sv2v_reg ,\nz.mem_1696_sv2v_reg ,\nz.mem_1695_sv2v_reg ,\nz.mem_1694_sv2v_reg ,
  \nz.mem_1693_sv2v_reg ,\nz.mem_1692_sv2v_reg ,\nz.mem_1691_sv2v_reg ,
  \nz.mem_1690_sv2v_reg ,\nz.mem_1689_sv2v_reg ,\nz.mem_1688_sv2v_reg ,\nz.mem_1687_sv2v_reg ,
  \nz.mem_1686_sv2v_reg ,\nz.mem_1685_sv2v_reg ,\nz.mem_1684_sv2v_reg ,
  \nz.mem_1683_sv2v_reg ,\nz.mem_1682_sv2v_reg ,\nz.mem_1681_sv2v_reg ,\nz.mem_1680_sv2v_reg ,
  \nz.mem_1679_sv2v_reg ,\nz.mem_1678_sv2v_reg ,\nz.mem_1677_sv2v_reg ,
  \nz.mem_1676_sv2v_reg ,\nz.mem_1675_sv2v_reg ,\nz.mem_1674_sv2v_reg ,
  \nz.mem_1673_sv2v_reg ,\nz.mem_1672_sv2v_reg ,\nz.mem_1671_sv2v_reg ,\nz.mem_1670_sv2v_reg ,
  \nz.mem_1669_sv2v_reg ,\nz.mem_1668_sv2v_reg ,\nz.mem_1667_sv2v_reg ,
  \nz.mem_1666_sv2v_reg ,\nz.mem_1665_sv2v_reg ,\nz.mem_1664_sv2v_reg ,\nz.mem_1663_sv2v_reg ,
  \nz.mem_1662_sv2v_reg ,\nz.mem_1661_sv2v_reg ,\nz.mem_1660_sv2v_reg ,
  \nz.mem_1659_sv2v_reg ,\nz.mem_1658_sv2v_reg ,\nz.mem_1657_sv2v_reg ,\nz.mem_1656_sv2v_reg ,
  \nz.mem_1655_sv2v_reg ,\nz.mem_1654_sv2v_reg ,\nz.mem_1653_sv2v_reg ,
  \nz.mem_1652_sv2v_reg ,\nz.mem_1651_sv2v_reg ,\nz.mem_1650_sv2v_reg ,\nz.mem_1649_sv2v_reg ,
  \nz.mem_1648_sv2v_reg ,\nz.mem_1647_sv2v_reg ,\nz.mem_1646_sv2v_reg ,
  \nz.mem_1645_sv2v_reg ,\nz.mem_1644_sv2v_reg ,\nz.mem_1643_sv2v_reg ,\nz.mem_1642_sv2v_reg ,
  \nz.mem_1641_sv2v_reg ,\nz.mem_1640_sv2v_reg ,\nz.mem_1639_sv2v_reg ,
  \nz.mem_1638_sv2v_reg ,\nz.mem_1637_sv2v_reg ,\nz.mem_1636_sv2v_reg ,\nz.mem_1635_sv2v_reg ,
  \nz.mem_1634_sv2v_reg ,\nz.mem_1633_sv2v_reg ,\nz.mem_1632_sv2v_reg ,
  \nz.mem_1631_sv2v_reg ,\nz.mem_1630_sv2v_reg ,\nz.mem_1629_sv2v_reg ,\nz.mem_1628_sv2v_reg ,
  \nz.mem_1627_sv2v_reg ,\nz.mem_1626_sv2v_reg ,\nz.mem_1625_sv2v_reg ,
  \nz.mem_1624_sv2v_reg ,\nz.mem_1623_sv2v_reg ,\nz.mem_1622_sv2v_reg ,\nz.mem_1621_sv2v_reg ,
  \nz.mem_1620_sv2v_reg ,\nz.mem_1619_sv2v_reg ,\nz.mem_1618_sv2v_reg ,
  \nz.mem_1617_sv2v_reg ,\nz.mem_1616_sv2v_reg ,\nz.mem_1615_sv2v_reg ,\nz.mem_1614_sv2v_reg ,
  \nz.mem_1613_sv2v_reg ,\nz.mem_1612_sv2v_reg ,\nz.mem_1611_sv2v_reg ,
  \nz.mem_1610_sv2v_reg ,\nz.mem_1609_sv2v_reg ,\nz.mem_1608_sv2v_reg ,\nz.mem_1607_sv2v_reg ,
  \nz.mem_1606_sv2v_reg ,\nz.mem_1605_sv2v_reg ,\nz.mem_1604_sv2v_reg ,
  \nz.mem_1603_sv2v_reg ,\nz.mem_1602_sv2v_reg ,\nz.mem_1601_sv2v_reg ,\nz.mem_1600_sv2v_reg ,
  \nz.mem_1599_sv2v_reg ,\nz.mem_1598_sv2v_reg ,\nz.mem_1597_sv2v_reg ,
  \nz.mem_1596_sv2v_reg ,\nz.mem_1595_sv2v_reg ,\nz.mem_1594_sv2v_reg ,
  \nz.mem_1593_sv2v_reg ,\nz.mem_1592_sv2v_reg ,\nz.mem_1591_sv2v_reg ,\nz.mem_1590_sv2v_reg ,
  \nz.mem_1589_sv2v_reg ,\nz.mem_1588_sv2v_reg ,\nz.mem_1587_sv2v_reg ,
  \nz.mem_1586_sv2v_reg ,\nz.mem_1585_sv2v_reg ,\nz.mem_1584_sv2v_reg ,\nz.mem_1583_sv2v_reg ,
  \nz.mem_1582_sv2v_reg ,\nz.mem_1581_sv2v_reg ,\nz.mem_1580_sv2v_reg ,
  \nz.mem_1579_sv2v_reg ,\nz.mem_1578_sv2v_reg ,\nz.mem_1577_sv2v_reg ,\nz.mem_1576_sv2v_reg ,
  \nz.mem_1575_sv2v_reg ,\nz.mem_1574_sv2v_reg ,\nz.mem_1573_sv2v_reg ,
  \nz.mem_1572_sv2v_reg ,\nz.mem_1571_sv2v_reg ,\nz.mem_1570_sv2v_reg ,\nz.mem_1569_sv2v_reg ,
  \nz.mem_1568_sv2v_reg ,\nz.mem_1567_sv2v_reg ,\nz.mem_1566_sv2v_reg ,
  \nz.mem_1565_sv2v_reg ,\nz.mem_1564_sv2v_reg ,\nz.mem_1563_sv2v_reg ,\nz.mem_1562_sv2v_reg ,
  \nz.mem_1561_sv2v_reg ,\nz.mem_1560_sv2v_reg ,\nz.mem_1559_sv2v_reg ,
  \nz.mem_1558_sv2v_reg ,\nz.mem_1557_sv2v_reg ,\nz.mem_1556_sv2v_reg ,\nz.mem_1555_sv2v_reg ,
  \nz.mem_1554_sv2v_reg ,\nz.mem_1553_sv2v_reg ,\nz.mem_1552_sv2v_reg ,
  \nz.mem_1551_sv2v_reg ,\nz.mem_1550_sv2v_reg ,\nz.mem_1549_sv2v_reg ,\nz.mem_1548_sv2v_reg ,
  \nz.mem_1547_sv2v_reg ,\nz.mem_1546_sv2v_reg ,\nz.mem_1545_sv2v_reg ,
  \nz.mem_1544_sv2v_reg ,\nz.mem_1543_sv2v_reg ,\nz.mem_1542_sv2v_reg ,\nz.mem_1541_sv2v_reg ,
  \nz.mem_1540_sv2v_reg ,\nz.mem_1539_sv2v_reg ,\nz.mem_1538_sv2v_reg ,
  \nz.mem_1537_sv2v_reg ,\nz.mem_1536_sv2v_reg ,\nz.mem_1535_sv2v_reg ,\nz.mem_1534_sv2v_reg ,
  \nz.mem_1533_sv2v_reg ,\nz.mem_1532_sv2v_reg ,\nz.mem_1531_sv2v_reg ,
  \nz.mem_1530_sv2v_reg ,\nz.mem_1529_sv2v_reg ,\nz.mem_1528_sv2v_reg ,\nz.mem_1527_sv2v_reg ,
  \nz.mem_1526_sv2v_reg ,\nz.mem_1525_sv2v_reg ,\nz.mem_1524_sv2v_reg ,
  \nz.mem_1523_sv2v_reg ,\nz.mem_1522_sv2v_reg ,\nz.mem_1521_sv2v_reg ,\nz.mem_1520_sv2v_reg ,
  \nz.mem_1519_sv2v_reg ,\nz.mem_1518_sv2v_reg ,\nz.mem_1517_sv2v_reg ,
  \nz.mem_1516_sv2v_reg ,\nz.mem_1515_sv2v_reg ,\nz.mem_1514_sv2v_reg ,
  \nz.mem_1513_sv2v_reg ,\nz.mem_1512_sv2v_reg ,\nz.mem_1511_sv2v_reg ,\nz.mem_1510_sv2v_reg ,
  \nz.mem_1509_sv2v_reg ,\nz.mem_1508_sv2v_reg ,\nz.mem_1507_sv2v_reg ,
  \nz.mem_1506_sv2v_reg ,\nz.mem_1505_sv2v_reg ,\nz.mem_1504_sv2v_reg ,\nz.mem_1503_sv2v_reg ,
  \nz.mem_1502_sv2v_reg ,\nz.mem_1501_sv2v_reg ,\nz.mem_1500_sv2v_reg ,
  \nz.mem_1499_sv2v_reg ,\nz.mem_1498_sv2v_reg ,\nz.mem_1497_sv2v_reg ,\nz.mem_1496_sv2v_reg ,
  \nz.mem_1495_sv2v_reg ,\nz.mem_1494_sv2v_reg ,\nz.mem_1493_sv2v_reg ,
  \nz.mem_1492_sv2v_reg ,\nz.mem_1491_sv2v_reg ,\nz.mem_1490_sv2v_reg ,\nz.mem_1489_sv2v_reg ,
  \nz.mem_1488_sv2v_reg ,\nz.mem_1487_sv2v_reg ,\nz.mem_1486_sv2v_reg ,
  \nz.mem_1485_sv2v_reg ,\nz.mem_1484_sv2v_reg ,\nz.mem_1483_sv2v_reg ,\nz.mem_1482_sv2v_reg ,
  \nz.mem_1481_sv2v_reg ,\nz.mem_1480_sv2v_reg ,\nz.mem_1479_sv2v_reg ,
  \nz.mem_1478_sv2v_reg ,\nz.mem_1477_sv2v_reg ,\nz.mem_1476_sv2v_reg ,\nz.mem_1475_sv2v_reg ,
  \nz.mem_1474_sv2v_reg ,\nz.mem_1473_sv2v_reg ,\nz.mem_1472_sv2v_reg ,
  \nz.mem_1471_sv2v_reg ,\nz.mem_1470_sv2v_reg ,\nz.mem_1469_sv2v_reg ,\nz.mem_1468_sv2v_reg ,
  \nz.mem_1467_sv2v_reg ,\nz.mem_1466_sv2v_reg ,\nz.mem_1465_sv2v_reg ,
  \nz.mem_1464_sv2v_reg ,\nz.mem_1463_sv2v_reg ,\nz.mem_1462_sv2v_reg ,\nz.mem_1461_sv2v_reg ,
  \nz.mem_1460_sv2v_reg ,\nz.mem_1459_sv2v_reg ,\nz.mem_1458_sv2v_reg ,
  \nz.mem_1457_sv2v_reg ,\nz.mem_1456_sv2v_reg ,\nz.mem_1455_sv2v_reg ,\nz.mem_1454_sv2v_reg ,
  \nz.mem_1453_sv2v_reg ,\nz.mem_1452_sv2v_reg ,\nz.mem_1451_sv2v_reg ,
  \nz.mem_1450_sv2v_reg ,\nz.mem_1449_sv2v_reg ,\nz.mem_1448_sv2v_reg ,\nz.mem_1447_sv2v_reg ,
  \nz.mem_1446_sv2v_reg ,\nz.mem_1445_sv2v_reg ,\nz.mem_1444_sv2v_reg ,
  \nz.mem_1443_sv2v_reg ,\nz.mem_1442_sv2v_reg ,\nz.mem_1441_sv2v_reg ,\nz.mem_1440_sv2v_reg ,
  \nz.mem_1439_sv2v_reg ,\nz.mem_1438_sv2v_reg ,\nz.mem_1437_sv2v_reg ,
  \nz.mem_1436_sv2v_reg ,\nz.mem_1435_sv2v_reg ,\nz.mem_1434_sv2v_reg ,
  \nz.mem_1433_sv2v_reg ,\nz.mem_1432_sv2v_reg ,\nz.mem_1431_sv2v_reg ,\nz.mem_1430_sv2v_reg ,
  \nz.mem_1429_sv2v_reg ,\nz.mem_1428_sv2v_reg ,\nz.mem_1427_sv2v_reg ,
  \nz.mem_1426_sv2v_reg ,\nz.mem_1425_sv2v_reg ,\nz.mem_1424_sv2v_reg ,\nz.mem_1423_sv2v_reg ,
  \nz.mem_1422_sv2v_reg ,\nz.mem_1421_sv2v_reg ,\nz.mem_1420_sv2v_reg ,
  \nz.mem_1419_sv2v_reg ,\nz.mem_1418_sv2v_reg ,\nz.mem_1417_sv2v_reg ,\nz.mem_1416_sv2v_reg ,
  \nz.mem_1415_sv2v_reg ,\nz.mem_1414_sv2v_reg ,\nz.mem_1413_sv2v_reg ,
  \nz.mem_1412_sv2v_reg ,\nz.mem_1411_sv2v_reg ,\nz.mem_1410_sv2v_reg ,\nz.mem_1409_sv2v_reg ,
  \nz.mem_1408_sv2v_reg ,\nz.mem_1407_sv2v_reg ,\nz.mem_1406_sv2v_reg ,
  \nz.mem_1405_sv2v_reg ,\nz.mem_1404_sv2v_reg ,\nz.mem_1403_sv2v_reg ,\nz.mem_1402_sv2v_reg ,
  \nz.mem_1401_sv2v_reg ,\nz.mem_1400_sv2v_reg ,\nz.mem_1399_sv2v_reg ,
  \nz.mem_1398_sv2v_reg ,\nz.mem_1397_sv2v_reg ,\nz.mem_1396_sv2v_reg ,\nz.mem_1395_sv2v_reg ,
  \nz.mem_1394_sv2v_reg ,\nz.mem_1393_sv2v_reg ,\nz.mem_1392_sv2v_reg ,
  \nz.mem_1391_sv2v_reg ,\nz.mem_1390_sv2v_reg ,\nz.mem_1389_sv2v_reg ,\nz.mem_1388_sv2v_reg ,
  \nz.mem_1387_sv2v_reg ,\nz.mem_1386_sv2v_reg ,\nz.mem_1385_sv2v_reg ,
  \nz.mem_1384_sv2v_reg ,\nz.mem_1383_sv2v_reg ,\nz.mem_1382_sv2v_reg ,\nz.mem_1381_sv2v_reg ,
  \nz.mem_1380_sv2v_reg ,\nz.mem_1379_sv2v_reg ,\nz.mem_1378_sv2v_reg ,
  \nz.mem_1377_sv2v_reg ,\nz.mem_1376_sv2v_reg ,\nz.mem_1375_sv2v_reg ,\nz.mem_1374_sv2v_reg ,
  \nz.mem_1373_sv2v_reg ,\nz.mem_1372_sv2v_reg ,\nz.mem_1371_sv2v_reg ,
  \nz.mem_1370_sv2v_reg ,\nz.mem_1369_sv2v_reg ,\nz.mem_1368_sv2v_reg ,\nz.mem_1367_sv2v_reg ,
  \nz.mem_1366_sv2v_reg ,\nz.mem_1365_sv2v_reg ,\nz.mem_1364_sv2v_reg ,
  \nz.mem_1363_sv2v_reg ,\nz.mem_1362_sv2v_reg ,\nz.mem_1361_sv2v_reg ,\nz.mem_1360_sv2v_reg ,
  \nz.mem_1359_sv2v_reg ,\nz.mem_1358_sv2v_reg ,\nz.mem_1357_sv2v_reg ,
  \nz.mem_1356_sv2v_reg ,\nz.mem_1355_sv2v_reg ,\nz.mem_1354_sv2v_reg ,
  \nz.mem_1353_sv2v_reg ,\nz.mem_1352_sv2v_reg ,\nz.mem_1351_sv2v_reg ,\nz.mem_1350_sv2v_reg ,
  \nz.mem_1349_sv2v_reg ,\nz.mem_1348_sv2v_reg ,\nz.mem_1347_sv2v_reg ,
  \nz.mem_1346_sv2v_reg ,\nz.mem_1345_sv2v_reg ,\nz.mem_1344_sv2v_reg ,\nz.mem_1343_sv2v_reg ,
  \nz.mem_1342_sv2v_reg ,\nz.mem_1341_sv2v_reg ,\nz.mem_1340_sv2v_reg ,
  \nz.mem_1339_sv2v_reg ,\nz.mem_1338_sv2v_reg ,\nz.mem_1337_sv2v_reg ,\nz.mem_1336_sv2v_reg ,
  \nz.mem_1335_sv2v_reg ,\nz.mem_1334_sv2v_reg ,\nz.mem_1333_sv2v_reg ,
  \nz.mem_1332_sv2v_reg ,\nz.mem_1331_sv2v_reg ,\nz.mem_1330_sv2v_reg ,\nz.mem_1329_sv2v_reg ,
  \nz.mem_1328_sv2v_reg ,\nz.mem_1327_sv2v_reg ,\nz.mem_1326_sv2v_reg ,
  \nz.mem_1325_sv2v_reg ,\nz.mem_1324_sv2v_reg ,\nz.mem_1323_sv2v_reg ,\nz.mem_1322_sv2v_reg ,
  \nz.mem_1321_sv2v_reg ,\nz.mem_1320_sv2v_reg ,\nz.mem_1319_sv2v_reg ,
  \nz.mem_1318_sv2v_reg ,\nz.mem_1317_sv2v_reg ,\nz.mem_1316_sv2v_reg ,\nz.mem_1315_sv2v_reg ,
  \nz.mem_1314_sv2v_reg ,\nz.mem_1313_sv2v_reg ,\nz.mem_1312_sv2v_reg ,
  \nz.mem_1311_sv2v_reg ,\nz.mem_1310_sv2v_reg ,\nz.mem_1309_sv2v_reg ,\nz.mem_1308_sv2v_reg ,
  \nz.mem_1307_sv2v_reg ,\nz.mem_1306_sv2v_reg ,\nz.mem_1305_sv2v_reg ,
  \nz.mem_1304_sv2v_reg ,\nz.mem_1303_sv2v_reg ,\nz.mem_1302_sv2v_reg ,\nz.mem_1301_sv2v_reg ,
  \nz.mem_1300_sv2v_reg ,\nz.mem_1299_sv2v_reg ,\nz.mem_1298_sv2v_reg ,
  \nz.mem_1297_sv2v_reg ,\nz.mem_1296_sv2v_reg ,\nz.mem_1295_sv2v_reg ,\nz.mem_1294_sv2v_reg ,
  \nz.mem_1293_sv2v_reg ,\nz.mem_1292_sv2v_reg ,\nz.mem_1291_sv2v_reg ,
  \nz.mem_1290_sv2v_reg ,\nz.mem_1289_sv2v_reg ,\nz.mem_1288_sv2v_reg ,\nz.mem_1287_sv2v_reg ,
  \nz.mem_1286_sv2v_reg ,\nz.mem_1285_sv2v_reg ,\nz.mem_1284_sv2v_reg ,
  \nz.mem_1283_sv2v_reg ,\nz.mem_1282_sv2v_reg ,\nz.mem_1281_sv2v_reg ,\nz.mem_1280_sv2v_reg ,
  \nz.mem_1279_sv2v_reg ,\nz.mem_1278_sv2v_reg ,\nz.mem_1277_sv2v_reg ,
  \nz.mem_1276_sv2v_reg ,\nz.mem_1275_sv2v_reg ,\nz.mem_1274_sv2v_reg ,
  \nz.mem_1273_sv2v_reg ,\nz.mem_1272_sv2v_reg ,\nz.mem_1271_sv2v_reg ,\nz.mem_1270_sv2v_reg ,
  \nz.mem_1269_sv2v_reg ,\nz.mem_1268_sv2v_reg ,\nz.mem_1267_sv2v_reg ,
  \nz.mem_1266_sv2v_reg ,\nz.mem_1265_sv2v_reg ,\nz.mem_1264_sv2v_reg ,\nz.mem_1263_sv2v_reg ,
  \nz.mem_1262_sv2v_reg ,\nz.mem_1261_sv2v_reg ,\nz.mem_1260_sv2v_reg ,
  \nz.mem_1259_sv2v_reg ,\nz.mem_1258_sv2v_reg ,\nz.mem_1257_sv2v_reg ,\nz.mem_1256_sv2v_reg ,
  \nz.mem_1255_sv2v_reg ,\nz.mem_1254_sv2v_reg ,\nz.mem_1253_sv2v_reg ,
  \nz.mem_1252_sv2v_reg ,\nz.mem_1251_sv2v_reg ,\nz.mem_1250_sv2v_reg ,\nz.mem_1249_sv2v_reg ,
  \nz.mem_1248_sv2v_reg ,\nz.mem_1247_sv2v_reg ,\nz.mem_1246_sv2v_reg ,
  \nz.mem_1245_sv2v_reg ,\nz.mem_1244_sv2v_reg ,\nz.mem_1243_sv2v_reg ,\nz.mem_1242_sv2v_reg ,
  \nz.mem_1241_sv2v_reg ,\nz.mem_1240_sv2v_reg ,\nz.mem_1239_sv2v_reg ,
  \nz.mem_1238_sv2v_reg ,\nz.mem_1237_sv2v_reg ,\nz.mem_1236_sv2v_reg ,\nz.mem_1235_sv2v_reg ,
  \nz.mem_1234_sv2v_reg ,\nz.mem_1233_sv2v_reg ,\nz.mem_1232_sv2v_reg ,
  \nz.mem_1231_sv2v_reg ,\nz.mem_1230_sv2v_reg ,\nz.mem_1229_sv2v_reg ,\nz.mem_1228_sv2v_reg ,
  \nz.mem_1227_sv2v_reg ,\nz.mem_1226_sv2v_reg ,\nz.mem_1225_sv2v_reg ,
  \nz.mem_1224_sv2v_reg ,\nz.mem_1223_sv2v_reg ,\nz.mem_1222_sv2v_reg ,\nz.mem_1221_sv2v_reg ,
  \nz.mem_1220_sv2v_reg ,\nz.mem_1219_sv2v_reg ,\nz.mem_1218_sv2v_reg ,
  \nz.mem_1217_sv2v_reg ,\nz.mem_1216_sv2v_reg ,\nz.mem_1215_sv2v_reg ,\nz.mem_1214_sv2v_reg ,
  \nz.mem_1213_sv2v_reg ,\nz.mem_1212_sv2v_reg ,\nz.mem_1211_sv2v_reg ,
  \nz.mem_1210_sv2v_reg ,\nz.mem_1209_sv2v_reg ,\nz.mem_1208_sv2v_reg ,\nz.mem_1207_sv2v_reg ,
  \nz.mem_1206_sv2v_reg ,\nz.mem_1205_sv2v_reg ,\nz.mem_1204_sv2v_reg ,
  \nz.mem_1203_sv2v_reg ,\nz.mem_1202_sv2v_reg ,\nz.mem_1201_sv2v_reg ,\nz.mem_1200_sv2v_reg ,
  \nz.mem_1199_sv2v_reg ,\nz.mem_1198_sv2v_reg ,\nz.mem_1197_sv2v_reg ,
  \nz.mem_1196_sv2v_reg ,\nz.mem_1195_sv2v_reg ,\nz.mem_1194_sv2v_reg ,
  \nz.mem_1193_sv2v_reg ,\nz.mem_1192_sv2v_reg ,\nz.mem_1191_sv2v_reg ,\nz.mem_1190_sv2v_reg ,
  \nz.mem_1189_sv2v_reg ,\nz.mem_1188_sv2v_reg ,\nz.mem_1187_sv2v_reg ,
  \nz.mem_1186_sv2v_reg ,\nz.mem_1185_sv2v_reg ,\nz.mem_1184_sv2v_reg ,\nz.mem_1183_sv2v_reg ,
  \nz.mem_1182_sv2v_reg ,\nz.mem_1181_sv2v_reg ,\nz.mem_1180_sv2v_reg ,
  \nz.mem_1179_sv2v_reg ,\nz.mem_1178_sv2v_reg ,\nz.mem_1177_sv2v_reg ,\nz.mem_1176_sv2v_reg ,
  \nz.mem_1175_sv2v_reg ,\nz.mem_1174_sv2v_reg ,\nz.mem_1173_sv2v_reg ,
  \nz.mem_1172_sv2v_reg ,\nz.mem_1171_sv2v_reg ,\nz.mem_1170_sv2v_reg ,\nz.mem_1169_sv2v_reg ,
  \nz.mem_1168_sv2v_reg ,\nz.mem_1167_sv2v_reg ,\nz.mem_1166_sv2v_reg ,
  \nz.mem_1165_sv2v_reg ,\nz.mem_1164_sv2v_reg ,\nz.mem_1163_sv2v_reg ,\nz.mem_1162_sv2v_reg ,
  \nz.mem_1161_sv2v_reg ,\nz.mem_1160_sv2v_reg ,\nz.mem_1159_sv2v_reg ,
  \nz.mem_1158_sv2v_reg ,\nz.mem_1157_sv2v_reg ,\nz.mem_1156_sv2v_reg ,\nz.mem_1155_sv2v_reg ,
  \nz.mem_1154_sv2v_reg ,\nz.mem_1153_sv2v_reg ,\nz.mem_1152_sv2v_reg ,
  \nz.mem_1151_sv2v_reg ,\nz.mem_1150_sv2v_reg ,\nz.mem_1149_sv2v_reg ,\nz.mem_1148_sv2v_reg ,
  \nz.mem_1147_sv2v_reg ,\nz.mem_1146_sv2v_reg ,\nz.mem_1145_sv2v_reg ,
  \nz.mem_1144_sv2v_reg ,\nz.mem_1143_sv2v_reg ,\nz.mem_1142_sv2v_reg ,\nz.mem_1141_sv2v_reg ,
  \nz.mem_1140_sv2v_reg ,\nz.mem_1139_sv2v_reg ,\nz.mem_1138_sv2v_reg ,
  \nz.mem_1137_sv2v_reg ,\nz.mem_1136_sv2v_reg ,\nz.mem_1135_sv2v_reg ,\nz.mem_1134_sv2v_reg ,
  \nz.mem_1133_sv2v_reg ,\nz.mem_1132_sv2v_reg ,\nz.mem_1131_sv2v_reg ,
  \nz.mem_1130_sv2v_reg ,\nz.mem_1129_sv2v_reg ,\nz.mem_1128_sv2v_reg ,\nz.mem_1127_sv2v_reg ,
  \nz.mem_1126_sv2v_reg ,\nz.mem_1125_sv2v_reg ,\nz.mem_1124_sv2v_reg ,
  \nz.mem_1123_sv2v_reg ,\nz.mem_1122_sv2v_reg ,\nz.mem_1121_sv2v_reg ,\nz.mem_1120_sv2v_reg ,
  \nz.mem_1119_sv2v_reg ,\nz.mem_1118_sv2v_reg ,\nz.mem_1117_sv2v_reg ,
  \nz.mem_1116_sv2v_reg ,\nz.mem_1115_sv2v_reg ,\nz.mem_1114_sv2v_reg ,
  \nz.mem_1113_sv2v_reg ,\nz.mem_1112_sv2v_reg ,\nz.mem_1111_sv2v_reg ,\nz.mem_1110_sv2v_reg ,
  \nz.mem_1109_sv2v_reg ,\nz.mem_1108_sv2v_reg ,\nz.mem_1107_sv2v_reg ,
  \nz.mem_1106_sv2v_reg ,\nz.mem_1105_sv2v_reg ,\nz.mem_1104_sv2v_reg ,\nz.mem_1103_sv2v_reg ,
  \nz.mem_1102_sv2v_reg ,\nz.mem_1101_sv2v_reg ,\nz.mem_1100_sv2v_reg ,
  \nz.mem_1099_sv2v_reg ,\nz.mem_1098_sv2v_reg ,\nz.mem_1097_sv2v_reg ,\nz.mem_1096_sv2v_reg ,
  \nz.mem_1095_sv2v_reg ,\nz.mem_1094_sv2v_reg ,\nz.mem_1093_sv2v_reg ,
  \nz.mem_1092_sv2v_reg ,\nz.mem_1091_sv2v_reg ,\nz.mem_1090_sv2v_reg ,\nz.mem_1089_sv2v_reg ,
  \nz.mem_1088_sv2v_reg ,\nz.mem_1087_sv2v_reg ,\nz.mem_1086_sv2v_reg ,
  \nz.mem_1085_sv2v_reg ,\nz.mem_1084_sv2v_reg ,\nz.mem_1083_sv2v_reg ,\nz.mem_1082_sv2v_reg ,
  \nz.mem_1081_sv2v_reg ,\nz.mem_1080_sv2v_reg ,\nz.mem_1079_sv2v_reg ,
  \nz.mem_1078_sv2v_reg ,\nz.mem_1077_sv2v_reg ,\nz.mem_1076_sv2v_reg ,\nz.mem_1075_sv2v_reg ,
  \nz.mem_1074_sv2v_reg ,\nz.mem_1073_sv2v_reg ,\nz.mem_1072_sv2v_reg ,
  \nz.mem_1071_sv2v_reg ,\nz.mem_1070_sv2v_reg ,\nz.mem_1069_sv2v_reg ,\nz.mem_1068_sv2v_reg ,
  \nz.mem_1067_sv2v_reg ,\nz.mem_1066_sv2v_reg ,\nz.mem_1065_sv2v_reg ,
  \nz.mem_1064_sv2v_reg ,\nz.mem_1063_sv2v_reg ,\nz.mem_1062_sv2v_reg ,\nz.mem_1061_sv2v_reg ,
  \nz.mem_1060_sv2v_reg ,\nz.mem_1059_sv2v_reg ,\nz.mem_1058_sv2v_reg ,
  \nz.mem_1057_sv2v_reg ,\nz.mem_1056_sv2v_reg ,\nz.mem_1055_sv2v_reg ,\nz.mem_1054_sv2v_reg ,
  \nz.mem_1053_sv2v_reg ,\nz.mem_1052_sv2v_reg ,\nz.mem_1051_sv2v_reg ,
  \nz.mem_1050_sv2v_reg ,\nz.mem_1049_sv2v_reg ,\nz.mem_1048_sv2v_reg ,\nz.mem_1047_sv2v_reg ,
  \nz.mem_1046_sv2v_reg ,\nz.mem_1045_sv2v_reg ,\nz.mem_1044_sv2v_reg ,
  \nz.mem_1043_sv2v_reg ,\nz.mem_1042_sv2v_reg ,\nz.mem_1041_sv2v_reg ,\nz.mem_1040_sv2v_reg ,
  \nz.mem_1039_sv2v_reg ,\nz.mem_1038_sv2v_reg ,\nz.mem_1037_sv2v_reg ,
  \nz.mem_1036_sv2v_reg ,\nz.mem_1035_sv2v_reg ,\nz.mem_1034_sv2v_reg ,
  \nz.mem_1033_sv2v_reg ,\nz.mem_1032_sv2v_reg ,\nz.mem_1031_sv2v_reg ,\nz.mem_1030_sv2v_reg ,
  \nz.mem_1029_sv2v_reg ,\nz.mem_1028_sv2v_reg ,\nz.mem_1027_sv2v_reg ,
  \nz.mem_1026_sv2v_reg ,\nz.mem_1025_sv2v_reg ,\nz.mem_1024_sv2v_reg ,\nz.mem_1023_sv2v_reg ,
  \nz.mem_1022_sv2v_reg ,\nz.mem_1021_sv2v_reg ,\nz.mem_1020_sv2v_reg ,
  \nz.mem_1019_sv2v_reg ,\nz.mem_1018_sv2v_reg ,\nz.mem_1017_sv2v_reg ,\nz.mem_1016_sv2v_reg ,
  \nz.mem_1015_sv2v_reg ,\nz.mem_1014_sv2v_reg ,\nz.mem_1013_sv2v_reg ,
  \nz.mem_1012_sv2v_reg ,\nz.mem_1011_sv2v_reg ,\nz.mem_1010_sv2v_reg ,\nz.mem_1009_sv2v_reg ,
  \nz.mem_1008_sv2v_reg ,\nz.mem_1007_sv2v_reg ,\nz.mem_1006_sv2v_reg ,
  \nz.mem_1005_sv2v_reg ,\nz.mem_1004_sv2v_reg ,\nz.mem_1003_sv2v_reg ,\nz.mem_1002_sv2v_reg ,
  \nz.mem_1001_sv2v_reg ,\nz.mem_1000_sv2v_reg ,\nz.mem_999_sv2v_reg ,
  \nz.mem_998_sv2v_reg ,\nz.mem_997_sv2v_reg ,\nz.mem_996_sv2v_reg ,\nz.mem_995_sv2v_reg ,
  \nz.mem_994_sv2v_reg ,\nz.mem_993_sv2v_reg ,\nz.mem_992_sv2v_reg ,\nz.mem_991_sv2v_reg ,
  \nz.mem_990_sv2v_reg ,\nz.mem_989_sv2v_reg ,\nz.mem_988_sv2v_reg ,
  \nz.mem_987_sv2v_reg ,\nz.mem_986_sv2v_reg ,\nz.mem_985_sv2v_reg ,\nz.mem_984_sv2v_reg ,
  \nz.mem_983_sv2v_reg ,\nz.mem_982_sv2v_reg ,\nz.mem_981_sv2v_reg ,\nz.mem_980_sv2v_reg ,
  \nz.mem_979_sv2v_reg ,\nz.mem_978_sv2v_reg ,\nz.mem_977_sv2v_reg ,
  \nz.mem_976_sv2v_reg ,\nz.mem_975_sv2v_reg ,\nz.mem_974_sv2v_reg ,\nz.mem_973_sv2v_reg ,
  \nz.mem_972_sv2v_reg ,\nz.mem_971_sv2v_reg ,\nz.mem_970_sv2v_reg ,
  \nz.mem_969_sv2v_reg ,\nz.mem_968_sv2v_reg ,\nz.mem_967_sv2v_reg ,\nz.mem_966_sv2v_reg ,
  \nz.mem_965_sv2v_reg ,\nz.mem_964_sv2v_reg ,\nz.mem_963_sv2v_reg ,\nz.mem_962_sv2v_reg ,
  \nz.mem_961_sv2v_reg ,\nz.mem_960_sv2v_reg ,\nz.mem_959_sv2v_reg ,
  \nz.mem_958_sv2v_reg ,\nz.mem_957_sv2v_reg ,\nz.mem_956_sv2v_reg ,\nz.mem_955_sv2v_reg ,
  \nz.mem_954_sv2v_reg ,\nz.mem_953_sv2v_reg ,\nz.mem_952_sv2v_reg ,\nz.mem_951_sv2v_reg ,
  \nz.mem_950_sv2v_reg ,\nz.mem_949_sv2v_reg ,\nz.mem_948_sv2v_reg ,
  \nz.mem_947_sv2v_reg ,\nz.mem_946_sv2v_reg ,\nz.mem_945_sv2v_reg ,\nz.mem_944_sv2v_reg ,
  \nz.mem_943_sv2v_reg ,\nz.mem_942_sv2v_reg ,\nz.mem_941_sv2v_reg ,\nz.mem_940_sv2v_reg ,
  \nz.mem_939_sv2v_reg ,\nz.mem_938_sv2v_reg ,\nz.mem_937_sv2v_reg ,
  \nz.mem_936_sv2v_reg ,\nz.mem_935_sv2v_reg ,\nz.mem_934_sv2v_reg ,\nz.mem_933_sv2v_reg ,
  \nz.mem_932_sv2v_reg ,\nz.mem_931_sv2v_reg ,\nz.mem_930_sv2v_reg ,
  \nz.mem_929_sv2v_reg ,\nz.mem_928_sv2v_reg ,\nz.mem_927_sv2v_reg ,\nz.mem_926_sv2v_reg ,
  \nz.mem_925_sv2v_reg ,\nz.mem_924_sv2v_reg ,\nz.mem_923_sv2v_reg ,\nz.mem_922_sv2v_reg ,
  \nz.mem_921_sv2v_reg ,\nz.mem_920_sv2v_reg ,\nz.mem_919_sv2v_reg ,
  \nz.mem_918_sv2v_reg ,\nz.mem_917_sv2v_reg ,\nz.mem_916_sv2v_reg ,\nz.mem_915_sv2v_reg ,
  \nz.mem_914_sv2v_reg ,\nz.mem_913_sv2v_reg ,\nz.mem_912_sv2v_reg ,\nz.mem_911_sv2v_reg ,
  \nz.mem_910_sv2v_reg ,\nz.mem_909_sv2v_reg ,\nz.mem_908_sv2v_reg ,
  \nz.mem_907_sv2v_reg ,\nz.mem_906_sv2v_reg ,\nz.mem_905_sv2v_reg ,\nz.mem_904_sv2v_reg ,
  \nz.mem_903_sv2v_reg ,\nz.mem_902_sv2v_reg ,\nz.mem_901_sv2v_reg ,\nz.mem_900_sv2v_reg ,
  \nz.mem_899_sv2v_reg ,\nz.mem_898_sv2v_reg ,\nz.mem_897_sv2v_reg ,
  \nz.mem_896_sv2v_reg ,\nz.mem_895_sv2v_reg ,\nz.mem_894_sv2v_reg ,\nz.mem_893_sv2v_reg ,
  \nz.mem_892_sv2v_reg ,\nz.mem_891_sv2v_reg ,\nz.mem_890_sv2v_reg ,
  \nz.mem_889_sv2v_reg ,\nz.mem_888_sv2v_reg ,\nz.mem_887_sv2v_reg ,\nz.mem_886_sv2v_reg ,
  \nz.mem_885_sv2v_reg ,\nz.mem_884_sv2v_reg ,\nz.mem_883_sv2v_reg ,\nz.mem_882_sv2v_reg ,
  \nz.mem_881_sv2v_reg ,\nz.mem_880_sv2v_reg ,\nz.mem_879_sv2v_reg ,
  \nz.mem_878_sv2v_reg ,\nz.mem_877_sv2v_reg ,\nz.mem_876_sv2v_reg ,\nz.mem_875_sv2v_reg ,
  \nz.mem_874_sv2v_reg ,\nz.mem_873_sv2v_reg ,\nz.mem_872_sv2v_reg ,\nz.mem_871_sv2v_reg ,
  \nz.mem_870_sv2v_reg ,\nz.mem_869_sv2v_reg ,\nz.mem_868_sv2v_reg ,
  \nz.mem_867_sv2v_reg ,\nz.mem_866_sv2v_reg ,\nz.mem_865_sv2v_reg ,\nz.mem_864_sv2v_reg ,
  \nz.mem_863_sv2v_reg ,\nz.mem_862_sv2v_reg ,\nz.mem_861_sv2v_reg ,\nz.mem_860_sv2v_reg ,
  \nz.mem_859_sv2v_reg ,\nz.mem_858_sv2v_reg ,\nz.mem_857_sv2v_reg ,
  \nz.mem_856_sv2v_reg ,\nz.mem_855_sv2v_reg ,\nz.mem_854_sv2v_reg ,\nz.mem_853_sv2v_reg ,
  \nz.mem_852_sv2v_reg ,\nz.mem_851_sv2v_reg ,\nz.mem_850_sv2v_reg ,
  \nz.mem_849_sv2v_reg ,\nz.mem_848_sv2v_reg ,\nz.mem_847_sv2v_reg ,\nz.mem_846_sv2v_reg ,
  \nz.mem_845_sv2v_reg ,\nz.mem_844_sv2v_reg ,\nz.mem_843_sv2v_reg ,\nz.mem_842_sv2v_reg ,
  \nz.mem_841_sv2v_reg ,\nz.mem_840_sv2v_reg ,\nz.mem_839_sv2v_reg ,
  \nz.mem_838_sv2v_reg ,\nz.mem_837_sv2v_reg ,\nz.mem_836_sv2v_reg ,\nz.mem_835_sv2v_reg ,
  \nz.mem_834_sv2v_reg ,\nz.mem_833_sv2v_reg ,\nz.mem_832_sv2v_reg ,\nz.mem_831_sv2v_reg ,
  \nz.mem_830_sv2v_reg ,\nz.mem_829_sv2v_reg ,\nz.mem_828_sv2v_reg ,
  \nz.mem_827_sv2v_reg ,\nz.mem_826_sv2v_reg ,\nz.mem_825_sv2v_reg ,\nz.mem_824_sv2v_reg ,
  \nz.mem_823_sv2v_reg ,\nz.mem_822_sv2v_reg ,\nz.mem_821_sv2v_reg ,\nz.mem_820_sv2v_reg ,
  \nz.mem_819_sv2v_reg ,\nz.mem_818_sv2v_reg ,\nz.mem_817_sv2v_reg ,
  \nz.mem_816_sv2v_reg ,\nz.mem_815_sv2v_reg ,\nz.mem_814_sv2v_reg ,\nz.mem_813_sv2v_reg ,
  \nz.mem_812_sv2v_reg ,\nz.mem_811_sv2v_reg ,\nz.mem_810_sv2v_reg ,
  \nz.mem_809_sv2v_reg ,\nz.mem_808_sv2v_reg ,\nz.mem_807_sv2v_reg ,\nz.mem_806_sv2v_reg ,
  \nz.mem_805_sv2v_reg ,\nz.mem_804_sv2v_reg ,\nz.mem_803_sv2v_reg ,\nz.mem_802_sv2v_reg ,
  \nz.mem_801_sv2v_reg ,\nz.mem_800_sv2v_reg ,\nz.mem_799_sv2v_reg ,
  \nz.mem_798_sv2v_reg ,\nz.mem_797_sv2v_reg ,\nz.mem_796_sv2v_reg ,\nz.mem_795_sv2v_reg ,
  \nz.mem_794_sv2v_reg ,\nz.mem_793_sv2v_reg ,\nz.mem_792_sv2v_reg ,\nz.mem_791_sv2v_reg ,
  \nz.mem_790_sv2v_reg ,\nz.mem_789_sv2v_reg ,\nz.mem_788_sv2v_reg ,
  \nz.mem_787_sv2v_reg ,\nz.mem_786_sv2v_reg ,\nz.mem_785_sv2v_reg ,\nz.mem_784_sv2v_reg ,
  \nz.mem_783_sv2v_reg ,\nz.mem_782_sv2v_reg ,\nz.mem_781_sv2v_reg ,\nz.mem_780_sv2v_reg ,
  \nz.mem_779_sv2v_reg ,\nz.mem_778_sv2v_reg ,\nz.mem_777_sv2v_reg ,
  \nz.mem_776_sv2v_reg ,\nz.mem_775_sv2v_reg ,\nz.mem_774_sv2v_reg ,\nz.mem_773_sv2v_reg ,
  \nz.mem_772_sv2v_reg ,\nz.mem_771_sv2v_reg ,\nz.mem_770_sv2v_reg ,
  \nz.mem_769_sv2v_reg ,\nz.mem_768_sv2v_reg ,\nz.mem_767_sv2v_reg ,\nz.mem_766_sv2v_reg ,
  \nz.mem_765_sv2v_reg ,\nz.mem_764_sv2v_reg ,\nz.mem_763_sv2v_reg ,\nz.mem_762_sv2v_reg ,
  \nz.mem_761_sv2v_reg ,\nz.mem_760_sv2v_reg ,\nz.mem_759_sv2v_reg ,
  \nz.mem_758_sv2v_reg ,\nz.mem_757_sv2v_reg ,\nz.mem_756_sv2v_reg ,\nz.mem_755_sv2v_reg ,
  \nz.mem_754_sv2v_reg ,\nz.mem_753_sv2v_reg ,\nz.mem_752_sv2v_reg ,\nz.mem_751_sv2v_reg ,
  \nz.mem_750_sv2v_reg ,\nz.mem_749_sv2v_reg ,\nz.mem_748_sv2v_reg ,
  \nz.mem_747_sv2v_reg ,\nz.mem_746_sv2v_reg ,\nz.mem_745_sv2v_reg ,\nz.mem_744_sv2v_reg ,
  \nz.mem_743_sv2v_reg ,\nz.mem_742_sv2v_reg ,\nz.mem_741_sv2v_reg ,\nz.mem_740_sv2v_reg ,
  \nz.mem_739_sv2v_reg ,\nz.mem_738_sv2v_reg ,\nz.mem_737_sv2v_reg ,
  \nz.mem_736_sv2v_reg ,\nz.mem_735_sv2v_reg ,\nz.mem_734_sv2v_reg ,\nz.mem_733_sv2v_reg ,
  \nz.mem_732_sv2v_reg ,\nz.mem_731_sv2v_reg ,\nz.mem_730_sv2v_reg ,
  \nz.mem_729_sv2v_reg ,\nz.mem_728_sv2v_reg ,\nz.mem_727_sv2v_reg ,\nz.mem_726_sv2v_reg ,
  \nz.mem_725_sv2v_reg ,\nz.mem_724_sv2v_reg ,\nz.mem_723_sv2v_reg ,\nz.mem_722_sv2v_reg ,
  \nz.mem_721_sv2v_reg ,\nz.mem_720_sv2v_reg ,\nz.mem_719_sv2v_reg ,
  \nz.mem_718_sv2v_reg ,\nz.mem_717_sv2v_reg ,\nz.mem_716_sv2v_reg ,\nz.mem_715_sv2v_reg ,
  \nz.mem_714_sv2v_reg ,\nz.mem_713_sv2v_reg ,\nz.mem_712_sv2v_reg ,\nz.mem_711_sv2v_reg ,
  \nz.mem_710_sv2v_reg ,\nz.mem_709_sv2v_reg ,\nz.mem_708_sv2v_reg ,
  \nz.mem_707_sv2v_reg ,\nz.mem_706_sv2v_reg ,\nz.mem_705_sv2v_reg ,\nz.mem_704_sv2v_reg ,
  \nz.mem_703_sv2v_reg ,\nz.mem_702_sv2v_reg ,\nz.mem_701_sv2v_reg ,\nz.mem_700_sv2v_reg ,
  \nz.mem_699_sv2v_reg ,\nz.mem_698_sv2v_reg ,\nz.mem_697_sv2v_reg ,
  \nz.mem_696_sv2v_reg ,\nz.mem_695_sv2v_reg ,\nz.mem_694_sv2v_reg ,\nz.mem_693_sv2v_reg ,
  \nz.mem_692_sv2v_reg ,\nz.mem_691_sv2v_reg ,\nz.mem_690_sv2v_reg ,
  \nz.mem_689_sv2v_reg ,\nz.mem_688_sv2v_reg ,\nz.mem_687_sv2v_reg ,\nz.mem_686_sv2v_reg ,
  \nz.mem_685_sv2v_reg ,\nz.mem_684_sv2v_reg ,\nz.mem_683_sv2v_reg ,\nz.mem_682_sv2v_reg ,
  \nz.mem_681_sv2v_reg ,\nz.mem_680_sv2v_reg ,\nz.mem_679_sv2v_reg ,
  \nz.mem_678_sv2v_reg ,\nz.mem_677_sv2v_reg ,\nz.mem_676_sv2v_reg ,\nz.mem_675_sv2v_reg ,
  \nz.mem_674_sv2v_reg ,\nz.mem_673_sv2v_reg ,\nz.mem_672_sv2v_reg ,\nz.mem_671_sv2v_reg ,
  \nz.mem_670_sv2v_reg ,\nz.mem_669_sv2v_reg ,\nz.mem_668_sv2v_reg ,
  \nz.mem_667_sv2v_reg ,\nz.mem_666_sv2v_reg ,\nz.mem_665_sv2v_reg ,\nz.mem_664_sv2v_reg ,
  \nz.mem_663_sv2v_reg ,\nz.mem_662_sv2v_reg ,\nz.mem_661_sv2v_reg ,\nz.mem_660_sv2v_reg ,
  \nz.mem_659_sv2v_reg ,\nz.mem_658_sv2v_reg ,\nz.mem_657_sv2v_reg ,
  \nz.mem_656_sv2v_reg ,\nz.mem_655_sv2v_reg ,\nz.mem_654_sv2v_reg ,\nz.mem_653_sv2v_reg ,
  \nz.mem_652_sv2v_reg ,\nz.mem_651_sv2v_reg ,\nz.mem_650_sv2v_reg ,
  \nz.mem_649_sv2v_reg ,\nz.mem_648_sv2v_reg ,\nz.mem_647_sv2v_reg ,\nz.mem_646_sv2v_reg ,
  \nz.mem_645_sv2v_reg ,\nz.mem_644_sv2v_reg ,\nz.mem_643_sv2v_reg ,\nz.mem_642_sv2v_reg ,
  \nz.mem_641_sv2v_reg ,\nz.mem_640_sv2v_reg ,\nz.mem_639_sv2v_reg ,
  \nz.mem_638_sv2v_reg ,\nz.mem_637_sv2v_reg ,\nz.mem_636_sv2v_reg ,\nz.mem_635_sv2v_reg ,
  \nz.mem_634_sv2v_reg ,\nz.mem_633_sv2v_reg ,\nz.mem_632_sv2v_reg ,\nz.mem_631_sv2v_reg ,
  \nz.mem_630_sv2v_reg ,\nz.mem_629_sv2v_reg ,\nz.mem_628_sv2v_reg ,
  \nz.mem_627_sv2v_reg ,\nz.mem_626_sv2v_reg ,\nz.mem_625_sv2v_reg ,\nz.mem_624_sv2v_reg ,
  \nz.mem_623_sv2v_reg ,\nz.mem_622_sv2v_reg ,\nz.mem_621_sv2v_reg ,\nz.mem_620_sv2v_reg ,
  \nz.mem_619_sv2v_reg ,\nz.mem_618_sv2v_reg ,\nz.mem_617_sv2v_reg ,
  \nz.mem_616_sv2v_reg ,\nz.mem_615_sv2v_reg ,\nz.mem_614_sv2v_reg ,\nz.mem_613_sv2v_reg ,
  \nz.mem_612_sv2v_reg ,\nz.mem_611_sv2v_reg ,\nz.mem_610_sv2v_reg ,
  \nz.mem_609_sv2v_reg ,\nz.mem_608_sv2v_reg ,\nz.mem_607_sv2v_reg ,\nz.mem_606_sv2v_reg ,
  \nz.mem_605_sv2v_reg ,\nz.mem_604_sv2v_reg ,\nz.mem_603_sv2v_reg ,\nz.mem_602_sv2v_reg ,
  \nz.mem_601_sv2v_reg ,\nz.mem_600_sv2v_reg ,\nz.mem_599_sv2v_reg ,
  \nz.mem_598_sv2v_reg ,\nz.mem_597_sv2v_reg ,\nz.mem_596_sv2v_reg ,\nz.mem_595_sv2v_reg ,
  \nz.mem_594_sv2v_reg ,\nz.mem_593_sv2v_reg ,\nz.mem_592_sv2v_reg ,\nz.mem_591_sv2v_reg ,
  \nz.mem_590_sv2v_reg ,\nz.mem_589_sv2v_reg ,\nz.mem_588_sv2v_reg ,
  \nz.mem_587_sv2v_reg ,\nz.mem_586_sv2v_reg ,\nz.mem_585_sv2v_reg ,\nz.mem_584_sv2v_reg ,
  \nz.mem_583_sv2v_reg ,\nz.mem_582_sv2v_reg ,\nz.mem_581_sv2v_reg ,\nz.mem_580_sv2v_reg ,
  \nz.mem_579_sv2v_reg ,\nz.mem_578_sv2v_reg ,\nz.mem_577_sv2v_reg ,
  \nz.mem_576_sv2v_reg ,\nz.mem_575_sv2v_reg ,\nz.mem_574_sv2v_reg ,\nz.mem_573_sv2v_reg ,
  \nz.mem_572_sv2v_reg ,\nz.mem_571_sv2v_reg ,\nz.mem_570_sv2v_reg ,
  \nz.mem_569_sv2v_reg ,\nz.mem_568_sv2v_reg ,\nz.mem_567_sv2v_reg ,\nz.mem_566_sv2v_reg ,
  \nz.mem_565_sv2v_reg ,\nz.mem_564_sv2v_reg ,\nz.mem_563_sv2v_reg ,\nz.mem_562_sv2v_reg ,
  \nz.mem_561_sv2v_reg ,\nz.mem_560_sv2v_reg ,\nz.mem_559_sv2v_reg ,
  \nz.mem_558_sv2v_reg ,\nz.mem_557_sv2v_reg ,\nz.mem_556_sv2v_reg ,\nz.mem_555_sv2v_reg ,
  \nz.mem_554_sv2v_reg ,\nz.mem_553_sv2v_reg ,\nz.mem_552_sv2v_reg ,\nz.mem_551_sv2v_reg ,
  \nz.mem_550_sv2v_reg ,\nz.mem_549_sv2v_reg ,\nz.mem_548_sv2v_reg ,
  \nz.mem_547_sv2v_reg ,\nz.mem_546_sv2v_reg ,\nz.mem_545_sv2v_reg ,\nz.mem_544_sv2v_reg ,
  \nz.mem_543_sv2v_reg ,\nz.mem_542_sv2v_reg ,\nz.mem_541_sv2v_reg ,\nz.mem_540_sv2v_reg ,
  \nz.mem_539_sv2v_reg ,\nz.mem_538_sv2v_reg ,\nz.mem_537_sv2v_reg ,
  \nz.mem_536_sv2v_reg ,\nz.mem_535_sv2v_reg ,\nz.mem_534_sv2v_reg ,\nz.mem_533_sv2v_reg ,
  \nz.mem_532_sv2v_reg ,\nz.mem_531_sv2v_reg ,\nz.mem_530_sv2v_reg ,
  \nz.mem_529_sv2v_reg ,\nz.mem_528_sv2v_reg ,\nz.mem_527_sv2v_reg ,\nz.mem_526_sv2v_reg ,
  \nz.mem_525_sv2v_reg ,\nz.mem_524_sv2v_reg ,\nz.mem_523_sv2v_reg ,\nz.mem_522_sv2v_reg ,
  \nz.mem_521_sv2v_reg ,\nz.mem_520_sv2v_reg ,\nz.mem_519_sv2v_reg ,
  \nz.mem_518_sv2v_reg ,\nz.mem_517_sv2v_reg ,\nz.mem_516_sv2v_reg ,\nz.mem_515_sv2v_reg ,
  \nz.mem_514_sv2v_reg ,\nz.mem_513_sv2v_reg ,\nz.mem_512_sv2v_reg ,\nz.mem_511_sv2v_reg ,
  \nz.mem_510_sv2v_reg ,\nz.mem_509_sv2v_reg ,\nz.mem_508_sv2v_reg ,
  \nz.mem_507_sv2v_reg ,\nz.mem_506_sv2v_reg ,\nz.mem_505_sv2v_reg ,\nz.mem_504_sv2v_reg ,
  \nz.mem_503_sv2v_reg ,\nz.mem_502_sv2v_reg ,\nz.mem_501_sv2v_reg ,\nz.mem_500_sv2v_reg ,
  \nz.mem_499_sv2v_reg ,\nz.mem_498_sv2v_reg ,\nz.mem_497_sv2v_reg ,
  \nz.mem_496_sv2v_reg ,\nz.mem_495_sv2v_reg ,\nz.mem_494_sv2v_reg ,\nz.mem_493_sv2v_reg ,
  \nz.mem_492_sv2v_reg ,\nz.mem_491_sv2v_reg ,\nz.mem_490_sv2v_reg ,
  \nz.mem_489_sv2v_reg ,\nz.mem_488_sv2v_reg ,\nz.mem_487_sv2v_reg ,\nz.mem_486_sv2v_reg ,
  \nz.mem_485_sv2v_reg ,\nz.mem_484_sv2v_reg ,\nz.mem_483_sv2v_reg ,\nz.mem_482_sv2v_reg ,
  \nz.mem_481_sv2v_reg ,\nz.mem_480_sv2v_reg ,\nz.mem_479_sv2v_reg ,
  \nz.mem_478_sv2v_reg ,\nz.mem_477_sv2v_reg ,\nz.mem_476_sv2v_reg ,\nz.mem_475_sv2v_reg ,
  \nz.mem_474_sv2v_reg ,\nz.mem_473_sv2v_reg ,\nz.mem_472_sv2v_reg ,\nz.mem_471_sv2v_reg ,
  \nz.mem_470_sv2v_reg ,\nz.mem_469_sv2v_reg ,\nz.mem_468_sv2v_reg ,
  \nz.mem_467_sv2v_reg ,\nz.mem_466_sv2v_reg ,\nz.mem_465_sv2v_reg ,\nz.mem_464_sv2v_reg ,
  \nz.mem_463_sv2v_reg ,\nz.mem_462_sv2v_reg ,\nz.mem_461_sv2v_reg ,\nz.mem_460_sv2v_reg ,
  \nz.mem_459_sv2v_reg ,\nz.mem_458_sv2v_reg ,\nz.mem_457_sv2v_reg ,
  \nz.mem_456_sv2v_reg ,\nz.mem_455_sv2v_reg ,\nz.mem_454_sv2v_reg ,\nz.mem_453_sv2v_reg ,
  \nz.mem_452_sv2v_reg ,\nz.mem_451_sv2v_reg ,\nz.mem_450_sv2v_reg ,
  \nz.mem_449_sv2v_reg ,\nz.mem_448_sv2v_reg ,\nz.mem_447_sv2v_reg ,\nz.mem_446_sv2v_reg ,
  \nz.mem_445_sv2v_reg ,\nz.mem_444_sv2v_reg ,\nz.mem_443_sv2v_reg ,\nz.mem_442_sv2v_reg ,
  \nz.mem_441_sv2v_reg ,\nz.mem_440_sv2v_reg ,\nz.mem_439_sv2v_reg ,
  \nz.mem_438_sv2v_reg ,\nz.mem_437_sv2v_reg ,\nz.mem_436_sv2v_reg ,\nz.mem_435_sv2v_reg ,
  \nz.mem_434_sv2v_reg ,\nz.mem_433_sv2v_reg ,\nz.mem_432_sv2v_reg ,\nz.mem_431_sv2v_reg ,
  \nz.mem_430_sv2v_reg ,\nz.mem_429_sv2v_reg ,\nz.mem_428_sv2v_reg ,
  \nz.mem_427_sv2v_reg ,\nz.mem_426_sv2v_reg ,\nz.mem_425_sv2v_reg ,\nz.mem_424_sv2v_reg ,
  \nz.mem_423_sv2v_reg ,\nz.mem_422_sv2v_reg ,\nz.mem_421_sv2v_reg ,\nz.mem_420_sv2v_reg ,
  \nz.mem_419_sv2v_reg ,\nz.mem_418_sv2v_reg ,\nz.mem_417_sv2v_reg ,
  \nz.mem_416_sv2v_reg ,\nz.mem_415_sv2v_reg ,\nz.mem_414_sv2v_reg ,\nz.mem_413_sv2v_reg ,
  \nz.mem_412_sv2v_reg ,\nz.mem_411_sv2v_reg ,\nz.mem_410_sv2v_reg ,
  \nz.mem_409_sv2v_reg ,\nz.mem_408_sv2v_reg ,\nz.mem_407_sv2v_reg ,\nz.mem_406_sv2v_reg ,
  \nz.mem_405_sv2v_reg ,\nz.mem_404_sv2v_reg ,\nz.mem_403_sv2v_reg ,\nz.mem_402_sv2v_reg ,
  \nz.mem_401_sv2v_reg ,\nz.mem_400_sv2v_reg ,\nz.mem_399_sv2v_reg ,
  \nz.mem_398_sv2v_reg ,\nz.mem_397_sv2v_reg ,\nz.mem_396_sv2v_reg ,\nz.mem_395_sv2v_reg ,
  \nz.mem_394_sv2v_reg ,\nz.mem_393_sv2v_reg ,\nz.mem_392_sv2v_reg ,\nz.mem_391_sv2v_reg ,
  \nz.mem_390_sv2v_reg ,\nz.mem_389_sv2v_reg ,\nz.mem_388_sv2v_reg ,
  \nz.mem_387_sv2v_reg ,\nz.mem_386_sv2v_reg ,\nz.mem_385_sv2v_reg ,\nz.mem_384_sv2v_reg ,
  \nz.mem_383_sv2v_reg ,\nz.mem_382_sv2v_reg ,\nz.mem_381_sv2v_reg ,\nz.mem_380_sv2v_reg ,
  \nz.mem_379_sv2v_reg ,\nz.mem_378_sv2v_reg ,\nz.mem_377_sv2v_reg ,
  \nz.mem_376_sv2v_reg ,\nz.mem_375_sv2v_reg ,\nz.mem_374_sv2v_reg ,\nz.mem_373_sv2v_reg ,
  \nz.mem_372_sv2v_reg ,\nz.mem_371_sv2v_reg ,\nz.mem_370_sv2v_reg ,
  \nz.mem_369_sv2v_reg ,\nz.mem_368_sv2v_reg ,\nz.mem_367_sv2v_reg ,\nz.mem_366_sv2v_reg ,
  \nz.mem_365_sv2v_reg ,\nz.mem_364_sv2v_reg ,\nz.mem_363_sv2v_reg ,\nz.mem_362_sv2v_reg ,
  \nz.mem_361_sv2v_reg ,\nz.mem_360_sv2v_reg ,\nz.mem_359_sv2v_reg ,
  \nz.mem_358_sv2v_reg ,\nz.mem_357_sv2v_reg ,\nz.mem_356_sv2v_reg ,\nz.mem_355_sv2v_reg ,
  \nz.mem_354_sv2v_reg ,\nz.mem_353_sv2v_reg ,\nz.mem_352_sv2v_reg ,\nz.mem_351_sv2v_reg ,
  \nz.mem_350_sv2v_reg ,\nz.mem_349_sv2v_reg ,\nz.mem_348_sv2v_reg ,
  \nz.mem_347_sv2v_reg ,\nz.mem_346_sv2v_reg ,\nz.mem_345_sv2v_reg ,\nz.mem_344_sv2v_reg ,
  \nz.mem_343_sv2v_reg ,\nz.mem_342_sv2v_reg ,\nz.mem_341_sv2v_reg ,\nz.mem_340_sv2v_reg ,
  \nz.mem_339_sv2v_reg ,\nz.mem_338_sv2v_reg ,\nz.mem_337_sv2v_reg ,
  \nz.mem_336_sv2v_reg ,\nz.mem_335_sv2v_reg ,\nz.mem_334_sv2v_reg ,\nz.mem_333_sv2v_reg ,
  \nz.mem_332_sv2v_reg ,\nz.mem_331_sv2v_reg ,\nz.mem_330_sv2v_reg ,
  \nz.mem_329_sv2v_reg ,\nz.mem_328_sv2v_reg ,\nz.mem_327_sv2v_reg ,\nz.mem_326_sv2v_reg ,
  \nz.mem_325_sv2v_reg ,\nz.mem_324_sv2v_reg ,\nz.mem_323_sv2v_reg ,\nz.mem_322_sv2v_reg ,
  \nz.mem_321_sv2v_reg ,\nz.mem_320_sv2v_reg ,\nz.mem_319_sv2v_reg ,
  \nz.mem_318_sv2v_reg ,\nz.mem_317_sv2v_reg ,\nz.mem_316_sv2v_reg ,\nz.mem_315_sv2v_reg ,
  \nz.mem_314_sv2v_reg ,\nz.mem_313_sv2v_reg ,\nz.mem_312_sv2v_reg ,\nz.mem_311_sv2v_reg ,
  \nz.mem_310_sv2v_reg ,\nz.mem_309_sv2v_reg ,\nz.mem_308_sv2v_reg ,
  \nz.mem_307_sv2v_reg ,\nz.mem_306_sv2v_reg ,\nz.mem_305_sv2v_reg ,\nz.mem_304_sv2v_reg ,
  \nz.mem_303_sv2v_reg ,\nz.mem_302_sv2v_reg ,\nz.mem_301_sv2v_reg ,\nz.mem_300_sv2v_reg ,
  \nz.mem_299_sv2v_reg ,\nz.mem_298_sv2v_reg ,\nz.mem_297_sv2v_reg ,
  \nz.mem_296_sv2v_reg ,\nz.mem_295_sv2v_reg ,\nz.mem_294_sv2v_reg ,\nz.mem_293_sv2v_reg ,
  \nz.mem_292_sv2v_reg ,\nz.mem_291_sv2v_reg ,\nz.mem_290_sv2v_reg ,
  \nz.mem_289_sv2v_reg ,\nz.mem_288_sv2v_reg ,\nz.mem_287_sv2v_reg ,\nz.mem_286_sv2v_reg ,
  \nz.mem_285_sv2v_reg ,\nz.mem_284_sv2v_reg ,\nz.mem_283_sv2v_reg ,\nz.mem_282_sv2v_reg ,
  \nz.mem_281_sv2v_reg ,\nz.mem_280_sv2v_reg ,\nz.mem_279_sv2v_reg ,
  \nz.mem_278_sv2v_reg ,\nz.mem_277_sv2v_reg ,\nz.mem_276_sv2v_reg ,\nz.mem_275_sv2v_reg ,
  \nz.mem_274_sv2v_reg ,\nz.mem_273_sv2v_reg ,\nz.mem_272_sv2v_reg ,\nz.mem_271_sv2v_reg ,
  \nz.mem_270_sv2v_reg ,\nz.mem_269_sv2v_reg ,\nz.mem_268_sv2v_reg ,
  \nz.mem_267_sv2v_reg ,\nz.mem_266_sv2v_reg ,\nz.mem_265_sv2v_reg ,\nz.mem_264_sv2v_reg ,
  \nz.mem_263_sv2v_reg ,\nz.mem_262_sv2v_reg ,\nz.mem_261_sv2v_reg ,\nz.mem_260_sv2v_reg ,
  \nz.mem_259_sv2v_reg ,\nz.mem_258_sv2v_reg ,\nz.mem_257_sv2v_reg ,
  \nz.mem_256_sv2v_reg ,\nz.mem_255_sv2v_reg ,\nz.mem_254_sv2v_reg ,\nz.mem_253_sv2v_reg ,
  \nz.mem_252_sv2v_reg ,\nz.mem_251_sv2v_reg ,\nz.mem_250_sv2v_reg ,
  \nz.mem_249_sv2v_reg ,\nz.mem_248_sv2v_reg ,\nz.mem_247_sv2v_reg ,\nz.mem_246_sv2v_reg ,
  \nz.mem_245_sv2v_reg ,\nz.mem_244_sv2v_reg ,\nz.mem_243_sv2v_reg ,\nz.mem_242_sv2v_reg ,
  \nz.mem_241_sv2v_reg ,\nz.mem_240_sv2v_reg ,\nz.mem_239_sv2v_reg ,
  \nz.mem_238_sv2v_reg ,\nz.mem_237_sv2v_reg ,\nz.mem_236_sv2v_reg ,\nz.mem_235_sv2v_reg ,
  \nz.mem_234_sv2v_reg ,\nz.mem_233_sv2v_reg ,\nz.mem_232_sv2v_reg ,\nz.mem_231_sv2v_reg ,
  \nz.mem_230_sv2v_reg ,\nz.mem_229_sv2v_reg ,\nz.mem_228_sv2v_reg ,
  \nz.mem_227_sv2v_reg ,\nz.mem_226_sv2v_reg ,\nz.mem_225_sv2v_reg ,\nz.mem_224_sv2v_reg ,
  \nz.mem_223_sv2v_reg ,\nz.mem_222_sv2v_reg ,\nz.mem_221_sv2v_reg ,\nz.mem_220_sv2v_reg ,
  \nz.mem_219_sv2v_reg ,\nz.mem_218_sv2v_reg ,\nz.mem_217_sv2v_reg ,
  \nz.mem_216_sv2v_reg ,\nz.mem_215_sv2v_reg ,\nz.mem_214_sv2v_reg ,\nz.mem_213_sv2v_reg ,
  \nz.mem_212_sv2v_reg ,\nz.mem_211_sv2v_reg ,\nz.mem_210_sv2v_reg ,
  \nz.mem_209_sv2v_reg ,\nz.mem_208_sv2v_reg ,\nz.mem_207_sv2v_reg ,\nz.mem_206_sv2v_reg ,
  \nz.mem_205_sv2v_reg ,\nz.mem_204_sv2v_reg ,\nz.mem_203_sv2v_reg ,\nz.mem_202_sv2v_reg ,
  \nz.mem_201_sv2v_reg ,\nz.mem_200_sv2v_reg ,\nz.mem_199_sv2v_reg ,
  \nz.mem_198_sv2v_reg ,\nz.mem_197_sv2v_reg ,\nz.mem_196_sv2v_reg ,\nz.mem_195_sv2v_reg ,
  \nz.mem_194_sv2v_reg ,\nz.mem_193_sv2v_reg ,\nz.mem_192_sv2v_reg ,\nz.mem_191_sv2v_reg ,
  \nz.mem_190_sv2v_reg ,\nz.mem_189_sv2v_reg ,\nz.mem_188_sv2v_reg ,
  \nz.mem_187_sv2v_reg ,\nz.mem_186_sv2v_reg ,\nz.mem_185_sv2v_reg ,\nz.mem_184_sv2v_reg ,
  \nz.mem_183_sv2v_reg ,\nz.mem_182_sv2v_reg ,\nz.mem_181_sv2v_reg ,\nz.mem_180_sv2v_reg ,
  \nz.mem_179_sv2v_reg ,\nz.mem_178_sv2v_reg ,\nz.mem_177_sv2v_reg ,
  \nz.mem_176_sv2v_reg ,\nz.mem_175_sv2v_reg ,\nz.mem_174_sv2v_reg ,\nz.mem_173_sv2v_reg ,
  \nz.mem_172_sv2v_reg ,\nz.mem_171_sv2v_reg ,\nz.mem_170_sv2v_reg ,
  \nz.mem_169_sv2v_reg ,\nz.mem_168_sv2v_reg ,\nz.mem_167_sv2v_reg ,\nz.mem_166_sv2v_reg ,
  \nz.mem_165_sv2v_reg ,\nz.mem_164_sv2v_reg ,\nz.mem_163_sv2v_reg ,\nz.mem_162_sv2v_reg ,
  \nz.mem_161_sv2v_reg ,\nz.mem_160_sv2v_reg ,\nz.mem_159_sv2v_reg ,
  \nz.mem_158_sv2v_reg ,\nz.mem_157_sv2v_reg ,\nz.mem_156_sv2v_reg ,\nz.mem_155_sv2v_reg ,
  \nz.mem_154_sv2v_reg ,\nz.mem_153_sv2v_reg ,\nz.mem_152_sv2v_reg ,\nz.mem_151_sv2v_reg ,
  \nz.mem_150_sv2v_reg ,\nz.mem_149_sv2v_reg ,\nz.mem_148_sv2v_reg ,
  \nz.mem_147_sv2v_reg ,\nz.mem_146_sv2v_reg ,\nz.mem_145_sv2v_reg ,\nz.mem_144_sv2v_reg ,
  \nz.mem_143_sv2v_reg ,\nz.mem_142_sv2v_reg ,\nz.mem_141_sv2v_reg ,\nz.mem_140_sv2v_reg ,
  \nz.mem_139_sv2v_reg ,\nz.mem_138_sv2v_reg ,\nz.mem_137_sv2v_reg ,
  \nz.mem_136_sv2v_reg ,\nz.mem_135_sv2v_reg ,\nz.mem_134_sv2v_reg ,\nz.mem_133_sv2v_reg ,
  \nz.mem_132_sv2v_reg ,\nz.mem_131_sv2v_reg ,\nz.mem_130_sv2v_reg ,
  \nz.mem_129_sv2v_reg ,\nz.mem_128_sv2v_reg ,\nz.mem_127_sv2v_reg ,\nz.mem_126_sv2v_reg ,
  \nz.mem_125_sv2v_reg ,\nz.mem_124_sv2v_reg ,\nz.mem_123_sv2v_reg ,\nz.mem_122_sv2v_reg ,
  \nz.mem_121_sv2v_reg ,\nz.mem_120_sv2v_reg ,\nz.mem_119_sv2v_reg ,
  \nz.mem_118_sv2v_reg ,\nz.mem_117_sv2v_reg ,\nz.mem_116_sv2v_reg ,\nz.mem_115_sv2v_reg ,
  \nz.mem_114_sv2v_reg ,\nz.mem_113_sv2v_reg ,\nz.mem_112_sv2v_reg ,\nz.mem_111_sv2v_reg ,
  \nz.mem_110_sv2v_reg ,\nz.mem_109_sv2v_reg ,\nz.mem_108_sv2v_reg ,
  \nz.mem_107_sv2v_reg ,\nz.mem_106_sv2v_reg ,\nz.mem_105_sv2v_reg ,\nz.mem_104_sv2v_reg ,
  \nz.mem_103_sv2v_reg ,\nz.mem_102_sv2v_reg ,\nz.mem_101_sv2v_reg ,\nz.mem_100_sv2v_reg ,
  \nz.mem_99_sv2v_reg ,\nz.mem_98_sv2v_reg ,\nz.mem_97_sv2v_reg ,
  \nz.mem_96_sv2v_reg ,\nz.mem_95_sv2v_reg ,\nz.mem_94_sv2v_reg ,\nz.mem_93_sv2v_reg ,
  \nz.mem_92_sv2v_reg ,\nz.mem_91_sv2v_reg ,\nz.mem_90_sv2v_reg ,\nz.mem_89_sv2v_reg ,
  \nz.mem_88_sv2v_reg ,\nz.mem_87_sv2v_reg ,\nz.mem_86_sv2v_reg ,\nz.mem_85_sv2v_reg ,
  \nz.mem_84_sv2v_reg ,\nz.mem_83_sv2v_reg ,\nz.mem_82_sv2v_reg ,\nz.mem_81_sv2v_reg ,
  \nz.mem_80_sv2v_reg ,\nz.mem_79_sv2v_reg ,\nz.mem_78_sv2v_reg ,
  \nz.mem_77_sv2v_reg ,\nz.mem_76_sv2v_reg ,\nz.mem_75_sv2v_reg ,\nz.mem_74_sv2v_reg ,
  \nz.mem_73_sv2v_reg ,\nz.mem_72_sv2v_reg ,\nz.mem_71_sv2v_reg ,\nz.mem_70_sv2v_reg ,
  \nz.mem_69_sv2v_reg ,\nz.mem_68_sv2v_reg ,\nz.mem_67_sv2v_reg ,\nz.mem_66_sv2v_reg ,
  \nz.mem_65_sv2v_reg ,\nz.mem_64_sv2v_reg ,\nz.mem_63_sv2v_reg ,\nz.mem_62_sv2v_reg ,
  \nz.mem_61_sv2v_reg ,\nz.mem_60_sv2v_reg ,\nz.mem_59_sv2v_reg ,
  \nz.mem_58_sv2v_reg ,\nz.mem_57_sv2v_reg ,\nz.mem_56_sv2v_reg ,\nz.mem_55_sv2v_reg ,
  \nz.mem_54_sv2v_reg ,\nz.mem_53_sv2v_reg ,\nz.mem_52_sv2v_reg ,\nz.mem_51_sv2v_reg ,
  \nz.mem_50_sv2v_reg ,\nz.mem_49_sv2v_reg ,\nz.mem_48_sv2v_reg ,\nz.mem_47_sv2v_reg ,
  \nz.mem_46_sv2v_reg ,\nz.mem_45_sv2v_reg ,\nz.mem_44_sv2v_reg ,\nz.mem_43_sv2v_reg ,
  \nz.mem_42_sv2v_reg ,\nz.mem_41_sv2v_reg ,\nz.mem_40_sv2v_reg ,
  \nz.mem_39_sv2v_reg ,\nz.mem_38_sv2v_reg ,\nz.mem_37_sv2v_reg ,\nz.mem_36_sv2v_reg ,
  \nz.mem_35_sv2v_reg ,\nz.mem_34_sv2v_reg ,\nz.mem_33_sv2v_reg ,\nz.mem_32_sv2v_reg ,
  \nz.mem_31_sv2v_reg ,\nz.mem_30_sv2v_reg ,\nz.mem_29_sv2v_reg ,\nz.mem_28_sv2v_reg ,
  \nz.mem_27_sv2v_reg ,\nz.mem_26_sv2v_reg ,\nz.mem_25_sv2v_reg ,\nz.mem_24_sv2v_reg ,
  \nz.mem_23_sv2v_reg ,\nz.mem_22_sv2v_reg ,\nz.mem_21_sv2v_reg ,\nz.mem_20_sv2v_reg ,
  \nz.mem_19_sv2v_reg ,\nz.mem_18_sv2v_reg ,\nz.mem_17_sv2v_reg ,
  \nz.mem_16_sv2v_reg ,\nz.mem_15_sv2v_reg ,\nz.mem_14_sv2v_reg ,\nz.mem_13_sv2v_reg ,
  \nz.mem_12_sv2v_reg ,\nz.mem_11_sv2v_reg ,\nz.mem_10_sv2v_reg ,\nz.mem_9_sv2v_reg ,
  \nz.mem_8_sv2v_reg ,\nz.mem_7_sv2v_reg ,\nz.mem_6_sv2v_reg ,\nz.mem_5_sv2v_reg ,
  \nz.mem_4_sv2v_reg ,\nz.mem_3_sv2v_reg ,\nz.mem_2_sv2v_reg ,\nz.mem_1_sv2v_reg ,
  \nz.mem_0_sv2v_reg ;
  assign \nz.mem [3199] = \nz.mem_3199_sv2v_reg ;
  assign \nz.mem [3198] = \nz.mem_3198_sv2v_reg ;
  assign \nz.mem [3197] = \nz.mem_3197_sv2v_reg ;
  assign \nz.mem [3196] = \nz.mem_3196_sv2v_reg ;
  assign \nz.mem [3195] = \nz.mem_3195_sv2v_reg ;
  assign \nz.mem [3194] = \nz.mem_3194_sv2v_reg ;
  assign \nz.mem [3193] = \nz.mem_3193_sv2v_reg ;
  assign \nz.mem [3192] = \nz.mem_3192_sv2v_reg ;
  assign \nz.mem [3191] = \nz.mem_3191_sv2v_reg ;
  assign \nz.mem [3190] = \nz.mem_3190_sv2v_reg ;
  assign \nz.mem [3189] = \nz.mem_3189_sv2v_reg ;
  assign \nz.mem [3188] = \nz.mem_3188_sv2v_reg ;
  assign \nz.mem [3187] = \nz.mem_3187_sv2v_reg ;
  assign \nz.mem [3186] = \nz.mem_3186_sv2v_reg ;
  assign \nz.mem [3185] = \nz.mem_3185_sv2v_reg ;
  assign \nz.mem [3184] = \nz.mem_3184_sv2v_reg ;
  assign \nz.mem [3183] = \nz.mem_3183_sv2v_reg ;
  assign \nz.mem [3182] = \nz.mem_3182_sv2v_reg ;
  assign \nz.mem [3181] = \nz.mem_3181_sv2v_reg ;
  assign \nz.mem [3180] = \nz.mem_3180_sv2v_reg ;
  assign \nz.mem [3179] = \nz.mem_3179_sv2v_reg ;
  assign \nz.mem [3178] = \nz.mem_3178_sv2v_reg ;
  assign \nz.mem [3177] = \nz.mem_3177_sv2v_reg ;
  assign \nz.mem [3176] = \nz.mem_3176_sv2v_reg ;
  assign \nz.mem [3175] = \nz.mem_3175_sv2v_reg ;
  assign \nz.mem [3174] = \nz.mem_3174_sv2v_reg ;
  assign \nz.mem [3173] = \nz.mem_3173_sv2v_reg ;
  assign \nz.mem [3172] = \nz.mem_3172_sv2v_reg ;
  assign \nz.mem [3171] = \nz.mem_3171_sv2v_reg ;
  assign \nz.mem [3170] = \nz.mem_3170_sv2v_reg ;
  assign \nz.mem [3169] = \nz.mem_3169_sv2v_reg ;
  assign \nz.mem [3168] = \nz.mem_3168_sv2v_reg ;
  assign \nz.mem [3167] = \nz.mem_3167_sv2v_reg ;
  assign \nz.mem [3166] = \nz.mem_3166_sv2v_reg ;
  assign \nz.mem [3165] = \nz.mem_3165_sv2v_reg ;
  assign \nz.mem [3164] = \nz.mem_3164_sv2v_reg ;
  assign \nz.mem [3163] = \nz.mem_3163_sv2v_reg ;
  assign \nz.mem [3162] = \nz.mem_3162_sv2v_reg ;
  assign \nz.mem [3161] = \nz.mem_3161_sv2v_reg ;
  assign \nz.mem [3160] = \nz.mem_3160_sv2v_reg ;
  assign \nz.mem [3159] = \nz.mem_3159_sv2v_reg ;
  assign \nz.mem [3158] = \nz.mem_3158_sv2v_reg ;
  assign \nz.mem [3157] = \nz.mem_3157_sv2v_reg ;
  assign \nz.mem [3156] = \nz.mem_3156_sv2v_reg ;
  assign \nz.mem [3155] = \nz.mem_3155_sv2v_reg ;
  assign \nz.mem [3154] = \nz.mem_3154_sv2v_reg ;
  assign \nz.mem [3153] = \nz.mem_3153_sv2v_reg ;
  assign \nz.mem [3152] = \nz.mem_3152_sv2v_reg ;
  assign \nz.mem [3151] = \nz.mem_3151_sv2v_reg ;
  assign \nz.mem [3150] = \nz.mem_3150_sv2v_reg ;
  assign \nz.mem [3149] = \nz.mem_3149_sv2v_reg ;
  assign \nz.mem [3148] = \nz.mem_3148_sv2v_reg ;
  assign \nz.mem [3147] = \nz.mem_3147_sv2v_reg ;
  assign \nz.mem [3146] = \nz.mem_3146_sv2v_reg ;
  assign \nz.mem [3145] = \nz.mem_3145_sv2v_reg ;
  assign \nz.mem [3144] = \nz.mem_3144_sv2v_reg ;
  assign \nz.mem [3143] = \nz.mem_3143_sv2v_reg ;
  assign \nz.mem [3142] = \nz.mem_3142_sv2v_reg ;
  assign \nz.mem [3141] = \nz.mem_3141_sv2v_reg ;
  assign \nz.mem [3140] = \nz.mem_3140_sv2v_reg ;
  assign \nz.mem [3139] = \nz.mem_3139_sv2v_reg ;
  assign \nz.mem [3138] = \nz.mem_3138_sv2v_reg ;
  assign \nz.mem [3137] = \nz.mem_3137_sv2v_reg ;
  assign \nz.mem [3136] = \nz.mem_3136_sv2v_reg ;
  assign \nz.mem [3135] = \nz.mem_3135_sv2v_reg ;
  assign \nz.mem [3134] = \nz.mem_3134_sv2v_reg ;
  assign \nz.mem [3133] = \nz.mem_3133_sv2v_reg ;
  assign \nz.mem [3132] = \nz.mem_3132_sv2v_reg ;
  assign \nz.mem [3131] = \nz.mem_3131_sv2v_reg ;
  assign \nz.mem [3130] = \nz.mem_3130_sv2v_reg ;
  assign \nz.mem [3129] = \nz.mem_3129_sv2v_reg ;
  assign \nz.mem [3128] = \nz.mem_3128_sv2v_reg ;
  assign \nz.mem [3127] = \nz.mem_3127_sv2v_reg ;
  assign \nz.mem [3126] = \nz.mem_3126_sv2v_reg ;
  assign \nz.mem [3125] = \nz.mem_3125_sv2v_reg ;
  assign \nz.mem [3124] = \nz.mem_3124_sv2v_reg ;
  assign \nz.mem [3123] = \nz.mem_3123_sv2v_reg ;
  assign \nz.mem [3122] = \nz.mem_3122_sv2v_reg ;
  assign \nz.mem [3121] = \nz.mem_3121_sv2v_reg ;
  assign \nz.mem [3120] = \nz.mem_3120_sv2v_reg ;
  assign \nz.mem [3119] = \nz.mem_3119_sv2v_reg ;
  assign \nz.mem [3118] = \nz.mem_3118_sv2v_reg ;
  assign \nz.mem [3117] = \nz.mem_3117_sv2v_reg ;
  assign \nz.mem [3116] = \nz.mem_3116_sv2v_reg ;
  assign \nz.mem [3115] = \nz.mem_3115_sv2v_reg ;
  assign \nz.mem [3114] = \nz.mem_3114_sv2v_reg ;
  assign \nz.mem [3113] = \nz.mem_3113_sv2v_reg ;
  assign \nz.mem [3112] = \nz.mem_3112_sv2v_reg ;
  assign \nz.mem [3111] = \nz.mem_3111_sv2v_reg ;
  assign \nz.mem [3110] = \nz.mem_3110_sv2v_reg ;
  assign \nz.mem [3109] = \nz.mem_3109_sv2v_reg ;
  assign \nz.mem [3108] = \nz.mem_3108_sv2v_reg ;
  assign \nz.mem [3107] = \nz.mem_3107_sv2v_reg ;
  assign \nz.mem [3106] = \nz.mem_3106_sv2v_reg ;
  assign \nz.mem [3105] = \nz.mem_3105_sv2v_reg ;
  assign \nz.mem [3104] = \nz.mem_3104_sv2v_reg ;
  assign \nz.mem [3103] = \nz.mem_3103_sv2v_reg ;
  assign \nz.mem [3102] = \nz.mem_3102_sv2v_reg ;
  assign \nz.mem [3101] = \nz.mem_3101_sv2v_reg ;
  assign \nz.mem [3100] = \nz.mem_3100_sv2v_reg ;
  assign \nz.mem [3099] = \nz.mem_3099_sv2v_reg ;
  assign \nz.mem [3098] = \nz.mem_3098_sv2v_reg ;
  assign \nz.mem [3097] = \nz.mem_3097_sv2v_reg ;
  assign \nz.mem [3096] = \nz.mem_3096_sv2v_reg ;
  assign \nz.mem [3095] = \nz.mem_3095_sv2v_reg ;
  assign \nz.mem [3094] = \nz.mem_3094_sv2v_reg ;
  assign \nz.mem [3093] = \nz.mem_3093_sv2v_reg ;
  assign \nz.mem [3092] = \nz.mem_3092_sv2v_reg ;
  assign \nz.mem [3091] = \nz.mem_3091_sv2v_reg ;
  assign \nz.mem [3090] = \nz.mem_3090_sv2v_reg ;
  assign \nz.mem [3089] = \nz.mem_3089_sv2v_reg ;
  assign \nz.mem [3088] = \nz.mem_3088_sv2v_reg ;
  assign \nz.mem [3087] = \nz.mem_3087_sv2v_reg ;
  assign \nz.mem [3086] = \nz.mem_3086_sv2v_reg ;
  assign \nz.mem [3085] = \nz.mem_3085_sv2v_reg ;
  assign \nz.mem [3084] = \nz.mem_3084_sv2v_reg ;
  assign \nz.mem [3083] = \nz.mem_3083_sv2v_reg ;
  assign \nz.mem [3082] = \nz.mem_3082_sv2v_reg ;
  assign \nz.mem [3081] = \nz.mem_3081_sv2v_reg ;
  assign \nz.mem [3080] = \nz.mem_3080_sv2v_reg ;
  assign \nz.mem [3079] = \nz.mem_3079_sv2v_reg ;
  assign \nz.mem [3078] = \nz.mem_3078_sv2v_reg ;
  assign \nz.mem [3077] = \nz.mem_3077_sv2v_reg ;
  assign \nz.mem [3076] = \nz.mem_3076_sv2v_reg ;
  assign \nz.mem [3075] = \nz.mem_3075_sv2v_reg ;
  assign \nz.mem [3074] = \nz.mem_3074_sv2v_reg ;
  assign \nz.mem [3073] = \nz.mem_3073_sv2v_reg ;
  assign \nz.mem [3072] = \nz.mem_3072_sv2v_reg ;
  assign \nz.mem [3071] = \nz.mem_3071_sv2v_reg ;
  assign \nz.mem [3070] = \nz.mem_3070_sv2v_reg ;
  assign \nz.mem [3069] = \nz.mem_3069_sv2v_reg ;
  assign \nz.mem [3068] = \nz.mem_3068_sv2v_reg ;
  assign \nz.mem [3067] = \nz.mem_3067_sv2v_reg ;
  assign \nz.mem [3066] = \nz.mem_3066_sv2v_reg ;
  assign \nz.mem [3065] = \nz.mem_3065_sv2v_reg ;
  assign \nz.mem [3064] = \nz.mem_3064_sv2v_reg ;
  assign \nz.mem [3063] = \nz.mem_3063_sv2v_reg ;
  assign \nz.mem [3062] = \nz.mem_3062_sv2v_reg ;
  assign \nz.mem [3061] = \nz.mem_3061_sv2v_reg ;
  assign \nz.mem [3060] = \nz.mem_3060_sv2v_reg ;
  assign \nz.mem [3059] = \nz.mem_3059_sv2v_reg ;
  assign \nz.mem [3058] = \nz.mem_3058_sv2v_reg ;
  assign \nz.mem [3057] = \nz.mem_3057_sv2v_reg ;
  assign \nz.mem [3056] = \nz.mem_3056_sv2v_reg ;
  assign \nz.mem [3055] = \nz.mem_3055_sv2v_reg ;
  assign \nz.mem [3054] = \nz.mem_3054_sv2v_reg ;
  assign \nz.mem [3053] = \nz.mem_3053_sv2v_reg ;
  assign \nz.mem [3052] = \nz.mem_3052_sv2v_reg ;
  assign \nz.mem [3051] = \nz.mem_3051_sv2v_reg ;
  assign \nz.mem [3050] = \nz.mem_3050_sv2v_reg ;
  assign \nz.mem [3049] = \nz.mem_3049_sv2v_reg ;
  assign \nz.mem [3048] = \nz.mem_3048_sv2v_reg ;
  assign \nz.mem [3047] = \nz.mem_3047_sv2v_reg ;
  assign \nz.mem [3046] = \nz.mem_3046_sv2v_reg ;
  assign \nz.mem [3045] = \nz.mem_3045_sv2v_reg ;
  assign \nz.mem [3044] = \nz.mem_3044_sv2v_reg ;
  assign \nz.mem [3043] = \nz.mem_3043_sv2v_reg ;
  assign \nz.mem [3042] = \nz.mem_3042_sv2v_reg ;
  assign \nz.mem [3041] = \nz.mem_3041_sv2v_reg ;
  assign \nz.mem [3040] = \nz.mem_3040_sv2v_reg ;
  assign \nz.mem [3039] = \nz.mem_3039_sv2v_reg ;
  assign \nz.mem [3038] = \nz.mem_3038_sv2v_reg ;
  assign \nz.mem [3037] = \nz.mem_3037_sv2v_reg ;
  assign \nz.mem [3036] = \nz.mem_3036_sv2v_reg ;
  assign \nz.mem [3035] = \nz.mem_3035_sv2v_reg ;
  assign \nz.mem [3034] = \nz.mem_3034_sv2v_reg ;
  assign \nz.mem [3033] = \nz.mem_3033_sv2v_reg ;
  assign \nz.mem [3032] = \nz.mem_3032_sv2v_reg ;
  assign \nz.mem [3031] = \nz.mem_3031_sv2v_reg ;
  assign \nz.mem [3030] = \nz.mem_3030_sv2v_reg ;
  assign \nz.mem [3029] = \nz.mem_3029_sv2v_reg ;
  assign \nz.mem [3028] = \nz.mem_3028_sv2v_reg ;
  assign \nz.mem [3027] = \nz.mem_3027_sv2v_reg ;
  assign \nz.mem [3026] = \nz.mem_3026_sv2v_reg ;
  assign \nz.mem [3025] = \nz.mem_3025_sv2v_reg ;
  assign \nz.mem [3024] = \nz.mem_3024_sv2v_reg ;
  assign \nz.mem [3023] = \nz.mem_3023_sv2v_reg ;
  assign \nz.mem [3022] = \nz.mem_3022_sv2v_reg ;
  assign \nz.mem [3021] = \nz.mem_3021_sv2v_reg ;
  assign \nz.mem [3020] = \nz.mem_3020_sv2v_reg ;
  assign \nz.mem [3019] = \nz.mem_3019_sv2v_reg ;
  assign \nz.mem [3018] = \nz.mem_3018_sv2v_reg ;
  assign \nz.mem [3017] = \nz.mem_3017_sv2v_reg ;
  assign \nz.mem [3016] = \nz.mem_3016_sv2v_reg ;
  assign \nz.mem [3015] = \nz.mem_3015_sv2v_reg ;
  assign \nz.mem [3014] = \nz.mem_3014_sv2v_reg ;
  assign \nz.mem [3013] = \nz.mem_3013_sv2v_reg ;
  assign \nz.mem [3012] = \nz.mem_3012_sv2v_reg ;
  assign \nz.mem [3011] = \nz.mem_3011_sv2v_reg ;
  assign \nz.mem [3010] = \nz.mem_3010_sv2v_reg ;
  assign \nz.mem [3009] = \nz.mem_3009_sv2v_reg ;
  assign \nz.mem [3008] = \nz.mem_3008_sv2v_reg ;
  assign \nz.mem [3007] = \nz.mem_3007_sv2v_reg ;
  assign \nz.mem [3006] = \nz.mem_3006_sv2v_reg ;
  assign \nz.mem [3005] = \nz.mem_3005_sv2v_reg ;
  assign \nz.mem [3004] = \nz.mem_3004_sv2v_reg ;
  assign \nz.mem [3003] = \nz.mem_3003_sv2v_reg ;
  assign \nz.mem [3002] = \nz.mem_3002_sv2v_reg ;
  assign \nz.mem [3001] = \nz.mem_3001_sv2v_reg ;
  assign \nz.mem [3000] = \nz.mem_3000_sv2v_reg ;
  assign \nz.mem [2999] = \nz.mem_2999_sv2v_reg ;
  assign \nz.mem [2998] = \nz.mem_2998_sv2v_reg ;
  assign \nz.mem [2997] = \nz.mem_2997_sv2v_reg ;
  assign \nz.mem [2996] = \nz.mem_2996_sv2v_reg ;
  assign \nz.mem [2995] = \nz.mem_2995_sv2v_reg ;
  assign \nz.mem [2994] = \nz.mem_2994_sv2v_reg ;
  assign \nz.mem [2993] = \nz.mem_2993_sv2v_reg ;
  assign \nz.mem [2992] = \nz.mem_2992_sv2v_reg ;
  assign \nz.mem [2991] = \nz.mem_2991_sv2v_reg ;
  assign \nz.mem [2990] = \nz.mem_2990_sv2v_reg ;
  assign \nz.mem [2989] = \nz.mem_2989_sv2v_reg ;
  assign \nz.mem [2988] = \nz.mem_2988_sv2v_reg ;
  assign \nz.mem [2987] = \nz.mem_2987_sv2v_reg ;
  assign \nz.mem [2986] = \nz.mem_2986_sv2v_reg ;
  assign \nz.mem [2985] = \nz.mem_2985_sv2v_reg ;
  assign \nz.mem [2984] = \nz.mem_2984_sv2v_reg ;
  assign \nz.mem [2983] = \nz.mem_2983_sv2v_reg ;
  assign \nz.mem [2982] = \nz.mem_2982_sv2v_reg ;
  assign \nz.mem [2981] = \nz.mem_2981_sv2v_reg ;
  assign \nz.mem [2980] = \nz.mem_2980_sv2v_reg ;
  assign \nz.mem [2979] = \nz.mem_2979_sv2v_reg ;
  assign \nz.mem [2978] = \nz.mem_2978_sv2v_reg ;
  assign \nz.mem [2977] = \nz.mem_2977_sv2v_reg ;
  assign \nz.mem [2976] = \nz.mem_2976_sv2v_reg ;
  assign \nz.mem [2975] = \nz.mem_2975_sv2v_reg ;
  assign \nz.mem [2974] = \nz.mem_2974_sv2v_reg ;
  assign \nz.mem [2973] = \nz.mem_2973_sv2v_reg ;
  assign \nz.mem [2972] = \nz.mem_2972_sv2v_reg ;
  assign \nz.mem [2971] = \nz.mem_2971_sv2v_reg ;
  assign \nz.mem [2970] = \nz.mem_2970_sv2v_reg ;
  assign \nz.mem [2969] = \nz.mem_2969_sv2v_reg ;
  assign \nz.mem [2968] = \nz.mem_2968_sv2v_reg ;
  assign \nz.mem [2967] = \nz.mem_2967_sv2v_reg ;
  assign \nz.mem [2966] = \nz.mem_2966_sv2v_reg ;
  assign \nz.mem [2965] = \nz.mem_2965_sv2v_reg ;
  assign \nz.mem [2964] = \nz.mem_2964_sv2v_reg ;
  assign \nz.mem [2963] = \nz.mem_2963_sv2v_reg ;
  assign \nz.mem [2962] = \nz.mem_2962_sv2v_reg ;
  assign \nz.mem [2961] = \nz.mem_2961_sv2v_reg ;
  assign \nz.mem [2960] = \nz.mem_2960_sv2v_reg ;
  assign \nz.mem [2959] = \nz.mem_2959_sv2v_reg ;
  assign \nz.mem [2958] = \nz.mem_2958_sv2v_reg ;
  assign \nz.mem [2957] = \nz.mem_2957_sv2v_reg ;
  assign \nz.mem [2956] = \nz.mem_2956_sv2v_reg ;
  assign \nz.mem [2955] = \nz.mem_2955_sv2v_reg ;
  assign \nz.mem [2954] = \nz.mem_2954_sv2v_reg ;
  assign \nz.mem [2953] = \nz.mem_2953_sv2v_reg ;
  assign \nz.mem [2952] = \nz.mem_2952_sv2v_reg ;
  assign \nz.mem [2951] = \nz.mem_2951_sv2v_reg ;
  assign \nz.mem [2950] = \nz.mem_2950_sv2v_reg ;
  assign \nz.mem [2949] = \nz.mem_2949_sv2v_reg ;
  assign \nz.mem [2948] = \nz.mem_2948_sv2v_reg ;
  assign \nz.mem [2947] = \nz.mem_2947_sv2v_reg ;
  assign \nz.mem [2946] = \nz.mem_2946_sv2v_reg ;
  assign \nz.mem [2945] = \nz.mem_2945_sv2v_reg ;
  assign \nz.mem [2944] = \nz.mem_2944_sv2v_reg ;
  assign \nz.mem [2943] = \nz.mem_2943_sv2v_reg ;
  assign \nz.mem [2942] = \nz.mem_2942_sv2v_reg ;
  assign \nz.mem [2941] = \nz.mem_2941_sv2v_reg ;
  assign \nz.mem [2940] = \nz.mem_2940_sv2v_reg ;
  assign \nz.mem [2939] = \nz.mem_2939_sv2v_reg ;
  assign \nz.mem [2938] = \nz.mem_2938_sv2v_reg ;
  assign \nz.mem [2937] = \nz.mem_2937_sv2v_reg ;
  assign \nz.mem [2936] = \nz.mem_2936_sv2v_reg ;
  assign \nz.mem [2935] = \nz.mem_2935_sv2v_reg ;
  assign \nz.mem [2934] = \nz.mem_2934_sv2v_reg ;
  assign \nz.mem [2933] = \nz.mem_2933_sv2v_reg ;
  assign \nz.mem [2932] = \nz.mem_2932_sv2v_reg ;
  assign \nz.mem [2931] = \nz.mem_2931_sv2v_reg ;
  assign \nz.mem [2930] = \nz.mem_2930_sv2v_reg ;
  assign \nz.mem [2929] = \nz.mem_2929_sv2v_reg ;
  assign \nz.mem [2928] = \nz.mem_2928_sv2v_reg ;
  assign \nz.mem [2927] = \nz.mem_2927_sv2v_reg ;
  assign \nz.mem [2926] = \nz.mem_2926_sv2v_reg ;
  assign \nz.mem [2925] = \nz.mem_2925_sv2v_reg ;
  assign \nz.mem [2924] = \nz.mem_2924_sv2v_reg ;
  assign \nz.mem [2923] = \nz.mem_2923_sv2v_reg ;
  assign \nz.mem [2922] = \nz.mem_2922_sv2v_reg ;
  assign \nz.mem [2921] = \nz.mem_2921_sv2v_reg ;
  assign \nz.mem [2920] = \nz.mem_2920_sv2v_reg ;
  assign \nz.mem [2919] = \nz.mem_2919_sv2v_reg ;
  assign \nz.mem [2918] = \nz.mem_2918_sv2v_reg ;
  assign \nz.mem [2917] = \nz.mem_2917_sv2v_reg ;
  assign \nz.mem [2916] = \nz.mem_2916_sv2v_reg ;
  assign \nz.mem [2915] = \nz.mem_2915_sv2v_reg ;
  assign \nz.mem [2914] = \nz.mem_2914_sv2v_reg ;
  assign \nz.mem [2913] = \nz.mem_2913_sv2v_reg ;
  assign \nz.mem [2912] = \nz.mem_2912_sv2v_reg ;
  assign \nz.mem [2911] = \nz.mem_2911_sv2v_reg ;
  assign \nz.mem [2910] = \nz.mem_2910_sv2v_reg ;
  assign \nz.mem [2909] = \nz.mem_2909_sv2v_reg ;
  assign \nz.mem [2908] = \nz.mem_2908_sv2v_reg ;
  assign \nz.mem [2907] = \nz.mem_2907_sv2v_reg ;
  assign \nz.mem [2906] = \nz.mem_2906_sv2v_reg ;
  assign \nz.mem [2905] = \nz.mem_2905_sv2v_reg ;
  assign \nz.mem [2904] = \nz.mem_2904_sv2v_reg ;
  assign \nz.mem [2903] = \nz.mem_2903_sv2v_reg ;
  assign \nz.mem [2902] = \nz.mem_2902_sv2v_reg ;
  assign \nz.mem [2901] = \nz.mem_2901_sv2v_reg ;
  assign \nz.mem [2900] = \nz.mem_2900_sv2v_reg ;
  assign \nz.mem [2899] = \nz.mem_2899_sv2v_reg ;
  assign \nz.mem [2898] = \nz.mem_2898_sv2v_reg ;
  assign \nz.mem [2897] = \nz.mem_2897_sv2v_reg ;
  assign \nz.mem [2896] = \nz.mem_2896_sv2v_reg ;
  assign \nz.mem [2895] = \nz.mem_2895_sv2v_reg ;
  assign \nz.mem [2894] = \nz.mem_2894_sv2v_reg ;
  assign \nz.mem [2893] = \nz.mem_2893_sv2v_reg ;
  assign \nz.mem [2892] = \nz.mem_2892_sv2v_reg ;
  assign \nz.mem [2891] = \nz.mem_2891_sv2v_reg ;
  assign \nz.mem [2890] = \nz.mem_2890_sv2v_reg ;
  assign \nz.mem [2889] = \nz.mem_2889_sv2v_reg ;
  assign \nz.mem [2888] = \nz.mem_2888_sv2v_reg ;
  assign \nz.mem [2887] = \nz.mem_2887_sv2v_reg ;
  assign \nz.mem [2886] = \nz.mem_2886_sv2v_reg ;
  assign \nz.mem [2885] = \nz.mem_2885_sv2v_reg ;
  assign \nz.mem [2884] = \nz.mem_2884_sv2v_reg ;
  assign \nz.mem [2883] = \nz.mem_2883_sv2v_reg ;
  assign \nz.mem [2882] = \nz.mem_2882_sv2v_reg ;
  assign \nz.mem [2881] = \nz.mem_2881_sv2v_reg ;
  assign \nz.mem [2880] = \nz.mem_2880_sv2v_reg ;
  assign \nz.mem [2879] = \nz.mem_2879_sv2v_reg ;
  assign \nz.mem [2878] = \nz.mem_2878_sv2v_reg ;
  assign \nz.mem [2877] = \nz.mem_2877_sv2v_reg ;
  assign \nz.mem [2876] = \nz.mem_2876_sv2v_reg ;
  assign \nz.mem [2875] = \nz.mem_2875_sv2v_reg ;
  assign \nz.mem [2874] = \nz.mem_2874_sv2v_reg ;
  assign \nz.mem [2873] = \nz.mem_2873_sv2v_reg ;
  assign \nz.mem [2872] = \nz.mem_2872_sv2v_reg ;
  assign \nz.mem [2871] = \nz.mem_2871_sv2v_reg ;
  assign \nz.mem [2870] = \nz.mem_2870_sv2v_reg ;
  assign \nz.mem [2869] = \nz.mem_2869_sv2v_reg ;
  assign \nz.mem [2868] = \nz.mem_2868_sv2v_reg ;
  assign \nz.mem [2867] = \nz.mem_2867_sv2v_reg ;
  assign \nz.mem [2866] = \nz.mem_2866_sv2v_reg ;
  assign \nz.mem [2865] = \nz.mem_2865_sv2v_reg ;
  assign \nz.mem [2864] = \nz.mem_2864_sv2v_reg ;
  assign \nz.mem [2863] = \nz.mem_2863_sv2v_reg ;
  assign \nz.mem [2862] = \nz.mem_2862_sv2v_reg ;
  assign \nz.mem [2861] = \nz.mem_2861_sv2v_reg ;
  assign \nz.mem [2860] = \nz.mem_2860_sv2v_reg ;
  assign \nz.mem [2859] = \nz.mem_2859_sv2v_reg ;
  assign \nz.mem [2858] = \nz.mem_2858_sv2v_reg ;
  assign \nz.mem [2857] = \nz.mem_2857_sv2v_reg ;
  assign \nz.mem [2856] = \nz.mem_2856_sv2v_reg ;
  assign \nz.mem [2855] = \nz.mem_2855_sv2v_reg ;
  assign \nz.mem [2854] = \nz.mem_2854_sv2v_reg ;
  assign \nz.mem [2853] = \nz.mem_2853_sv2v_reg ;
  assign \nz.mem [2852] = \nz.mem_2852_sv2v_reg ;
  assign \nz.mem [2851] = \nz.mem_2851_sv2v_reg ;
  assign \nz.mem [2850] = \nz.mem_2850_sv2v_reg ;
  assign \nz.mem [2849] = \nz.mem_2849_sv2v_reg ;
  assign \nz.mem [2848] = \nz.mem_2848_sv2v_reg ;
  assign \nz.mem [2847] = \nz.mem_2847_sv2v_reg ;
  assign \nz.mem [2846] = \nz.mem_2846_sv2v_reg ;
  assign \nz.mem [2845] = \nz.mem_2845_sv2v_reg ;
  assign \nz.mem [2844] = \nz.mem_2844_sv2v_reg ;
  assign \nz.mem [2843] = \nz.mem_2843_sv2v_reg ;
  assign \nz.mem [2842] = \nz.mem_2842_sv2v_reg ;
  assign \nz.mem [2841] = \nz.mem_2841_sv2v_reg ;
  assign \nz.mem [2840] = \nz.mem_2840_sv2v_reg ;
  assign \nz.mem [2839] = \nz.mem_2839_sv2v_reg ;
  assign \nz.mem [2838] = \nz.mem_2838_sv2v_reg ;
  assign \nz.mem [2837] = \nz.mem_2837_sv2v_reg ;
  assign \nz.mem [2836] = \nz.mem_2836_sv2v_reg ;
  assign \nz.mem [2835] = \nz.mem_2835_sv2v_reg ;
  assign \nz.mem [2834] = \nz.mem_2834_sv2v_reg ;
  assign \nz.mem [2833] = \nz.mem_2833_sv2v_reg ;
  assign \nz.mem [2832] = \nz.mem_2832_sv2v_reg ;
  assign \nz.mem [2831] = \nz.mem_2831_sv2v_reg ;
  assign \nz.mem [2830] = \nz.mem_2830_sv2v_reg ;
  assign \nz.mem [2829] = \nz.mem_2829_sv2v_reg ;
  assign \nz.mem [2828] = \nz.mem_2828_sv2v_reg ;
  assign \nz.mem [2827] = \nz.mem_2827_sv2v_reg ;
  assign \nz.mem [2826] = \nz.mem_2826_sv2v_reg ;
  assign \nz.mem [2825] = \nz.mem_2825_sv2v_reg ;
  assign \nz.mem [2824] = \nz.mem_2824_sv2v_reg ;
  assign \nz.mem [2823] = \nz.mem_2823_sv2v_reg ;
  assign \nz.mem [2822] = \nz.mem_2822_sv2v_reg ;
  assign \nz.mem [2821] = \nz.mem_2821_sv2v_reg ;
  assign \nz.mem [2820] = \nz.mem_2820_sv2v_reg ;
  assign \nz.mem [2819] = \nz.mem_2819_sv2v_reg ;
  assign \nz.mem [2818] = \nz.mem_2818_sv2v_reg ;
  assign \nz.mem [2817] = \nz.mem_2817_sv2v_reg ;
  assign \nz.mem [2816] = \nz.mem_2816_sv2v_reg ;
  assign \nz.mem [2815] = \nz.mem_2815_sv2v_reg ;
  assign \nz.mem [2814] = \nz.mem_2814_sv2v_reg ;
  assign \nz.mem [2813] = \nz.mem_2813_sv2v_reg ;
  assign \nz.mem [2812] = \nz.mem_2812_sv2v_reg ;
  assign \nz.mem [2811] = \nz.mem_2811_sv2v_reg ;
  assign \nz.mem [2810] = \nz.mem_2810_sv2v_reg ;
  assign \nz.mem [2809] = \nz.mem_2809_sv2v_reg ;
  assign \nz.mem [2808] = \nz.mem_2808_sv2v_reg ;
  assign \nz.mem [2807] = \nz.mem_2807_sv2v_reg ;
  assign \nz.mem [2806] = \nz.mem_2806_sv2v_reg ;
  assign \nz.mem [2805] = \nz.mem_2805_sv2v_reg ;
  assign \nz.mem [2804] = \nz.mem_2804_sv2v_reg ;
  assign \nz.mem [2803] = \nz.mem_2803_sv2v_reg ;
  assign \nz.mem [2802] = \nz.mem_2802_sv2v_reg ;
  assign \nz.mem [2801] = \nz.mem_2801_sv2v_reg ;
  assign \nz.mem [2800] = \nz.mem_2800_sv2v_reg ;
  assign \nz.mem [2799] = \nz.mem_2799_sv2v_reg ;
  assign \nz.mem [2798] = \nz.mem_2798_sv2v_reg ;
  assign \nz.mem [2797] = \nz.mem_2797_sv2v_reg ;
  assign \nz.mem [2796] = \nz.mem_2796_sv2v_reg ;
  assign \nz.mem [2795] = \nz.mem_2795_sv2v_reg ;
  assign \nz.mem [2794] = \nz.mem_2794_sv2v_reg ;
  assign \nz.mem [2793] = \nz.mem_2793_sv2v_reg ;
  assign \nz.mem [2792] = \nz.mem_2792_sv2v_reg ;
  assign \nz.mem [2791] = \nz.mem_2791_sv2v_reg ;
  assign \nz.mem [2790] = \nz.mem_2790_sv2v_reg ;
  assign \nz.mem [2789] = \nz.mem_2789_sv2v_reg ;
  assign \nz.mem [2788] = \nz.mem_2788_sv2v_reg ;
  assign \nz.mem [2787] = \nz.mem_2787_sv2v_reg ;
  assign \nz.mem [2786] = \nz.mem_2786_sv2v_reg ;
  assign \nz.mem [2785] = \nz.mem_2785_sv2v_reg ;
  assign \nz.mem [2784] = \nz.mem_2784_sv2v_reg ;
  assign \nz.mem [2783] = \nz.mem_2783_sv2v_reg ;
  assign \nz.mem [2782] = \nz.mem_2782_sv2v_reg ;
  assign \nz.mem [2781] = \nz.mem_2781_sv2v_reg ;
  assign \nz.mem [2780] = \nz.mem_2780_sv2v_reg ;
  assign \nz.mem [2779] = \nz.mem_2779_sv2v_reg ;
  assign \nz.mem [2778] = \nz.mem_2778_sv2v_reg ;
  assign \nz.mem [2777] = \nz.mem_2777_sv2v_reg ;
  assign \nz.mem [2776] = \nz.mem_2776_sv2v_reg ;
  assign \nz.mem [2775] = \nz.mem_2775_sv2v_reg ;
  assign \nz.mem [2774] = \nz.mem_2774_sv2v_reg ;
  assign \nz.mem [2773] = \nz.mem_2773_sv2v_reg ;
  assign \nz.mem [2772] = \nz.mem_2772_sv2v_reg ;
  assign \nz.mem [2771] = \nz.mem_2771_sv2v_reg ;
  assign \nz.mem [2770] = \nz.mem_2770_sv2v_reg ;
  assign \nz.mem [2769] = \nz.mem_2769_sv2v_reg ;
  assign \nz.mem [2768] = \nz.mem_2768_sv2v_reg ;
  assign \nz.mem [2767] = \nz.mem_2767_sv2v_reg ;
  assign \nz.mem [2766] = \nz.mem_2766_sv2v_reg ;
  assign \nz.mem [2765] = \nz.mem_2765_sv2v_reg ;
  assign \nz.mem [2764] = \nz.mem_2764_sv2v_reg ;
  assign \nz.mem [2763] = \nz.mem_2763_sv2v_reg ;
  assign \nz.mem [2762] = \nz.mem_2762_sv2v_reg ;
  assign \nz.mem [2761] = \nz.mem_2761_sv2v_reg ;
  assign \nz.mem [2760] = \nz.mem_2760_sv2v_reg ;
  assign \nz.mem [2759] = \nz.mem_2759_sv2v_reg ;
  assign \nz.mem [2758] = \nz.mem_2758_sv2v_reg ;
  assign \nz.mem [2757] = \nz.mem_2757_sv2v_reg ;
  assign \nz.mem [2756] = \nz.mem_2756_sv2v_reg ;
  assign \nz.mem [2755] = \nz.mem_2755_sv2v_reg ;
  assign \nz.mem [2754] = \nz.mem_2754_sv2v_reg ;
  assign \nz.mem [2753] = \nz.mem_2753_sv2v_reg ;
  assign \nz.mem [2752] = \nz.mem_2752_sv2v_reg ;
  assign \nz.mem [2751] = \nz.mem_2751_sv2v_reg ;
  assign \nz.mem [2750] = \nz.mem_2750_sv2v_reg ;
  assign \nz.mem [2749] = \nz.mem_2749_sv2v_reg ;
  assign \nz.mem [2748] = \nz.mem_2748_sv2v_reg ;
  assign \nz.mem [2747] = \nz.mem_2747_sv2v_reg ;
  assign \nz.mem [2746] = \nz.mem_2746_sv2v_reg ;
  assign \nz.mem [2745] = \nz.mem_2745_sv2v_reg ;
  assign \nz.mem [2744] = \nz.mem_2744_sv2v_reg ;
  assign \nz.mem [2743] = \nz.mem_2743_sv2v_reg ;
  assign \nz.mem [2742] = \nz.mem_2742_sv2v_reg ;
  assign \nz.mem [2741] = \nz.mem_2741_sv2v_reg ;
  assign \nz.mem [2740] = \nz.mem_2740_sv2v_reg ;
  assign \nz.mem [2739] = \nz.mem_2739_sv2v_reg ;
  assign \nz.mem [2738] = \nz.mem_2738_sv2v_reg ;
  assign \nz.mem [2737] = \nz.mem_2737_sv2v_reg ;
  assign \nz.mem [2736] = \nz.mem_2736_sv2v_reg ;
  assign \nz.mem [2735] = \nz.mem_2735_sv2v_reg ;
  assign \nz.mem [2734] = \nz.mem_2734_sv2v_reg ;
  assign \nz.mem [2733] = \nz.mem_2733_sv2v_reg ;
  assign \nz.mem [2732] = \nz.mem_2732_sv2v_reg ;
  assign \nz.mem [2731] = \nz.mem_2731_sv2v_reg ;
  assign \nz.mem [2730] = \nz.mem_2730_sv2v_reg ;
  assign \nz.mem [2729] = \nz.mem_2729_sv2v_reg ;
  assign \nz.mem [2728] = \nz.mem_2728_sv2v_reg ;
  assign \nz.mem [2727] = \nz.mem_2727_sv2v_reg ;
  assign \nz.mem [2726] = \nz.mem_2726_sv2v_reg ;
  assign \nz.mem [2725] = \nz.mem_2725_sv2v_reg ;
  assign \nz.mem [2724] = \nz.mem_2724_sv2v_reg ;
  assign \nz.mem [2723] = \nz.mem_2723_sv2v_reg ;
  assign \nz.mem [2722] = \nz.mem_2722_sv2v_reg ;
  assign \nz.mem [2721] = \nz.mem_2721_sv2v_reg ;
  assign \nz.mem [2720] = \nz.mem_2720_sv2v_reg ;
  assign \nz.mem [2719] = \nz.mem_2719_sv2v_reg ;
  assign \nz.mem [2718] = \nz.mem_2718_sv2v_reg ;
  assign \nz.mem [2717] = \nz.mem_2717_sv2v_reg ;
  assign \nz.mem [2716] = \nz.mem_2716_sv2v_reg ;
  assign \nz.mem [2715] = \nz.mem_2715_sv2v_reg ;
  assign \nz.mem [2714] = \nz.mem_2714_sv2v_reg ;
  assign \nz.mem [2713] = \nz.mem_2713_sv2v_reg ;
  assign \nz.mem [2712] = \nz.mem_2712_sv2v_reg ;
  assign \nz.mem [2711] = \nz.mem_2711_sv2v_reg ;
  assign \nz.mem [2710] = \nz.mem_2710_sv2v_reg ;
  assign \nz.mem [2709] = \nz.mem_2709_sv2v_reg ;
  assign \nz.mem [2708] = \nz.mem_2708_sv2v_reg ;
  assign \nz.mem [2707] = \nz.mem_2707_sv2v_reg ;
  assign \nz.mem [2706] = \nz.mem_2706_sv2v_reg ;
  assign \nz.mem [2705] = \nz.mem_2705_sv2v_reg ;
  assign \nz.mem [2704] = \nz.mem_2704_sv2v_reg ;
  assign \nz.mem [2703] = \nz.mem_2703_sv2v_reg ;
  assign \nz.mem [2702] = \nz.mem_2702_sv2v_reg ;
  assign \nz.mem [2701] = \nz.mem_2701_sv2v_reg ;
  assign \nz.mem [2700] = \nz.mem_2700_sv2v_reg ;
  assign \nz.mem [2699] = \nz.mem_2699_sv2v_reg ;
  assign \nz.mem [2698] = \nz.mem_2698_sv2v_reg ;
  assign \nz.mem [2697] = \nz.mem_2697_sv2v_reg ;
  assign \nz.mem [2696] = \nz.mem_2696_sv2v_reg ;
  assign \nz.mem [2695] = \nz.mem_2695_sv2v_reg ;
  assign \nz.mem [2694] = \nz.mem_2694_sv2v_reg ;
  assign \nz.mem [2693] = \nz.mem_2693_sv2v_reg ;
  assign \nz.mem [2692] = \nz.mem_2692_sv2v_reg ;
  assign \nz.mem [2691] = \nz.mem_2691_sv2v_reg ;
  assign \nz.mem [2690] = \nz.mem_2690_sv2v_reg ;
  assign \nz.mem [2689] = \nz.mem_2689_sv2v_reg ;
  assign \nz.mem [2688] = \nz.mem_2688_sv2v_reg ;
  assign \nz.mem [2687] = \nz.mem_2687_sv2v_reg ;
  assign \nz.mem [2686] = \nz.mem_2686_sv2v_reg ;
  assign \nz.mem [2685] = \nz.mem_2685_sv2v_reg ;
  assign \nz.mem [2684] = \nz.mem_2684_sv2v_reg ;
  assign \nz.mem [2683] = \nz.mem_2683_sv2v_reg ;
  assign \nz.mem [2682] = \nz.mem_2682_sv2v_reg ;
  assign \nz.mem [2681] = \nz.mem_2681_sv2v_reg ;
  assign \nz.mem [2680] = \nz.mem_2680_sv2v_reg ;
  assign \nz.mem [2679] = \nz.mem_2679_sv2v_reg ;
  assign \nz.mem [2678] = \nz.mem_2678_sv2v_reg ;
  assign \nz.mem [2677] = \nz.mem_2677_sv2v_reg ;
  assign \nz.mem [2676] = \nz.mem_2676_sv2v_reg ;
  assign \nz.mem [2675] = \nz.mem_2675_sv2v_reg ;
  assign \nz.mem [2674] = \nz.mem_2674_sv2v_reg ;
  assign \nz.mem [2673] = \nz.mem_2673_sv2v_reg ;
  assign \nz.mem [2672] = \nz.mem_2672_sv2v_reg ;
  assign \nz.mem [2671] = \nz.mem_2671_sv2v_reg ;
  assign \nz.mem [2670] = \nz.mem_2670_sv2v_reg ;
  assign \nz.mem [2669] = \nz.mem_2669_sv2v_reg ;
  assign \nz.mem [2668] = \nz.mem_2668_sv2v_reg ;
  assign \nz.mem [2667] = \nz.mem_2667_sv2v_reg ;
  assign \nz.mem [2666] = \nz.mem_2666_sv2v_reg ;
  assign \nz.mem [2665] = \nz.mem_2665_sv2v_reg ;
  assign \nz.mem [2664] = \nz.mem_2664_sv2v_reg ;
  assign \nz.mem [2663] = \nz.mem_2663_sv2v_reg ;
  assign \nz.mem [2662] = \nz.mem_2662_sv2v_reg ;
  assign \nz.mem [2661] = \nz.mem_2661_sv2v_reg ;
  assign \nz.mem [2660] = \nz.mem_2660_sv2v_reg ;
  assign \nz.mem [2659] = \nz.mem_2659_sv2v_reg ;
  assign \nz.mem [2658] = \nz.mem_2658_sv2v_reg ;
  assign \nz.mem [2657] = \nz.mem_2657_sv2v_reg ;
  assign \nz.mem [2656] = \nz.mem_2656_sv2v_reg ;
  assign \nz.mem [2655] = \nz.mem_2655_sv2v_reg ;
  assign \nz.mem [2654] = \nz.mem_2654_sv2v_reg ;
  assign \nz.mem [2653] = \nz.mem_2653_sv2v_reg ;
  assign \nz.mem [2652] = \nz.mem_2652_sv2v_reg ;
  assign \nz.mem [2651] = \nz.mem_2651_sv2v_reg ;
  assign \nz.mem [2650] = \nz.mem_2650_sv2v_reg ;
  assign \nz.mem [2649] = \nz.mem_2649_sv2v_reg ;
  assign \nz.mem [2648] = \nz.mem_2648_sv2v_reg ;
  assign \nz.mem [2647] = \nz.mem_2647_sv2v_reg ;
  assign \nz.mem [2646] = \nz.mem_2646_sv2v_reg ;
  assign \nz.mem [2645] = \nz.mem_2645_sv2v_reg ;
  assign \nz.mem [2644] = \nz.mem_2644_sv2v_reg ;
  assign \nz.mem [2643] = \nz.mem_2643_sv2v_reg ;
  assign \nz.mem [2642] = \nz.mem_2642_sv2v_reg ;
  assign \nz.mem [2641] = \nz.mem_2641_sv2v_reg ;
  assign \nz.mem [2640] = \nz.mem_2640_sv2v_reg ;
  assign \nz.mem [2639] = \nz.mem_2639_sv2v_reg ;
  assign \nz.mem [2638] = \nz.mem_2638_sv2v_reg ;
  assign \nz.mem [2637] = \nz.mem_2637_sv2v_reg ;
  assign \nz.mem [2636] = \nz.mem_2636_sv2v_reg ;
  assign \nz.mem [2635] = \nz.mem_2635_sv2v_reg ;
  assign \nz.mem [2634] = \nz.mem_2634_sv2v_reg ;
  assign \nz.mem [2633] = \nz.mem_2633_sv2v_reg ;
  assign \nz.mem [2632] = \nz.mem_2632_sv2v_reg ;
  assign \nz.mem [2631] = \nz.mem_2631_sv2v_reg ;
  assign \nz.mem [2630] = \nz.mem_2630_sv2v_reg ;
  assign \nz.mem [2629] = \nz.mem_2629_sv2v_reg ;
  assign \nz.mem [2628] = \nz.mem_2628_sv2v_reg ;
  assign \nz.mem [2627] = \nz.mem_2627_sv2v_reg ;
  assign \nz.mem [2626] = \nz.mem_2626_sv2v_reg ;
  assign \nz.mem [2625] = \nz.mem_2625_sv2v_reg ;
  assign \nz.mem [2624] = \nz.mem_2624_sv2v_reg ;
  assign \nz.mem [2623] = \nz.mem_2623_sv2v_reg ;
  assign \nz.mem [2622] = \nz.mem_2622_sv2v_reg ;
  assign \nz.mem [2621] = \nz.mem_2621_sv2v_reg ;
  assign \nz.mem [2620] = \nz.mem_2620_sv2v_reg ;
  assign \nz.mem [2619] = \nz.mem_2619_sv2v_reg ;
  assign \nz.mem [2618] = \nz.mem_2618_sv2v_reg ;
  assign \nz.mem [2617] = \nz.mem_2617_sv2v_reg ;
  assign \nz.mem [2616] = \nz.mem_2616_sv2v_reg ;
  assign \nz.mem [2615] = \nz.mem_2615_sv2v_reg ;
  assign \nz.mem [2614] = \nz.mem_2614_sv2v_reg ;
  assign \nz.mem [2613] = \nz.mem_2613_sv2v_reg ;
  assign \nz.mem [2612] = \nz.mem_2612_sv2v_reg ;
  assign \nz.mem [2611] = \nz.mem_2611_sv2v_reg ;
  assign \nz.mem [2610] = \nz.mem_2610_sv2v_reg ;
  assign \nz.mem [2609] = \nz.mem_2609_sv2v_reg ;
  assign \nz.mem [2608] = \nz.mem_2608_sv2v_reg ;
  assign \nz.mem [2607] = \nz.mem_2607_sv2v_reg ;
  assign \nz.mem [2606] = \nz.mem_2606_sv2v_reg ;
  assign \nz.mem [2605] = \nz.mem_2605_sv2v_reg ;
  assign \nz.mem [2604] = \nz.mem_2604_sv2v_reg ;
  assign \nz.mem [2603] = \nz.mem_2603_sv2v_reg ;
  assign \nz.mem [2602] = \nz.mem_2602_sv2v_reg ;
  assign \nz.mem [2601] = \nz.mem_2601_sv2v_reg ;
  assign \nz.mem [2600] = \nz.mem_2600_sv2v_reg ;
  assign \nz.mem [2599] = \nz.mem_2599_sv2v_reg ;
  assign \nz.mem [2598] = \nz.mem_2598_sv2v_reg ;
  assign \nz.mem [2597] = \nz.mem_2597_sv2v_reg ;
  assign \nz.mem [2596] = \nz.mem_2596_sv2v_reg ;
  assign \nz.mem [2595] = \nz.mem_2595_sv2v_reg ;
  assign \nz.mem [2594] = \nz.mem_2594_sv2v_reg ;
  assign \nz.mem [2593] = \nz.mem_2593_sv2v_reg ;
  assign \nz.mem [2592] = \nz.mem_2592_sv2v_reg ;
  assign \nz.mem [2591] = \nz.mem_2591_sv2v_reg ;
  assign \nz.mem [2590] = \nz.mem_2590_sv2v_reg ;
  assign \nz.mem [2589] = \nz.mem_2589_sv2v_reg ;
  assign \nz.mem [2588] = \nz.mem_2588_sv2v_reg ;
  assign \nz.mem [2587] = \nz.mem_2587_sv2v_reg ;
  assign \nz.mem [2586] = \nz.mem_2586_sv2v_reg ;
  assign \nz.mem [2585] = \nz.mem_2585_sv2v_reg ;
  assign \nz.mem [2584] = \nz.mem_2584_sv2v_reg ;
  assign \nz.mem [2583] = \nz.mem_2583_sv2v_reg ;
  assign \nz.mem [2582] = \nz.mem_2582_sv2v_reg ;
  assign \nz.mem [2581] = \nz.mem_2581_sv2v_reg ;
  assign \nz.mem [2580] = \nz.mem_2580_sv2v_reg ;
  assign \nz.mem [2579] = \nz.mem_2579_sv2v_reg ;
  assign \nz.mem [2578] = \nz.mem_2578_sv2v_reg ;
  assign \nz.mem [2577] = \nz.mem_2577_sv2v_reg ;
  assign \nz.mem [2576] = \nz.mem_2576_sv2v_reg ;
  assign \nz.mem [2575] = \nz.mem_2575_sv2v_reg ;
  assign \nz.mem [2574] = \nz.mem_2574_sv2v_reg ;
  assign \nz.mem [2573] = \nz.mem_2573_sv2v_reg ;
  assign \nz.mem [2572] = \nz.mem_2572_sv2v_reg ;
  assign \nz.mem [2571] = \nz.mem_2571_sv2v_reg ;
  assign \nz.mem [2570] = \nz.mem_2570_sv2v_reg ;
  assign \nz.mem [2569] = \nz.mem_2569_sv2v_reg ;
  assign \nz.mem [2568] = \nz.mem_2568_sv2v_reg ;
  assign \nz.mem [2567] = \nz.mem_2567_sv2v_reg ;
  assign \nz.mem [2566] = \nz.mem_2566_sv2v_reg ;
  assign \nz.mem [2565] = \nz.mem_2565_sv2v_reg ;
  assign \nz.mem [2564] = \nz.mem_2564_sv2v_reg ;
  assign \nz.mem [2563] = \nz.mem_2563_sv2v_reg ;
  assign \nz.mem [2562] = \nz.mem_2562_sv2v_reg ;
  assign \nz.mem [2561] = \nz.mem_2561_sv2v_reg ;
  assign \nz.mem [2560] = \nz.mem_2560_sv2v_reg ;
  assign \nz.mem [2559] = \nz.mem_2559_sv2v_reg ;
  assign \nz.mem [2558] = \nz.mem_2558_sv2v_reg ;
  assign \nz.mem [2557] = \nz.mem_2557_sv2v_reg ;
  assign \nz.mem [2556] = \nz.mem_2556_sv2v_reg ;
  assign \nz.mem [2555] = \nz.mem_2555_sv2v_reg ;
  assign \nz.mem [2554] = \nz.mem_2554_sv2v_reg ;
  assign \nz.mem [2553] = \nz.mem_2553_sv2v_reg ;
  assign \nz.mem [2552] = \nz.mem_2552_sv2v_reg ;
  assign \nz.mem [2551] = \nz.mem_2551_sv2v_reg ;
  assign \nz.mem [2550] = \nz.mem_2550_sv2v_reg ;
  assign \nz.mem [2549] = \nz.mem_2549_sv2v_reg ;
  assign \nz.mem [2548] = \nz.mem_2548_sv2v_reg ;
  assign \nz.mem [2547] = \nz.mem_2547_sv2v_reg ;
  assign \nz.mem [2546] = \nz.mem_2546_sv2v_reg ;
  assign \nz.mem [2545] = \nz.mem_2545_sv2v_reg ;
  assign \nz.mem [2544] = \nz.mem_2544_sv2v_reg ;
  assign \nz.mem [2543] = \nz.mem_2543_sv2v_reg ;
  assign \nz.mem [2542] = \nz.mem_2542_sv2v_reg ;
  assign \nz.mem [2541] = \nz.mem_2541_sv2v_reg ;
  assign \nz.mem [2540] = \nz.mem_2540_sv2v_reg ;
  assign \nz.mem [2539] = \nz.mem_2539_sv2v_reg ;
  assign \nz.mem [2538] = \nz.mem_2538_sv2v_reg ;
  assign \nz.mem [2537] = \nz.mem_2537_sv2v_reg ;
  assign \nz.mem [2536] = \nz.mem_2536_sv2v_reg ;
  assign \nz.mem [2535] = \nz.mem_2535_sv2v_reg ;
  assign \nz.mem [2534] = \nz.mem_2534_sv2v_reg ;
  assign \nz.mem [2533] = \nz.mem_2533_sv2v_reg ;
  assign \nz.mem [2532] = \nz.mem_2532_sv2v_reg ;
  assign \nz.mem [2531] = \nz.mem_2531_sv2v_reg ;
  assign \nz.mem [2530] = \nz.mem_2530_sv2v_reg ;
  assign \nz.mem [2529] = \nz.mem_2529_sv2v_reg ;
  assign \nz.mem [2528] = \nz.mem_2528_sv2v_reg ;
  assign \nz.mem [2527] = \nz.mem_2527_sv2v_reg ;
  assign \nz.mem [2526] = \nz.mem_2526_sv2v_reg ;
  assign \nz.mem [2525] = \nz.mem_2525_sv2v_reg ;
  assign \nz.mem [2524] = \nz.mem_2524_sv2v_reg ;
  assign \nz.mem [2523] = \nz.mem_2523_sv2v_reg ;
  assign \nz.mem [2522] = \nz.mem_2522_sv2v_reg ;
  assign \nz.mem [2521] = \nz.mem_2521_sv2v_reg ;
  assign \nz.mem [2520] = \nz.mem_2520_sv2v_reg ;
  assign \nz.mem [2519] = \nz.mem_2519_sv2v_reg ;
  assign \nz.mem [2518] = \nz.mem_2518_sv2v_reg ;
  assign \nz.mem [2517] = \nz.mem_2517_sv2v_reg ;
  assign \nz.mem [2516] = \nz.mem_2516_sv2v_reg ;
  assign \nz.mem [2515] = \nz.mem_2515_sv2v_reg ;
  assign \nz.mem [2514] = \nz.mem_2514_sv2v_reg ;
  assign \nz.mem [2513] = \nz.mem_2513_sv2v_reg ;
  assign \nz.mem [2512] = \nz.mem_2512_sv2v_reg ;
  assign \nz.mem [2511] = \nz.mem_2511_sv2v_reg ;
  assign \nz.mem [2510] = \nz.mem_2510_sv2v_reg ;
  assign \nz.mem [2509] = \nz.mem_2509_sv2v_reg ;
  assign \nz.mem [2508] = \nz.mem_2508_sv2v_reg ;
  assign \nz.mem [2507] = \nz.mem_2507_sv2v_reg ;
  assign \nz.mem [2506] = \nz.mem_2506_sv2v_reg ;
  assign \nz.mem [2505] = \nz.mem_2505_sv2v_reg ;
  assign \nz.mem [2504] = \nz.mem_2504_sv2v_reg ;
  assign \nz.mem [2503] = \nz.mem_2503_sv2v_reg ;
  assign \nz.mem [2502] = \nz.mem_2502_sv2v_reg ;
  assign \nz.mem [2501] = \nz.mem_2501_sv2v_reg ;
  assign \nz.mem [2500] = \nz.mem_2500_sv2v_reg ;
  assign \nz.mem [2499] = \nz.mem_2499_sv2v_reg ;
  assign \nz.mem [2498] = \nz.mem_2498_sv2v_reg ;
  assign \nz.mem [2497] = \nz.mem_2497_sv2v_reg ;
  assign \nz.mem [2496] = \nz.mem_2496_sv2v_reg ;
  assign \nz.mem [2495] = \nz.mem_2495_sv2v_reg ;
  assign \nz.mem [2494] = \nz.mem_2494_sv2v_reg ;
  assign \nz.mem [2493] = \nz.mem_2493_sv2v_reg ;
  assign \nz.mem [2492] = \nz.mem_2492_sv2v_reg ;
  assign \nz.mem [2491] = \nz.mem_2491_sv2v_reg ;
  assign \nz.mem [2490] = \nz.mem_2490_sv2v_reg ;
  assign \nz.mem [2489] = \nz.mem_2489_sv2v_reg ;
  assign \nz.mem [2488] = \nz.mem_2488_sv2v_reg ;
  assign \nz.mem [2487] = \nz.mem_2487_sv2v_reg ;
  assign \nz.mem [2486] = \nz.mem_2486_sv2v_reg ;
  assign \nz.mem [2485] = \nz.mem_2485_sv2v_reg ;
  assign \nz.mem [2484] = \nz.mem_2484_sv2v_reg ;
  assign \nz.mem [2483] = \nz.mem_2483_sv2v_reg ;
  assign \nz.mem [2482] = \nz.mem_2482_sv2v_reg ;
  assign \nz.mem [2481] = \nz.mem_2481_sv2v_reg ;
  assign \nz.mem [2480] = \nz.mem_2480_sv2v_reg ;
  assign \nz.mem [2479] = \nz.mem_2479_sv2v_reg ;
  assign \nz.mem [2478] = \nz.mem_2478_sv2v_reg ;
  assign \nz.mem [2477] = \nz.mem_2477_sv2v_reg ;
  assign \nz.mem [2476] = \nz.mem_2476_sv2v_reg ;
  assign \nz.mem [2475] = \nz.mem_2475_sv2v_reg ;
  assign \nz.mem [2474] = \nz.mem_2474_sv2v_reg ;
  assign \nz.mem [2473] = \nz.mem_2473_sv2v_reg ;
  assign \nz.mem [2472] = \nz.mem_2472_sv2v_reg ;
  assign \nz.mem [2471] = \nz.mem_2471_sv2v_reg ;
  assign \nz.mem [2470] = \nz.mem_2470_sv2v_reg ;
  assign \nz.mem [2469] = \nz.mem_2469_sv2v_reg ;
  assign \nz.mem [2468] = \nz.mem_2468_sv2v_reg ;
  assign \nz.mem [2467] = \nz.mem_2467_sv2v_reg ;
  assign \nz.mem [2466] = \nz.mem_2466_sv2v_reg ;
  assign \nz.mem [2465] = \nz.mem_2465_sv2v_reg ;
  assign \nz.mem [2464] = \nz.mem_2464_sv2v_reg ;
  assign \nz.mem [2463] = \nz.mem_2463_sv2v_reg ;
  assign \nz.mem [2462] = \nz.mem_2462_sv2v_reg ;
  assign \nz.mem [2461] = \nz.mem_2461_sv2v_reg ;
  assign \nz.mem [2460] = \nz.mem_2460_sv2v_reg ;
  assign \nz.mem [2459] = \nz.mem_2459_sv2v_reg ;
  assign \nz.mem [2458] = \nz.mem_2458_sv2v_reg ;
  assign \nz.mem [2457] = \nz.mem_2457_sv2v_reg ;
  assign \nz.mem [2456] = \nz.mem_2456_sv2v_reg ;
  assign \nz.mem [2455] = \nz.mem_2455_sv2v_reg ;
  assign \nz.mem [2454] = \nz.mem_2454_sv2v_reg ;
  assign \nz.mem [2453] = \nz.mem_2453_sv2v_reg ;
  assign \nz.mem [2452] = \nz.mem_2452_sv2v_reg ;
  assign \nz.mem [2451] = \nz.mem_2451_sv2v_reg ;
  assign \nz.mem [2450] = \nz.mem_2450_sv2v_reg ;
  assign \nz.mem [2449] = \nz.mem_2449_sv2v_reg ;
  assign \nz.mem [2448] = \nz.mem_2448_sv2v_reg ;
  assign \nz.mem [2447] = \nz.mem_2447_sv2v_reg ;
  assign \nz.mem [2446] = \nz.mem_2446_sv2v_reg ;
  assign \nz.mem [2445] = \nz.mem_2445_sv2v_reg ;
  assign \nz.mem [2444] = \nz.mem_2444_sv2v_reg ;
  assign \nz.mem [2443] = \nz.mem_2443_sv2v_reg ;
  assign \nz.mem [2442] = \nz.mem_2442_sv2v_reg ;
  assign \nz.mem [2441] = \nz.mem_2441_sv2v_reg ;
  assign \nz.mem [2440] = \nz.mem_2440_sv2v_reg ;
  assign \nz.mem [2439] = \nz.mem_2439_sv2v_reg ;
  assign \nz.mem [2438] = \nz.mem_2438_sv2v_reg ;
  assign \nz.mem [2437] = \nz.mem_2437_sv2v_reg ;
  assign \nz.mem [2436] = \nz.mem_2436_sv2v_reg ;
  assign \nz.mem [2435] = \nz.mem_2435_sv2v_reg ;
  assign \nz.mem [2434] = \nz.mem_2434_sv2v_reg ;
  assign \nz.mem [2433] = \nz.mem_2433_sv2v_reg ;
  assign \nz.mem [2432] = \nz.mem_2432_sv2v_reg ;
  assign \nz.mem [2431] = \nz.mem_2431_sv2v_reg ;
  assign \nz.mem [2430] = \nz.mem_2430_sv2v_reg ;
  assign \nz.mem [2429] = \nz.mem_2429_sv2v_reg ;
  assign \nz.mem [2428] = \nz.mem_2428_sv2v_reg ;
  assign \nz.mem [2427] = \nz.mem_2427_sv2v_reg ;
  assign \nz.mem [2426] = \nz.mem_2426_sv2v_reg ;
  assign \nz.mem [2425] = \nz.mem_2425_sv2v_reg ;
  assign \nz.mem [2424] = \nz.mem_2424_sv2v_reg ;
  assign \nz.mem [2423] = \nz.mem_2423_sv2v_reg ;
  assign \nz.mem [2422] = \nz.mem_2422_sv2v_reg ;
  assign \nz.mem [2421] = \nz.mem_2421_sv2v_reg ;
  assign \nz.mem [2420] = \nz.mem_2420_sv2v_reg ;
  assign \nz.mem [2419] = \nz.mem_2419_sv2v_reg ;
  assign \nz.mem [2418] = \nz.mem_2418_sv2v_reg ;
  assign \nz.mem [2417] = \nz.mem_2417_sv2v_reg ;
  assign \nz.mem [2416] = \nz.mem_2416_sv2v_reg ;
  assign \nz.mem [2415] = \nz.mem_2415_sv2v_reg ;
  assign \nz.mem [2414] = \nz.mem_2414_sv2v_reg ;
  assign \nz.mem [2413] = \nz.mem_2413_sv2v_reg ;
  assign \nz.mem [2412] = \nz.mem_2412_sv2v_reg ;
  assign \nz.mem [2411] = \nz.mem_2411_sv2v_reg ;
  assign \nz.mem [2410] = \nz.mem_2410_sv2v_reg ;
  assign \nz.mem [2409] = \nz.mem_2409_sv2v_reg ;
  assign \nz.mem [2408] = \nz.mem_2408_sv2v_reg ;
  assign \nz.mem [2407] = \nz.mem_2407_sv2v_reg ;
  assign \nz.mem [2406] = \nz.mem_2406_sv2v_reg ;
  assign \nz.mem [2405] = \nz.mem_2405_sv2v_reg ;
  assign \nz.mem [2404] = \nz.mem_2404_sv2v_reg ;
  assign \nz.mem [2403] = \nz.mem_2403_sv2v_reg ;
  assign \nz.mem [2402] = \nz.mem_2402_sv2v_reg ;
  assign \nz.mem [2401] = \nz.mem_2401_sv2v_reg ;
  assign \nz.mem [2400] = \nz.mem_2400_sv2v_reg ;
  assign \nz.mem [2399] = \nz.mem_2399_sv2v_reg ;
  assign \nz.mem [2398] = \nz.mem_2398_sv2v_reg ;
  assign \nz.mem [2397] = \nz.mem_2397_sv2v_reg ;
  assign \nz.mem [2396] = \nz.mem_2396_sv2v_reg ;
  assign \nz.mem [2395] = \nz.mem_2395_sv2v_reg ;
  assign \nz.mem [2394] = \nz.mem_2394_sv2v_reg ;
  assign \nz.mem [2393] = \nz.mem_2393_sv2v_reg ;
  assign \nz.mem [2392] = \nz.mem_2392_sv2v_reg ;
  assign \nz.mem [2391] = \nz.mem_2391_sv2v_reg ;
  assign \nz.mem [2390] = \nz.mem_2390_sv2v_reg ;
  assign \nz.mem [2389] = \nz.mem_2389_sv2v_reg ;
  assign \nz.mem [2388] = \nz.mem_2388_sv2v_reg ;
  assign \nz.mem [2387] = \nz.mem_2387_sv2v_reg ;
  assign \nz.mem [2386] = \nz.mem_2386_sv2v_reg ;
  assign \nz.mem [2385] = \nz.mem_2385_sv2v_reg ;
  assign \nz.mem [2384] = \nz.mem_2384_sv2v_reg ;
  assign \nz.mem [2383] = \nz.mem_2383_sv2v_reg ;
  assign \nz.mem [2382] = \nz.mem_2382_sv2v_reg ;
  assign \nz.mem [2381] = \nz.mem_2381_sv2v_reg ;
  assign \nz.mem [2380] = \nz.mem_2380_sv2v_reg ;
  assign \nz.mem [2379] = \nz.mem_2379_sv2v_reg ;
  assign \nz.mem [2378] = \nz.mem_2378_sv2v_reg ;
  assign \nz.mem [2377] = \nz.mem_2377_sv2v_reg ;
  assign \nz.mem [2376] = \nz.mem_2376_sv2v_reg ;
  assign \nz.mem [2375] = \nz.mem_2375_sv2v_reg ;
  assign \nz.mem [2374] = \nz.mem_2374_sv2v_reg ;
  assign \nz.mem [2373] = \nz.mem_2373_sv2v_reg ;
  assign \nz.mem [2372] = \nz.mem_2372_sv2v_reg ;
  assign \nz.mem [2371] = \nz.mem_2371_sv2v_reg ;
  assign \nz.mem [2370] = \nz.mem_2370_sv2v_reg ;
  assign \nz.mem [2369] = \nz.mem_2369_sv2v_reg ;
  assign \nz.mem [2368] = \nz.mem_2368_sv2v_reg ;
  assign \nz.mem [2367] = \nz.mem_2367_sv2v_reg ;
  assign \nz.mem [2366] = \nz.mem_2366_sv2v_reg ;
  assign \nz.mem [2365] = \nz.mem_2365_sv2v_reg ;
  assign \nz.mem [2364] = \nz.mem_2364_sv2v_reg ;
  assign \nz.mem [2363] = \nz.mem_2363_sv2v_reg ;
  assign \nz.mem [2362] = \nz.mem_2362_sv2v_reg ;
  assign \nz.mem [2361] = \nz.mem_2361_sv2v_reg ;
  assign \nz.mem [2360] = \nz.mem_2360_sv2v_reg ;
  assign \nz.mem [2359] = \nz.mem_2359_sv2v_reg ;
  assign \nz.mem [2358] = \nz.mem_2358_sv2v_reg ;
  assign \nz.mem [2357] = \nz.mem_2357_sv2v_reg ;
  assign \nz.mem [2356] = \nz.mem_2356_sv2v_reg ;
  assign \nz.mem [2355] = \nz.mem_2355_sv2v_reg ;
  assign \nz.mem [2354] = \nz.mem_2354_sv2v_reg ;
  assign \nz.mem [2353] = \nz.mem_2353_sv2v_reg ;
  assign \nz.mem [2352] = \nz.mem_2352_sv2v_reg ;
  assign \nz.mem [2351] = \nz.mem_2351_sv2v_reg ;
  assign \nz.mem [2350] = \nz.mem_2350_sv2v_reg ;
  assign \nz.mem [2349] = \nz.mem_2349_sv2v_reg ;
  assign \nz.mem [2348] = \nz.mem_2348_sv2v_reg ;
  assign \nz.mem [2347] = \nz.mem_2347_sv2v_reg ;
  assign \nz.mem [2346] = \nz.mem_2346_sv2v_reg ;
  assign \nz.mem [2345] = \nz.mem_2345_sv2v_reg ;
  assign \nz.mem [2344] = \nz.mem_2344_sv2v_reg ;
  assign \nz.mem [2343] = \nz.mem_2343_sv2v_reg ;
  assign \nz.mem [2342] = \nz.mem_2342_sv2v_reg ;
  assign \nz.mem [2341] = \nz.mem_2341_sv2v_reg ;
  assign \nz.mem [2340] = \nz.mem_2340_sv2v_reg ;
  assign \nz.mem [2339] = \nz.mem_2339_sv2v_reg ;
  assign \nz.mem [2338] = \nz.mem_2338_sv2v_reg ;
  assign \nz.mem [2337] = \nz.mem_2337_sv2v_reg ;
  assign \nz.mem [2336] = \nz.mem_2336_sv2v_reg ;
  assign \nz.mem [2335] = \nz.mem_2335_sv2v_reg ;
  assign \nz.mem [2334] = \nz.mem_2334_sv2v_reg ;
  assign \nz.mem [2333] = \nz.mem_2333_sv2v_reg ;
  assign \nz.mem [2332] = \nz.mem_2332_sv2v_reg ;
  assign \nz.mem [2331] = \nz.mem_2331_sv2v_reg ;
  assign \nz.mem [2330] = \nz.mem_2330_sv2v_reg ;
  assign \nz.mem [2329] = \nz.mem_2329_sv2v_reg ;
  assign \nz.mem [2328] = \nz.mem_2328_sv2v_reg ;
  assign \nz.mem [2327] = \nz.mem_2327_sv2v_reg ;
  assign \nz.mem [2326] = \nz.mem_2326_sv2v_reg ;
  assign \nz.mem [2325] = \nz.mem_2325_sv2v_reg ;
  assign \nz.mem [2324] = \nz.mem_2324_sv2v_reg ;
  assign \nz.mem [2323] = \nz.mem_2323_sv2v_reg ;
  assign \nz.mem [2322] = \nz.mem_2322_sv2v_reg ;
  assign \nz.mem [2321] = \nz.mem_2321_sv2v_reg ;
  assign \nz.mem [2320] = \nz.mem_2320_sv2v_reg ;
  assign \nz.mem [2319] = \nz.mem_2319_sv2v_reg ;
  assign \nz.mem [2318] = \nz.mem_2318_sv2v_reg ;
  assign \nz.mem [2317] = \nz.mem_2317_sv2v_reg ;
  assign \nz.mem [2316] = \nz.mem_2316_sv2v_reg ;
  assign \nz.mem [2315] = \nz.mem_2315_sv2v_reg ;
  assign \nz.mem [2314] = \nz.mem_2314_sv2v_reg ;
  assign \nz.mem [2313] = \nz.mem_2313_sv2v_reg ;
  assign \nz.mem [2312] = \nz.mem_2312_sv2v_reg ;
  assign \nz.mem [2311] = \nz.mem_2311_sv2v_reg ;
  assign \nz.mem [2310] = \nz.mem_2310_sv2v_reg ;
  assign \nz.mem [2309] = \nz.mem_2309_sv2v_reg ;
  assign \nz.mem [2308] = \nz.mem_2308_sv2v_reg ;
  assign \nz.mem [2307] = \nz.mem_2307_sv2v_reg ;
  assign \nz.mem [2306] = \nz.mem_2306_sv2v_reg ;
  assign \nz.mem [2305] = \nz.mem_2305_sv2v_reg ;
  assign \nz.mem [2304] = \nz.mem_2304_sv2v_reg ;
  assign \nz.mem [2303] = \nz.mem_2303_sv2v_reg ;
  assign \nz.mem [2302] = \nz.mem_2302_sv2v_reg ;
  assign \nz.mem [2301] = \nz.mem_2301_sv2v_reg ;
  assign \nz.mem [2300] = \nz.mem_2300_sv2v_reg ;
  assign \nz.mem [2299] = \nz.mem_2299_sv2v_reg ;
  assign \nz.mem [2298] = \nz.mem_2298_sv2v_reg ;
  assign \nz.mem [2297] = \nz.mem_2297_sv2v_reg ;
  assign \nz.mem [2296] = \nz.mem_2296_sv2v_reg ;
  assign \nz.mem [2295] = \nz.mem_2295_sv2v_reg ;
  assign \nz.mem [2294] = \nz.mem_2294_sv2v_reg ;
  assign \nz.mem [2293] = \nz.mem_2293_sv2v_reg ;
  assign \nz.mem [2292] = \nz.mem_2292_sv2v_reg ;
  assign \nz.mem [2291] = \nz.mem_2291_sv2v_reg ;
  assign \nz.mem [2290] = \nz.mem_2290_sv2v_reg ;
  assign \nz.mem [2289] = \nz.mem_2289_sv2v_reg ;
  assign \nz.mem [2288] = \nz.mem_2288_sv2v_reg ;
  assign \nz.mem [2287] = \nz.mem_2287_sv2v_reg ;
  assign \nz.mem [2286] = \nz.mem_2286_sv2v_reg ;
  assign \nz.mem [2285] = \nz.mem_2285_sv2v_reg ;
  assign \nz.mem [2284] = \nz.mem_2284_sv2v_reg ;
  assign \nz.mem [2283] = \nz.mem_2283_sv2v_reg ;
  assign \nz.mem [2282] = \nz.mem_2282_sv2v_reg ;
  assign \nz.mem [2281] = \nz.mem_2281_sv2v_reg ;
  assign \nz.mem [2280] = \nz.mem_2280_sv2v_reg ;
  assign \nz.mem [2279] = \nz.mem_2279_sv2v_reg ;
  assign \nz.mem [2278] = \nz.mem_2278_sv2v_reg ;
  assign \nz.mem [2277] = \nz.mem_2277_sv2v_reg ;
  assign \nz.mem [2276] = \nz.mem_2276_sv2v_reg ;
  assign \nz.mem [2275] = \nz.mem_2275_sv2v_reg ;
  assign \nz.mem [2274] = \nz.mem_2274_sv2v_reg ;
  assign \nz.mem [2273] = \nz.mem_2273_sv2v_reg ;
  assign \nz.mem [2272] = \nz.mem_2272_sv2v_reg ;
  assign \nz.mem [2271] = \nz.mem_2271_sv2v_reg ;
  assign \nz.mem [2270] = \nz.mem_2270_sv2v_reg ;
  assign \nz.mem [2269] = \nz.mem_2269_sv2v_reg ;
  assign \nz.mem [2268] = \nz.mem_2268_sv2v_reg ;
  assign \nz.mem [2267] = \nz.mem_2267_sv2v_reg ;
  assign \nz.mem [2266] = \nz.mem_2266_sv2v_reg ;
  assign \nz.mem [2265] = \nz.mem_2265_sv2v_reg ;
  assign \nz.mem [2264] = \nz.mem_2264_sv2v_reg ;
  assign \nz.mem [2263] = \nz.mem_2263_sv2v_reg ;
  assign \nz.mem [2262] = \nz.mem_2262_sv2v_reg ;
  assign \nz.mem [2261] = \nz.mem_2261_sv2v_reg ;
  assign \nz.mem [2260] = \nz.mem_2260_sv2v_reg ;
  assign \nz.mem [2259] = \nz.mem_2259_sv2v_reg ;
  assign \nz.mem [2258] = \nz.mem_2258_sv2v_reg ;
  assign \nz.mem [2257] = \nz.mem_2257_sv2v_reg ;
  assign \nz.mem [2256] = \nz.mem_2256_sv2v_reg ;
  assign \nz.mem [2255] = \nz.mem_2255_sv2v_reg ;
  assign \nz.mem [2254] = \nz.mem_2254_sv2v_reg ;
  assign \nz.mem [2253] = \nz.mem_2253_sv2v_reg ;
  assign \nz.mem [2252] = \nz.mem_2252_sv2v_reg ;
  assign \nz.mem [2251] = \nz.mem_2251_sv2v_reg ;
  assign \nz.mem [2250] = \nz.mem_2250_sv2v_reg ;
  assign \nz.mem [2249] = \nz.mem_2249_sv2v_reg ;
  assign \nz.mem [2248] = \nz.mem_2248_sv2v_reg ;
  assign \nz.mem [2247] = \nz.mem_2247_sv2v_reg ;
  assign \nz.mem [2246] = \nz.mem_2246_sv2v_reg ;
  assign \nz.mem [2245] = \nz.mem_2245_sv2v_reg ;
  assign \nz.mem [2244] = \nz.mem_2244_sv2v_reg ;
  assign \nz.mem [2243] = \nz.mem_2243_sv2v_reg ;
  assign \nz.mem [2242] = \nz.mem_2242_sv2v_reg ;
  assign \nz.mem [2241] = \nz.mem_2241_sv2v_reg ;
  assign \nz.mem [2240] = \nz.mem_2240_sv2v_reg ;
  assign \nz.mem [2239] = \nz.mem_2239_sv2v_reg ;
  assign \nz.mem [2238] = \nz.mem_2238_sv2v_reg ;
  assign \nz.mem [2237] = \nz.mem_2237_sv2v_reg ;
  assign \nz.mem [2236] = \nz.mem_2236_sv2v_reg ;
  assign \nz.mem [2235] = \nz.mem_2235_sv2v_reg ;
  assign \nz.mem [2234] = \nz.mem_2234_sv2v_reg ;
  assign \nz.mem [2233] = \nz.mem_2233_sv2v_reg ;
  assign \nz.mem [2232] = \nz.mem_2232_sv2v_reg ;
  assign \nz.mem [2231] = \nz.mem_2231_sv2v_reg ;
  assign \nz.mem [2230] = \nz.mem_2230_sv2v_reg ;
  assign \nz.mem [2229] = \nz.mem_2229_sv2v_reg ;
  assign \nz.mem [2228] = \nz.mem_2228_sv2v_reg ;
  assign \nz.mem [2227] = \nz.mem_2227_sv2v_reg ;
  assign \nz.mem [2226] = \nz.mem_2226_sv2v_reg ;
  assign \nz.mem [2225] = \nz.mem_2225_sv2v_reg ;
  assign \nz.mem [2224] = \nz.mem_2224_sv2v_reg ;
  assign \nz.mem [2223] = \nz.mem_2223_sv2v_reg ;
  assign \nz.mem [2222] = \nz.mem_2222_sv2v_reg ;
  assign \nz.mem [2221] = \nz.mem_2221_sv2v_reg ;
  assign \nz.mem [2220] = \nz.mem_2220_sv2v_reg ;
  assign \nz.mem [2219] = \nz.mem_2219_sv2v_reg ;
  assign \nz.mem [2218] = \nz.mem_2218_sv2v_reg ;
  assign \nz.mem [2217] = \nz.mem_2217_sv2v_reg ;
  assign \nz.mem [2216] = \nz.mem_2216_sv2v_reg ;
  assign \nz.mem [2215] = \nz.mem_2215_sv2v_reg ;
  assign \nz.mem [2214] = \nz.mem_2214_sv2v_reg ;
  assign \nz.mem [2213] = \nz.mem_2213_sv2v_reg ;
  assign \nz.mem [2212] = \nz.mem_2212_sv2v_reg ;
  assign \nz.mem [2211] = \nz.mem_2211_sv2v_reg ;
  assign \nz.mem [2210] = \nz.mem_2210_sv2v_reg ;
  assign \nz.mem [2209] = \nz.mem_2209_sv2v_reg ;
  assign \nz.mem [2208] = \nz.mem_2208_sv2v_reg ;
  assign \nz.mem [2207] = \nz.mem_2207_sv2v_reg ;
  assign \nz.mem [2206] = \nz.mem_2206_sv2v_reg ;
  assign \nz.mem [2205] = \nz.mem_2205_sv2v_reg ;
  assign \nz.mem [2204] = \nz.mem_2204_sv2v_reg ;
  assign \nz.mem [2203] = \nz.mem_2203_sv2v_reg ;
  assign \nz.mem [2202] = \nz.mem_2202_sv2v_reg ;
  assign \nz.mem [2201] = \nz.mem_2201_sv2v_reg ;
  assign \nz.mem [2200] = \nz.mem_2200_sv2v_reg ;
  assign \nz.mem [2199] = \nz.mem_2199_sv2v_reg ;
  assign \nz.mem [2198] = \nz.mem_2198_sv2v_reg ;
  assign \nz.mem [2197] = \nz.mem_2197_sv2v_reg ;
  assign \nz.mem [2196] = \nz.mem_2196_sv2v_reg ;
  assign \nz.mem [2195] = \nz.mem_2195_sv2v_reg ;
  assign \nz.mem [2194] = \nz.mem_2194_sv2v_reg ;
  assign \nz.mem [2193] = \nz.mem_2193_sv2v_reg ;
  assign \nz.mem [2192] = \nz.mem_2192_sv2v_reg ;
  assign \nz.mem [2191] = \nz.mem_2191_sv2v_reg ;
  assign \nz.mem [2190] = \nz.mem_2190_sv2v_reg ;
  assign \nz.mem [2189] = \nz.mem_2189_sv2v_reg ;
  assign \nz.mem [2188] = \nz.mem_2188_sv2v_reg ;
  assign \nz.mem [2187] = \nz.mem_2187_sv2v_reg ;
  assign \nz.mem [2186] = \nz.mem_2186_sv2v_reg ;
  assign \nz.mem [2185] = \nz.mem_2185_sv2v_reg ;
  assign \nz.mem [2184] = \nz.mem_2184_sv2v_reg ;
  assign \nz.mem [2183] = \nz.mem_2183_sv2v_reg ;
  assign \nz.mem [2182] = \nz.mem_2182_sv2v_reg ;
  assign \nz.mem [2181] = \nz.mem_2181_sv2v_reg ;
  assign \nz.mem [2180] = \nz.mem_2180_sv2v_reg ;
  assign \nz.mem [2179] = \nz.mem_2179_sv2v_reg ;
  assign \nz.mem [2178] = \nz.mem_2178_sv2v_reg ;
  assign \nz.mem [2177] = \nz.mem_2177_sv2v_reg ;
  assign \nz.mem [2176] = \nz.mem_2176_sv2v_reg ;
  assign \nz.mem [2175] = \nz.mem_2175_sv2v_reg ;
  assign \nz.mem [2174] = \nz.mem_2174_sv2v_reg ;
  assign \nz.mem [2173] = \nz.mem_2173_sv2v_reg ;
  assign \nz.mem [2172] = \nz.mem_2172_sv2v_reg ;
  assign \nz.mem [2171] = \nz.mem_2171_sv2v_reg ;
  assign \nz.mem [2170] = \nz.mem_2170_sv2v_reg ;
  assign \nz.mem [2169] = \nz.mem_2169_sv2v_reg ;
  assign \nz.mem [2168] = \nz.mem_2168_sv2v_reg ;
  assign \nz.mem [2167] = \nz.mem_2167_sv2v_reg ;
  assign \nz.mem [2166] = \nz.mem_2166_sv2v_reg ;
  assign \nz.mem [2165] = \nz.mem_2165_sv2v_reg ;
  assign \nz.mem [2164] = \nz.mem_2164_sv2v_reg ;
  assign \nz.mem [2163] = \nz.mem_2163_sv2v_reg ;
  assign \nz.mem [2162] = \nz.mem_2162_sv2v_reg ;
  assign \nz.mem [2161] = \nz.mem_2161_sv2v_reg ;
  assign \nz.mem [2160] = \nz.mem_2160_sv2v_reg ;
  assign \nz.mem [2159] = \nz.mem_2159_sv2v_reg ;
  assign \nz.mem [2158] = \nz.mem_2158_sv2v_reg ;
  assign \nz.mem [2157] = \nz.mem_2157_sv2v_reg ;
  assign \nz.mem [2156] = \nz.mem_2156_sv2v_reg ;
  assign \nz.mem [2155] = \nz.mem_2155_sv2v_reg ;
  assign \nz.mem [2154] = \nz.mem_2154_sv2v_reg ;
  assign \nz.mem [2153] = \nz.mem_2153_sv2v_reg ;
  assign \nz.mem [2152] = \nz.mem_2152_sv2v_reg ;
  assign \nz.mem [2151] = \nz.mem_2151_sv2v_reg ;
  assign \nz.mem [2150] = \nz.mem_2150_sv2v_reg ;
  assign \nz.mem [2149] = \nz.mem_2149_sv2v_reg ;
  assign \nz.mem [2148] = \nz.mem_2148_sv2v_reg ;
  assign \nz.mem [2147] = \nz.mem_2147_sv2v_reg ;
  assign \nz.mem [2146] = \nz.mem_2146_sv2v_reg ;
  assign \nz.mem [2145] = \nz.mem_2145_sv2v_reg ;
  assign \nz.mem [2144] = \nz.mem_2144_sv2v_reg ;
  assign \nz.mem [2143] = \nz.mem_2143_sv2v_reg ;
  assign \nz.mem [2142] = \nz.mem_2142_sv2v_reg ;
  assign \nz.mem [2141] = \nz.mem_2141_sv2v_reg ;
  assign \nz.mem [2140] = \nz.mem_2140_sv2v_reg ;
  assign \nz.mem [2139] = \nz.mem_2139_sv2v_reg ;
  assign \nz.mem [2138] = \nz.mem_2138_sv2v_reg ;
  assign \nz.mem [2137] = \nz.mem_2137_sv2v_reg ;
  assign \nz.mem [2136] = \nz.mem_2136_sv2v_reg ;
  assign \nz.mem [2135] = \nz.mem_2135_sv2v_reg ;
  assign \nz.mem [2134] = \nz.mem_2134_sv2v_reg ;
  assign \nz.mem [2133] = \nz.mem_2133_sv2v_reg ;
  assign \nz.mem [2132] = \nz.mem_2132_sv2v_reg ;
  assign \nz.mem [2131] = \nz.mem_2131_sv2v_reg ;
  assign \nz.mem [2130] = \nz.mem_2130_sv2v_reg ;
  assign \nz.mem [2129] = \nz.mem_2129_sv2v_reg ;
  assign \nz.mem [2128] = \nz.mem_2128_sv2v_reg ;
  assign \nz.mem [2127] = \nz.mem_2127_sv2v_reg ;
  assign \nz.mem [2126] = \nz.mem_2126_sv2v_reg ;
  assign \nz.mem [2125] = \nz.mem_2125_sv2v_reg ;
  assign \nz.mem [2124] = \nz.mem_2124_sv2v_reg ;
  assign \nz.mem [2123] = \nz.mem_2123_sv2v_reg ;
  assign \nz.mem [2122] = \nz.mem_2122_sv2v_reg ;
  assign \nz.mem [2121] = \nz.mem_2121_sv2v_reg ;
  assign \nz.mem [2120] = \nz.mem_2120_sv2v_reg ;
  assign \nz.mem [2119] = \nz.mem_2119_sv2v_reg ;
  assign \nz.mem [2118] = \nz.mem_2118_sv2v_reg ;
  assign \nz.mem [2117] = \nz.mem_2117_sv2v_reg ;
  assign \nz.mem [2116] = \nz.mem_2116_sv2v_reg ;
  assign \nz.mem [2115] = \nz.mem_2115_sv2v_reg ;
  assign \nz.mem [2114] = \nz.mem_2114_sv2v_reg ;
  assign \nz.mem [2113] = \nz.mem_2113_sv2v_reg ;
  assign \nz.mem [2112] = \nz.mem_2112_sv2v_reg ;
  assign \nz.mem [2111] = \nz.mem_2111_sv2v_reg ;
  assign \nz.mem [2110] = \nz.mem_2110_sv2v_reg ;
  assign \nz.mem [2109] = \nz.mem_2109_sv2v_reg ;
  assign \nz.mem [2108] = \nz.mem_2108_sv2v_reg ;
  assign \nz.mem [2107] = \nz.mem_2107_sv2v_reg ;
  assign \nz.mem [2106] = \nz.mem_2106_sv2v_reg ;
  assign \nz.mem [2105] = \nz.mem_2105_sv2v_reg ;
  assign \nz.mem [2104] = \nz.mem_2104_sv2v_reg ;
  assign \nz.mem [2103] = \nz.mem_2103_sv2v_reg ;
  assign \nz.mem [2102] = \nz.mem_2102_sv2v_reg ;
  assign \nz.mem [2101] = \nz.mem_2101_sv2v_reg ;
  assign \nz.mem [2100] = \nz.mem_2100_sv2v_reg ;
  assign \nz.mem [2099] = \nz.mem_2099_sv2v_reg ;
  assign \nz.mem [2098] = \nz.mem_2098_sv2v_reg ;
  assign \nz.mem [2097] = \nz.mem_2097_sv2v_reg ;
  assign \nz.mem [2096] = \nz.mem_2096_sv2v_reg ;
  assign \nz.mem [2095] = \nz.mem_2095_sv2v_reg ;
  assign \nz.mem [2094] = \nz.mem_2094_sv2v_reg ;
  assign \nz.mem [2093] = \nz.mem_2093_sv2v_reg ;
  assign \nz.mem [2092] = \nz.mem_2092_sv2v_reg ;
  assign \nz.mem [2091] = \nz.mem_2091_sv2v_reg ;
  assign \nz.mem [2090] = \nz.mem_2090_sv2v_reg ;
  assign \nz.mem [2089] = \nz.mem_2089_sv2v_reg ;
  assign \nz.mem [2088] = \nz.mem_2088_sv2v_reg ;
  assign \nz.mem [2087] = \nz.mem_2087_sv2v_reg ;
  assign \nz.mem [2086] = \nz.mem_2086_sv2v_reg ;
  assign \nz.mem [2085] = \nz.mem_2085_sv2v_reg ;
  assign \nz.mem [2084] = \nz.mem_2084_sv2v_reg ;
  assign \nz.mem [2083] = \nz.mem_2083_sv2v_reg ;
  assign \nz.mem [2082] = \nz.mem_2082_sv2v_reg ;
  assign \nz.mem [2081] = \nz.mem_2081_sv2v_reg ;
  assign \nz.mem [2080] = \nz.mem_2080_sv2v_reg ;
  assign \nz.mem [2079] = \nz.mem_2079_sv2v_reg ;
  assign \nz.mem [2078] = \nz.mem_2078_sv2v_reg ;
  assign \nz.mem [2077] = \nz.mem_2077_sv2v_reg ;
  assign \nz.mem [2076] = \nz.mem_2076_sv2v_reg ;
  assign \nz.mem [2075] = \nz.mem_2075_sv2v_reg ;
  assign \nz.mem [2074] = \nz.mem_2074_sv2v_reg ;
  assign \nz.mem [2073] = \nz.mem_2073_sv2v_reg ;
  assign \nz.mem [2072] = \nz.mem_2072_sv2v_reg ;
  assign \nz.mem [2071] = \nz.mem_2071_sv2v_reg ;
  assign \nz.mem [2070] = \nz.mem_2070_sv2v_reg ;
  assign \nz.mem [2069] = \nz.mem_2069_sv2v_reg ;
  assign \nz.mem [2068] = \nz.mem_2068_sv2v_reg ;
  assign \nz.mem [2067] = \nz.mem_2067_sv2v_reg ;
  assign \nz.mem [2066] = \nz.mem_2066_sv2v_reg ;
  assign \nz.mem [2065] = \nz.mem_2065_sv2v_reg ;
  assign \nz.mem [2064] = \nz.mem_2064_sv2v_reg ;
  assign \nz.mem [2063] = \nz.mem_2063_sv2v_reg ;
  assign \nz.mem [2062] = \nz.mem_2062_sv2v_reg ;
  assign \nz.mem [2061] = \nz.mem_2061_sv2v_reg ;
  assign \nz.mem [2060] = \nz.mem_2060_sv2v_reg ;
  assign \nz.mem [2059] = \nz.mem_2059_sv2v_reg ;
  assign \nz.mem [2058] = \nz.mem_2058_sv2v_reg ;
  assign \nz.mem [2057] = \nz.mem_2057_sv2v_reg ;
  assign \nz.mem [2056] = \nz.mem_2056_sv2v_reg ;
  assign \nz.mem [2055] = \nz.mem_2055_sv2v_reg ;
  assign \nz.mem [2054] = \nz.mem_2054_sv2v_reg ;
  assign \nz.mem [2053] = \nz.mem_2053_sv2v_reg ;
  assign \nz.mem [2052] = \nz.mem_2052_sv2v_reg ;
  assign \nz.mem [2051] = \nz.mem_2051_sv2v_reg ;
  assign \nz.mem [2050] = \nz.mem_2050_sv2v_reg ;
  assign \nz.mem [2049] = \nz.mem_2049_sv2v_reg ;
  assign \nz.mem [2048] = \nz.mem_2048_sv2v_reg ;
  assign \nz.mem [2047] = \nz.mem_2047_sv2v_reg ;
  assign \nz.mem [2046] = \nz.mem_2046_sv2v_reg ;
  assign \nz.mem [2045] = \nz.mem_2045_sv2v_reg ;
  assign \nz.mem [2044] = \nz.mem_2044_sv2v_reg ;
  assign \nz.mem [2043] = \nz.mem_2043_sv2v_reg ;
  assign \nz.mem [2042] = \nz.mem_2042_sv2v_reg ;
  assign \nz.mem [2041] = \nz.mem_2041_sv2v_reg ;
  assign \nz.mem [2040] = \nz.mem_2040_sv2v_reg ;
  assign \nz.mem [2039] = \nz.mem_2039_sv2v_reg ;
  assign \nz.mem [2038] = \nz.mem_2038_sv2v_reg ;
  assign \nz.mem [2037] = \nz.mem_2037_sv2v_reg ;
  assign \nz.mem [2036] = \nz.mem_2036_sv2v_reg ;
  assign \nz.mem [2035] = \nz.mem_2035_sv2v_reg ;
  assign \nz.mem [2034] = \nz.mem_2034_sv2v_reg ;
  assign \nz.mem [2033] = \nz.mem_2033_sv2v_reg ;
  assign \nz.mem [2032] = \nz.mem_2032_sv2v_reg ;
  assign \nz.mem [2031] = \nz.mem_2031_sv2v_reg ;
  assign \nz.mem [2030] = \nz.mem_2030_sv2v_reg ;
  assign \nz.mem [2029] = \nz.mem_2029_sv2v_reg ;
  assign \nz.mem [2028] = \nz.mem_2028_sv2v_reg ;
  assign \nz.mem [2027] = \nz.mem_2027_sv2v_reg ;
  assign \nz.mem [2026] = \nz.mem_2026_sv2v_reg ;
  assign \nz.mem [2025] = \nz.mem_2025_sv2v_reg ;
  assign \nz.mem [2024] = \nz.mem_2024_sv2v_reg ;
  assign \nz.mem [2023] = \nz.mem_2023_sv2v_reg ;
  assign \nz.mem [2022] = \nz.mem_2022_sv2v_reg ;
  assign \nz.mem [2021] = \nz.mem_2021_sv2v_reg ;
  assign \nz.mem [2020] = \nz.mem_2020_sv2v_reg ;
  assign \nz.mem [2019] = \nz.mem_2019_sv2v_reg ;
  assign \nz.mem [2018] = \nz.mem_2018_sv2v_reg ;
  assign \nz.mem [2017] = \nz.mem_2017_sv2v_reg ;
  assign \nz.mem [2016] = \nz.mem_2016_sv2v_reg ;
  assign \nz.mem [2015] = \nz.mem_2015_sv2v_reg ;
  assign \nz.mem [2014] = \nz.mem_2014_sv2v_reg ;
  assign \nz.mem [2013] = \nz.mem_2013_sv2v_reg ;
  assign \nz.mem [2012] = \nz.mem_2012_sv2v_reg ;
  assign \nz.mem [2011] = \nz.mem_2011_sv2v_reg ;
  assign \nz.mem [2010] = \nz.mem_2010_sv2v_reg ;
  assign \nz.mem [2009] = \nz.mem_2009_sv2v_reg ;
  assign \nz.mem [2008] = \nz.mem_2008_sv2v_reg ;
  assign \nz.mem [2007] = \nz.mem_2007_sv2v_reg ;
  assign \nz.mem [2006] = \nz.mem_2006_sv2v_reg ;
  assign \nz.mem [2005] = \nz.mem_2005_sv2v_reg ;
  assign \nz.mem [2004] = \nz.mem_2004_sv2v_reg ;
  assign \nz.mem [2003] = \nz.mem_2003_sv2v_reg ;
  assign \nz.mem [2002] = \nz.mem_2002_sv2v_reg ;
  assign \nz.mem [2001] = \nz.mem_2001_sv2v_reg ;
  assign \nz.mem [2000] = \nz.mem_2000_sv2v_reg ;
  assign \nz.mem [1999] = \nz.mem_1999_sv2v_reg ;
  assign \nz.mem [1998] = \nz.mem_1998_sv2v_reg ;
  assign \nz.mem [1997] = \nz.mem_1997_sv2v_reg ;
  assign \nz.mem [1996] = \nz.mem_1996_sv2v_reg ;
  assign \nz.mem [1995] = \nz.mem_1995_sv2v_reg ;
  assign \nz.mem [1994] = \nz.mem_1994_sv2v_reg ;
  assign \nz.mem [1993] = \nz.mem_1993_sv2v_reg ;
  assign \nz.mem [1992] = \nz.mem_1992_sv2v_reg ;
  assign \nz.mem [1991] = \nz.mem_1991_sv2v_reg ;
  assign \nz.mem [1990] = \nz.mem_1990_sv2v_reg ;
  assign \nz.mem [1989] = \nz.mem_1989_sv2v_reg ;
  assign \nz.mem [1988] = \nz.mem_1988_sv2v_reg ;
  assign \nz.mem [1987] = \nz.mem_1987_sv2v_reg ;
  assign \nz.mem [1986] = \nz.mem_1986_sv2v_reg ;
  assign \nz.mem [1985] = \nz.mem_1985_sv2v_reg ;
  assign \nz.mem [1984] = \nz.mem_1984_sv2v_reg ;
  assign \nz.mem [1983] = \nz.mem_1983_sv2v_reg ;
  assign \nz.mem [1982] = \nz.mem_1982_sv2v_reg ;
  assign \nz.mem [1981] = \nz.mem_1981_sv2v_reg ;
  assign \nz.mem [1980] = \nz.mem_1980_sv2v_reg ;
  assign \nz.mem [1979] = \nz.mem_1979_sv2v_reg ;
  assign \nz.mem [1978] = \nz.mem_1978_sv2v_reg ;
  assign \nz.mem [1977] = \nz.mem_1977_sv2v_reg ;
  assign \nz.mem [1976] = \nz.mem_1976_sv2v_reg ;
  assign \nz.mem [1975] = \nz.mem_1975_sv2v_reg ;
  assign \nz.mem [1974] = \nz.mem_1974_sv2v_reg ;
  assign \nz.mem [1973] = \nz.mem_1973_sv2v_reg ;
  assign \nz.mem [1972] = \nz.mem_1972_sv2v_reg ;
  assign \nz.mem [1971] = \nz.mem_1971_sv2v_reg ;
  assign \nz.mem [1970] = \nz.mem_1970_sv2v_reg ;
  assign \nz.mem [1969] = \nz.mem_1969_sv2v_reg ;
  assign \nz.mem [1968] = \nz.mem_1968_sv2v_reg ;
  assign \nz.mem [1967] = \nz.mem_1967_sv2v_reg ;
  assign \nz.mem [1966] = \nz.mem_1966_sv2v_reg ;
  assign \nz.mem [1965] = \nz.mem_1965_sv2v_reg ;
  assign \nz.mem [1964] = \nz.mem_1964_sv2v_reg ;
  assign \nz.mem [1963] = \nz.mem_1963_sv2v_reg ;
  assign \nz.mem [1962] = \nz.mem_1962_sv2v_reg ;
  assign \nz.mem [1961] = \nz.mem_1961_sv2v_reg ;
  assign \nz.mem [1960] = \nz.mem_1960_sv2v_reg ;
  assign \nz.mem [1959] = \nz.mem_1959_sv2v_reg ;
  assign \nz.mem [1958] = \nz.mem_1958_sv2v_reg ;
  assign \nz.mem [1957] = \nz.mem_1957_sv2v_reg ;
  assign \nz.mem [1956] = \nz.mem_1956_sv2v_reg ;
  assign \nz.mem [1955] = \nz.mem_1955_sv2v_reg ;
  assign \nz.mem [1954] = \nz.mem_1954_sv2v_reg ;
  assign \nz.mem [1953] = \nz.mem_1953_sv2v_reg ;
  assign \nz.mem [1952] = \nz.mem_1952_sv2v_reg ;
  assign \nz.mem [1951] = \nz.mem_1951_sv2v_reg ;
  assign \nz.mem [1950] = \nz.mem_1950_sv2v_reg ;
  assign \nz.mem [1949] = \nz.mem_1949_sv2v_reg ;
  assign \nz.mem [1948] = \nz.mem_1948_sv2v_reg ;
  assign \nz.mem [1947] = \nz.mem_1947_sv2v_reg ;
  assign \nz.mem [1946] = \nz.mem_1946_sv2v_reg ;
  assign \nz.mem [1945] = \nz.mem_1945_sv2v_reg ;
  assign \nz.mem [1944] = \nz.mem_1944_sv2v_reg ;
  assign \nz.mem [1943] = \nz.mem_1943_sv2v_reg ;
  assign \nz.mem [1942] = \nz.mem_1942_sv2v_reg ;
  assign \nz.mem [1941] = \nz.mem_1941_sv2v_reg ;
  assign \nz.mem [1940] = \nz.mem_1940_sv2v_reg ;
  assign \nz.mem [1939] = \nz.mem_1939_sv2v_reg ;
  assign \nz.mem [1938] = \nz.mem_1938_sv2v_reg ;
  assign \nz.mem [1937] = \nz.mem_1937_sv2v_reg ;
  assign \nz.mem [1936] = \nz.mem_1936_sv2v_reg ;
  assign \nz.mem [1935] = \nz.mem_1935_sv2v_reg ;
  assign \nz.mem [1934] = \nz.mem_1934_sv2v_reg ;
  assign \nz.mem [1933] = \nz.mem_1933_sv2v_reg ;
  assign \nz.mem [1932] = \nz.mem_1932_sv2v_reg ;
  assign \nz.mem [1931] = \nz.mem_1931_sv2v_reg ;
  assign \nz.mem [1930] = \nz.mem_1930_sv2v_reg ;
  assign \nz.mem [1929] = \nz.mem_1929_sv2v_reg ;
  assign \nz.mem [1928] = \nz.mem_1928_sv2v_reg ;
  assign \nz.mem [1927] = \nz.mem_1927_sv2v_reg ;
  assign \nz.mem [1926] = \nz.mem_1926_sv2v_reg ;
  assign \nz.mem [1925] = \nz.mem_1925_sv2v_reg ;
  assign \nz.mem [1924] = \nz.mem_1924_sv2v_reg ;
  assign \nz.mem [1923] = \nz.mem_1923_sv2v_reg ;
  assign \nz.mem [1922] = \nz.mem_1922_sv2v_reg ;
  assign \nz.mem [1921] = \nz.mem_1921_sv2v_reg ;
  assign \nz.mem [1920] = \nz.mem_1920_sv2v_reg ;
  assign \nz.mem [1919] = \nz.mem_1919_sv2v_reg ;
  assign \nz.mem [1918] = \nz.mem_1918_sv2v_reg ;
  assign \nz.mem [1917] = \nz.mem_1917_sv2v_reg ;
  assign \nz.mem [1916] = \nz.mem_1916_sv2v_reg ;
  assign \nz.mem [1915] = \nz.mem_1915_sv2v_reg ;
  assign \nz.mem [1914] = \nz.mem_1914_sv2v_reg ;
  assign \nz.mem [1913] = \nz.mem_1913_sv2v_reg ;
  assign \nz.mem [1912] = \nz.mem_1912_sv2v_reg ;
  assign \nz.mem [1911] = \nz.mem_1911_sv2v_reg ;
  assign \nz.mem [1910] = \nz.mem_1910_sv2v_reg ;
  assign \nz.mem [1909] = \nz.mem_1909_sv2v_reg ;
  assign \nz.mem [1908] = \nz.mem_1908_sv2v_reg ;
  assign \nz.mem [1907] = \nz.mem_1907_sv2v_reg ;
  assign \nz.mem [1906] = \nz.mem_1906_sv2v_reg ;
  assign \nz.mem [1905] = \nz.mem_1905_sv2v_reg ;
  assign \nz.mem [1904] = \nz.mem_1904_sv2v_reg ;
  assign \nz.mem [1903] = \nz.mem_1903_sv2v_reg ;
  assign \nz.mem [1902] = \nz.mem_1902_sv2v_reg ;
  assign \nz.mem [1901] = \nz.mem_1901_sv2v_reg ;
  assign \nz.mem [1900] = \nz.mem_1900_sv2v_reg ;
  assign \nz.mem [1899] = \nz.mem_1899_sv2v_reg ;
  assign \nz.mem [1898] = \nz.mem_1898_sv2v_reg ;
  assign \nz.mem [1897] = \nz.mem_1897_sv2v_reg ;
  assign \nz.mem [1896] = \nz.mem_1896_sv2v_reg ;
  assign \nz.mem [1895] = \nz.mem_1895_sv2v_reg ;
  assign \nz.mem [1894] = \nz.mem_1894_sv2v_reg ;
  assign \nz.mem [1893] = \nz.mem_1893_sv2v_reg ;
  assign \nz.mem [1892] = \nz.mem_1892_sv2v_reg ;
  assign \nz.mem [1891] = \nz.mem_1891_sv2v_reg ;
  assign \nz.mem [1890] = \nz.mem_1890_sv2v_reg ;
  assign \nz.mem [1889] = \nz.mem_1889_sv2v_reg ;
  assign \nz.mem [1888] = \nz.mem_1888_sv2v_reg ;
  assign \nz.mem [1887] = \nz.mem_1887_sv2v_reg ;
  assign \nz.mem [1886] = \nz.mem_1886_sv2v_reg ;
  assign \nz.mem [1885] = \nz.mem_1885_sv2v_reg ;
  assign \nz.mem [1884] = \nz.mem_1884_sv2v_reg ;
  assign \nz.mem [1883] = \nz.mem_1883_sv2v_reg ;
  assign \nz.mem [1882] = \nz.mem_1882_sv2v_reg ;
  assign \nz.mem [1881] = \nz.mem_1881_sv2v_reg ;
  assign \nz.mem [1880] = \nz.mem_1880_sv2v_reg ;
  assign \nz.mem [1879] = \nz.mem_1879_sv2v_reg ;
  assign \nz.mem [1878] = \nz.mem_1878_sv2v_reg ;
  assign \nz.mem [1877] = \nz.mem_1877_sv2v_reg ;
  assign \nz.mem [1876] = \nz.mem_1876_sv2v_reg ;
  assign \nz.mem [1875] = \nz.mem_1875_sv2v_reg ;
  assign \nz.mem [1874] = \nz.mem_1874_sv2v_reg ;
  assign \nz.mem [1873] = \nz.mem_1873_sv2v_reg ;
  assign \nz.mem [1872] = \nz.mem_1872_sv2v_reg ;
  assign \nz.mem [1871] = \nz.mem_1871_sv2v_reg ;
  assign \nz.mem [1870] = \nz.mem_1870_sv2v_reg ;
  assign \nz.mem [1869] = \nz.mem_1869_sv2v_reg ;
  assign \nz.mem [1868] = \nz.mem_1868_sv2v_reg ;
  assign \nz.mem [1867] = \nz.mem_1867_sv2v_reg ;
  assign \nz.mem [1866] = \nz.mem_1866_sv2v_reg ;
  assign \nz.mem [1865] = \nz.mem_1865_sv2v_reg ;
  assign \nz.mem [1864] = \nz.mem_1864_sv2v_reg ;
  assign \nz.mem [1863] = \nz.mem_1863_sv2v_reg ;
  assign \nz.mem [1862] = \nz.mem_1862_sv2v_reg ;
  assign \nz.mem [1861] = \nz.mem_1861_sv2v_reg ;
  assign \nz.mem [1860] = \nz.mem_1860_sv2v_reg ;
  assign \nz.mem [1859] = \nz.mem_1859_sv2v_reg ;
  assign \nz.mem [1858] = \nz.mem_1858_sv2v_reg ;
  assign \nz.mem [1857] = \nz.mem_1857_sv2v_reg ;
  assign \nz.mem [1856] = \nz.mem_1856_sv2v_reg ;
  assign \nz.mem [1855] = \nz.mem_1855_sv2v_reg ;
  assign \nz.mem [1854] = \nz.mem_1854_sv2v_reg ;
  assign \nz.mem [1853] = \nz.mem_1853_sv2v_reg ;
  assign \nz.mem [1852] = \nz.mem_1852_sv2v_reg ;
  assign \nz.mem [1851] = \nz.mem_1851_sv2v_reg ;
  assign \nz.mem [1850] = \nz.mem_1850_sv2v_reg ;
  assign \nz.mem [1849] = \nz.mem_1849_sv2v_reg ;
  assign \nz.mem [1848] = \nz.mem_1848_sv2v_reg ;
  assign \nz.mem [1847] = \nz.mem_1847_sv2v_reg ;
  assign \nz.mem [1846] = \nz.mem_1846_sv2v_reg ;
  assign \nz.mem [1845] = \nz.mem_1845_sv2v_reg ;
  assign \nz.mem [1844] = \nz.mem_1844_sv2v_reg ;
  assign \nz.mem [1843] = \nz.mem_1843_sv2v_reg ;
  assign \nz.mem [1842] = \nz.mem_1842_sv2v_reg ;
  assign \nz.mem [1841] = \nz.mem_1841_sv2v_reg ;
  assign \nz.mem [1840] = \nz.mem_1840_sv2v_reg ;
  assign \nz.mem [1839] = \nz.mem_1839_sv2v_reg ;
  assign \nz.mem [1838] = \nz.mem_1838_sv2v_reg ;
  assign \nz.mem [1837] = \nz.mem_1837_sv2v_reg ;
  assign \nz.mem [1836] = \nz.mem_1836_sv2v_reg ;
  assign \nz.mem [1835] = \nz.mem_1835_sv2v_reg ;
  assign \nz.mem [1834] = \nz.mem_1834_sv2v_reg ;
  assign \nz.mem [1833] = \nz.mem_1833_sv2v_reg ;
  assign \nz.mem [1832] = \nz.mem_1832_sv2v_reg ;
  assign \nz.mem [1831] = \nz.mem_1831_sv2v_reg ;
  assign \nz.mem [1830] = \nz.mem_1830_sv2v_reg ;
  assign \nz.mem [1829] = \nz.mem_1829_sv2v_reg ;
  assign \nz.mem [1828] = \nz.mem_1828_sv2v_reg ;
  assign \nz.mem [1827] = \nz.mem_1827_sv2v_reg ;
  assign \nz.mem [1826] = \nz.mem_1826_sv2v_reg ;
  assign \nz.mem [1825] = \nz.mem_1825_sv2v_reg ;
  assign \nz.mem [1824] = \nz.mem_1824_sv2v_reg ;
  assign \nz.mem [1823] = \nz.mem_1823_sv2v_reg ;
  assign \nz.mem [1822] = \nz.mem_1822_sv2v_reg ;
  assign \nz.mem [1821] = \nz.mem_1821_sv2v_reg ;
  assign \nz.mem [1820] = \nz.mem_1820_sv2v_reg ;
  assign \nz.mem [1819] = \nz.mem_1819_sv2v_reg ;
  assign \nz.mem [1818] = \nz.mem_1818_sv2v_reg ;
  assign \nz.mem [1817] = \nz.mem_1817_sv2v_reg ;
  assign \nz.mem [1816] = \nz.mem_1816_sv2v_reg ;
  assign \nz.mem [1815] = \nz.mem_1815_sv2v_reg ;
  assign \nz.mem [1814] = \nz.mem_1814_sv2v_reg ;
  assign \nz.mem [1813] = \nz.mem_1813_sv2v_reg ;
  assign \nz.mem [1812] = \nz.mem_1812_sv2v_reg ;
  assign \nz.mem [1811] = \nz.mem_1811_sv2v_reg ;
  assign \nz.mem [1810] = \nz.mem_1810_sv2v_reg ;
  assign \nz.mem [1809] = \nz.mem_1809_sv2v_reg ;
  assign \nz.mem [1808] = \nz.mem_1808_sv2v_reg ;
  assign \nz.mem [1807] = \nz.mem_1807_sv2v_reg ;
  assign \nz.mem [1806] = \nz.mem_1806_sv2v_reg ;
  assign \nz.mem [1805] = \nz.mem_1805_sv2v_reg ;
  assign \nz.mem [1804] = \nz.mem_1804_sv2v_reg ;
  assign \nz.mem [1803] = \nz.mem_1803_sv2v_reg ;
  assign \nz.mem [1802] = \nz.mem_1802_sv2v_reg ;
  assign \nz.mem [1801] = \nz.mem_1801_sv2v_reg ;
  assign \nz.mem [1800] = \nz.mem_1800_sv2v_reg ;
  assign \nz.mem [1799] = \nz.mem_1799_sv2v_reg ;
  assign \nz.mem [1798] = \nz.mem_1798_sv2v_reg ;
  assign \nz.mem [1797] = \nz.mem_1797_sv2v_reg ;
  assign \nz.mem [1796] = \nz.mem_1796_sv2v_reg ;
  assign \nz.mem [1795] = \nz.mem_1795_sv2v_reg ;
  assign \nz.mem [1794] = \nz.mem_1794_sv2v_reg ;
  assign \nz.mem [1793] = \nz.mem_1793_sv2v_reg ;
  assign \nz.mem [1792] = \nz.mem_1792_sv2v_reg ;
  assign \nz.mem [1791] = \nz.mem_1791_sv2v_reg ;
  assign \nz.mem [1790] = \nz.mem_1790_sv2v_reg ;
  assign \nz.mem [1789] = \nz.mem_1789_sv2v_reg ;
  assign \nz.mem [1788] = \nz.mem_1788_sv2v_reg ;
  assign \nz.mem [1787] = \nz.mem_1787_sv2v_reg ;
  assign \nz.mem [1786] = \nz.mem_1786_sv2v_reg ;
  assign \nz.mem [1785] = \nz.mem_1785_sv2v_reg ;
  assign \nz.mem [1784] = \nz.mem_1784_sv2v_reg ;
  assign \nz.mem [1783] = \nz.mem_1783_sv2v_reg ;
  assign \nz.mem [1782] = \nz.mem_1782_sv2v_reg ;
  assign \nz.mem [1781] = \nz.mem_1781_sv2v_reg ;
  assign \nz.mem [1780] = \nz.mem_1780_sv2v_reg ;
  assign \nz.mem [1779] = \nz.mem_1779_sv2v_reg ;
  assign \nz.mem [1778] = \nz.mem_1778_sv2v_reg ;
  assign \nz.mem [1777] = \nz.mem_1777_sv2v_reg ;
  assign \nz.mem [1776] = \nz.mem_1776_sv2v_reg ;
  assign \nz.mem [1775] = \nz.mem_1775_sv2v_reg ;
  assign \nz.mem [1774] = \nz.mem_1774_sv2v_reg ;
  assign \nz.mem [1773] = \nz.mem_1773_sv2v_reg ;
  assign \nz.mem [1772] = \nz.mem_1772_sv2v_reg ;
  assign \nz.mem [1771] = \nz.mem_1771_sv2v_reg ;
  assign \nz.mem [1770] = \nz.mem_1770_sv2v_reg ;
  assign \nz.mem [1769] = \nz.mem_1769_sv2v_reg ;
  assign \nz.mem [1768] = \nz.mem_1768_sv2v_reg ;
  assign \nz.mem [1767] = \nz.mem_1767_sv2v_reg ;
  assign \nz.mem [1766] = \nz.mem_1766_sv2v_reg ;
  assign \nz.mem [1765] = \nz.mem_1765_sv2v_reg ;
  assign \nz.mem [1764] = \nz.mem_1764_sv2v_reg ;
  assign \nz.mem [1763] = \nz.mem_1763_sv2v_reg ;
  assign \nz.mem [1762] = \nz.mem_1762_sv2v_reg ;
  assign \nz.mem [1761] = \nz.mem_1761_sv2v_reg ;
  assign \nz.mem [1760] = \nz.mem_1760_sv2v_reg ;
  assign \nz.mem [1759] = \nz.mem_1759_sv2v_reg ;
  assign \nz.mem [1758] = \nz.mem_1758_sv2v_reg ;
  assign \nz.mem [1757] = \nz.mem_1757_sv2v_reg ;
  assign \nz.mem [1756] = \nz.mem_1756_sv2v_reg ;
  assign \nz.mem [1755] = \nz.mem_1755_sv2v_reg ;
  assign \nz.mem [1754] = \nz.mem_1754_sv2v_reg ;
  assign \nz.mem [1753] = \nz.mem_1753_sv2v_reg ;
  assign \nz.mem [1752] = \nz.mem_1752_sv2v_reg ;
  assign \nz.mem [1751] = \nz.mem_1751_sv2v_reg ;
  assign \nz.mem [1750] = \nz.mem_1750_sv2v_reg ;
  assign \nz.mem [1749] = \nz.mem_1749_sv2v_reg ;
  assign \nz.mem [1748] = \nz.mem_1748_sv2v_reg ;
  assign \nz.mem [1747] = \nz.mem_1747_sv2v_reg ;
  assign \nz.mem [1746] = \nz.mem_1746_sv2v_reg ;
  assign \nz.mem [1745] = \nz.mem_1745_sv2v_reg ;
  assign \nz.mem [1744] = \nz.mem_1744_sv2v_reg ;
  assign \nz.mem [1743] = \nz.mem_1743_sv2v_reg ;
  assign \nz.mem [1742] = \nz.mem_1742_sv2v_reg ;
  assign \nz.mem [1741] = \nz.mem_1741_sv2v_reg ;
  assign \nz.mem [1740] = \nz.mem_1740_sv2v_reg ;
  assign \nz.mem [1739] = \nz.mem_1739_sv2v_reg ;
  assign \nz.mem [1738] = \nz.mem_1738_sv2v_reg ;
  assign \nz.mem [1737] = \nz.mem_1737_sv2v_reg ;
  assign \nz.mem [1736] = \nz.mem_1736_sv2v_reg ;
  assign \nz.mem [1735] = \nz.mem_1735_sv2v_reg ;
  assign \nz.mem [1734] = \nz.mem_1734_sv2v_reg ;
  assign \nz.mem [1733] = \nz.mem_1733_sv2v_reg ;
  assign \nz.mem [1732] = \nz.mem_1732_sv2v_reg ;
  assign \nz.mem [1731] = \nz.mem_1731_sv2v_reg ;
  assign \nz.mem [1730] = \nz.mem_1730_sv2v_reg ;
  assign \nz.mem [1729] = \nz.mem_1729_sv2v_reg ;
  assign \nz.mem [1728] = \nz.mem_1728_sv2v_reg ;
  assign \nz.mem [1727] = \nz.mem_1727_sv2v_reg ;
  assign \nz.mem [1726] = \nz.mem_1726_sv2v_reg ;
  assign \nz.mem [1725] = \nz.mem_1725_sv2v_reg ;
  assign \nz.mem [1724] = \nz.mem_1724_sv2v_reg ;
  assign \nz.mem [1723] = \nz.mem_1723_sv2v_reg ;
  assign \nz.mem [1722] = \nz.mem_1722_sv2v_reg ;
  assign \nz.mem [1721] = \nz.mem_1721_sv2v_reg ;
  assign \nz.mem [1720] = \nz.mem_1720_sv2v_reg ;
  assign \nz.mem [1719] = \nz.mem_1719_sv2v_reg ;
  assign \nz.mem [1718] = \nz.mem_1718_sv2v_reg ;
  assign \nz.mem [1717] = \nz.mem_1717_sv2v_reg ;
  assign \nz.mem [1716] = \nz.mem_1716_sv2v_reg ;
  assign \nz.mem [1715] = \nz.mem_1715_sv2v_reg ;
  assign \nz.mem [1714] = \nz.mem_1714_sv2v_reg ;
  assign \nz.mem [1713] = \nz.mem_1713_sv2v_reg ;
  assign \nz.mem [1712] = \nz.mem_1712_sv2v_reg ;
  assign \nz.mem [1711] = \nz.mem_1711_sv2v_reg ;
  assign \nz.mem [1710] = \nz.mem_1710_sv2v_reg ;
  assign \nz.mem [1709] = \nz.mem_1709_sv2v_reg ;
  assign \nz.mem [1708] = \nz.mem_1708_sv2v_reg ;
  assign \nz.mem [1707] = \nz.mem_1707_sv2v_reg ;
  assign \nz.mem [1706] = \nz.mem_1706_sv2v_reg ;
  assign \nz.mem [1705] = \nz.mem_1705_sv2v_reg ;
  assign \nz.mem [1704] = \nz.mem_1704_sv2v_reg ;
  assign \nz.mem [1703] = \nz.mem_1703_sv2v_reg ;
  assign \nz.mem [1702] = \nz.mem_1702_sv2v_reg ;
  assign \nz.mem [1701] = \nz.mem_1701_sv2v_reg ;
  assign \nz.mem [1700] = \nz.mem_1700_sv2v_reg ;
  assign \nz.mem [1699] = \nz.mem_1699_sv2v_reg ;
  assign \nz.mem [1698] = \nz.mem_1698_sv2v_reg ;
  assign \nz.mem [1697] = \nz.mem_1697_sv2v_reg ;
  assign \nz.mem [1696] = \nz.mem_1696_sv2v_reg ;
  assign \nz.mem [1695] = \nz.mem_1695_sv2v_reg ;
  assign \nz.mem [1694] = \nz.mem_1694_sv2v_reg ;
  assign \nz.mem [1693] = \nz.mem_1693_sv2v_reg ;
  assign \nz.mem [1692] = \nz.mem_1692_sv2v_reg ;
  assign \nz.mem [1691] = \nz.mem_1691_sv2v_reg ;
  assign \nz.mem [1690] = \nz.mem_1690_sv2v_reg ;
  assign \nz.mem [1689] = \nz.mem_1689_sv2v_reg ;
  assign \nz.mem [1688] = \nz.mem_1688_sv2v_reg ;
  assign \nz.mem [1687] = \nz.mem_1687_sv2v_reg ;
  assign \nz.mem [1686] = \nz.mem_1686_sv2v_reg ;
  assign \nz.mem [1685] = \nz.mem_1685_sv2v_reg ;
  assign \nz.mem [1684] = \nz.mem_1684_sv2v_reg ;
  assign \nz.mem [1683] = \nz.mem_1683_sv2v_reg ;
  assign \nz.mem [1682] = \nz.mem_1682_sv2v_reg ;
  assign \nz.mem [1681] = \nz.mem_1681_sv2v_reg ;
  assign \nz.mem [1680] = \nz.mem_1680_sv2v_reg ;
  assign \nz.mem [1679] = \nz.mem_1679_sv2v_reg ;
  assign \nz.mem [1678] = \nz.mem_1678_sv2v_reg ;
  assign \nz.mem [1677] = \nz.mem_1677_sv2v_reg ;
  assign \nz.mem [1676] = \nz.mem_1676_sv2v_reg ;
  assign \nz.mem [1675] = \nz.mem_1675_sv2v_reg ;
  assign \nz.mem [1674] = \nz.mem_1674_sv2v_reg ;
  assign \nz.mem [1673] = \nz.mem_1673_sv2v_reg ;
  assign \nz.mem [1672] = \nz.mem_1672_sv2v_reg ;
  assign \nz.mem [1671] = \nz.mem_1671_sv2v_reg ;
  assign \nz.mem [1670] = \nz.mem_1670_sv2v_reg ;
  assign \nz.mem [1669] = \nz.mem_1669_sv2v_reg ;
  assign \nz.mem [1668] = \nz.mem_1668_sv2v_reg ;
  assign \nz.mem [1667] = \nz.mem_1667_sv2v_reg ;
  assign \nz.mem [1666] = \nz.mem_1666_sv2v_reg ;
  assign \nz.mem [1665] = \nz.mem_1665_sv2v_reg ;
  assign \nz.mem [1664] = \nz.mem_1664_sv2v_reg ;
  assign \nz.mem [1663] = \nz.mem_1663_sv2v_reg ;
  assign \nz.mem [1662] = \nz.mem_1662_sv2v_reg ;
  assign \nz.mem [1661] = \nz.mem_1661_sv2v_reg ;
  assign \nz.mem [1660] = \nz.mem_1660_sv2v_reg ;
  assign \nz.mem [1659] = \nz.mem_1659_sv2v_reg ;
  assign \nz.mem [1658] = \nz.mem_1658_sv2v_reg ;
  assign \nz.mem [1657] = \nz.mem_1657_sv2v_reg ;
  assign \nz.mem [1656] = \nz.mem_1656_sv2v_reg ;
  assign \nz.mem [1655] = \nz.mem_1655_sv2v_reg ;
  assign \nz.mem [1654] = \nz.mem_1654_sv2v_reg ;
  assign \nz.mem [1653] = \nz.mem_1653_sv2v_reg ;
  assign \nz.mem [1652] = \nz.mem_1652_sv2v_reg ;
  assign \nz.mem [1651] = \nz.mem_1651_sv2v_reg ;
  assign \nz.mem [1650] = \nz.mem_1650_sv2v_reg ;
  assign \nz.mem [1649] = \nz.mem_1649_sv2v_reg ;
  assign \nz.mem [1648] = \nz.mem_1648_sv2v_reg ;
  assign \nz.mem [1647] = \nz.mem_1647_sv2v_reg ;
  assign \nz.mem [1646] = \nz.mem_1646_sv2v_reg ;
  assign \nz.mem [1645] = \nz.mem_1645_sv2v_reg ;
  assign \nz.mem [1644] = \nz.mem_1644_sv2v_reg ;
  assign \nz.mem [1643] = \nz.mem_1643_sv2v_reg ;
  assign \nz.mem [1642] = \nz.mem_1642_sv2v_reg ;
  assign \nz.mem [1641] = \nz.mem_1641_sv2v_reg ;
  assign \nz.mem [1640] = \nz.mem_1640_sv2v_reg ;
  assign \nz.mem [1639] = \nz.mem_1639_sv2v_reg ;
  assign \nz.mem [1638] = \nz.mem_1638_sv2v_reg ;
  assign \nz.mem [1637] = \nz.mem_1637_sv2v_reg ;
  assign \nz.mem [1636] = \nz.mem_1636_sv2v_reg ;
  assign \nz.mem [1635] = \nz.mem_1635_sv2v_reg ;
  assign \nz.mem [1634] = \nz.mem_1634_sv2v_reg ;
  assign \nz.mem [1633] = \nz.mem_1633_sv2v_reg ;
  assign \nz.mem [1632] = \nz.mem_1632_sv2v_reg ;
  assign \nz.mem [1631] = \nz.mem_1631_sv2v_reg ;
  assign \nz.mem [1630] = \nz.mem_1630_sv2v_reg ;
  assign \nz.mem [1629] = \nz.mem_1629_sv2v_reg ;
  assign \nz.mem [1628] = \nz.mem_1628_sv2v_reg ;
  assign \nz.mem [1627] = \nz.mem_1627_sv2v_reg ;
  assign \nz.mem [1626] = \nz.mem_1626_sv2v_reg ;
  assign \nz.mem [1625] = \nz.mem_1625_sv2v_reg ;
  assign \nz.mem [1624] = \nz.mem_1624_sv2v_reg ;
  assign \nz.mem [1623] = \nz.mem_1623_sv2v_reg ;
  assign \nz.mem [1622] = \nz.mem_1622_sv2v_reg ;
  assign \nz.mem [1621] = \nz.mem_1621_sv2v_reg ;
  assign \nz.mem [1620] = \nz.mem_1620_sv2v_reg ;
  assign \nz.mem [1619] = \nz.mem_1619_sv2v_reg ;
  assign \nz.mem [1618] = \nz.mem_1618_sv2v_reg ;
  assign \nz.mem [1617] = \nz.mem_1617_sv2v_reg ;
  assign \nz.mem [1616] = \nz.mem_1616_sv2v_reg ;
  assign \nz.mem [1615] = \nz.mem_1615_sv2v_reg ;
  assign \nz.mem [1614] = \nz.mem_1614_sv2v_reg ;
  assign \nz.mem [1613] = \nz.mem_1613_sv2v_reg ;
  assign \nz.mem [1612] = \nz.mem_1612_sv2v_reg ;
  assign \nz.mem [1611] = \nz.mem_1611_sv2v_reg ;
  assign \nz.mem [1610] = \nz.mem_1610_sv2v_reg ;
  assign \nz.mem [1609] = \nz.mem_1609_sv2v_reg ;
  assign \nz.mem [1608] = \nz.mem_1608_sv2v_reg ;
  assign \nz.mem [1607] = \nz.mem_1607_sv2v_reg ;
  assign \nz.mem [1606] = \nz.mem_1606_sv2v_reg ;
  assign \nz.mem [1605] = \nz.mem_1605_sv2v_reg ;
  assign \nz.mem [1604] = \nz.mem_1604_sv2v_reg ;
  assign \nz.mem [1603] = \nz.mem_1603_sv2v_reg ;
  assign \nz.mem [1602] = \nz.mem_1602_sv2v_reg ;
  assign \nz.mem [1601] = \nz.mem_1601_sv2v_reg ;
  assign \nz.mem [1600] = \nz.mem_1600_sv2v_reg ;
  assign \nz.mem [1599] = \nz.mem_1599_sv2v_reg ;
  assign \nz.mem [1598] = \nz.mem_1598_sv2v_reg ;
  assign \nz.mem [1597] = \nz.mem_1597_sv2v_reg ;
  assign \nz.mem [1596] = \nz.mem_1596_sv2v_reg ;
  assign \nz.mem [1595] = \nz.mem_1595_sv2v_reg ;
  assign \nz.mem [1594] = \nz.mem_1594_sv2v_reg ;
  assign \nz.mem [1593] = \nz.mem_1593_sv2v_reg ;
  assign \nz.mem [1592] = \nz.mem_1592_sv2v_reg ;
  assign \nz.mem [1591] = \nz.mem_1591_sv2v_reg ;
  assign \nz.mem [1590] = \nz.mem_1590_sv2v_reg ;
  assign \nz.mem [1589] = \nz.mem_1589_sv2v_reg ;
  assign \nz.mem [1588] = \nz.mem_1588_sv2v_reg ;
  assign \nz.mem [1587] = \nz.mem_1587_sv2v_reg ;
  assign \nz.mem [1586] = \nz.mem_1586_sv2v_reg ;
  assign \nz.mem [1585] = \nz.mem_1585_sv2v_reg ;
  assign \nz.mem [1584] = \nz.mem_1584_sv2v_reg ;
  assign \nz.mem [1583] = \nz.mem_1583_sv2v_reg ;
  assign \nz.mem [1582] = \nz.mem_1582_sv2v_reg ;
  assign \nz.mem [1581] = \nz.mem_1581_sv2v_reg ;
  assign \nz.mem [1580] = \nz.mem_1580_sv2v_reg ;
  assign \nz.mem [1579] = \nz.mem_1579_sv2v_reg ;
  assign \nz.mem [1578] = \nz.mem_1578_sv2v_reg ;
  assign \nz.mem [1577] = \nz.mem_1577_sv2v_reg ;
  assign \nz.mem [1576] = \nz.mem_1576_sv2v_reg ;
  assign \nz.mem [1575] = \nz.mem_1575_sv2v_reg ;
  assign \nz.mem [1574] = \nz.mem_1574_sv2v_reg ;
  assign \nz.mem [1573] = \nz.mem_1573_sv2v_reg ;
  assign \nz.mem [1572] = \nz.mem_1572_sv2v_reg ;
  assign \nz.mem [1571] = \nz.mem_1571_sv2v_reg ;
  assign \nz.mem [1570] = \nz.mem_1570_sv2v_reg ;
  assign \nz.mem [1569] = \nz.mem_1569_sv2v_reg ;
  assign \nz.mem [1568] = \nz.mem_1568_sv2v_reg ;
  assign \nz.mem [1567] = \nz.mem_1567_sv2v_reg ;
  assign \nz.mem [1566] = \nz.mem_1566_sv2v_reg ;
  assign \nz.mem [1565] = \nz.mem_1565_sv2v_reg ;
  assign \nz.mem [1564] = \nz.mem_1564_sv2v_reg ;
  assign \nz.mem [1563] = \nz.mem_1563_sv2v_reg ;
  assign \nz.mem [1562] = \nz.mem_1562_sv2v_reg ;
  assign \nz.mem [1561] = \nz.mem_1561_sv2v_reg ;
  assign \nz.mem [1560] = \nz.mem_1560_sv2v_reg ;
  assign \nz.mem [1559] = \nz.mem_1559_sv2v_reg ;
  assign \nz.mem [1558] = \nz.mem_1558_sv2v_reg ;
  assign \nz.mem [1557] = \nz.mem_1557_sv2v_reg ;
  assign \nz.mem [1556] = \nz.mem_1556_sv2v_reg ;
  assign \nz.mem [1555] = \nz.mem_1555_sv2v_reg ;
  assign \nz.mem [1554] = \nz.mem_1554_sv2v_reg ;
  assign \nz.mem [1553] = \nz.mem_1553_sv2v_reg ;
  assign \nz.mem [1552] = \nz.mem_1552_sv2v_reg ;
  assign \nz.mem [1551] = \nz.mem_1551_sv2v_reg ;
  assign \nz.mem [1550] = \nz.mem_1550_sv2v_reg ;
  assign \nz.mem [1549] = \nz.mem_1549_sv2v_reg ;
  assign \nz.mem [1548] = \nz.mem_1548_sv2v_reg ;
  assign \nz.mem [1547] = \nz.mem_1547_sv2v_reg ;
  assign \nz.mem [1546] = \nz.mem_1546_sv2v_reg ;
  assign \nz.mem [1545] = \nz.mem_1545_sv2v_reg ;
  assign \nz.mem [1544] = \nz.mem_1544_sv2v_reg ;
  assign \nz.mem [1543] = \nz.mem_1543_sv2v_reg ;
  assign \nz.mem [1542] = \nz.mem_1542_sv2v_reg ;
  assign \nz.mem [1541] = \nz.mem_1541_sv2v_reg ;
  assign \nz.mem [1540] = \nz.mem_1540_sv2v_reg ;
  assign \nz.mem [1539] = \nz.mem_1539_sv2v_reg ;
  assign \nz.mem [1538] = \nz.mem_1538_sv2v_reg ;
  assign \nz.mem [1537] = \nz.mem_1537_sv2v_reg ;
  assign \nz.mem [1536] = \nz.mem_1536_sv2v_reg ;
  assign \nz.mem [1535] = \nz.mem_1535_sv2v_reg ;
  assign \nz.mem [1534] = \nz.mem_1534_sv2v_reg ;
  assign \nz.mem [1533] = \nz.mem_1533_sv2v_reg ;
  assign \nz.mem [1532] = \nz.mem_1532_sv2v_reg ;
  assign \nz.mem [1531] = \nz.mem_1531_sv2v_reg ;
  assign \nz.mem [1530] = \nz.mem_1530_sv2v_reg ;
  assign \nz.mem [1529] = \nz.mem_1529_sv2v_reg ;
  assign \nz.mem [1528] = \nz.mem_1528_sv2v_reg ;
  assign \nz.mem [1527] = \nz.mem_1527_sv2v_reg ;
  assign \nz.mem [1526] = \nz.mem_1526_sv2v_reg ;
  assign \nz.mem [1525] = \nz.mem_1525_sv2v_reg ;
  assign \nz.mem [1524] = \nz.mem_1524_sv2v_reg ;
  assign \nz.mem [1523] = \nz.mem_1523_sv2v_reg ;
  assign \nz.mem [1522] = \nz.mem_1522_sv2v_reg ;
  assign \nz.mem [1521] = \nz.mem_1521_sv2v_reg ;
  assign \nz.mem [1520] = \nz.mem_1520_sv2v_reg ;
  assign \nz.mem [1519] = \nz.mem_1519_sv2v_reg ;
  assign \nz.mem [1518] = \nz.mem_1518_sv2v_reg ;
  assign \nz.mem [1517] = \nz.mem_1517_sv2v_reg ;
  assign \nz.mem [1516] = \nz.mem_1516_sv2v_reg ;
  assign \nz.mem [1515] = \nz.mem_1515_sv2v_reg ;
  assign \nz.mem [1514] = \nz.mem_1514_sv2v_reg ;
  assign \nz.mem [1513] = \nz.mem_1513_sv2v_reg ;
  assign \nz.mem [1512] = \nz.mem_1512_sv2v_reg ;
  assign \nz.mem [1511] = \nz.mem_1511_sv2v_reg ;
  assign \nz.mem [1510] = \nz.mem_1510_sv2v_reg ;
  assign \nz.mem [1509] = \nz.mem_1509_sv2v_reg ;
  assign \nz.mem [1508] = \nz.mem_1508_sv2v_reg ;
  assign \nz.mem [1507] = \nz.mem_1507_sv2v_reg ;
  assign \nz.mem [1506] = \nz.mem_1506_sv2v_reg ;
  assign \nz.mem [1505] = \nz.mem_1505_sv2v_reg ;
  assign \nz.mem [1504] = \nz.mem_1504_sv2v_reg ;
  assign \nz.mem [1503] = \nz.mem_1503_sv2v_reg ;
  assign \nz.mem [1502] = \nz.mem_1502_sv2v_reg ;
  assign \nz.mem [1501] = \nz.mem_1501_sv2v_reg ;
  assign \nz.mem [1500] = \nz.mem_1500_sv2v_reg ;
  assign \nz.mem [1499] = \nz.mem_1499_sv2v_reg ;
  assign \nz.mem [1498] = \nz.mem_1498_sv2v_reg ;
  assign \nz.mem [1497] = \nz.mem_1497_sv2v_reg ;
  assign \nz.mem [1496] = \nz.mem_1496_sv2v_reg ;
  assign \nz.mem [1495] = \nz.mem_1495_sv2v_reg ;
  assign \nz.mem [1494] = \nz.mem_1494_sv2v_reg ;
  assign \nz.mem [1493] = \nz.mem_1493_sv2v_reg ;
  assign \nz.mem [1492] = \nz.mem_1492_sv2v_reg ;
  assign \nz.mem [1491] = \nz.mem_1491_sv2v_reg ;
  assign \nz.mem [1490] = \nz.mem_1490_sv2v_reg ;
  assign \nz.mem [1489] = \nz.mem_1489_sv2v_reg ;
  assign \nz.mem [1488] = \nz.mem_1488_sv2v_reg ;
  assign \nz.mem [1487] = \nz.mem_1487_sv2v_reg ;
  assign \nz.mem [1486] = \nz.mem_1486_sv2v_reg ;
  assign \nz.mem [1485] = \nz.mem_1485_sv2v_reg ;
  assign \nz.mem [1484] = \nz.mem_1484_sv2v_reg ;
  assign \nz.mem [1483] = \nz.mem_1483_sv2v_reg ;
  assign \nz.mem [1482] = \nz.mem_1482_sv2v_reg ;
  assign \nz.mem [1481] = \nz.mem_1481_sv2v_reg ;
  assign \nz.mem [1480] = \nz.mem_1480_sv2v_reg ;
  assign \nz.mem [1479] = \nz.mem_1479_sv2v_reg ;
  assign \nz.mem [1478] = \nz.mem_1478_sv2v_reg ;
  assign \nz.mem [1477] = \nz.mem_1477_sv2v_reg ;
  assign \nz.mem [1476] = \nz.mem_1476_sv2v_reg ;
  assign \nz.mem [1475] = \nz.mem_1475_sv2v_reg ;
  assign \nz.mem [1474] = \nz.mem_1474_sv2v_reg ;
  assign \nz.mem [1473] = \nz.mem_1473_sv2v_reg ;
  assign \nz.mem [1472] = \nz.mem_1472_sv2v_reg ;
  assign \nz.mem [1471] = \nz.mem_1471_sv2v_reg ;
  assign \nz.mem [1470] = \nz.mem_1470_sv2v_reg ;
  assign \nz.mem [1469] = \nz.mem_1469_sv2v_reg ;
  assign \nz.mem [1468] = \nz.mem_1468_sv2v_reg ;
  assign \nz.mem [1467] = \nz.mem_1467_sv2v_reg ;
  assign \nz.mem [1466] = \nz.mem_1466_sv2v_reg ;
  assign \nz.mem [1465] = \nz.mem_1465_sv2v_reg ;
  assign \nz.mem [1464] = \nz.mem_1464_sv2v_reg ;
  assign \nz.mem [1463] = \nz.mem_1463_sv2v_reg ;
  assign \nz.mem [1462] = \nz.mem_1462_sv2v_reg ;
  assign \nz.mem [1461] = \nz.mem_1461_sv2v_reg ;
  assign \nz.mem [1460] = \nz.mem_1460_sv2v_reg ;
  assign \nz.mem [1459] = \nz.mem_1459_sv2v_reg ;
  assign \nz.mem [1458] = \nz.mem_1458_sv2v_reg ;
  assign \nz.mem [1457] = \nz.mem_1457_sv2v_reg ;
  assign \nz.mem [1456] = \nz.mem_1456_sv2v_reg ;
  assign \nz.mem [1455] = \nz.mem_1455_sv2v_reg ;
  assign \nz.mem [1454] = \nz.mem_1454_sv2v_reg ;
  assign \nz.mem [1453] = \nz.mem_1453_sv2v_reg ;
  assign \nz.mem [1452] = \nz.mem_1452_sv2v_reg ;
  assign \nz.mem [1451] = \nz.mem_1451_sv2v_reg ;
  assign \nz.mem [1450] = \nz.mem_1450_sv2v_reg ;
  assign \nz.mem [1449] = \nz.mem_1449_sv2v_reg ;
  assign \nz.mem [1448] = \nz.mem_1448_sv2v_reg ;
  assign \nz.mem [1447] = \nz.mem_1447_sv2v_reg ;
  assign \nz.mem [1446] = \nz.mem_1446_sv2v_reg ;
  assign \nz.mem [1445] = \nz.mem_1445_sv2v_reg ;
  assign \nz.mem [1444] = \nz.mem_1444_sv2v_reg ;
  assign \nz.mem [1443] = \nz.mem_1443_sv2v_reg ;
  assign \nz.mem [1442] = \nz.mem_1442_sv2v_reg ;
  assign \nz.mem [1441] = \nz.mem_1441_sv2v_reg ;
  assign \nz.mem [1440] = \nz.mem_1440_sv2v_reg ;
  assign \nz.mem [1439] = \nz.mem_1439_sv2v_reg ;
  assign \nz.mem [1438] = \nz.mem_1438_sv2v_reg ;
  assign \nz.mem [1437] = \nz.mem_1437_sv2v_reg ;
  assign \nz.mem [1436] = \nz.mem_1436_sv2v_reg ;
  assign \nz.mem [1435] = \nz.mem_1435_sv2v_reg ;
  assign \nz.mem [1434] = \nz.mem_1434_sv2v_reg ;
  assign \nz.mem [1433] = \nz.mem_1433_sv2v_reg ;
  assign \nz.mem [1432] = \nz.mem_1432_sv2v_reg ;
  assign \nz.mem [1431] = \nz.mem_1431_sv2v_reg ;
  assign \nz.mem [1430] = \nz.mem_1430_sv2v_reg ;
  assign \nz.mem [1429] = \nz.mem_1429_sv2v_reg ;
  assign \nz.mem [1428] = \nz.mem_1428_sv2v_reg ;
  assign \nz.mem [1427] = \nz.mem_1427_sv2v_reg ;
  assign \nz.mem [1426] = \nz.mem_1426_sv2v_reg ;
  assign \nz.mem [1425] = \nz.mem_1425_sv2v_reg ;
  assign \nz.mem [1424] = \nz.mem_1424_sv2v_reg ;
  assign \nz.mem [1423] = \nz.mem_1423_sv2v_reg ;
  assign \nz.mem [1422] = \nz.mem_1422_sv2v_reg ;
  assign \nz.mem [1421] = \nz.mem_1421_sv2v_reg ;
  assign \nz.mem [1420] = \nz.mem_1420_sv2v_reg ;
  assign \nz.mem [1419] = \nz.mem_1419_sv2v_reg ;
  assign \nz.mem [1418] = \nz.mem_1418_sv2v_reg ;
  assign \nz.mem [1417] = \nz.mem_1417_sv2v_reg ;
  assign \nz.mem [1416] = \nz.mem_1416_sv2v_reg ;
  assign \nz.mem [1415] = \nz.mem_1415_sv2v_reg ;
  assign \nz.mem [1414] = \nz.mem_1414_sv2v_reg ;
  assign \nz.mem [1413] = \nz.mem_1413_sv2v_reg ;
  assign \nz.mem [1412] = \nz.mem_1412_sv2v_reg ;
  assign \nz.mem [1411] = \nz.mem_1411_sv2v_reg ;
  assign \nz.mem [1410] = \nz.mem_1410_sv2v_reg ;
  assign \nz.mem [1409] = \nz.mem_1409_sv2v_reg ;
  assign \nz.mem [1408] = \nz.mem_1408_sv2v_reg ;
  assign \nz.mem [1407] = \nz.mem_1407_sv2v_reg ;
  assign \nz.mem [1406] = \nz.mem_1406_sv2v_reg ;
  assign \nz.mem [1405] = \nz.mem_1405_sv2v_reg ;
  assign \nz.mem [1404] = \nz.mem_1404_sv2v_reg ;
  assign \nz.mem [1403] = \nz.mem_1403_sv2v_reg ;
  assign \nz.mem [1402] = \nz.mem_1402_sv2v_reg ;
  assign \nz.mem [1401] = \nz.mem_1401_sv2v_reg ;
  assign \nz.mem [1400] = \nz.mem_1400_sv2v_reg ;
  assign \nz.mem [1399] = \nz.mem_1399_sv2v_reg ;
  assign \nz.mem [1398] = \nz.mem_1398_sv2v_reg ;
  assign \nz.mem [1397] = \nz.mem_1397_sv2v_reg ;
  assign \nz.mem [1396] = \nz.mem_1396_sv2v_reg ;
  assign \nz.mem [1395] = \nz.mem_1395_sv2v_reg ;
  assign \nz.mem [1394] = \nz.mem_1394_sv2v_reg ;
  assign \nz.mem [1393] = \nz.mem_1393_sv2v_reg ;
  assign \nz.mem [1392] = \nz.mem_1392_sv2v_reg ;
  assign \nz.mem [1391] = \nz.mem_1391_sv2v_reg ;
  assign \nz.mem [1390] = \nz.mem_1390_sv2v_reg ;
  assign \nz.mem [1389] = \nz.mem_1389_sv2v_reg ;
  assign \nz.mem [1388] = \nz.mem_1388_sv2v_reg ;
  assign \nz.mem [1387] = \nz.mem_1387_sv2v_reg ;
  assign \nz.mem [1386] = \nz.mem_1386_sv2v_reg ;
  assign \nz.mem [1385] = \nz.mem_1385_sv2v_reg ;
  assign \nz.mem [1384] = \nz.mem_1384_sv2v_reg ;
  assign \nz.mem [1383] = \nz.mem_1383_sv2v_reg ;
  assign \nz.mem [1382] = \nz.mem_1382_sv2v_reg ;
  assign \nz.mem [1381] = \nz.mem_1381_sv2v_reg ;
  assign \nz.mem [1380] = \nz.mem_1380_sv2v_reg ;
  assign \nz.mem [1379] = \nz.mem_1379_sv2v_reg ;
  assign \nz.mem [1378] = \nz.mem_1378_sv2v_reg ;
  assign \nz.mem [1377] = \nz.mem_1377_sv2v_reg ;
  assign \nz.mem [1376] = \nz.mem_1376_sv2v_reg ;
  assign \nz.mem [1375] = \nz.mem_1375_sv2v_reg ;
  assign \nz.mem [1374] = \nz.mem_1374_sv2v_reg ;
  assign \nz.mem [1373] = \nz.mem_1373_sv2v_reg ;
  assign \nz.mem [1372] = \nz.mem_1372_sv2v_reg ;
  assign \nz.mem [1371] = \nz.mem_1371_sv2v_reg ;
  assign \nz.mem [1370] = \nz.mem_1370_sv2v_reg ;
  assign \nz.mem [1369] = \nz.mem_1369_sv2v_reg ;
  assign \nz.mem [1368] = \nz.mem_1368_sv2v_reg ;
  assign \nz.mem [1367] = \nz.mem_1367_sv2v_reg ;
  assign \nz.mem [1366] = \nz.mem_1366_sv2v_reg ;
  assign \nz.mem [1365] = \nz.mem_1365_sv2v_reg ;
  assign \nz.mem [1364] = \nz.mem_1364_sv2v_reg ;
  assign \nz.mem [1363] = \nz.mem_1363_sv2v_reg ;
  assign \nz.mem [1362] = \nz.mem_1362_sv2v_reg ;
  assign \nz.mem [1361] = \nz.mem_1361_sv2v_reg ;
  assign \nz.mem [1360] = \nz.mem_1360_sv2v_reg ;
  assign \nz.mem [1359] = \nz.mem_1359_sv2v_reg ;
  assign \nz.mem [1358] = \nz.mem_1358_sv2v_reg ;
  assign \nz.mem [1357] = \nz.mem_1357_sv2v_reg ;
  assign \nz.mem [1356] = \nz.mem_1356_sv2v_reg ;
  assign \nz.mem [1355] = \nz.mem_1355_sv2v_reg ;
  assign \nz.mem [1354] = \nz.mem_1354_sv2v_reg ;
  assign \nz.mem [1353] = \nz.mem_1353_sv2v_reg ;
  assign \nz.mem [1352] = \nz.mem_1352_sv2v_reg ;
  assign \nz.mem [1351] = \nz.mem_1351_sv2v_reg ;
  assign \nz.mem [1350] = \nz.mem_1350_sv2v_reg ;
  assign \nz.mem [1349] = \nz.mem_1349_sv2v_reg ;
  assign \nz.mem [1348] = \nz.mem_1348_sv2v_reg ;
  assign \nz.mem [1347] = \nz.mem_1347_sv2v_reg ;
  assign \nz.mem [1346] = \nz.mem_1346_sv2v_reg ;
  assign \nz.mem [1345] = \nz.mem_1345_sv2v_reg ;
  assign \nz.mem [1344] = \nz.mem_1344_sv2v_reg ;
  assign \nz.mem [1343] = \nz.mem_1343_sv2v_reg ;
  assign \nz.mem [1342] = \nz.mem_1342_sv2v_reg ;
  assign \nz.mem [1341] = \nz.mem_1341_sv2v_reg ;
  assign \nz.mem [1340] = \nz.mem_1340_sv2v_reg ;
  assign \nz.mem [1339] = \nz.mem_1339_sv2v_reg ;
  assign \nz.mem [1338] = \nz.mem_1338_sv2v_reg ;
  assign \nz.mem [1337] = \nz.mem_1337_sv2v_reg ;
  assign \nz.mem [1336] = \nz.mem_1336_sv2v_reg ;
  assign \nz.mem [1335] = \nz.mem_1335_sv2v_reg ;
  assign \nz.mem [1334] = \nz.mem_1334_sv2v_reg ;
  assign \nz.mem [1333] = \nz.mem_1333_sv2v_reg ;
  assign \nz.mem [1332] = \nz.mem_1332_sv2v_reg ;
  assign \nz.mem [1331] = \nz.mem_1331_sv2v_reg ;
  assign \nz.mem [1330] = \nz.mem_1330_sv2v_reg ;
  assign \nz.mem [1329] = \nz.mem_1329_sv2v_reg ;
  assign \nz.mem [1328] = \nz.mem_1328_sv2v_reg ;
  assign \nz.mem [1327] = \nz.mem_1327_sv2v_reg ;
  assign \nz.mem [1326] = \nz.mem_1326_sv2v_reg ;
  assign \nz.mem [1325] = \nz.mem_1325_sv2v_reg ;
  assign \nz.mem [1324] = \nz.mem_1324_sv2v_reg ;
  assign \nz.mem [1323] = \nz.mem_1323_sv2v_reg ;
  assign \nz.mem [1322] = \nz.mem_1322_sv2v_reg ;
  assign \nz.mem [1321] = \nz.mem_1321_sv2v_reg ;
  assign \nz.mem [1320] = \nz.mem_1320_sv2v_reg ;
  assign \nz.mem [1319] = \nz.mem_1319_sv2v_reg ;
  assign \nz.mem [1318] = \nz.mem_1318_sv2v_reg ;
  assign \nz.mem [1317] = \nz.mem_1317_sv2v_reg ;
  assign \nz.mem [1316] = \nz.mem_1316_sv2v_reg ;
  assign \nz.mem [1315] = \nz.mem_1315_sv2v_reg ;
  assign \nz.mem [1314] = \nz.mem_1314_sv2v_reg ;
  assign \nz.mem [1313] = \nz.mem_1313_sv2v_reg ;
  assign \nz.mem [1312] = \nz.mem_1312_sv2v_reg ;
  assign \nz.mem [1311] = \nz.mem_1311_sv2v_reg ;
  assign \nz.mem [1310] = \nz.mem_1310_sv2v_reg ;
  assign \nz.mem [1309] = \nz.mem_1309_sv2v_reg ;
  assign \nz.mem [1308] = \nz.mem_1308_sv2v_reg ;
  assign \nz.mem [1307] = \nz.mem_1307_sv2v_reg ;
  assign \nz.mem [1306] = \nz.mem_1306_sv2v_reg ;
  assign \nz.mem [1305] = \nz.mem_1305_sv2v_reg ;
  assign \nz.mem [1304] = \nz.mem_1304_sv2v_reg ;
  assign \nz.mem [1303] = \nz.mem_1303_sv2v_reg ;
  assign \nz.mem [1302] = \nz.mem_1302_sv2v_reg ;
  assign \nz.mem [1301] = \nz.mem_1301_sv2v_reg ;
  assign \nz.mem [1300] = \nz.mem_1300_sv2v_reg ;
  assign \nz.mem [1299] = \nz.mem_1299_sv2v_reg ;
  assign \nz.mem [1298] = \nz.mem_1298_sv2v_reg ;
  assign \nz.mem [1297] = \nz.mem_1297_sv2v_reg ;
  assign \nz.mem [1296] = \nz.mem_1296_sv2v_reg ;
  assign \nz.mem [1295] = \nz.mem_1295_sv2v_reg ;
  assign \nz.mem [1294] = \nz.mem_1294_sv2v_reg ;
  assign \nz.mem [1293] = \nz.mem_1293_sv2v_reg ;
  assign \nz.mem [1292] = \nz.mem_1292_sv2v_reg ;
  assign \nz.mem [1291] = \nz.mem_1291_sv2v_reg ;
  assign \nz.mem [1290] = \nz.mem_1290_sv2v_reg ;
  assign \nz.mem [1289] = \nz.mem_1289_sv2v_reg ;
  assign \nz.mem [1288] = \nz.mem_1288_sv2v_reg ;
  assign \nz.mem [1287] = \nz.mem_1287_sv2v_reg ;
  assign \nz.mem [1286] = \nz.mem_1286_sv2v_reg ;
  assign \nz.mem [1285] = \nz.mem_1285_sv2v_reg ;
  assign \nz.mem [1284] = \nz.mem_1284_sv2v_reg ;
  assign \nz.mem [1283] = \nz.mem_1283_sv2v_reg ;
  assign \nz.mem [1282] = \nz.mem_1282_sv2v_reg ;
  assign \nz.mem [1281] = \nz.mem_1281_sv2v_reg ;
  assign \nz.mem [1280] = \nz.mem_1280_sv2v_reg ;
  assign \nz.mem [1279] = \nz.mem_1279_sv2v_reg ;
  assign \nz.mem [1278] = \nz.mem_1278_sv2v_reg ;
  assign \nz.mem [1277] = \nz.mem_1277_sv2v_reg ;
  assign \nz.mem [1276] = \nz.mem_1276_sv2v_reg ;
  assign \nz.mem [1275] = \nz.mem_1275_sv2v_reg ;
  assign \nz.mem [1274] = \nz.mem_1274_sv2v_reg ;
  assign \nz.mem [1273] = \nz.mem_1273_sv2v_reg ;
  assign \nz.mem [1272] = \nz.mem_1272_sv2v_reg ;
  assign \nz.mem [1271] = \nz.mem_1271_sv2v_reg ;
  assign \nz.mem [1270] = \nz.mem_1270_sv2v_reg ;
  assign \nz.mem [1269] = \nz.mem_1269_sv2v_reg ;
  assign \nz.mem [1268] = \nz.mem_1268_sv2v_reg ;
  assign \nz.mem [1267] = \nz.mem_1267_sv2v_reg ;
  assign \nz.mem [1266] = \nz.mem_1266_sv2v_reg ;
  assign \nz.mem [1265] = \nz.mem_1265_sv2v_reg ;
  assign \nz.mem [1264] = \nz.mem_1264_sv2v_reg ;
  assign \nz.mem [1263] = \nz.mem_1263_sv2v_reg ;
  assign \nz.mem [1262] = \nz.mem_1262_sv2v_reg ;
  assign \nz.mem [1261] = \nz.mem_1261_sv2v_reg ;
  assign \nz.mem [1260] = \nz.mem_1260_sv2v_reg ;
  assign \nz.mem [1259] = \nz.mem_1259_sv2v_reg ;
  assign \nz.mem [1258] = \nz.mem_1258_sv2v_reg ;
  assign \nz.mem [1257] = \nz.mem_1257_sv2v_reg ;
  assign \nz.mem [1256] = \nz.mem_1256_sv2v_reg ;
  assign \nz.mem [1255] = \nz.mem_1255_sv2v_reg ;
  assign \nz.mem [1254] = \nz.mem_1254_sv2v_reg ;
  assign \nz.mem [1253] = \nz.mem_1253_sv2v_reg ;
  assign \nz.mem [1252] = \nz.mem_1252_sv2v_reg ;
  assign \nz.mem [1251] = \nz.mem_1251_sv2v_reg ;
  assign \nz.mem [1250] = \nz.mem_1250_sv2v_reg ;
  assign \nz.mem [1249] = \nz.mem_1249_sv2v_reg ;
  assign \nz.mem [1248] = \nz.mem_1248_sv2v_reg ;
  assign \nz.mem [1247] = \nz.mem_1247_sv2v_reg ;
  assign \nz.mem [1246] = \nz.mem_1246_sv2v_reg ;
  assign \nz.mem [1245] = \nz.mem_1245_sv2v_reg ;
  assign \nz.mem [1244] = \nz.mem_1244_sv2v_reg ;
  assign \nz.mem [1243] = \nz.mem_1243_sv2v_reg ;
  assign \nz.mem [1242] = \nz.mem_1242_sv2v_reg ;
  assign \nz.mem [1241] = \nz.mem_1241_sv2v_reg ;
  assign \nz.mem [1240] = \nz.mem_1240_sv2v_reg ;
  assign \nz.mem [1239] = \nz.mem_1239_sv2v_reg ;
  assign \nz.mem [1238] = \nz.mem_1238_sv2v_reg ;
  assign \nz.mem [1237] = \nz.mem_1237_sv2v_reg ;
  assign \nz.mem [1236] = \nz.mem_1236_sv2v_reg ;
  assign \nz.mem [1235] = \nz.mem_1235_sv2v_reg ;
  assign \nz.mem [1234] = \nz.mem_1234_sv2v_reg ;
  assign \nz.mem [1233] = \nz.mem_1233_sv2v_reg ;
  assign \nz.mem [1232] = \nz.mem_1232_sv2v_reg ;
  assign \nz.mem [1231] = \nz.mem_1231_sv2v_reg ;
  assign \nz.mem [1230] = \nz.mem_1230_sv2v_reg ;
  assign \nz.mem [1229] = \nz.mem_1229_sv2v_reg ;
  assign \nz.mem [1228] = \nz.mem_1228_sv2v_reg ;
  assign \nz.mem [1227] = \nz.mem_1227_sv2v_reg ;
  assign \nz.mem [1226] = \nz.mem_1226_sv2v_reg ;
  assign \nz.mem [1225] = \nz.mem_1225_sv2v_reg ;
  assign \nz.mem [1224] = \nz.mem_1224_sv2v_reg ;
  assign \nz.mem [1223] = \nz.mem_1223_sv2v_reg ;
  assign \nz.mem [1222] = \nz.mem_1222_sv2v_reg ;
  assign \nz.mem [1221] = \nz.mem_1221_sv2v_reg ;
  assign \nz.mem [1220] = \nz.mem_1220_sv2v_reg ;
  assign \nz.mem [1219] = \nz.mem_1219_sv2v_reg ;
  assign \nz.mem [1218] = \nz.mem_1218_sv2v_reg ;
  assign \nz.mem [1217] = \nz.mem_1217_sv2v_reg ;
  assign \nz.mem [1216] = \nz.mem_1216_sv2v_reg ;
  assign \nz.mem [1215] = \nz.mem_1215_sv2v_reg ;
  assign \nz.mem [1214] = \nz.mem_1214_sv2v_reg ;
  assign \nz.mem [1213] = \nz.mem_1213_sv2v_reg ;
  assign \nz.mem [1212] = \nz.mem_1212_sv2v_reg ;
  assign \nz.mem [1211] = \nz.mem_1211_sv2v_reg ;
  assign \nz.mem [1210] = \nz.mem_1210_sv2v_reg ;
  assign \nz.mem [1209] = \nz.mem_1209_sv2v_reg ;
  assign \nz.mem [1208] = \nz.mem_1208_sv2v_reg ;
  assign \nz.mem [1207] = \nz.mem_1207_sv2v_reg ;
  assign \nz.mem [1206] = \nz.mem_1206_sv2v_reg ;
  assign \nz.mem [1205] = \nz.mem_1205_sv2v_reg ;
  assign \nz.mem [1204] = \nz.mem_1204_sv2v_reg ;
  assign \nz.mem [1203] = \nz.mem_1203_sv2v_reg ;
  assign \nz.mem [1202] = \nz.mem_1202_sv2v_reg ;
  assign \nz.mem [1201] = \nz.mem_1201_sv2v_reg ;
  assign \nz.mem [1200] = \nz.mem_1200_sv2v_reg ;
  assign \nz.mem [1199] = \nz.mem_1199_sv2v_reg ;
  assign \nz.mem [1198] = \nz.mem_1198_sv2v_reg ;
  assign \nz.mem [1197] = \nz.mem_1197_sv2v_reg ;
  assign \nz.mem [1196] = \nz.mem_1196_sv2v_reg ;
  assign \nz.mem [1195] = \nz.mem_1195_sv2v_reg ;
  assign \nz.mem [1194] = \nz.mem_1194_sv2v_reg ;
  assign \nz.mem [1193] = \nz.mem_1193_sv2v_reg ;
  assign \nz.mem [1192] = \nz.mem_1192_sv2v_reg ;
  assign \nz.mem [1191] = \nz.mem_1191_sv2v_reg ;
  assign \nz.mem [1190] = \nz.mem_1190_sv2v_reg ;
  assign \nz.mem [1189] = \nz.mem_1189_sv2v_reg ;
  assign \nz.mem [1188] = \nz.mem_1188_sv2v_reg ;
  assign \nz.mem [1187] = \nz.mem_1187_sv2v_reg ;
  assign \nz.mem [1186] = \nz.mem_1186_sv2v_reg ;
  assign \nz.mem [1185] = \nz.mem_1185_sv2v_reg ;
  assign \nz.mem [1184] = \nz.mem_1184_sv2v_reg ;
  assign \nz.mem [1183] = \nz.mem_1183_sv2v_reg ;
  assign \nz.mem [1182] = \nz.mem_1182_sv2v_reg ;
  assign \nz.mem [1181] = \nz.mem_1181_sv2v_reg ;
  assign \nz.mem [1180] = \nz.mem_1180_sv2v_reg ;
  assign \nz.mem [1179] = \nz.mem_1179_sv2v_reg ;
  assign \nz.mem [1178] = \nz.mem_1178_sv2v_reg ;
  assign \nz.mem [1177] = \nz.mem_1177_sv2v_reg ;
  assign \nz.mem [1176] = \nz.mem_1176_sv2v_reg ;
  assign \nz.mem [1175] = \nz.mem_1175_sv2v_reg ;
  assign \nz.mem [1174] = \nz.mem_1174_sv2v_reg ;
  assign \nz.mem [1173] = \nz.mem_1173_sv2v_reg ;
  assign \nz.mem [1172] = \nz.mem_1172_sv2v_reg ;
  assign \nz.mem [1171] = \nz.mem_1171_sv2v_reg ;
  assign \nz.mem [1170] = \nz.mem_1170_sv2v_reg ;
  assign \nz.mem [1169] = \nz.mem_1169_sv2v_reg ;
  assign \nz.mem [1168] = \nz.mem_1168_sv2v_reg ;
  assign \nz.mem [1167] = \nz.mem_1167_sv2v_reg ;
  assign \nz.mem [1166] = \nz.mem_1166_sv2v_reg ;
  assign \nz.mem [1165] = \nz.mem_1165_sv2v_reg ;
  assign \nz.mem [1164] = \nz.mem_1164_sv2v_reg ;
  assign \nz.mem [1163] = \nz.mem_1163_sv2v_reg ;
  assign \nz.mem [1162] = \nz.mem_1162_sv2v_reg ;
  assign \nz.mem [1161] = \nz.mem_1161_sv2v_reg ;
  assign \nz.mem [1160] = \nz.mem_1160_sv2v_reg ;
  assign \nz.mem [1159] = \nz.mem_1159_sv2v_reg ;
  assign \nz.mem [1158] = \nz.mem_1158_sv2v_reg ;
  assign \nz.mem [1157] = \nz.mem_1157_sv2v_reg ;
  assign \nz.mem [1156] = \nz.mem_1156_sv2v_reg ;
  assign \nz.mem [1155] = \nz.mem_1155_sv2v_reg ;
  assign \nz.mem [1154] = \nz.mem_1154_sv2v_reg ;
  assign \nz.mem [1153] = \nz.mem_1153_sv2v_reg ;
  assign \nz.mem [1152] = \nz.mem_1152_sv2v_reg ;
  assign \nz.mem [1151] = \nz.mem_1151_sv2v_reg ;
  assign \nz.mem [1150] = \nz.mem_1150_sv2v_reg ;
  assign \nz.mem [1149] = \nz.mem_1149_sv2v_reg ;
  assign \nz.mem [1148] = \nz.mem_1148_sv2v_reg ;
  assign \nz.mem [1147] = \nz.mem_1147_sv2v_reg ;
  assign \nz.mem [1146] = \nz.mem_1146_sv2v_reg ;
  assign \nz.mem [1145] = \nz.mem_1145_sv2v_reg ;
  assign \nz.mem [1144] = \nz.mem_1144_sv2v_reg ;
  assign \nz.mem [1143] = \nz.mem_1143_sv2v_reg ;
  assign \nz.mem [1142] = \nz.mem_1142_sv2v_reg ;
  assign \nz.mem [1141] = \nz.mem_1141_sv2v_reg ;
  assign \nz.mem [1140] = \nz.mem_1140_sv2v_reg ;
  assign \nz.mem [1139] = \nz.mem_1139_sv2v_reg ;
  assign \nz.mem [1138] = \nz.mem_1138_sv2v_reg ;
  assign \nz.mem [1137] = \nz.mem_1137_sv2v_reg ;
  assign \nz.mem [1136] = \nz.mem_1136_sv2v_reg ;
  assign \nz.mem [1135] = \nz.mem_1135_sv2v_reg ;
  assign \nz.mem [1134] = \nz.mem_1134_sv2v_reg ;
  assign \nz.mem [1133] = \nz.mem_1133_sv2v_reg ;
  assign \nz.mem [1132] = \nz.mem_1132_sv2v_reg ;
  assign \nz.mem [1131] = \nz.mem_1131_sv2v_reg ;
  assign \nz.mem [1130] = \nz.mem_1130_sv2v_reg ;
  assign \nz.mem [1129] = \nz.mem_1129_sv2v_reg ;
  assign \nz.mem [1128] = \nz.mem_1128_sv2v_reg ;
  assign \nz.mem [1127] = \nz.mem_1127_sv2v_reg ;
  assign \nz.mem [1126] = \nz.mem_1126_sv2v_reg ;
  assign \nz.mem [1125] = \nz.mem_1125_sv2v_reg ;
  assign \nz.mem [1124] = \nz.mem_1124_sv2v_reg ;
  assign \nz.mem [1123] = \nz.mem_1123_sv2v_reg ;
  assign \nz.mem [1122] = \nz.mem_1122_sv2v_reg ;
  assign \nz.mem [1121] = \nz.mem_1121_sv2v_reg ;
  assign \nz.mem [1120] = \nz.mem_1120_sv2v_reg ;
  assign \nz.mem [1119] = \nz.mem_1119_sv2v_reg ;
  assign \nz.mem [1118] = \nz.mem_1118_sv2v_reg ;
  assign \nz.mem [1117] = \nz.mem_1117_sv2v_reg ;
  assign \nz.mem [1116] = \nz.mem_1116_sv2v_reg ;
  assign \nz.mem [1115] = \nz.mem_1115_sv2v_reg ;
  assign \nz.mem [1114] = \nz.mem_1114_sv2v_reg ;
  assign \nz.mem [1113] = \nz.mem_1113_sv2v_reg ;
  assign \nz.mem [1112] = \nz.mem_1112_sv2v_reg ;
  assign \nz.mem [1111] = \nz.mem_1111_sv2v_reg ;
  assign \nz.mem [1110] = \nz.mem_1110_sv2v_reg ;
  assign \nz.mem [1109] = \nz.mem_1109_sv2v_reg ;
  assign \nz.mem [1108] = \nz.mem_1108_sv2v_reg ;
  assign \nz.mem [1107] = \nz.mem_1107_sv2v_reg ;
  assign \nz.mem [1106] = \nz.mem_1106_sv2v_reg ;
  assign \nz.mem [1105] = \nz.mem_1105_sv2v_reg ;
  assign \nz.mem [1104] = \nz.mem_1104_sv2v_reg ;
  assign \nz.mem [1103] = \nz.mem_1103_sv2v_reg ;
  assign \nz.mem [1102] = \nz.mem_1102_sv2v_reg ;
  assign \nz.mem [1101] = \nz.mem_1101_sv2v_reg ;
  assign \nz.mem [1100] = \nz.mem_1100_sv2v_reg ;
  assign \nz.mem [1099] = \nz.mem_1099_sv2v_reg ;
  assign \nz.mem [1098] = \nz.mem_1098_sv2v_reg ;
  assign \nz.mem [1097] = \nz.mem_1097_sv2v_reg ;
  assign \nz.mem [1096] = \nz.mem_1096_sv2v_reg ;
  assign \nz.mem [1095] = \nz.mem_1095_sv2v_reg ;
  assign \nz.mem [1094] = \nz.mem_1094_sv2v_reg ;
  assign \nz.mem [1093] = \nz.mem_1093_sv2v_reg ;
  assign \nz.mem [1092] = \nz.mem_1092_sv2v_reg ;
  assign \nz.mem [1091] = \nz.mem_1091_sv2v_reg ;
  assign \nz.mem [1090] = \nz.mem_1090_sv2v_reg ;
  assign \nz.mem [1089] = \nz.mem_1089_sv2v_reg ;
  assign \nz.mem [1088] = \nz.mem_1088_sv2v_reg ;
  assign \nz.mem [1087] = \nz.mem_1087_sv2v_reg ;
  assign \nz.mem [1086] = \nz.mem_1086_sv2v_reg ;
  assign \nz.mem [1085] = \nz.mem_1085_sv2v_reg ;
  assign \nz.mem [1084] = \nz.mem_1084_sv2v_reg ;
  assign \nz.mem [1083] = \nz.mem_1083_sv2v_reg ;
  assign \nz.mem [1082] = \nz.mem_1082_sv2v_reg ;
  assign \nz.mem [1081] = \nz.mem_1081_sv2v_reg ;
  assign \nz.mem [1080] = \nz.mem_1080_sv2v_reg ;
  assign \nz.mem [1079] = \nz.mem_1079_sv2v_reg ;
  assign \nz.mem [1078] = \nz.mem_1078_sv2v_reg ;
  assign \nz.mem [1077] = \nz.mem_1077_sv2v_reg ;
  assign \nz.mem [1076] = \nz.mem_1076_sv2v_reg ;
  assign \nz.mem [1075] = \nz.mem_1075_sv2v_reg ;
  assign \nz.mem [1074] = \nz.mem_1074_sv2v_reg ;
  assign \nz.mem [1073] = \nz.mem_1073_sv2v_reg ;
  assign \nz.mem [1072] = \nz.mem_1072_sv2v_reg ;
  assign \nz.mem [1071] = \nz.mem_1071_sv2v_reg ;
  assign \nz.mem [1070] = \nz.mem_1070_sv2v_reg ;
  assign \nz.mem [1069] = \nz.mem_1069_sv2v_reg ;
  assign \nz.mem [1068] = \nz.mem_1068_sv2v_reg ;
  assign \nz.mem [1067] = \nz.mem_1067_sv2v_reg ;
  assign \nz.mem [1066] = \nz.mem_1066_sv2v_reg ;
  assign \nz.mem [1065] = \nz.mem_1065_sv2v_reg ;
  assign \nz.mem [1064] = \nz.mem_1064_sv2v_reg ;
  assign \nz.mem [1063] = \nz.mem_1063_sv2v_reg ;
  assign \nz.mem [1062] = \nz.mem_1062_sv2v_reg ;
  assign \nz.mem [1061] = \nz.mem_1061_sv2v_reg ;
  assign \nz.mem [1060] = \nz.mem_1060_sv2v_reg ;
  assign \nz.mem [1059] = \nz.mem_1059_sv2v_reg ;
  assign \nz.mem [1058] = \nz.mem_1058_sv2v_reg ;
  assign \nz.mem [1057] = \nz.mem_1057_sv2v_reg ;
  assign \nz.mem [1056] = \nz.mem_1056_sv2v_reg ;
  assign \nz.mem [1055] = \nz.mem_1055_sv2v_reg ;
  assign \nz.mem [1054] = \nz.mem_1054_sv2v_reg ;
  assign \nz.mem [1053] = \nz.mem_1053_sv2v_reg ;
  assign \nz.mem [1052] = \nz.mem_1052_sv2v_reg ;
  assign \nz.mem [1051] = \nz.mem_1051_sv2v_reg ;
  assign \nz.mem [1050] = \nz.mem_1050_sv2v_reg ;
  assign \nz.mem [1049] = \nz.mem_1049_sv2v_reg ;
  assign \nz.mem [1048] = \nz.mem_1048_sv2v_reg ;
  assign \nz.mem [1047] = \nz.mem_1047_sv2v_reg ;
  assign \nz.mem [1046] = \nz.mem_1046_sv2v_reg ;
  assign \nz.mem [1045] = \nz.mem_1045_sv2v_reg ;
  assign \nz.mem [1044] = \nz.mem_1044_sv2v_reg ;
  assign \nz.mem [1043] = \nz.mem_1043_sv2v_reg ;
  assign \nz.mem [1042] = \nz.mem_1042_sv2v_reg ;
  assign \nz.mem [1041] = \nz.mem_1041_sv2v_reg ;
  assign \nz.mem [1040] = \nz.mem_1040_sv2v_reg ;
  assign \nz.mem [1039] = \nz.mem_1039_sv2v_reg ;
  assign \nz.mem [1038] = \nz.mem_1038_sv2v_reg ;
  assign \nz.mem [1037] = \nz.mem_1037_sv2v_reg ;
  assign \nz.mem [1036] = \nz.mem_1036_sv2v_reg ;
  assign \nz.mem [1035] = \nz.mem_1035_sv2v_reg ;
  assign \nz.mem [1034] = \nz.mem_1034_sv2v_reg ;
  assign \nz.mem [1033] = \nz.mem_1033_sv2v_reg ;
  assign \nz.mem [1032] = \nz.mem_1032_sv2v_reg ;
  assign \nz.mem [1031] = \nz.mem_1031_sv2v_reg ;
  assign \nz.mem [1030] = \nz.mem_1030_sv2v_reg ;
  assign \nz.mem [1029] = \nz.mem_1029_sv2v_reg ;
  assign \nz.mem [1028] = \nz.mem_1028_sv2v_reg ;
  assign \nz.mem [1027] = \nz.mem_1027_sv2v_reg ;
  assign \nz.mem [1026] = \nz.mem_1026_sv2v_reg ;
  assign \nz.mem [1025] = \nz.mem_1025_sv2v_reg ;
  assign \nz.mem [1024] = \nz.mem_1024_sv2v_reg ;
  assign \nz.mem [1023] = \nz.mem_1023_sv2v_reg ;
  assign \nz.mem [1022] = \nz.mem_1022_sv2v_reg ;
  assign \nz.mem [1021] = \nz.mem_1021_sv2v_reg ;
  assign \nz.mem [1020] = \nz.mem_1020_sv2v_reg ;
  assign \nz.mem [1019] = \nz.mem_1019_sv2v_reg ;
  assign \nz.mem [1018] = \nz.mem_1018_sv2v_reg ;
  assign \nz.mem [1017] = \nz.mem_1017_sv2v_reg ;
  assign \nz.mem [1016] = \nz.mem_1016_sv2v_reg ;
  assign \nz.mem [1015] = \nz.mem_1015_sv2v_reg ;
  assign \nz.mem [1014] = \nz.mem_1014_sv2v_reg ;
  assign \nz.mem [1013] = \nz.mem_1013_sv2v_reg ;
  assign \nz.mem [1012] = \nz.mem_1012_sv2v_reg ;
  assign \nz.mem [1011] = \nz.mem_1011_sv2v_reg ;
  assign \nz.mem [1010] = \nz.mem_1010_sv2v_reg ;
  assign \nz.mem [1009] = \nz.mem_1009_sv2v_reg ;
  assign \nz.mem [1008] = \nz.mem_1008_sv2v_reg ;
  assign \nz.mem [1007] = \nz.mem_1007_sv2v_reg ;
  assign \nz.mem [1006] = \nz.mem_1006_sv2v_reg ;
  assign \nz.mem [1005] = \nz.mem_1005_sv2v_reg ;
  assign \nz.mem [1004] = \nz.mem_1004_sv2v_reg ;
  assign \nz.mem [1003] = \nz.mem_1003_sv2v_reg ;
  assign \nz.mem [1002] = \nz.mem_1002_sv2v_reg ;
  assign \nz.mem [1001] = \nz.mem_1001_sv2v_reg ;
  assign \nz.mem [1000] = \nz.mem_1000_sv2v_reg ;
  assign \nz.mem [999] = \nz.mem_999_sv2v_reg ;
  assign \nz.mem [998] = \nz.mem_998_sv2v_reg ;
  assign \nz.mem [997] = \nz.mem_997_sv2v_reg ;
  assign \nz.mem [996] = \nz.mem_996_sv2v_reg ;
  assign \nz.mem [995] = \nz.mem_995_sv2v_reg ;
  assign \nz.mem [994] = \nz.mem_994_sv2v_reg ;
  assign \nz.mem [993] = \nz.mem_993_sv2v_reg ;
  assign \nz.mem [992] = \nz.mem_992_sv2v_reg ;
  assign \nz.mem [991] = \nz.mem_991_sv2v_reg ;
  assign \nz.mem [990] = \nz.mem_990_sv2v_reg ;
  assign \nz.mem [989] = \nz.mem_989_sv2v_reg ;
  assign \nz.mem [988] = \nz.mem_988_sv2v_reg ;
  assign \nz.mem [987] = \nz.mem_987_sv2v_reg ;
  assign \nz.mem [986] = \nz.mem_986_sv2v_reg ;
  assign \nz.mem [985] = \nz.mem_985_sv2v_reg ;
  assign \nz.mem [984] = \nz.mem_984_sv2v_reg ;
  assign \nz.mem [983] = \nz.mem_983_sv2v_reg ;
  assign \nz.mem [982] = \nz.mem_982_sv2v_reg ;
  assign \nz.mem [981] = \nz.mem_981_sv2v_reg ;
  assign \nz.mem [980] = \nz.mem_980_sv2v_reg ;
  assign \nz.mem [979] = \nz.mem_979_sv2v_reg ;
  assign \nz.mem [978] = \nz.mem_978_sv2v_reg ;
  assign \nz.mem [977] = \nz.mem_977_sv2v_reg ;
  assign \nz.mem [976] = \nz.mem_976_sv2v_reg ;
  assign \nz.mem [975] = \nz.mem_975_sv2v_reg ;
  assign \nz.mem [974] = \nz.mem_974_sv2v_reg ;
  assign \nz.mem [973] = \nz.mem_973_sv2v_reg ;
  assign \nz.mem [972] = \nz.mem_972_sv2v_reg ;
  assign \nz.mem [971] = \nz.mem_971_sv2v_reg ;
  assign \nz.mem [970] = \nz.mem_970_sv2v_reg ;
  assign \nz.mem [969] = \nz.mem_969_sv2v_reg ;
  assign \nz.mem [968] = \nz.mem_968_sv2v_reg ;
  assign \nz.mem [967] = \nz.mem_967_sv2v_reg ;
  assign \nz.mem [966] = \nz.mem_966_sv2v_reg ;
  assign \nz.mem [965] = \nz.mem_965_sv2v_reg ;
  assign \nz.mem [964] = \nz.mem_964_sv2v_reg ;
  assign \nz.mem [963] = \nz.mem_963_sv2v_reg ;
  assign \nz.mem [962] = \nz.mem_962_sv2v_reg ;
  assign \nz.mem [961] = \nz.mem_961_sv2v_reg ;
  assign \nz.mem [960] = \nz.mem_960_sv2v_reg ;
  assign \nz.mem [959] = \nz.mem_959_sv2v_reg ;
  assign \nz.mem [958] = \nz.mem_958_sv2v_reg ;
  assign \nz.mem [957] = \nz.mem_957_sv2v_reg ;
  assign \nz.mem [956] = \nz.mem_956_sv2v_reg ;
  assign \nz.mem [955] = \nz.mem_955_sv2v_reg ;
  assign \nz.mem [954] = \nz.mem_954_sv2v_reg ;
  assign \nz.mem [953] = \nz.mem_953_sv2v_reg ;
  assign \nz.mem [952] = \nz.mem_952_sv2v_reg ;
  assign \nz.mem [951] = \nz.mem_951_sv2v_reg ;
  assign \nz.mem [950] = \nz.mem_950_sv2v_reg ;
  assign \nz.mem [949] = \nz.mem_949_sv2v_reg ;
  assign \nz.mem [948] = \nz.mem_948_sv2v_reg ;
  assign \nz.mem [947] = \nz.mem_947_sv2v_reg ;
  assign \nz.mem [946] = \nz.mem_946_sv2v_reg ;
  assign \nz.mem [945] = \nz.mem_945_sv2v_reg ;
  assign \nz.mem [944] = \nz.mem_944_sv2v_reg ;
  assign \nz.mem [943] = \nz.mem_943_sv2v_reg ;
  assign \nz.mem [942] = \nz.mem_942_sv2v_reg ;
  assign \nz.mem [941] = \nz.mem_941_sv2v_reg ;
  assign \nz.mem [940] = \nz.mem_940_sv2v_reg ;
  assign \nz.mem [939] = \nz.mem_939_sv2v_reg ;
  assign \nz.mem [938] = \nz.mem_938_sv2v_reg ;
  assign \nz.mem [937] = \nz.mem_937_sv2v_reg ;
  assign \nz.mem [936] = \nz.mem_936_sv2v_reg ;
  assign \nz.mem [935] = \nz.mem_935_sv2v_reg ;
  assign \nz.mem [934] = \nz.mem_934_sv2v_reg ;
  assign \nz.mem [933] = \nz.mem_933_sv2v_reg ;
  assign \nz.mem [932] = \nz.mem_932_sv2v_reg ;
  assign \nz.mem [931] = \nz.mem_931_sv2v_reg ;
  assign \nz.mem [930] = \nz.mem_930_sv2v_reg ;
  assign \nz.mem [929] = \nz.mem_929_sv2v_reg ;
  assign \nz.mem [928] = \nz.mem_928_sv2v_reg ;
  assign \nz.mem [927] = \nz.mem_927_sv2v_reg ;
  assign \nz.mem [926] = \nz.mem_926_sv2v_reg ;
  assign \nz.mem [925] = \nz.mem_925_sv2v_reg ;
  assign \nz.mem [924] = \nz.mem_924_sv2v_reg ;
  assign \nz.mem [923] = \nz.mem_923_sv2v_reg ;
  assign \nz.mem [922] = \nz.mem_922_sv2v_reg ;
  assign \nz.mem [921] = \nz.mem_921_sv2v_reg ;
  assign \nz.mem [920] = \nz.mem_920_sv2v_reg ;
  assign \nz.mem [919] = \nz.mem_919_sv2v_reg ;
  assign \nz.mem [918] = \nz.mem_918_sv2v_reg ;
  assign \nz.mem [917] = \nz.mem_917_sv2v_reg ;
  assign \nz.mem [916] = \nz.mem_916_sv2v_reg ;
  assign \nz.mem [915] = \nz.mem_915_sv2v_reg ;
  assign \nz.mem [914] = \nz.mem_914_sv2v_reg ;
  assign \nz.mem [913] = \nz.mem_913_sv2v_reg ;
  assign \nz.mem [912] = \nz.mem_912_sv2v_reg ;
  assign \nz.mem [911] = \nz.mem_911_sv2v_reg ;
  assign \nz.mem [910] = \nz.mem_910_sv2v_reg ;
  assign \nz.mem [909] = \nz.mem_909_sv2v_reg ;
  assign \nz.mem [908] = \nz.mem_908_sv2v_reg ;
  assign \nz.mem [907] = \nz.mem_907_sv2v_reg ;
  assign \nz.mem [906] = \nz.mem_906_sv2v_reg ;
  assign \nz.mem [905] = \nz.mem_905_sv2v_reg ;
  assign \nz.mem [904] = \nz.mem_904_sv2v_reg ;
  assign \nz.mem [903] = \nz.mem_903_sv2v_reg ;
  assign \nz.mem [902] = \nz.mem_902_sv2v_reg ;
  assign \nz.mem [901] = \nz.mem_901_sv2v_reg ;
  assign \nz.mem [900] = \nz.mem_900_sv2v_reg ;
  assign \nz.mem [899] = \nz.mem_899_sv2v_reg ;
  assign \nz.mem [898] = \nz.mem_898_sv2v_reg ;
  assign \nz.mem [897] = \nz.mem_897_sv2v_reg ;
  assign \nz.mem [896] = \nz.mem_896_sv2v_reg ;
  assign \nz.mem [895] = \nz.mem_895_sv2v_reg ;
  assign \nz.mem [894] = \nz.mem_894_sv2v_reg ;
  assign \nz.mem [893] = \nz.mem_893_sv2v_reg ;
  assign \nz.mem [892] = \nz.mem_892_sv2v_reg ;
  assign \nz.mem [891] = \nz.mem_891_sv2v_reg ;
  assign \nz.mem [890] = \nz.mem_890_sv2v_reg ;
  assign \nz.mem [889] = \nz.mem_889_sv2v_reg ;
  assign \nz.mem [888] = \nz.mem_888_sv2v_reg ;
  assign \nz.mem [887] = \nz.mem_887_sv2v_reg ;
  assign \nz.mem [886] = \nz.mem_886_sv2v_reg ;
  assign \nz.mem [885] = \nz.mem_885_sv2v_reg ;
  assign \nz.mem [884] = \nz.mem_884_sv2v_reg ;
  assign \nz.mem [883] = \nz.mem_883_sv2v_reg ;
  assign \nz.mem [882] = \nz.mem_882_sv2v_reg ;
  assign \nz.mem [881] = \nz.mem_881_sv2v_reg ;
  assign \nz.mem [880] = \nz.mem_880_sv2v_reg ;
  assign \nz.mem [879] = \nz.mem_879_sv2v_reg ;
  assign \nz.mem [878] = \nz.mem_878_sv2v_reg ;
  assign \nz.mem [877] = \nz.mem_877_sv2v_reg ;
  assign \nz.mem [876] = \nz.mem_876_sv2v_reg ;
  assign \nz.mem [875] = \nz.mem_875_sv2v_reg ;
  assign \nz.mem [874] = \nz.mem_874_sv2v_reg ;
  assign \nz.mem [873] = \nz.mem_873_sv2v_reg ;
  assign \nz.mem [872] = \nz.mem_872_sv2v_reg ;
  assign \nz.mem [871] = \nz.mem_871_sv2v_reg ;
  assign \nz.mem [870] = \nz.mem_870_sv2v_reg ;
  assign \nz.mem [869] = \nz.mem_869_sv2v_reg ;
  assign \nz.mem [868] = \nz.mem_868_sv2v_reg ;
  assign \nz.mem [867] = \nz.mem_867_sv2v_reg ;
  assign \nz.mem [866] = \nz.mem_866_sv2v_reg ;
  assign \nz.mem [865] = \nz.mem_865_sv2v_reg ;
  assign \nz.mem [864] = \nz.mem_864_sv2v_reg ;
  assign \nz.mem [863] = \nz.mem_863_sv2v_reg ;
  assign \nz.mem [862] = \nz.mem_862_sv2v_reg ;
  assign \nz.mem [861] = \nz.mem_861_sv2v_reg ;
  assign \nz.mem [860] = \nz.mem_860_sv2v_reg ;
  assign \nz.mem [859] = \nz.mem_859_sv2v_reg ;
  assign \nz.mem [858] = \nz.mem_858_sv2v_reg ;
  assign \nz.mem [857] = \nz.mem_857_sv2v_reg ;
  assign \nz.mem [856] = \nz.mem_856_sv2v_reg ;
  assign \nz.mem [855] = \nz.mem_855_sv2v_reg ;
  assign \nz.mem [854] = \nz.mem_854_sv2v_reg ;
  assign \nz.mem [853] = \nz.mem_853_sv2v_reg ;
  assign \nz.mem [852] = \nz.mem_852_sv2v_reg ;
  assign \nz.mem [851] = \nz.mem_851_sv2v_reg ;
  assign \nz.mem [850] = \nz.mem_850_sv2v_reg ;
  assign \nz.mem [849] = \nz.mem_849_sv2v_reg ;
  assign \nz.mem [848] = \nz.mem_848_sv2v_reg ;
  assign \nz.mem [847] = \nz.mem_847_sv2v_reg ;
  assign \nz.mem [846] = \nz.mem_846_sv2v_reg ;
  assign \nz.mem [845] = \nz.mem_845_sv2v_reg ;
  assign \nz.mem [844] = \nz.mem_844_sv2v_reg ;
  assign \nz.mem [843] = \nz.mem_843_sv2v_reg ;
  assign \nz.mem [842] = \nz.mem_842_sv2v_reg ;
  assign \nz.mem [841] = \nz.mem_841_sv2v_reg ;
  assign \nz.mem [840] = \nz.mem_840_sv2v_reg ;
  assign \nz.mem [839] = \nz.mem_839_sv2v_reg ;
  assign \nz.mem [838] = \nz.mem_838_sv2v_reg ;
  assign \nz.mem [837] = \nz.mem_837_sv2v_reg ;
  assign \nz.mem [836] = \nz.mem_836_sv2v_reg ;
  assign \nz.mem [835] = \nz.mem_835_sv2v_reg ;
  assign \nz.mem [834] = \nz.mem_834_sv2v_reg ;
  assign \nz.mem [833] = \nz.mem_833_sv2v_reg ;
  assign \nz.mem [832] = \nz.mem_832_sv2v_reg ;
  assign \nz.mem [831] = \nz.mem_831_sv2v_reg ;
  assign \nz.mem [830] = \nz.mem_830_sv2v_reg ;
  assign \nz.mem [829] = \nz.mem_829_sv2v_reg ;
  assign \nz.mem [828] = \nz.mem_828_sv2v_reg ;
  assign \nz.mem [827] = \nz.mem_827_sv2v_reg ;
  assign \nz.mem [826] = \nz.mem_826_sv2v_reg ;
  assign \nz.mem [825] = \nz.mem_825_sv2v_reg ;
  assign \nz.mem [824] = \nz.mem_824_sv2v_reg ;
  assign \nz.mem [823] = \nz.mem_823_sv2v_reg ;
  assign \nz.mem [822] = \nz.mem_822_sv2v_reg ;
  assign \nz.mem [821] = \nz.mem_821_sv2v_reg ;
  assign \nz.mem [820] = \nz.mem_820_sv2v_reg ;
  assign \nz.mem [819] = \nz.mem_819_sv2v_reg ;
  assign \nz.mem [818] = \nz.mem_818_sv2v_reg ;
  assign \nz.mem [817] = \nz.mem_817_sv2v_reg ;
  assign \nz.mem [816] = \nz.mem_816_sv2v_reg ;
  assign \nz.mem [815] = \nz.mem_815_sv2v_reg ;
  assign \nz.mem [814] = \nz.mem_814_sv2v_reg ;
  assign \nz.mem [813] = \nz.mem_813_sv2v_reg ;
  assign \nz.mem [812] = \nz.mem_812_sv2v_reg ;
  assign \nz.mem [811] = \nz.mem_811_sv2v_reg ;
  assign \nz.mem [810] = \nz.mem_810_sv2v_reg ;
  assign \nz.mem [809] = \nz.mem_809_sv2v_reg ;
  assign \nz.mem [808] = \nz.mem_808_sv2v_reg ;
  assign \nz.mem [807] = \nz.mem_807_sv2v_reg ;
  assign \nz.mem [806] = \nz.mem_806_sv2v_reg ;
  assign \nz.mem [805] = \nz.mem_805_sv2v_reg ;
  assign \nz.mem [804] = \nz.mem_804_sv2v_reg ;
  assign \nz.mem [803] = \nz.mem_803_sv2v_reg ;
  assign \nz.mem [802] = \nz.mem_802_sv2v_reg ;
  assign \nz.mem [801] = \nz.mem_801_sv2v_reg ;
  assign \nz.mem [800] = \nz.mem_800_sv2v_reg ;
  assign \nz.mem [799] = \nz.mem_799_sv2v_reg ;
  assign \nz.mem [798] = \nz.mem_798_sv2v_reg ;
  assign \nz.mem [797] = \nz.mem_797_sv2v_reg ;
  assign \nz.mem [796] = \nz.mem_796_sv2v_reg ;
  assign \nz.mem [795] = \nz.mem_795_sv2v_reg ;
  assign \nz.mem [794] = \nz.mem_794_sv2v_reg ;
  assign \nz.mem [793] = \nz.mem_793_sv2v_reg ;
  assign \nz.mem [792] = \nz.mem_792_sv2v_reg ;
  assign \nz.mem [791] = \nz.mem_791_sv2v_reg ;
  assign \nz.mem [790] = \nz.mem_790_sv2v_reg ;
  assign \nz.mem [789] = \nz.mem_789_sv2v_reg ;
  assign \nz.mem [788] = \nz.mem_788_sv2v_reg ;
  assign \nz.mem [787] = \nz.mem_787_sv2v_reg ;
  assign \nz.mem [786] = \nz.mem_786_sv2v_reg ;
  assign \nz.mem [785] = \nz.mem_785_sv2v_reg ;
  assign \nz.mem [784] = \nz.mem_784_sv2v_reg ;
  assign \nz.mem [783] = \nz.mem_783_sv2v_reg ;
  assign \nz.mem [782] = \nz.mem_782_sv2v_reg ;
  assign \nz.mem [781] = \nz.mem_781_sv2v_reg ;
  assign \nz.mem [780] = \nz.mem_780_sv2v_reg ;
  assign \nz.mem [779] = \nz.mem_779_sv2v_reg ;
  assign \nz.mem [778] = \nz.mem_778_sv2v_reg ;
  assign \nz.mem [777] = \nz.mem_777_sv2v_reg ;
  assign \nz.mem [776] = \nz.mem_776_sv2v_reg ;
  assign \nz.mem [775] = \nz.mem_775_sv2v_reg ;
  assign \nz.mem [774] = \nz.mem_774_sv2v_reg ;
  assign \nz.mem [773] = \nz.mem_773_sv2v_reg ;
  assign \nz.mem [772] = \nz.mem_772_sv2v_reg ;
  assign \nz.mem [771] = \nz.mem_771_sv2v_reg ;
  assign \nz.mem [770] = \nz.mem_770_sv2v_reg ;
  assign \nz.mem [769] = \nz.mem_769_sv2v_reg ;
  assign \nz.mem [768] = \nz.mem_768_sv2v_reg ;
  assign \nz.mem [767] = \nz.mem_767_sv2v_reg ;
  assign \nz.mem [766] = \nz.mem_766_sv2v_reg ;
  assign \nz.mem [765] = \nz.mem_765_sv2v_reg ;
  assign \nz.mem [764] = \nz.mem_764_sv2v_reg ;
  assign \nz.mem [763] = \nz.mem_763_sv2v_reg ;
  assign \nz.mem [762] = \nz.mem_762_sv2v_reg ;
  assign \nz.mem [761] = \nz.mem_761_sv2v_reg ;
  assign \nz.mem [760] = \nz.mem_760_sv2v_reg ;
  assign \nz.mem [759] = \nz.mem_759_sv2v_reg ;
  assign \nz.mem [758] = \nz.mem_758_sv2v_reg ;
  assign \nz.mem [757] = \nz.mem_757_sv2v_reg ;
  assign \nz.mem [756] = \nz.mem_756_sv2v_reg ;
  assign \nz.mem [755] = \nz.mem_755_sv2v_reg ;
  assign \nz.mem [754] = \nz.mem_754_sv2v_reg ;
  assign \nz.mem [753] = \nz.mem_753_sv2v_reg ;
  assign \nz.mem [752] = \nz.mem_752_sv2v_reg ;
  assign \nz.mem [751] = \nz.mem_751_sv2v_reg ;
  assign \nz.mem [750] = \nz.mem_750_sv2v_reg ;
  assign \nz.mem [749] = \nz.mem_749_sv2v_reg ;
  assign \nz.mem [748] = \nz.mem_748_sv2v_reg ;
  assign \nz.mem [747] = \nz.mem_747_sv2v_reg ;
  assign \nz.mem [746] = \nz.mem_746_sv2v_reg ;
  assign \nz.mem [745] = \nz.mem_745_sv2v_reg ;
  assign \nz.mem [744] = \nz.mem_744_sv2v_reg ;
  assign \nz.mem [743] = \nz.mem_743_sv2v_reg ;
  assign \nz.mem [742] = \nz.mem_742_sv2v_reg ;
  assign \nz.mem [741] = \nz.mem_741_sv2v_reg ;
  assign \nz.mem [740] = \nz.mem_740_sv2v_reg ;
  assign \nz.mem [739] = \nz.mem_739_sv2v_reg ;
  assign \nz.mem [738] = \nz.mem_738_sv2v_reg ;
  assign \nz.mem [737] = \nz.mem_737_sv2v_reg ;
  assign \nz.mem [736] = \nz.mem_736_sv2v_reg ;
  assign \nz.mem [735] = \nz.mem_735_sv2v_reg ;
  assign \nz.mem [734] = \nz.mem_734_sv2v_reg ;
  assign \nz.mem [733] = \nz.mem_733_sv2v_reg ;
  assign \nz.mem [732] = \nz.mem_732_sv2v_reg ;
  assign \nz.mem [731] = \nz.mem_731_sv2v_reg ;
  assign \nz.mem [730] = \nz.mem_730_sv2v_reg ;
  assign \nz.mem [729] = \nz.mem_729_sv2v_reg ;
  assign \nz.mem [728] = \nz.mem_728_sv2v_reg ;
  assign \nz.mem [727] = \nz.mem_727_sv2v_reg ;
  assign \nz.mem [726] = \nz.mem_726_sv2v_reg ;
  assign \nz.mem [725] = \nz.mem_725_sv2v_reg ;
  assign \nz.mem [724] = \nz.mem_724_sv2v_reg ;
  assign \nz.mem [723] = \nz.mem_723_sv2v_reg ;
  assign \nz.mem [722] = \nz.mem_722_sv2v_reg ;
  assign \nz.mem [721] = \nz.mem_721_sv2v_reg ;
  assign \nz.mem [720] = \nz.mem_720_sv2v_reg ;
  assign \nz.mem [719] = \nz.mem_719_sv2v_reg ;
  assign \nz.mem [718] = \nz.mem_718_sv2v_reg ;
  assign \nz.mem [717] = \nz.mem_717_sv2v_reg ;
  assign \nz.mem [716] = \nz.mem_716_sv2v_reg ;
  assign \nz.mem [715] = \nz.mem_715_sv2v_reg ;
  assign \nz.mem [714] = \nz.mem_714_sv2v_reg ;
  assign \nz.mem [713] = \nz.mem_713_sv2v_reg ;
  assign \nz.mem [712] = \nz.mem_712_sv2v_reg ;
  assign \nz.mem [711] = \nz.mem_711_sv2v_reg ;
  assign \nz.mem [710] = \nz.mem_710_sv2v_reg ;
  assign \nz.mem [709] = \nz.mem_709_sv2v_reg ;
  assign \nz.mem [708] = \nz.mem_708_sv2v_reg ;
  assign \nz.mem [707] = \nz.mem_707_sv2v_reg ;
  assign \nz.mem [706] = \nz.mem_706_sv2v_reg ;
  assign \nz.mem [705] = \nz.mem_705_sv2v_reg ;
  assign \nz.mem [704] = \nz.mem_704_sv2v_reg ;
  assign \nz.mem [703] = \nz.mem_703_sv2v_reg ;
  assign \nz.mem [702] = \nz.mem_702_sv2v_reg ;
  assign \nz.mem [701] = \nz.mem_701_sv2v_reg ;
  assign \nz.mem [700] = \nz.mem_700_sv2v_reg ;
  assign \nz.mem [699] = \nz.mem_699_sv2v_reg ;
  assign \nz.mem [698] = \nz.mem_698_sv2v_reg ;
  assign \nz.mem [697] = \nz.mem_697_sv2v_reg ;
  assign \nz.mem [696] = \nz.mem_696_sv2v_reg ;
  assign \nz.mem [695] = \nz.mem_695_sv2v_reg ;
  assign \nz.mem [694] = \nz.mem_694_sv2v_reg ;
  assign \nz.mem [693] = \nz.mem_693_sv2v_reg ;
  assign \nz.mem [692] = \nz.mem_692_sv2v_reg ;
  assign \nz.mem [691] = \nz.mem_691_sv2v_reg ;
  assign \nz.mem [690] = \nz.mem_690_sv2v_reg ;
  assign \nz.mem [689] = \nz.mem_689_sv2v_reg ;
  assign \nz.mem [688] = \nz.mem_688_sv2v_reg ;
  assign \nz.mem [687] = \nz.mem_687_sv2v_reg ;
  assign \nz.mem [686] = \nz.mem_686_sv2v_reg ;
  assign \nz.mem [685] = \nz.mem_685_sv2v_reg ;
  assign \nz.mem [684] = \nz.mem_684_sv2v_reg ;
  assign \nz.mem [683] = \nz.mem_683_sv2v_reg ;
  assign \nz.mem [682] = \nz.mem_682_sv2v_reg ;
  assign \nz.mem [681] = \nz.mem_681_sv2v_reg ;
  assign \nz.mem [680] = \nz.mem_680_sv2v_reg ;
  assign \nz.mem [679] = \nz.mem_679_sv2v_reg ;
  assign \nz.mem [678] = \nz.mem_678_sv2v_reg ;
  assign \nz.mem [677] = \nz.mem_677_sv2v_reg ;
  assign \nz.mem [676] = \nz.mem_676_sv2v_reg ;
  assign \nz.mem [675] = \nz.mem_675_sv2v_reg ;
  assign \nz.mem [674] = \nz.mem_674_sv2v_reg ;
  assign \nz.mem [673] = \nz.mem_673_sv2v_reg ;
  assign \nz.mem [672] = \nz.mem_672_sv2v_reg ;
  assign \nz.mem [671] = \nz.mem_671_sv2v_reg ;
  assign \nz.mem [670] = \nz.mem_670_sv2v_reg ;
  assign \nz.mem [669] = \nz.mem_669_sv2v_reg ;
  assign \nz.mem [668] = \nz.mem_668_sv2v_reg ;
  assign \nz.mem [667] = \nz.mem_667_sv2v_reg ;
  assign \nz.mem [666] = \nz.mem_666_sv2v_reg ;
  assign \nz.mem [665] = \nz.mem_665_sv2v_reg ;
  assign \nz.mem [664] = \nz.mem_664_sv2v_reg ;
  assign \nz.mem [663] = \nz.mem_663_sv2v_reg ;
  assign \nz.mem [662] = \nz.mem_662_sv2v_reg ;
  assign \nz.mem [661] = \nz.mem_661_sv2v_reg ;
  assign \nz.mem [660] = \nz.mem_660_sv2v_reg ;
  assign \nz.mem [659] = \nz.mem_659_sv2v_reg ;
  assign \nz.mem [658] = \nz.mem_658_sv2v_reg ;
  assign \nz.mem [657] = \nz.mem_657_sv2v_reg ;
  assign \nz.mem [656] = \nz.mem_656_sv2v_reg ;
  assign \nz.mem [655] = \nz.mem_655_sv2v_reg ;
  assign \nz.mem [654] = \nz.mem_654_sv2v_reg ;
  assign \nz.mem [653] = \nz.mem_653_sv2v_reg ;
  assign \nz.mem [652] = \nz.mem_652_sv2v_reg ;
  assign \nz.mem [651] = \nz.mem_651_sv2v_reg ;
  assign \nz.mem [650] = \nz.mem_650_sv2v_reg ;
  assign \nz.mem [649] = \nz.mem_649_sv2v_reg ;
  assign \nz.mem [648] = \nz.mem_648_sv2v_reg ;
  assign \nz.mem [647] = \nz.mem_647_sv2v_reg ;
  assign \nz.mem [646] = \nz.mem_646_sv2v_reg ;
  assign \nz.mem [645] = \nz.mem_645_sv2v_reg ;
  assign \nz.mem [644] = \nz.mem_644_sv2v_reg ;
  assign \nz.mem [643] = \nz.mem_643_sv2v_reg ;
  assign \nz.mem [642] = \nz.mem_642_sv2v_reg ;
  assign \nz.mem [641] = \nz.mem_641_sv2v_reg ;
  assign \nz.mem [640] = \nz.mem_640_sv2v_reg ;
  assign \nz.mem [639] = \nz.mem_639_sv2v_reg ;
  assign \nz.mem [638] = \nz.mem_638_sv2v_reg ;
  assign \nz.mem [637] = \nz.mem_637_sv2v_reg ;
  assign \nz.mem [636] = \nz.mem_636_sv2v_reg ;
  assign \nz.mem [635] = \nz.mem_635_sv2v_reg ;
  assign \nz.mem [634] = \nz.mem_634_sv2v_reg ;
  assign \nz.mem [633] = \nz.mem_633_sv2v_reg ;
  assign \nz.mem [632] = \nz.mem_632_sv2v_reg ;
  assign \nz.mem [631] = \nz.mem_631_sv2v_reg ;
  assign \nz.mem [630] = \nz.mem_630_sv2v_reg ;
  assign \nz.mem [629] = \nz.mem_629_sv2v_reg ;
  assign \nz.mem [628] = \nz.mem_628_sv2v_reg ;
  assign \nz.mem [627] = \nz.mem_627_sv2v_reg ;
  assign \nz.mem [626] = \nz.mem_626_sv2v_reg ;
  assign \nz.mem [625] = \nz.mem_625_sv2v_reg ;
  assign \nz.mem [624] = \nz.mem_624_sv2v_reg ;
  assign \nz.mem [623] = \nz.mem_623_sv2v_reg ;
  assign \nz.mem [622] = \nz.mem_622_sv2v_reg ;
  assign \nz.mem [621] = \nz.mem_621_sv2v_reg ;
  assign \nz.mem [620] = \nz.mem_620_sv2v_reg ;
  assign \nz.mem [619] = \nz.mem_619_sv2v_reg ;
  assign \nz.mem [618] = \nz.mem_618_sv2v_reg ;
  assign \nz.mem [617] = \nz.mem_617_sv2v_reg ;
  assign \nz.mem [616] = \nz.mem_616_sv2v_reg ;
  assign \nz.mem [615] = \nz.mem_615_sv2v_reg ;
  assign \nz.mem [614] = \nz.mem_614_sv2v_reg ;
  assign \nz.mem [613] = \nz.mem_613_sv2v_reg ;
  assign \nz.mem [612] = \nz.mem_612_sv2v_reg ;
  assign \nz.mem [611] = \nz.mem_611_sv2v_reg ;
  assign \nz.mem [610] = \nz.mem_610_sv2v_reg ;
  assign \nz.mem [609] = \nz.mem_609_sv2v_reg ;
  assign \nz.mem [608] = \nz.mem_608_sv2v_reg ;
  assign \nz.mem [607] = \nz.mem_607_sv2v_reg ;
  assign \nz.mem [606] = \nz.mem_606_sv2v_reg ;
  assign \nz.mem [605] = \nz.mem_605_sv2v_reg ;
  assign \nz.mem [604] = \nz.mem_604_sv2v_reg ;
  assign \nz.mem [603] = \nz.mem_603_sv2v_reg ;
  assign \nz.mem [602] = \nz.mem_602_sv2v_reg ;
  assign \nz.mem [601] = \nz.mem_601_sv2v_reg ;
  assign \nz.mem [600] = \nz.mem_600_sv2v_reg ;
  assign \nz.mem [599] = \nz.mem_599_sv2v_reg ;
  assign \nz.mem [598] = \nz.mem_598_sv2v_reg ;
  assign \nz.mem [597] = \nz.mem_597_sv2v_reg ;
  assign \nz.mem [596] = \nz.mem_596_sv2v_reg ;
  assign \nz.mem [595] = \nz.mem_595_sv2v_reg ;
  assign \nz.mem [594] = \nz.mem_594_sv2v_reg ;
  assign \nz.mem [593] = \nz.mem_593_sv2v_reg ;
  assign \nz.mem [592] = \nz.mem_592_sv2v_reg ;
  assign \nz.mem [591] = \nz.mem_591_sv2v_reg ;
  assign \nz.mem [590] = \nz.mem_590_sv2v_reg ;
  assign \nz.mem [589] = \nz.mem_589_sv2v_reg ;
  assign \nz.mem [588] = \nz.mem_588_sv2v_reg ;
  assign \nz.mem [587] = \nz.mem_587_sv2v_reg ;
  assign \nz.mem [586] = \nz.mem_586_sv2v_reg ;
  assign \nz.mem [585] = \nz.mem_585_sv2v_reg ;
  assign \nz.mem [584] = \nz.mem_584_sv2v_reg ;
  assign \nz.mem [583] = \nz.mem_583_sv2v_reg ;
  assign \nz.mem [582] = \nz.mem_582_sv2v_reg ;
  assign \nz.mem [581] = \nz.mem_581_sv2v_reg ;
  assign \nz.mem [580] = \nz.mem_580_sv2v_reg ;
  assign \nz.mem [579] = \nz.mem_579_sv2v_reg ;
  assign \nz.mem [578] = \nz.mem_578_sv2v_reg ;
  assign \nz.mem [577] = \nz.mem_577_sv2v_reg ;
  assign \nz.mem [576] = \nz.mem_576_sv2v_reg ;
  assign \nz.mem [575] = \nz.mem_575_sv2v_reg ;
  assign \nz.mem [574] = \nz.mem_574_sv2v_reg ;
  assign \nz.mem [573] = \nz.mem_573_sv2v_reg ;
  assign \nz.mem [572] = \nz.mem_572_sv2v_reg ;
  assign \nz.mem [571] = \nz.mem_571_sv2v_reg ;
  assign \nz.mem [570] = \nz.mem_570_sv2v_reg ;
  assign \nz.mem [569] = \nz.mem_569_sv2v_reg ;
  assign \nz.mem [568] = \nz.mem_568_sv2v_reg ;
  assign \nz.mem [567] = \nz.mem_567_sv2v_reg ;
  assign \nz.mem [566] = \nz.mem_566_sv2v_reg ;
  assign \nz.mem [565] = \nz.mem_565_sv2v_reg ;
  assign \nz.mem [564] = \nz.mem_564_sv2v_reg ;
  assign \nz.mem [563] = \nz.mem_563_sv2v_reg ;
  assign \nz.mem [562] = \nz.mem_562_sv2v_reg ;
  assign \nz.mem [561] = \nz.mem_561_sv2v_reg ;
  assign \nz.mem [560] = \nz.mem_560_sv2v_reg ;
  assign \nz.mem [559] = \nz.mem_559_sv2v_reg ;
  assign \nz.mem [558] = \nz.mem_558_sv2v_reg ;
  assign \nz.mem [557] = \nz.mem_557_sv2v_reg ;
  assign \nz.mem [556] = \nz.mem_556_sv2v_reg ;
  assign \nz.mem [555] = \nz.mem_555_sv2v_reg ;
  assign \nz.mem [554] = \nz.mem_554_sv2v_reg ;
  assign \nz.mem [553] = \nz.mem_553_sv2v_reg ;
  assign \nz.mem [552] = \nz.mem_552_sv2v_reg ;
  assign \nz.mem [551] = \nz.mem_551_sv2v_reg ;
  assign \nz.mem [550] = \nz.mem_550_sv2v_reg ;
  assign \nz.mem [549] = \nz.mem_549_sv2v_reg ;
  assign \nz.mem [548] = \nz.mem_548_sv2v_reg ;
  assign \nz.mem [547] = \nz.mem_547_sv2v_reg ;
  assign \nz.mem [546] = \nz.mem_546_sv2v_reg ;
  assign \nz.mem [545] = \nz.mem_545_sv2v_reg ;
  assign \nz.mem [544] = \nz.mem_544_sv2v_reg ;
  assign \nz.mem [543] = \nz.mem_543_sv2v_reg ;
  assign \nz.mem [542] = \nz.mem_542_sv2v_reg ;
  assign \nz.mem [541] = \nz.mem_541_sv2v_reg ;
  assign \nz.mem [540] = \nz.mem_540_sv2v_reg ;
  assign \nz.mem [539] = \nz.mem_539_sv2v_reg ;
  assign \nz.mem [538] = \nz.mem_538_sv2v_reg ;
  assign \nz.mem [537] = \nz.mem_537_sv2v_reg ;
  assign \nz.mem [536] = \nz.mem_536_sv2v_reg ;
  assign \nz.mem [535] = \nz.mem_535_sv2v_reg ;
  assign \nz.mem [534] = \nz.mem_534_sv2v_reg ;
  assign \nz.mem [533] = \nz.mem_533_sv2v_reg ;
  assign \nz.mem [532] = \nz.mem_532_sv2v_reg ;
  assign \nz.mem [531] = \nz.mem_531_sv2v_reg ;
  assign \nz.mem [530] = \nz.mem_530_sv2v_reg ;
  assign \nz.mem [529] = \nz.mem_529_sv2v_reg ;
  assign \nz.mem [528] = \nz.mem_528_sv2v_reg ;
  assign \nz.mem [527] = \nz.mem_527_sv2v_reg ;
  assign \nz.mem [526] = \nz.mem_526_sv2v_reg ;
  assign \nz.mem [525] = \nz.mem_525_sv2v_reg ;
  assign \nz.mem [524] = \nz.mem_524_sv2v_reg ;
  assign \nz.mem [523] = \nz.mem_523_sv2v_reg ;
  assign \nz.mem [522] = \nz.mem_522_sv2v_reg ;
  assign \nz.mem [521] = \nz.mem_521_sv2v_reg ;
  assign \nz.mem [520] = \nz.mem_520_sv2v_reg ;
  assign \nz.mem [519] = \nz.mem_519_sv2v_reg ;
  assign \nz.mem [518] = \nz.mem_518_sv2v_reg ;
  assign \nz.mem [517] = \nz.mem_517_sv2v_reg ;
  assign \nz.mem [516] = \nz.mem_516_sv2v_reg ;
  assign \nz.mem [515] = \nz.mem_515_sv2v_reg ;
  assign \nz.mem [514] = \nz.mem_514_sv2v_reg ;
  assign \nz.mem [513] = \nz.mem_513_sv2v_reg ;
  assign \nz.mem [512] = \nz.mem_512_sv2v_reg ;
  assign \nz.mem [511] = \nz.mem_511_sv2v_reg ;
  assign \nz.mem [510] = \nz.mem_510_sv2v_reg ;
  assign \nz.mem [509] = \nz.mem_509_sv2v_reg ;
  assign \nz.mem [508] = \nz.mem_508_sv2v_reg ;
  assign \nz.mem [507] = \nz.mem_507_sv2v_reg ;
  assign \nz.mem [506] = \nz.mem_506_sv2v_reg ;
  assign \nz.mem [505] = \nz.mem_505_sv2v_reg ;
  assign \nz.mem [504] = \nz.mem_504_sv2v_reg ;
  assign \nz.mem [503] = \nz.mem_503_sv2v_reg ;
  assign \nz.mem [502] = \nz.mem_502_sv2v_reg ;
  assign \nz.mem [501] = \nz.mem_501_sv2v_reg ;
  assign \nz.mem [500] = \nz.mem_500_sv2v_reg ;
  assign \nz.mem [499] = \nz.mem_499_sv2v_reg ;
  assign \nz.mem [498] = \nz.mem_498_sv2v_reg ;
  assign \nz.mem [497] = \nz.mem_497_sv2v_reg ;
  assign \nz.mem [496] = \nz.mem_496_sv2v_reg ;
  assign \nz.mem [495] = \nz.mem_495_sv2v_reg ;
  assign \nz.mem [494] = \nz.mem_494_sv2v_reg ;
  assign \nz.mem [493] = \nz.mem_493_sv2v_reg ;
  assign \nz.mem [492] = \nz.mem_492_sv2v_reg ;
  assign \nz.mem [491] = \nz.mem_491_sv2v_reg ;
  assign \nz.mem [490] = \nz.mem_490_sv2v_reg ;
  assign \nz.mem [489] = \nz.mem_489_sv2v_reg ;
  assign \nz.mem [488] = \nz.mem_488_sv2v_reg ;
  assign \nz.mem [487] = \nz.mem_487_sv2v_reg ;
  assign \nz.mem [486] = \nz.mem_486_sv2v_reg ;
  assign \nz.mem [485] = \nz.mem_485_sv2v_reg ;
  assign \nz.mem [484] = \nz.mem_484_sv2v_reg ;
  assign \nz.mem [483] = \nz.mem_483_sv2v_reg ;
  assign \nz.mem [482] = \nz.mem_482_sv2v_reg ;
  assign \nz.mem [481] = \nz.mem_481_sv2v_reg ;
  assign \nz.mem [480] = \nz.mem_480_sv2v_reg ;
  assign \nz.mem [479] = \nz.mem_479_sv2v_reg ;
  assign \nz.mem [478] = \nz.mem_478_sv2v_reg ;
  assign \nz.mem [477] = \nz.mem_477_sv2v_reg ;
  assign \nz.mem [476] = \nz.mem_476_sv2v_reg ;
  assign \nz.mem [475] = \nz.mem_475_sv2v_reg ;
  assign \nz.mem [474] = \nz.mem_474_sv2v_reg ;
  assign \nz.mem [473] = \nz.mem_473_sv2v_reg ;
  assign \nz.mem [472] = \nz.mem_472_sv2v_reg ;
  assign \nz.mem [471] = \nz.mem_471_sv2v_reg ;
  assign \nz.mem [470] = \nz.mem_470_sv2v_reg ;
  assign \nz.mem [469] = \nz.mem_469_sv2v_reg ;
  assign \nz.mem [468] = \nz.mem_468_sv2v_reg ;
  assign \nz.mem [467] = \nz.mem_467_sv2v_reg ;
  assign \nz.mem [466] = \nz.mem_466_sv2v_reg ;
  assign \nz.mem [465] = \nz.mem_465_sv2v_reg ;
  assign \nz.mem [464] = \nz.mem_464_sv2v_reg ;
  assign \nz.mem [463] = \nz.mem_463_sv2v_reg ;
  assign \nz.mem [462] = \nz.mem_462_sv2v_reg ;
  assign \nz.mem [461] = \nz.mem_461_sv2v_reg ;
  assign \nz.mem [460] = \nz.mem_460_sv2v_reg ;
  assign \nz.mem [459] = \nz.mem_459_sv2v_reg ;
  assign \nz.mem [458] = \nz.mem_458_sv2v_reg ;
  assign \nz.mem [457] = \nz.mem_457_sv2v_reg ;
  assign \nz.mem [456] = \nz.mem_456_sv2v_reg ;
  assign \nz.mem [455] = \nz.mem_455_sv2v_reg ;
  assign \nz.mem [454] = \nz.mem_454_sv2v_reg ;
  assign \nz.mem [453] = \nz.mem_453_sv2v_reg ;
  assign \nz.mem [452] = \nz.mem_452_sv2v_reg ;
  assign \nz.mem [451] = \nz.mem_451_sv2v_reg ;
  assign \nz.mem [450] = \nz.mem_450_sv2v_reg ;
  assign \nz.mem [449] = \nz.mem_449_sv2v_reg ;
  assign \nz.mem [448] = \nz.mem_448_sv2v_reg ;
  assign \nz.mem [447] = \nz.mem_447_sv2v_reg ;
  assign \nz.mem [446] = \nz.mem_446_sv2v_reg ;
  assign \nz.mem [445] = \nz.mem_445_sv2v_reg ;
  assign \nz.mem [444] = \nz.mem_444_sv2v_reg ;
  assign \nz.mem [443] = \nz.mem_443_sv2v_reg ;
  assign \nz.mem [442] = \nz.mem_442_sv2v_reg ;
  assign \nz.mem [441] = \nz.mem_441_sv2v_reg ;
  assign \nz.mem [440] = \nz.mem_440_sv2v_reg ;
  assign \nz.mem [439] = \nz.mem_439_sv2v_reg ;
  assign \nz.mem [438] = \nz.mem_438_sv2v_reg ;
  assign \nz.mem [437] = \nz.mem_437_sv2v_reg ;
  assign \nz.mem [436] = \nz.mem_436_sv2v_reg ;
  assign \nz.mem [435] = \nz.mem_435_sv2v_reg ;
  assign \nz.mem [434] = \nz.mem_434_sv2v_reg ;
  assign \nz.mem [433] = \nz.mem_433_sv2v_reg ;
  assign \nz.mem [432] = \nz.mem_432_sv2v_reg ;
  assign \nz.mem [431] = \nz.mem_431_sv2v_reg ;
  assign \nz.mem [430] = \nz.mem_430_sv2v_reg ;
  assign \nz.mem [429] = \nz.mem_429_sv2v_reg ;
  assign \nz.mem [428] = \nz.mem_428_sv2v_reg ;
  assign \nz.mem [427] = \nz.mem_427_sv2v_reg ;
  assign \nz.mem [426] = \nz.mem_426_sv2v_reg ;
  assign \nz.mem [425] = \nz.mem_425_sv2v_reg ;
  assign \nz.mem [424] = \nz.mem_424_sv2v_reg ;
  assign \nz.mem [423] = \nz.mem_423_sv2v_reg ;
  assign \nz.mem [422] = \nz.mem_422_sv2v_reg ;
  assign \nz.mem [421] = \nz.mem_421_sv2v_reg ;
  assign \nz.mem [420] = \nz.mem_420_sv2v_reg ;
  assign \nz.mem [419] = \nz.mem_419_sv2v_reg ;
  assign \nz.mem [418] = \nz.mem_418_sv2v_reg ;
  assign \nz.mem [417] = \nz.mem_417_sv2v_reg ;
  assign \nz.mem [416] = \nz.mem_416_sv2v_reg ;
  assign \nz.mem [415] = \nz.mem_415_sv2v_reg ;
  assign \nz.mem [414] = \nz.mem_414_sv2v_reg ;
  assign \nz.mem [413] = \nz.mem_413_sv2v_reg ;
  assign \nz.mem [412] = \nz.mem_412_sv2v_reg ;
  assign \nz.mem [411] = \nz.mem_411_sv2v_reg ;
  assign \nz.mem [410] = \nz.mem_410_sv2v_reg ;
  assign \nz.mem [409] = \nz.mem_409_sv2v_reg ;
  assign \nz.mem [408] = \nz.mem_408_sv2v_reg ;
  assign \nz.mem [407] = \nz.mem_407_sv2v_reg ;
  assign \nz.mem [406] = \nz.mem_406_sv2v_reg ;
  assign \nz.mem [405] = \nz.mem_405_sv2v_reg ;
  assign \nz.mem [404] = \nz.mem_404_sv2v_reg ;
  assign \nz.mem [403] = \nz.mem_403_sv2v_reg ;
  assign \nz.mem [402] = \nz.mem_402_sv2v_reg ;
  assign \nz.mem [401] = \nz.mem_401_sv2v_reg ;
  assign \nz.mem [400] = \nz.mem_400_sv2v_reg ;
  assign \nz.mem [399] = \nz.mem_399_sv2v_reg ;
  assign \nz.mem [398] = \nz.mem_398_sv2v_reg ;
  assign \nz.mem [397] = \nz.mem_397_sv2v_reg ;
  assign \nz.mem [396] = \nz.mem_396_sv2v_reg ;
  assign \nz.mem [395] = \nz.mem_395_sv2v_reg ;
  assign \nz.mem [394] = \nz.mem_394_sv2v_reg ;
  assign \nz.mem [393] = \nz.mem_393_sv2v_reg ;
  assign \nz.mem [392] = \nz.mem_392_sv2v_reg ;
  assign \nz.mem [391] = \nz.mem_391_sv2v_reg ;
  assign \nz.mem [390] = \nz.mem_390_sv2v_reg ;
  assign \nz.mem [389] = \nz.mem_389_sv2v_reg ;
  assign \nz.mem [388] = \nz.mem_388_sv2v_reg ;
  assign \nz.mem [387] = \nz.mem_387_sv2v_reg ;
  assign \nz.mem [386] = \nz.mem_386_sv2v_reg ;
  assign \nz.mem [385] = \nz.mem_385_sv2v_reg ;
  assign \nz.mem [384] = \nz.mem_384_sv2v_reg ;
  assign \nz.mem [383] = \nz.mem_383_sv2v_reg ;
  assign \nz.mem [382] = \nz.mem_382_sv2v_reg ;
  assign \nz.mem [381] = \nz.mem_381_sv2v_reg ;
  assign \nz.mem [380] = \nz.mem_380_sv2v_reg ;
  assign \nz.mem [379] = \nz.mem_379_sv2v_reg ;
  assign \nz.mem [378] = \nz.mem_378_sv2v_reg ;
  assign \nz.mem [377] = \nz.mem_377_sv2v_reg ;
  assign \nz.mem [376] = \nz.mem_376_sv2v_reg ;
  assign \nz.mem [375] = \nz.mem_375_sv2v_reg ;
  assign \nz.mem [374] = \nz.mem_374_sv2v_reg ;
  assign \nz.mem [373] = \nz.mem_373_sv2v_reg ;
  assign \nz.mem [372] = \nz.mem_372_sv2v_reg ;
  assign \nz.mem [371] = \nz.mem_371_sv2v_reg ;
  assign \nz.mem [370] = \nz.mem_370_sv2v_reg ;
  assign \nz.mem [369] = \nz.mem_369_sv2v_reg ;
  assign \nz.mem [368] = \nz.mem_368_sv2v_reg ;
  assign \nz.mem [367] = \nz.mem_367_sv2v_reg ;
  assign \nz.mem [366] = \nz.mem_366_sv2v_reg ;
  assign \nz.mem [365] = \nz.mem_365_sv2v_reg ;
  assign \nz.mem [364] = \nz.mem_364_sv2v_reg ;
  assign \nz.mem [363] = \nz.mem_363_sv2v_reg ;
  assign \nz.mem [362] = \nz.mem_362_sv2v_reg ;
  assign \nz.mem [361] = \nz.mem_361_sv2v_reg ;
  assign \nz.mem [360] = \nz.mem_360_sv2v_reg ;
  assign \nz.mem [359] = \nz.mem_359_sv2v_reg ;
  assign \nz.mem [358] = \nz.mem_358_sv2v_reg ;
  assign \nz.mem [357] = \nz.mem_357_sv2v_reg ;
  assign \nz.mem [356] = \nz.mem_356_sv2v_reg ;
  assign \nz.mem [355] = \nz.mem_355_sv2v_reg ;
  assign \nz.mem [354] = \nz.mem_354_sv2v_reg ;
  assign \nz.mem [353] = \nz.mem_353_sv2v_reg ;
  assign \nz.mem [352] = \nz.mem_352_sv2v_reg ;
  assign \nz.mem [351] = \nz.mem_351_sv2v_reg ;
  assign \nz.mem [350] = \nz.mem_350_sv2v_reg ;
  assign \nz.mem [349] = \nz.mem_349_sv2v_reg ;
  assign \nz.mem [348] = \nz.mem_348_sv2v_reg ;
  assign \nz.mem [347] = \nz.mem_347_sv2v_reg ;
  assign \nz.mem [346] = \nz.mem_346_sv2v_reg ;
  assign \nz.mem [345] = \nz.mem_345_sv2v_reg ;
  assign \nz.mem [344] = \nz.mem_344_sv2v_reg ;
  assign \nz.mem [343] = \nz.mem_343_sv2v_reg ;
  assign \nz.mem [342] = \nz.mem_342_sv2v_reg ;
  assign \nz.mem [341] = \nz.mem_341_sv2v_reg ;
  assign \nz.mem [340] = \nz.mem_340_sv2v_reg ;
  assign \nz.mem [339] = \nz.mem_339_sv2v_reg ;
  assign \nz.mem [338] = \nz.mem_338_sv2v_reg ;
  assign \nz.mem [337] = \nz.mem_337_sv2v_reg ;
  assign \nz.mem [336] = \nz.mem_336_sv2v_reg ;
  assign \nz.mem [335] = \nz.mem_335_sv2v_reg ;
  assign \nz.mem [334] = \nz.mem_334_sv2v_reg ;
  assign \nz.mem [333] = \nz.mem_333_sv2v_reg ;
  assign \nz.mem [332] = \nz.mem_332_sv2v_reg ;
  assign \nz.mem [331] = \nz.mem_331_sv2v_reg ;
  assign \nz.mem [330] = \nz.mem_330_sv2v_reg ;
  assign \nz.mem [329] = \nz.mem_329_sv2v_reg ;
  assign \nz.mem [328] = \nz.mem_328_sv2v_reg ;
  assign \nz.mem [327] = \nz.mem_327_sv2v_reg ;
  assign \nz.mem [326] = \nz.mem_326_sv2v_reg ;
  assign \nz.mem [325] = \nz.mem_325_sv2v_reg ;
  assign \nz.mem [324] = \nz.mem_324_sv2v_reg ;
  assign \nz.mem [323] = \nz.mem_323_sv2v_reg ;
  assign \nz.mem [322] = \nz.mem_322_sv2v_reg ;
  assign \nz.mem [321] = \nz.mem_321_sv2v_reg ;
  assign \nz.mem [320] = \nz.mem_320_sv2v_reg ;
  assign \nz.mem [319] = \nz.mem_319_sv2v_reg ;
  assign \nz.mem [318] = \nz.mem_318_sv2v_reg ;
  assign \nz.mem [317] = \nz.mem_317_sv2v_reg ;
  assign \nz.mem [316] = \nz.mem_316_sv2v_reg ;
  assign \nz.mem [315] = \nz.mem_315_sv2v_reg ;
  assign \nz.mem [314] = \nz.mem_314_sv2v_reg ;
  assign \nz.mem [313] = \nz.mem_313_sv2v_reg ;
  assign \nz.mem [312] = \nz.mem_312_sv2v_reg ;
  assign \nz.mem [311] = \nz.mem_311_sv2v_reg ;
  assign \nz.mem [310] = \nz.mem_310_sv2v_reg ;
  assign \nz.mem [309] = \nz.mem_309_sv2v_reg ;
  assign \nz.mem [308] = \nz.mem_308_sv2v_reg ;
  assign \nz.mem [307] = \nz.mem_307_sv2v_reg ;
  assign \nz.mem [306] = \nz.mem_306_sv2v_reg ;
  assign \nz.mem [305] = \nz.mem_305_sv2v_reg ;
  assign \nz.mem [304] = \nz.mem_304_sv2v_reg ;
  assign \nz.mem [303] = \nz.mem_303_sv2v_reg ;
  assign \nz.mem [302] = \nz.mem_302_sv2v_reg ;
  assign \nz.mem [301] = \nz.mem_301_sv2v_reg ;
  assign \nz.mem [300] = \nz.mem_300_sv2v_reg ;
  assign \nz.mem [299] = \nz.mem_299_sv2v_reg ;
  assign \nz.mem [298] = \nz.mem_298_sv2v_reg ;
  assign \nz.mem [297] = \nz.mem_297_sv2v_reg ;
  assign \nz.mem [296] = \nz.mem_296_sv2v_reg ;
  assign \nz.mem [295] = \nz.mem_295_sv2v_reg ;
  assign \nz.mem [294] = \nz.mem_294_sv2v_reg ;
  assign \nz.mem [293] = \nz.mem_293_sv2v_reg ;
  assign \nz.mem [292] = \nz.mem_292_sv2v_reg ;
  assign \nz.mem [291] = \nz.mem_291_sv2v_reg ;
  assign \nz.mem [290] = \nz.mem_290_sv2v_reg ;
  assign \nz.mem [289] = \nz.mem_289_sv2v_reg ;
  assign \nz.mem [288] = \nz.mem_288_sv2v_reg ;
  assign \nz.mem [287] = \nz.mem_287_sv2v_reg ;
  assign \nz.mem [286] = \nz.mem_286_sv2v_reg ;
  assign \nz.mem [285] = \nz.mem_285_sv2v_reg ;
  assign \nz.mem [284] = \nz.mem_284_sv2v_reg ;
  assign \nz.mem [283] = \nz.mem_283_sv2v_reg ;
  assign \nz.mem [282] = \nz.mem_282_sv2v_reg ;
  assign \nz.mem [281] = \nz.mem_281_sv2v_reg ;
  assign \nz.mem [280] = \nz.mem_280_sv2v_reg ;
  assign \nz.mem [279] = \nz.mem_279_sv2v_reg ;
  assign \nz.mem [278] = \nz.mem_278_sv2v_reg ;
  assign \nz.mem [277] = \nz.mem_277_sv2v_reg ;
  assign \nz.mem [276] = \nz.mem_276_sv2v_reg ;
  assign \nz.mem [275] = \nz.mem_275_sv2v_reg ;
  assign \nz.mem [274] = \nz.mem_274_sv2v_reg ;
  assign \nz.mem [273] = \nz.mem_273_sv2v_reg ;
  assign \nz.mem [272] = \nz.mem_272_sv2v_reg ;
  assign \nz.mem [271] = \nz.mem_271_sv2v_reg ;
  assign \nz.mem [270] = \nz.mem_270_sv2v_reg ;
  assign \nz.mem [269] = \nz.mem_269_sv2v_reg ;
  assign \nz.mem [268] = \nz.mem_268_sv2v_reg ;
  assign \nz.mem [267] = \nz.mem_267_sv2v_reg ;
  assign \nz.mem [266] = \nz.mem_266_sv2v_reg ;
  assign \nz.mem [265] = \nz.mem_265_sv2v_reg ;
  assign \nz.mem [264] = \nz.mem_264_sv2v_reg ;
  assign \nz.mem [263] = \nz.mem_263_sv2v_reg ;
  assign \nz.mem [262] = \nz.mem_262_sv2v_reg ;
  assign \nz.mem [261] = \nz.mem_261_sv2v_reg ;
  assign \nz.mem [260] = \nz.mem_260_sv2v_reg ;
  assign \nz.mem [259] = \nz.mem_259_sv2v_reg ;
  assign \nz.mem [258] = \nz.mem_258_sv2v_reg ;
  assign \nz.mem [257] = \nz.mem_257_sv2v_reg ;
  assign \nz.mem [256] = \nz.mem_256_sv2v_reg ;
  assign \nz.mem [255] = \nz.mem_255_sv2v_reg ;
  assign \nz.mem [254] = \nz.mem_254_sv2v_reg ;
  assign \nz.mem [253] = \nz.mem_253_sv2v_reg ;
  assign \nz.mem [252] = \nz.mem_252_sv2v_reg ;
  assign \nz.mem [251] = \nz.mem_251_sv2v_reg ;
  assign \nz.mem [250] = \nz.mem_250_sv2v_reg ;
  assign \nz.mem [249] = \nz.mem_249_sv2v_reg ;
  assign \nz.mem [248] = \nz.mem_248_sv2v_reg ;
  assign \nz.mem [247] = \nz.mem_247_sv2v_reg ;
  assign \nz.mem [246] = \nz.mem_246_sv2v_reg ;
  assign \nz.mem [245] = \nz.mem_245_sv2v_reg ;
  assign \nz.mem [244] = \nz.mem_244_sv2v_reg ;
  assign \nz.mem [243] = \nz.mem_243_sv2v_reg ;
  assign \nz.mem [242] = \nz.mem_242_sv2v_reg ;
  assign \nz.mem [241] = \nz.mem_241_sv2v_reg ;
  assign \nz.mem [240] = \nz.mem_240_sv2v_reg ;
  assign \nz.mem [239] = \nz.mem_239_sv2v_reg ;
  assign \nz.mem [238] = \nz.mem_238_sv2v_reg ;
  assign \nz.mem [237] = \nz.mem_237_sv2v_reg ;
  assign \nz.mem [236] = \nz.mem_236_sv2v_reg ;
  assign \nz.mem [235] = \nz.mem_235_sv2v_reg ;
  assign \nz.mem [234] = \nz.mem_234_sv2v_reg ;
  assign \nz.mem [233] = \nz.mem_233_sv2v_reg ;
  assign \nz.mem [232] = \nz.mem_232_sv2v_reg ;
  assign \nz.mem [231] = \nz.mem_231_sv2v_reg ;
  assign \nz.mem [230] = \nz.mem_230_sv2v_reg ;
  assign \nz.mem [229] = \nz.mem_229_sv2v_reg ;
  assign \nz.mem [228] = \nz.mem_228_sv2v_reg ;
  assign \nz.mem [227] = \nz.mem_227_sv2v_reg ;
  assign \nz.mem [226] = \nz.mem_226_sv2v_reg ;
  assign \nz.mem [225] = \nz.mem_225_sv2v_reg ;
  assign \nz.mem [224] = \nz.mem_224_sv2v_reg ;
  assign \nz.mem [223] = \nz.mem_223_sv2v_reg ;
  assign \nz.mem [222] = \nz.mem_222_sv2v_reg ;
  assign \nz.mem [221] = \nz.mem_221_sv2v_reg ;
  assign \nz.mem [220] = \nz.mem_220_sv2v_reg ;
  assign \nz.mem [219] = \nz.mem_219_sv2v_reg ;
  assign \nz.mem [218] = \nz.mem_218_sv2v_reg ;
  assign \nz.mem [217] = \nz.mem_217_sv2v_reg ;
  assign \nz.mem [216] = \nz.mem_216_sv2v_reg ;
  assign \nz.mem [215] = \nz.mem_215_sv2v_reg ;
  assign \nz.mem [214] = \nz.mem_214_sv2v_reg ;
  assign \nz.mem [213] = \nz.mem_213_sv2v_reg ;
  assign \nz.mem [212] = \nz.mem_212_sv2v_reg ;
  assign \nz.mem [211] = \nz.mem_211_sv2v_reg ;
  assign \nz.mem [210] = \nz.mem_210_sv2v_reg ;
  assign \nz.mem [209] = \nz.mem_209_sv2v_reg ;
  assign \nz.mem [208] = \nz.mem_208_sv2v_reg ;
  assign \nz.mem [207] = \nz.mem_207_sv2v_reg ;
  assign \nz.mem [206] = \nz.mem_206_sv2v_reg ;
  assign \nz.mem [205] = \nz.mem_205_sv2v_reg ;
  assign \nz.mem [204] = \nz.mem_204_sv2v_reg ;
  assign \nz.mem [203] = \nz.mem_203_sv2v_reg ;
  assign \nz.mem [202] = \nz.mem_202_sv2v_reg ;
  assign \nz.mem [201] = \nz.mem_201_sv2v_reg ;
  assign \nz.mem [200] = \nz.mem_200_sv2v_reg ;
  assign \nz.mem [199] = \nz.mem_199_sv2v_reg ;
  assign \nz.mem [198] = \nz.mem_198_sv2v_reg ;
  assign \nz.mem [197] = \nz.mem_197_sv2v_reg ;
  assign \nz.mem [196] = \nz.mem_196_sv2v_reg ;
  assign \nz.mem [195] = \nz.mem_195_sv2v_reg ;
  assign \nz.mem [194] = \nz.mem_194_sv2v_reg ;
  assign \nz.mem [193] = \nz.mem_193_sv2v_reg ;
  assign \nz.mem [192] = \nz.mem_192_sv2v_reg ;
  assign \nz.mem [191] = \nz.mem_191_sv2v_reg ;
  assign \nz.mem [190] = \nz.mem_190_sv2v_reg ;
  assign \nz.mem [189] = \nz.mem_189_sv2v_reg ;
  assign \nz.mem [188] = \nz.mem_188_sv2v_reg ;
  assign \nz.mem [187] = \nz.mem_187_sv2v_reg ;
  assign \nz.mem [186] = \nz.mem_186_sv2v_reg ;
  assign \nz.mem [185] = \nz.mem_185_sv2v_reg ;
  assign \nz.mem [184] = \nz.mem_184_sv2v_reg ;
  assign \nz.mem [183] = \nz.mem_183_sv2v_reg ;
  assign \nz.mem [182] = \nz.mem_182_sv2v_reg ;
  assign \nz.mem [181] = \nz.mem_181_sv2v_reg ;
  assign \nz.mem [180] = \nz.mem_180_sv2v_reg ;
  assign \nz.mem [179] = \nz.mem_179_sv2v_reg ;
  assign \nz.mem [178] = \nz.mem_178_sv2v_reg ;
  assign \nz.mem [177] = \nz.mem_177_sv2v_reg ;
  assign \nz.mem [176] = \nz.mem_176_sv2v_reg ;
  assign \nz.mem [175] = \nz.mem_175_sv2v_reg ;
  assign \nz.mem [174] = \nz.mem_174_sv2v_reg ;
  assign \nz.mem [173] = \nz.mem_173_sv2v_reg ;
  assign \nz.mem [172] = \nz.mem_172_sv2v_reg ;
  assign \nz.mem [171] = \nz.mem_171_sv2v_reg ;
  assign \nz.mem [170] = \nz.mem_170_sv2v_reg ;
  assign \nz.mem [169] = \nz.mem_169_sv2v_reg ;
  assign \nz.mem [168] = \nz.mem_168_sv2v_reg ;
  assign \nz.mem [167] = \nz.mem_167_sv2v_reg ;
  assign \nz.mem [166] = \nz.mem_166_sv2v_reg ;
  assign \nz.mem [165] = \nz.mem_165_sv2v_reg ;
  assign \nz.mem [164] = \nz.mem_164_sv2v_reg ;
  assign \nz.mem [163] = \nz.mem_163_sv2v_reg ;
  assign \nz.mem [162] = \nz.mem_162_sv2v_reg ;
  assign \nz.mem [161] = \nz.mem_161_sv2v_reg ;
  assign \nz.mem [160] = \nz.mem_160_sv2v_reg ;
  assign \nz.mem [159] = \nz.mem_159_sv2v_reg ;
  assign \nz.mem [158] = \nz.mem_158_sv2v_reg ;
  assign \nz.mem [157] = \nz.mem_157_sv2v_reg ;
  assign \nz.mem [156] = \nz.mem_156_sv2v_reg ;
  assign \nz.mem [155] = \nz.mem_155_sv2v_reg ;
  assign \nz.mem [154] = \nz.mem_154_sv2v_reg ;
  assign \nz.mem [153] = \nz.mem_153_sv2v_reg ;
  assign \nz.mem [152] = \nz.mem_152_sv2v_reg ;
  assign \nz.mem [151] = \nz.mem_151_sv2v_reg ;
  assign \nz.mem [150] = \nz.mem_150_sv2v_reg ;
  assign \nz.mem [149] = \nz.mem_149_sv2v_reg ;
  assign \nz.mem [148] = \nz.mem_148_sv2v_reg ;
  assign \nz.mem [147] = \nz.mem_147_sv2v_reg ;
  assign \nz.mem [146] = \nz.mem_146_sv2v_reg ;
  assign \nz.mem [145] = \nz.mem_145_sv2v_reg ;
  assign \nz.mem [144] = \nz.mem_144_sv2v_reg ;
  assign \nz.mem [143] = \nz.mem_143_sv2v_reg ;
  assign \nz.mem [142] = \nz.mem_142_sv2v_reg ;
  assign \nz.mem [141] = \nz.mem_141_sv2v_reg ;
  assign \nz.mem [140] = \nz.mem_140_sv2v_reg ;
  assign \nz.mem [139] = \nz.mem_139_sv2v_reg ;
  assign \nz.mem [138] = \nz.mem_138_sv2v_reg ;
  assign \nz.mem [137] = \nz.mem_137_sv2v_reg ;
  assign \nz.mem [136] = \nz.mem_136_sv2v_reg ;
  assign \nz.mem [135] = \nz.mem_135_sv2v_reg ;
  assign \nz.mem [134] = \nz.mem_134_sv2v_reg ;
  assign \nz.mem [133] = \nz.mem_133_sv2v_reg ;
  assign \nz.mem [132] = \nz.mem_132_sv2v_reg ;
  assign \nz.mem [131] = \nz.mem_131_sv2v_reg ;
  assign \nz.mem [130] = \nz.mem_130_sv2v_reg ;
  assign \nz.mem [129] = \nz.mem_129_sv2v_reg ;
  assign \nz.mem [128] = \nz.mem_128_sv2v_reg ;
  assign \nz.mem [127] = \nz.mem_127_sv2v_reg ;
  assign \nz.mem [126] = \nz.mem_126_sv2v_reg ;
  assign \nz.mem [125] = \nz.mem_125_sv2v_reg ;
  assign \nz.mem [124] = \nz.mem_124_sv2v_reg ;
  assign \nz.mem [123] = \nz.mem_123_sv2v_reg ;
  assign \nz.mem [122] = \nz.mem_122_sv2v_reg ;
  assign \nz.mem [121] = \nz.mem_121_sv2v_reg ;
  assign \nz.mem [120] = \nz.mem_120_sv2v_reg ;
  assign \nz.mem [119] = \nz.mem_119_sv2v_reg ;
  assign \nz.mem [118] = \nz.mem_118_sv2v_reg ;
  assign \nz.mem [117] = \nz.mem_117_sv2v_reg ;
  assign \nz.mem [116] = \nz.mem_116_sv2v_reg ;
  assign \nz.mem [115] = \nz.mem_115_sv2v_reg ;
  assign \nz.mem [114] = \nz.mem_114_sv2v_reg ;
  assign \nz.mem [113] = \nz.mem_113_sv2v_reg ;
  assign \nz.mem [112] = \nz.mem_112_sv2v_reg ;
  assign \nz.mem [111] = \nz.mem_111_sv2v_reg ;
  assign \nz.mem [110] = \nz.mem_110_sv2v_reg ;
  assign \nz.mem [109] = \nz.mem_109_sv2v_reg ;
  assign \nz.mem [108] = \nz.mem_108_sv2v_reg ;
  assign \nz.mem [107] = \nz.mem_107_sv2v_reg ;
  assign \nz.mem [106] = \nz.mem_106_sv2v_reg ;
  assign \nz.mem [105] = \nz.mem_105_sv2v_reg ;
  assign \nz.mem [104] = \nz.mem_104_sv2v_reg ;
  assign \nz.mem [103] = \nz.mem_103_sv2v_reg ;
  assign \nz.mem [102] = \nz.mem_102_sv2v_reg ;
  assign \nz.mem [101] = \nz.mem_101_sv2v_reg ;
  assign \nz.mem [100] = \nz.mem_100_sv2v_reg ;
  assign \nz.mem [99] = \nz.mem_99_sv2v_reg ;
  assign \nz.mem [98] = \nz.mem_98_sv2v_reg ;
  assign \nz.mem [97] = \nz.mem_97_sv2v_reg ;
  assign \nz.mem [96] = \nz.mem_96_sv2v_reg ;
  assign \nz.mem [95] = \nz.mem_95_sv2v_reg ;
  assign \nz.mem [94] = \nz.mem_94_sv2v_reg ;
  assign \nz.mem [93] = \nz.mem_93_sv2v_reg ;
  assign \nz.mem [92] = \nz.mem_92_sv2v_reg ;
  assign \nz.mem [91] = \nz.mem_91_sv2v_reg ;
  assign \nz.mem [90] = \nz.mem_90_sv2v_reg ;
  assign \nz.mem [89] = \nz.mem_89_sv2v_reg ;
  assign \nz.mem [88] = \nz.mem_88_sv2v_reg ;
  assign \nz.mem [87] = \nz.mem_87_sv2v_reg ;
  assign \nz.mem [86] = \nz.mem_86_sv2v_reg ;
  assign \nz.mem [85] = \nz.mem_85_sv2v_reg ;
  assign \nz.mem [84] = \nz.mem_84_sv2v_reg ;
  assign \nz.mem [83] = \nz.mem_83_sv2v_reg ;
  assign \nz.mem [82] = \nz.mem_82_sv2v_reg ;
  assign \nz.mem [81] = \nz.mem_81_sv2v_reg ;
  assign \nz.mem [80] = \nz.mem_80_sv2v_reg ;
  assign \nz.mem [79] = \nz.mem_79_sv2v_reg ;
  assign \nz.mem [78] = \nz.mem_78_sv2v_reg ;
  assign \nz.mem [77] = \nz.mem_77_sv2v_reg ;
  assign \nz.mem [76] = \nz.mem_76_sv2v_reg ;
  assign \nz.mem [75] = \nz.mem_75_sv2v_reg ;
  assign \nz.mem [74] = \nz.mem_74_sv2v_reg ;
  assign \nz.mem [73] = \nz.mem_73_sv2v_reg ;
  assign \nz.mem [72] = \nz.mem_72_sv2v_reg ;
  assign \nz.mem [71] = \nz.mem_71_sv2v_reg ;
  assign \nz.mem [70] = \nz.mem_70_sv2v_reg ;
  assign \nz.mem [69] = \nz.mem_69_sv2v_reg ;
  assign \nz.mem [68] = \nz.mem_68_sv2v_reg ;
  assign \nz.mem [67] = \nz.mem_67_sv2v_reg ;
  assign \nz.mem [66] = \nz.mem_66_sv2v_reg ;
  assign \nz.mem [65] = \nz.mem_65_sv2v_reg ;
  assign \nz.mem [64] = \nz.mem_64_sv2v_reg ;
  assign \nz.mem [63] = \nz.mem_63_sv2v_reg ;
  assign \nz.mem [62] = \nz.mem_62_sv2v_reg ;
  assign \nz.mem [61] = \nz.mem_61_sv2v_reg ;
  assign \nz.mem [60] = \nz.mem_60_sv2v_reg ;
  assign \nz.mem [59] = \nz.mem_59_sv2v_reg ;
  assign \nz.mem [58] = \nz.mem_58_sv2v_reg ;
  assign \nz.mem [57] = \nz.mem_57_sv2v_reg ;
  assign \nz.mem [56] = \nz.mem_56_sv2v_reg ;
  assign \nz.mem [55] = \nz.mem_55_sv2v_reg ;
  assign \nz.mem [54] = \nz.mem_54_sv2v_reg ;
  assign \nz.mem [53] = \nz.mem_53_sv2v_reg ;
  assign \nz.mem [52] = \nz.mem_52_sv2v_reg ;
  assign \nz.mem [51] = \nz.mem_51_sv2v_reg ;
  assign \nz.mem [50] = \nz.mem_50_sv2v_reg ;
  assign \nz.mem [49] = \nz.mem_49_sv2v_reg ;
  assign \nz.mem [48] = \nz.mem_48_sv2v_reg ;
  assign \nz.mem [47] = \nz.mem_47_sv2v_reg ;
  assign \nz.mem [46] = \nz.mem_46_sv2v_reg ;
  assign \nz.mem [45] = \nz.mem_45_sv2v_reg ;
  assign \nz.mem [44] = \nz.mem_44_sv2v_reg ;
  assign \nz.mem [43] = \nz.mem_43_sv2v_reg ;
  assign \nz.mem [42] = \nz.mem_42_sv2v_reg ;
  assign \nz.mem [41] = \nz.mem_41_sv2v_reg ;
  assign \nz.mem [40] = \nz.mem_40_sv2v_reg ;
  assign \nz.mem [39] = \nz.mem_39_sv2v_reg ;
  assign \nz.mem [38] = \nz.mem_38_sv2v_reg ;
  assign \nz.mem [37] = \nz.mem_37_sv2v_reg ;
  assign \nz.mem [36] = \nz.mem_36_sv2v_reg ;
  assign \nz.mem [35] = \nz.mem_35_sv2v_reg ;
  assign \nz.mem [34] = \nz.mem_34_sv2v_reg ;
  assign \nz.mem [33] = \nz.mem_33_sv2v_reg ;
  assign \nz.mem [32] = \nz.mem_32_sv2v_reg ;
  assign \nz.mem [31] = \nz.mem_31_sv2v_reg ;
  assign \nz.mem [30] = \nz.mem_30_sv2v_reg ;
  assign \nz.mem [29] = \nz.mem_29_sv2v_reg ;
  assign \nz.mem [28] = \nz.mem_28_sv2v_reg ;
  assign \nz.mem [27] = \nz.mem_27_sv2v_reg ;
  assign \nz.mem [26] = \nz.mem_26_sv2v_reg ;
  assign \nz.mem [25] = \nz.mem_25_sv2v_reg ;
  assign \nz.mem [24] = \nz.mem_24_sv2v_reg ;
  assign \nz.mem [23] = \nz.mem_23_sv2v_reg ;
  assign \nz.mem [22] = \nz.mem_22_sv2v_reg ;
  assign \nz.mem [21] = \nz.mem_21_sv2v_reg ;
  assign \nz.mem [20] = \nz.mem_20_sv2v_reg ;
  assign \nz.mem [19] = \nz.mem_19_sv2v_reg ;
  assign \nz.mem [18] = \nz.mem_18_sv2v_reg ;
  assign \nz.mem [17] = \nz.mem_17_sv2v_reg ;
  assign \nz.mem [16] = \nz.mem_16_sv2v_reg ;
  assign \nz.mem [15] = \nz.mem_15_sv2v_reg ;
  assign \nz.mem [14] = \nz.mem_14_sv2v_reg ;
  assign \nz.mem [13] = \nz.mem_13_sv2v_reg ;
  assign \nz.mem [12] = \nz.mem_12_sv2v_reg ;
  assign \nz.mem [11] = \nz.mem_11_sv2v_reg ;
  assign \nz.mem [10] = \nz.mem_10_sv2v_reg ;
  assign \nz.mem [9] = \nz.mem_9_sv2v_reg ;
  assign \nz.mem [8] = \nz.mem_8_sv2v_reg ;
  assign \nz.mem [7] = \nz.mem_7_sv2v_reg ;
  assign \nz.mem [6] = \nz.mem_6_sv2v_reg ;
  assign \nz.mem [5] = \nz.mem_5_sv2v_reg ;
  assign \nz.mem [4] = \nz.mem_4_sv2v_reg ;
  assign \nz.mem [3] = \nz.mem_3_sv2v_reg ;
  assign \nz.mem [2] = \nz.mem_2_sv2v_reg ;
  assign \nz.mem [1] = \nz.mem_1_sv2v_reg ;
  assign \nz.mem [0] = \nz.mem_0_sv2v_reg ;
  assign r_data_o[49] = (N76)? \nz.mem [49] : 
                        (N78)? \nz.mem [99] : 
                        (N80)? \nz.mem [149] : 
                        (N82)? \nz.mem [199] : 
                        (N84)? \nz.mem [249] : 
                        (N86)? \nz.mem [299] : 
                        (N88)? \nz.mem [349] : 
                        (N90)? \nz.mem [399] : 
                        (N92)? \nz.mem [449] : 
                        (N94)? \nz.mem [499] : 
                        (N96)? \nz.mem [549] : 
                        (N98)? \nz.mem [599] : 
                        (N100)? \nz.mem [649] : 
                        (N102)? \nz.mem [699] : 
                        (N104)? \nz.mem [749] : 
                        (N106)? \nz.mem [799] : 
                        (N108)? \nz.mem [849] : 
                        (N110)? \nz.mem [899] : 
                        (N112)? \nz.mem [949] : 
                        (N114)? \nz.mem [999] : 
                        (N116)? \nz.mem [1049] : 
                        (N118)? \nz.mem [1099] : 
                        (N120)? \nz.mem [1149] : 
                        (N122)? \nz.mem [1199] : 
                        (N124)? \nz.mem [1249] : 
                        (N126)? \nz.mem [1299] : 
                        (N128)? \nz.mem [1349] : 
                        (N130)? \nz.mem [1399] : 
                        (N132)? \nz.mem [1449] : 
                        (N134)? \nz.mem [1499] : 
                        (N136)? \nz.mem [1549] : 
                        (N138)? \nz.mem [1599] : 
                        (N77)? \nz.mem [1649] : 
                        (N79)? \nz.mem [1699] : 
                        (N81)? \nz.mem [1749] : 
                        (N83)? \nz.mem [1799] : 
                        (N85)? \nz.mem [1849] : 
                        (N87)? \nz.mem [1899] : 
                        (N89)? \nz.mem [1949] : 
                        (N91)? \nz.mem [1999] : 
                        (N93)? \nz.mem [2049] : 
                        (N95)? \nz.mem [2099] : 
                        (N97)? \nz.mem [2149] : 
                        (N99)? \nz.mem [2199] : 
                        (N101)? \nz.mem [2249] : 
                        (N103)? \nz.mem [2299] : 
                        (N105)? \nz.mem [2349] : 
                        (N107)? \nz.mem [2399] : 
                        (N109)? \nz.mem [2449] : 
                        (N111)? \nz.mem [2499] : 
                        (N113)? \nz.mem [2549] : 
                        (N115)? \nz.mem [2599] : 
                        (N117)? \nz.mem [2649] : 
                        (N119)? \nz.mem [2699] : 
                        (N121)? \nz.mem [2749] : 
                        (N123)? \nz.mem [2799] : 
                        (N125)? \nz.mem [2849] : 
                        (N127)? \nz.mem [2899] : 
                        (N129)? \nz.mem [2949] : 
                        (N131)? \nz.mem [2999] : 
                        (N133)? \nz.mem [3049] : 
                        (N135)? \nz.mem [3099] : 
                        (N137)? \nz.mem [3149] : 
                        (N139)? \nz.mem [3199] : 1'b0;
  assign r_data_o[48] = (N76)? \nz.mem [48] : 
                        (N78)? \nz.mem [98] : 
                        (N80)? \nz.mem [148] : 
                        (N82)? \nz.mem [198] : 
                        (N84)? \nz.mem [248] : 
                        (N86)? \nz.mem [298] : 
                        (N88)? \nz.mem [348] : 
                        (N90)? \nz.mem [398] : 
                        (N92)? \nz.mem [448] : 
                        (N94)? \nz.mem [498] : 
                        (N96)? \nz.mem [548] : 
                        (N98)? \nz.mem [598] : 
                        (N100)? \nz.mem [648] : 
                        (N102)? \nz.mem [698] : 
                        (N104)? \nz.mem [748] : 
                        (N106)? \nz.mem [798] : 
                        (N108)? \nz.mem [848] : 
                        (N110)? \nz.mem [898] : 
                        (N112)? \nz.mem [948] : 
                        (N114)? \nz.mem [998] : 
                        (N116)? \nz.mem [1048] : 
                        (N118)? \nz.mem [1098] : 
                        (N120)? \nz.mem [1148] : 
                        (N122)? \nz.mem [1198] : 
                        (N124)? \nz.mem [1248] : 
                        (N126)? \nz.mem [1298] : 
                        (N128)? \nz.mem [1348] : 
                        (N130)? \nz.mem [1398] : 
                        (N132)? \nz.mem [1448] : 
                        (N134)? \nz.mem [1498] : 
                        (N136)? \nz.mem [1548] : 
                        (N138)? \nz.mem [1598] : 
                        (N77)? \nz.mem [1648] : 
                        (N79)? \nz.mem [1698] : 
                        (N81)? \nz.mem [1748] : 
                        (N83)? \nz.mem [1798] : 
                        (N85)? \nz.mem [1848] : 
                        (N87)? \nz.mem [1898] : 
                        (N89)? \nz.mem [1948] : 
                        (N91)? \nz.mem [1998] : 
                        (N93)? \nz.mem [2048] : 
                        (N95)? \nz.mem [2098] : 
                        (N97)? \nz.mem [2148] : 
                        (N99)? \nz.mem [2198] : 
                        (N101)? \nz.mem [2248] : 
                        (N103)? \nz.mem [2298] : 
                        (N105)? \nz.mem [2348] : 
                        (N107)? \nz.mem [2398] : 
                        (N109)? \nz.mem [2448] : 
                        (N111)? \nz.mem [2498] : 
                        (N113)? \nz.mem [2548] : 
                        (N115)? \nz.mem [2598] : 
                        (N117)? \nz.mem [2648] : 
                        (N119)? \nz.mem [2698] : 
                        (N121)? \nz.mem [2748] : 
                        (N123)? \nz.mem [2798] : 
                        (N125)? \nz.mem [2848] : 
                        (N127)? \nz.mem [2898] : 
                        (N129)? \nz.mem [2948] : 
                        (N131)? \nz.mem [2998] : 
                        (N133)? \nz.mem [3048] : 
                        (N135)? \nz.mem [3098] : 
                        (N137)? \nz.mem [3148] : 
                        (N139)? \nz.mem [3198] : 1'b0;
  assign r_data_o[47] = (N76)? \nz.mem [47] : 
                        (N78)? \nz.mem [97] : 
                        (N80)? \nz.mem [147] : 
                        (N82)? \nz.mem [197] : 
                        (N84)? \nz.mem [247] : 
                        (N86)? \nz.mem [297] : 
                        (N88)? \nz.mem [347] : 
                        (N90)? \nz.mem [397] : 
                        (N92)? \nz.mem [447] : 
                        (N94)? \nz.mem [497] : 
                        (N96)? \nz.mem [547] : 
                        (N98)? \nz.mem [597] : 
                        (N100)? \nz.mem [647] : 
                        (N102)? \nz.mem [697] : 
                        (N104)? \nz.mem [747] : 
                        (N106)? \nz.mem [797] : 
                        (N108)? \nz.mem [847] : 
                        (N110)? \nz.mem [897] : 
                        (N112)? \nz.mem [947] : 
                        (N114)? \nz.mem [997] : 
                        (N116)? \nz.mem [1047] : 
                        (N118)? \nz.mem [1097] : 
                        (N120)? \nz.mem [1147] : 
                        (N122)? \nz.mem [1197] : 
                        (N124)? \nz.mem [1247] : 
                        (N126)? \nz.mem [1297] : 
                        (N128)? \nz.mem [1347] : 
                        (N130)? \nz.mem [1397] : 
                        (N132)? \nz.mem [1447] : 
                        (N134)? \nz.mem [1497] : 
                        (N136)? \nz.mem [1547] : 
                        (N138)? \nz.mem [1597] : 
                        (N77)? \nz.mem [1647] : 
                        (N79)? \nz.mem [1697] : 
                        (N81)? \nz.mem [1747] : 
                        (N83)? \nz.mem [1797] : 
                        (N85)? \nz.mem [1847] : 
                        (N87)? \nz.mem [1897] : 
                        (N89)? \nz.mem [1947] : 
                        (N91)? \nz.mem [1997] : 
                        (N93)? \nz.mem [2047] : 
                        (N95)? \nz.mem [2097] : 
                        (N97)? \nz.mem [2147] : 
                        (N99)? \nz.mem [2197] : 
                        (N101)? \nz.mem [2247] : 
                        (N103)? \nz.mem [2297] : 
                        (N105)? \nz.mem [2347] : 
                        (N107)? \nz.mem [2397] : 
                        (N109)? \nz.mem [2447] : 
                        (N111)? \nz.mem [2497] : 
                        (N113)? \nz.mem [2547] : 
                        (N115)? \nz.mem [2597] : 
                        (N117)? \nz.mem [2647] : 
                        (N119)? \nz.mem [2697] : 
                        (N121)? \nz.mem [2747] : 
                        (N123)? \nz.mem [2797] : 
                        (N125)? \nz.mem [2847] : 
                        (N127)? \nz.mem [2897] : 
                        (N129)? \nz.mem [2947] : 
                        (N131)? \nz.mem [2997] : 
                        (N133)? \nz.mem [3047] : 
                        (N135)? \nz.mem [3097] : 
                        (N137)? \nz.mem [3147] : 
                        (N139)? \nz.mem [3197] : 1'b0;
  assign r_data_o[46] = (N76)? \nz.mem [46] : 
                        (N78)? \nz.mem [96] : 
                        (N80)? \nz.mem [146] : 
                        (N82)? \nz.mem [196] : 
                        (N84)? \nz.mem [246] : 
                        (N86)? \nz.mem [296] : 
                        (N88)? \nz.mem [346] : 
                        (N90)? \nz.mem [396] : 
                        (N92)? \nz.mem [446] : 
                        (N94)? \nz.mem [496] : 
                        (N96)? \nz.mem [546] : 
                        (N98)? \nz.mem [596] : 
                        (N100)? \nz.mem [646] : 
                        (N102)? \nz.mem [696] : 
                        (N104)? \nz.mem [746] : 
                        (N106)? \nz.mem [796] : 
                        (N108)? \nz.mem [846] : 
                        (N110)? \nz.mem [896] : 
                        (N112)? \nz.mem [946] : 
                        (N114)? \nz.mem [996] : 
                        (N116)? \nz.mem [1046] : 
                        (N118)? \nz.mem [1096] : 
                        (N120)? \nz.mem [1146] : 
                        (N122)? \nz.mem [1196] : 
                        (N124)? \nz.mem [1246] : 
                        (N126)? \nz.mem [1296] : 
                        (N128)? \nz.mem [1346] : 
                        (N130)? \nz.mem [1396] : 
                        (N132)? \nz.mem [1446] : 
                        (N134)? \nz.mem [1496] : 
                        (N136)? \nz.mem [1546] : 
                        (N138)? \nz.mem [1596] : 
                        (N77)? \nz.mem [1646] : 
                        (N79)? \nz.mem [1696] : 
                        (N81)? \nz.mem [1746] : 
                        (N83)? \nz.mem [1796] : 
                        (N85)? \nz.mem [1846] : 
                        (N87)? \nz.mem [1896] : 
                        (N89)? \nz.mem [1946] : 
                        (N91)? \nz.mem [1996] : 
                        (N93)? \nz.mem [2046] : 
                        (N95)? \nz.mem [2096] : 
                        (N97)? \nz.mem [2146] : 
                        (N99)? \nz.mem [2196] : 
                        (N101)? \nz.mem [2246] : 
                        (N103)? \nz.mem [2296] : 
                        (N105)? \nz.mem [2346] : 
                        (N107)? \nz.mem [2396] : 
                        (N109)? \nz.mem [2446] : 
                        (N111)? \nz.mem [2496] : 
                        (N113)? \nz.mem [2546] : 
                        (N115)? \nz.mem [2596] : 
                        (N117)? \nz.mem [2646] : 
                        (N119)? \nz.mem [2696] : 
                        (N121)? \nz.mem [2746] : 
                        (N123)? \nz.mem [2796] : 
                        (N125)? \nz.mem [2846] : 
                        (N127)? \nz.mem [2896] : 
                        (N129)? \nz.mem [2946] : 
                        (N131)? \nz.mem [2996] : 
                        (N133)? \nz.mem [3046] : 
                        (N135)? \nz.mem [3096] : 
                        (N137)? \nz.mem [3146] : 
                        (N139)? \nz.mem [3196] : 1'b0;
  assign r_data_o[45] = (N76)? \nz.mem [45] : 
                        (N78)? \nz.mem [95] : 
                        (N80)? \nz.mem [145] : 
                        (N82)? \nz.mem [195] : 
                        (N84)? \nz.mem [245] : 
                        (N86)? \nz.mem [295] : 
                        (N88)? \nz.mem [345] : 
                        (N90)? \nz.mem [395] : 
                        (N92)? \nz.mem [445] : 
                        (N94)? \nz.mem [495] : 
                        (N96)? \nz.mem [545] : 
                        (N98)? \nz.mem [595] : 
                        (N100)? \nz.mem [645] : 
                        (N102)? \nz.mem [695] : 
                        (N104)? \nz.mem [745] : 
                        (N106)? \nz.mem [795] : 
                        (N108)? \nz.mem [845] : 
                        (N110)? \nz.mem [895] : 
                        (N112)? \nz.mem [945] : 
                        (N114)? \nz.mem [995] : 
                        (N116)? \nz.mem [1045] : 
                        (N118)? \nz.mem [1095] : 
                        (N120)? \nz.mem [1145] : 
                        (N122)? \nz.mem [1195] : 
                        (N124)? \nz.mem [1245] : 
                        (N126)? \nz.mem [1295] : 
                        (N128)? \nz.mem [1345] : 
                        (N130)? \nz.mem [1395] : 
                        (N132)? \nz.mem [1445] : 
                        (N134)? \nz.mem [1495] : 
                        (N136)? \nz.mem [1545] : 
                        (N138)? \nz.mem [1595] : 
                        (N77)? \nz.mem [1645] : 
                        (N79)? \nz.mem [1695] : 
                        (N81)? \nz.mem [1745] : 
                        (N83)? \nz.mem [1795] : 
                        (N85)? \nz.mem [1845] : 
                        (N87)? \nz.mem [1895] : 
                        (N89)? \nz.mem [1945] : 
                        (N91)? \nz.mem [1995] : 
                        (N93)? \nz.mem [2045] : 
                        (N95)? \nz.mem [2095] : 
                        (N97)? \nz.mem [2145] : 
                        (N99)? \nz.mem [2195] : 
                        (N101)? \nz.mem [2245] : 
                        (N103)? \nz.mem [2295] : 
                        (N105)? \nz.mem [2345] : 
                        (N107)? \nz.mem [2395] : 
                        (N109)? \nz.mem [2445] : 
                        (N111)? \nz.mem [2495] : 
                        (N113)? \nz.mem [2545] : 
                        (N115)? \nz.mem [2595] : 
                        (N117)? \nz.mem [2645] : 
                        (N119)? \nz.mem [2695] : 
                        (N121)? \nz.mem [2745] : 
                        (N123)? \nz.mem [2795] : 
                        (N125)? \nz.mem [2845] : 
                        (N127)? \nz.mem [2895] : 
                        (N129)? \nz.mem [2945] : 
                        (N131)? \nz.mem [2995] : 
                        (N133)? \nz.mem [3045] : 
                        (N135)? \nz.mem [3095] : 
                        (N137)? \nz.mem [3145] : 
                        (N139)? \nz.mem [3195] : 1'b0;
  assign r_data_o[44] = (N76)? \nz.mem [44] : 
                        (N78)? \nz.mem [94] : 
                        (N80)? \nz.mem [144] : 
                        (N82)? \nz.mem [194] : 
                        (N84)? \nz.mem [244] : 
                        (N86)? \nz.mem [294] : 
                        (N88)? \nz.mem [344] : 
                        (N90)? \nz.mem [394] : 
                        (N92)? \nz.mem [444] : 
                        (N94)? \nz.mem [494] : 
                        (N96)? \nz.mem [544] : 
                        (N98)? \nz.mem [594] : 
                        (N100)? \nz.mem [644] : 
                        (N102)? \nz.mem [694] : 
                        (N104)? \nz.mem [744] : 
                        (N106)? \nz.mem [794] : 
                        (N108)? \nz.mem [844] : 
                        (N110)? \nz.mem [894] : 
                        (N112)? \nz.mem [944] : 
                        (N114)? \nz.mem [994] : 
                        (N116)? \nz.mem [1044] : 
                        (N118)? \nz.mem [1094] : 
                        (N120)? \nz.mem [1144] : 
                        (N122)? \nz.mem [1194] : 
                        (N124)? \nz.mem [1244] : 
                        (N126)? \nz.mem [1294] : 
                        (N128)? \nz.mem [1344] : 
                        (N130)? \nz.mem [1394] : 
                        (N132)? \nz.mem [1444] : 
                        (N134)? \nz.mem [1494] : 
                        (N136)? \nz.mem [1544] : 
                        (N138)? \nz.mem [1594] : 
                        (N77)? \nz.mem [1644] : 
                        (N79)? \nz.mem [1694] : 
                        (N81)? \nz.mem [1744] : 
                        (N83)? \nz.mem [1794] : 
                        (N85)? \nz.mem [1844] : 
                        (N87)? \nz.mem [1894] : 
                        (N89)? \nz.mem [1944] : 
                        (N91)? \nz.mem [1994] : 
                        (N93)? \nz.mem [2044] : 
                        (N95)? \nz.mem [2094] : 
                        (N97)? \nz.mem [2144] : 
                        (N99)? \nz.mem [2194] : 
                        (N101)? \nz.mem [2244] : 
                        (N103)? \nz.mem [2294] : 
                        (N105)? \nz.mem [2344] : 
                        (N107)? \nz.mem [2394] : 
                        (N109)? \nz.mem [2444] : 
                        (N111)? \nz.mem [2494] : 
                        (N113)? \nz.mem [2544] : 
                        (N115)? \nz.mem [2594] : 
                        (N117)? \nz.mem [2644] : 
                        (N119)? \nz.mem [2694] : 
                        (N121)? \nz.mem [2744] : 
                        (N123)? \nz.mem [2794] : 
                        (N125)? \nz.mem [2844] : 
                        (N127)? \nz.mem [2894] : 
                        (N129)? \nz.mem [2944] : 
                        (N131)? \nz.mem [2994] : 
                        (N133)? \nz.mem [3044] : 
                        (N135)? \nz.mem [3094] : 
                        (N137)? \nz.mem [3144] : 
                        (N139)? \nz.mem [3194] : 1'b0;
  assign r_data_o[43] = (N76)? \nz.mem [43] : 
                        (N78)? \nz.mem [93] : 
                        (N80)? \nz.mem [143] : 
                        (N82)? \nz.mem [193] : 
                        (N84)? \nz.mem [243] : 
                        (N86)? \nz.mem [293] : 
                        (N88)? \nz.mem [343] : 
                        (N90)? \nz.mem [393] : 
                        (N92)? \nz.mem [443] : 
                        (N94)? \nz.mem [493] : 
                        (N96)? \nz.mem [543] : 
                        (N98)? \nz.mem [593] : 
                        (N100)? \nz.mem [643] : 
                        (N102)? \nz.mem [693] : 
                        (N104)? \nz.mem [743] : 
                        (N106)? \nz.mem [793] : 
                        (N108)? \nz.mem [843] : 
                        (N110)? \nz.mem [893] : 
                        (N112)? \nz.mem [943] : 
                        (N114)? \nz.mem [993] : 
                        (N116)? \nz.mem [1043] : 
                        (N118)? \nz.mem [1093] : 
                        (N120)? \nz.mem [1143] : 
                        (N122)? \nz.mem [1193] : 
                        (N124)? \nz.mem [1243] : 
                        (N126)? \nz.mem [1293] : 
                        (N128)? \nz.mem [1343] : 
                        (N130)? \nz.mem [1393] : 
                        (N132)? \nz.mem [1443] : 
                        (N134)? \nz.mem [1493] : 
                        (N136)? \nz.mem [1543] : 
                        (N138)? \nz.mem [1593] : 
                        (N77)? \nz.mem [1643] : 
                        (N79)? \nz.mem [1693] : 
                        (N81)? \nz.mem [1743] : 
                        (N83)? \nz.mem [1793] : 
                        (N85)? \nz.mem [1843] : 
                        (N87)? \nz.mem [1893] : 
                        (N89)? \nz.mem [1943] : 
                        (N91)? \nz.mem [1993] : 
                        (N93)? \nz.mem [2043] : 
                        (N95)? \nz.mem [2093] : 
                        (N97)? \nz.mem [2143] : 
                        (N99)? \nz.mem [2193] : 
                        (N101)? \nz.mem [2243] : 
                        (N103)? \nz.mem [2293] : 
                        (N105)? \nz.mem [2343] : 
                        (N107)? \nz.mem [2393] : 
                        (N109)? \nz.mem [2443] : 
                        (N111)? \nz.mem [2493] : 
                        (N113)? \nz.mem [2543] : 
                        (N115)? \nz.mem [2593] : 
                        (N117)? \nz.mem [2643] : 
                        (N119)? \nz.mem [2693] : 
                        (N121)? \nz.mem [2743] : 
                        (N123)? \nz.mem [2793] : 
                        (N125)? \nz.mem [2843] : 
                        (N127)? \nz.mem [2893] : 
                        (N129)? \nz.mem [2943] : 
                        (N131)? \nz.mem [2993] : 
                        (N133)? \nz.mem [3043] : 
                        (N135)? \nz.mem [3093] : 
                        (N137)? \nz.mem [3143] : 
                        (N139)? \nz.mem [3193] : 1'b0;
  assign r_data_o[42] = (N76)? \nz.mem [42] : 
                        (N78)? \nz.mem [92] : 
                        (N80)? \nz.mem [142] : 
                        (N82)? \nz.mem [192] : 
                        (N84)? \nz.mem [242] : 
                        (N86)? \nz.mem [292] : 
                        (N88)? \nz.mem [342] : 
                        (N90)? \nz.mem [392] : 
                        (N92)? \nz.mem [442] : 
                        (N94)? \nz.mem [492] : 
                        (N96)? \nz.mem [542] : 
                        (N98)? \nz.mem [592] : 
                        (N100)? \nz.mem [642] : 
                        (N102)? \nz.mem [692] : 
                        (N104)? \nz.mem [742] : 
                        (N106)? \nz.mem [792] : 
                        (N108)? \nz.mem [842] : 
                        (N110)? \nz.mem [892] : 
                        (N112)? \nz.mem [942] : 
                        (N114)? \nz.mem [992] : 
                        (N116)? \nz.mem [1042] : 
                        (N118)? \nz.mem [1092] : 
                        (N120)? \nz.mem [1142] : 
                        (N122)? \nz.mem [1192] : 
                        (N124)? \nz.mem [1242] : 
                        (N126)? \nz.mem [1292] : 
                        (N128)? \nz.mem [1342] : 
                        (N130)? \nz.mem [1392] : 
                        (N132)? \nz.mem [1442] : 
                        (N134)? \nz.mem [1492] : 
                        (N136)? \nz.mem [1542] : 
                        (N138)? \nz.mem [1592] : 
                        (N77)? \nz.mem [1642] : 
                        (N79)? \nz.mem [1692] : 
                        (N81)? \nz.mem [1742] : 
                        (N83)? \nz.mem [1792] : 
                        (N85)? \nz.mem [1842] : 
                        (N87)? \nz.mem [1892] : 
                        (N89)? \nz.mem [1942] : 
                        (N91)? \nz.mem [1992] : 
                        (N93)? \nz.mem [2042] : 
                        (N95)? \nz.mem [2092] : 
                        (N97)? \nz.mem [2142] : 
                        (N99)? \nz.mem [2192] : 
                        (N101)? \nz.mem [2242] : 
                        (N103)? \nz.mem [2292] : 
                        (N105)? \nz.mem [2342] : 
                        (N107)? \nz.mem [2392] : 
                        (N109)? \nz.mem [2442] : 
                        (N111)? \nz.mem [2492] : 
                        (N113)? \nz.mem [2542] : 
                        (N115)? \nz.mem [2592] : 
                        (N117)? \nz.mem [2642] : 
                        (N119)? \nz.mem [2692] : 
                        (N121)? \nz.mem [2742] : 
                        (N123)? \nz.mem [2792] : 
                        (N125)? \nz.mem [2842] : 
                        (N127)? \nz.mem [2892] : 
                        (N129)? \nz.mem [2942] : 
                        (N131)? \nz.mem [2992] : 
                        (N133)? \nz.mem [3042] : 
                        (N135)? \nz.mem [3092] : 
                        (N137)? \nz.mem [3142] : 
                        (N139)? \nz.mem [3192] : 1'b0;
  assign r_data_o[41] = (N76)? \nz.mem [41] : 
                        (N78)? \nz.mem [91] : 
                        (N80)? \nz.mem [141] : 
                        (N82)? \nz.mem [191] : 
                        (N84)? \nz.mem [241] : 
                        (N86)? \nz.mem [291] : 
                        (N88)? \nz.mem [341] : 
                        (N90)? \nz.mem [391] : 
                        (N92)? \nz.mem [441] : 
                        (N94)? \nz.mem [491] : 
                        (N96)? \nz.mem [541] : 
                        (N98)? \nz.mem [591] : 
                        (N100)? \nz.mem [641] : 
                        (N102)? \nz.mem [691] : 
                        (N104)? \nz.mem [741] : 
                        (N106)? \nz.mem [791] : 
                        (N108)? \nz.mem [841] : 
                        (N110)? \nz.mem [891] : 
                        (N112)? \nz.mem [941] : 
                        (N114)? \nz.mem [991] : 
                        (N116)? \nz.mem [1041] : 
                        (N118)? \nz.mem [1091] : 
                        (N120)? \nz.mem [1141] : 
                        (N122)? \nz.mem [1191] : 
                        (N124)? \nz.mem [1241] : 
                        (N126)? \nz.mem [1291] : 
                        (N128)? \nz.mem [1341] : 
                        (N130)? \nz.mem [1391] : 
                        (N132)? \nz.mem [1441] : 
                        (N134)? \nz.mem [1491] : 
                        (N136)? \nz.mem [1541] : 
                        (N138)? \nz.mem [1591] : 
                        (N77)? \nz.mem [1641] : 
                        (N79)? \nz.mem [1691] : 
                        (N81)? \nz.mem [1741] : 
                        (N83)? \nz.mem [1791] : 
                        (N85)? \nz.mem [1841] : 
                        (N87)? \nz.mem [1891] : 
                        (N89)? \nz.mem [1941] : 
                        (N91)? \nz.mem [1991] : 
                        (N93)? \nz.mem [2041] : 
                        (N95)? \nz.mem [2091] : 
                        (N97)? \nz.mem [2141] : 
                        (N99)? \nz.mem [2191] : 
                        (N101)? \nz.mem [2241] : 
                        (N103)? \nz.mem [2291] : 
                        (N105)? \nz.mem [2341] : 
                        (N107)? \nz.mem [2391] : 
                        (N109)? \nz.mem [2441] : 
                        (N111)? \nz.mem [2491] : 
                        (N113)? \nz.mem [2541] : 
                        (N115)? \nz.mem [2591] : 
                        (N117)? \nz.mem [2641] : 
                        (N119)? \nz.mem [2691] : 
                        (N121)? \nz.mem [2741] : 
                        (N123)? \nz.mem [2791] : 
                        (N125)? \nz.mem [2841] : 
                        (N127)? \nz.mem [2891] : 
                        (N129)? \nz.mem [2941] : 
                        (N131)? \nz.mem [2991] : 
                        (N133)? \nz.mem [3041] : 
                        (N135)? \nz.mem [3091] : 
                        (N137)? \nz.mem [3141] : 
                        (N139)? \nz.mem [3191] : 1'b0;
  assign r_data_o[40] = (N76)? \nz.mem [40] : 
                        (N78)? \nz.mem [90] : 
                        (N80)? \nz.mem [140] : 
                        (N82)? \nz.mem [190] : 
                        (N84)? \nz.mem [240] : 
                        (N86)? \nz.mem [290] : 
                        (N88)? \nz.mem [340] : 
                        (N90)? \nz.mem [390] : 
                        (N92)? \nz.mem [440] : 
                        (N94)? \nz.mem [490] : 
                        (N96)? \nz.mem [540] : 
                        (N98)? \nz.mem [590] : 
                        (N100)? \nz.mem [640] : 
                        (N102)? \nz.mem [690] : 
                        (N104)? \nz.mem [740] : 
                        (N106)? \nz.mem [790] : 
                        (N108)? \nz.mem [840] : 
                        (N110)? \nz.mem [890] : 
                        (N112)? \nz.mem [940] : 
                        (N114)? \nz.mem [990] : 
                        (N116)? \nz.mem [1040] : 
                        (N118)? \nz.mem [1090] : 
                        (N120)? \nz.mem [1140] : 
                        (N122)? \nz.mem [1190] : 
                        (N124)? \nz.mem [1240] : 
                        (N126)? \nz.mem [1290] : 
                        (N128)? \nz.mem [1340] : 
                        (N130)? \nz.mem [1390] : 
                        (N132)? \nz.mem [1440] : 
                        (N134)? \nz.mem [1490] : 
                        (N136)? \nz.mem [1540] : 
                        (N138)? \nz.mem [1590] : 
                        (N77)? \nz.mem [1640] : 
                        (N79)? \nz.mem [1690] : 
                        (N81)? \nz.mem [1740] : 
                        (N83)? \nz.mem [1790] : 
                        (N85)? \nz.mem [1840] : 
                        (N87)? \nz.mem [1890] : 
                        (N89)? \nz.mem [1940] : 
                        (N91)? \nz.mem [1990] : 
                        (N93)? \nz.mem [2040] : 
                        (N95)? \nz.mem [2090] : 
                        (N97)? \nz.mem [2140] : 
                        (N99)? \nz.mem [2190] : 
                        (N101)? \nz.mem [2240] : 
                        (N103)? \nz.mem [2290] : 
                        (N105)? \nz.mem [2340] : 
                        (N107)? \nz.mem [2390] : 
                        (N109)? \nz.mem [2440] : 
                        (N111)? \nz.mem [2490] : 
                        (N113)? \nz.mem [2540] : 
                        (N115)? \nz.mem [2590] : 
                        (N117)? \nz.mem [2640] : 
                        (N119)? \nz.mem [2690] : 
                        (N121)? \nz.mem [2740] : 
                        (N123)? \nz.mem [2790] : 
                        (N125)? \nz.mem [2840] : 
                        (N127)? \nz.mem [2890] : 
                        (N129)? \nz.mem [2940] : 
                        (N131)? \nz.mem [2990] : 
                        (N133)? \nz.mem [3040] : 
                        (N135)? \nz.mem [3090] : 
                        (N137)? \nz.mem [3140] : 
                        (N139)? \nz.mem [3190] : 1'b0;
  assign r_data_o[39] = (N76)? \nz.mem [39] : 
                        (N78)? \nz.mem [89] : 
                        (N80)? \nz.mem [139] : 
                        (N82)? \nz.mem [189] : 
                        (N84)? \nz.mem [239] : 
                        (N86)? \nz.mem [289] : 
                        (N88)? \nz.mem [339] : 
                        (N90)? \nz.mem [389] : 
                        (N92)? \nz.mem [439] : 
                        (N94)? \nz.mem [489] : 
                        (N96)? \nz.mem [539] : 
                        (N98)? \nz.mem [589] : 
                        (N100)? \nz.mem [639] : 
                        (N102)? \nz.mem [689] : 
                        (N104)? \nz.mem [739] : 
                        (N106)? \nz.mem [789] : 
                        (N108)? \nz.mem [839] : 
                        (N110)? \nz.mem [889] : 
                        (N112)? \nz.mem [939] : 
                        (N114)? \nz.mem [989] : 
                        (N116)? \nz.mem [1039] : 
                        (N118)? \nz.mem [1089] : 
                        (N120)? \nz.mem [1139] : 
                        (N122)? \nz.mem [1189] : 
                        (N124)? \nz.mem [1239] : 
                        (N126)? \nz.mem [1289] : 
                        (N128)? \nz.mem [1339] : 
                        (N130)? \nz.mem [1389] : 
                        (N132)? \nz.mem [1439] : 
                        (N134)? \nz.mem [1489] : 
                        (N136)? \nz.mem [1539] : 
                        (N138)? \nz.mem [1589] : 
                        (N77)? \nz.mem [1639] : 
                        (N79)? \nz.mem [1689] : 
                        (N81)? \nz.mem [1739] : 
                        (N83)? \nz.mem [1789] : 
                        (N85)? \nz.mem [1839] : 
                        (N87)? \nz.mem [1889] : 
                        (N89)? \nz.mem [1939] : 
                        (N91)? \nz.mem [1989] : 
                        (N93)? \nz.mem [2039] : 
                        (N95)? \nz.mem [2089] : 
                        (N97)? \nz.mem [2139] : 
                        (N99)? \nz.mem [2189] : 
                        (N101)? \nz.mem [2239] : 
                        (N103)? \nz.mem [2289] : 
                        (N105)? \nz.mem [2339] : 
                        (N107)? \nz.mem [2389] : 
                        (N109)? \nz.mem [2439] : 
                        (N111)? \nz.mem [2489] : 
                        (N113)? \nz.mem [2539] : 
                        (N115)? \nz.mem [2589] : 
                        (N117)? \nz.mem [2639] : 
                        (N119)? \nz.mem [2689] : 
                        (N121)? \nz.mem [2739] : 
                        (N123)? \nz.mem [2789] : 
                        (N125)? \nz.mem [2839] : 
                        (N127)? \nz.mem [2889] : 
                        (N129)? \nz.mem [2939] : 
                        (N131)? \nz.mem [2989] : 
                        (N133)? \nz.mem [3039] : 
                        (N135)? \nz.mem [3089] : 
                        (N137)? \nz.mem [3139] : 
                        (N139)? \nz.mem [3189] : 1'b0;
  assign r_data_o[38] = (N76)? \nz.mem [38] : 
                        (N78)? \nz.mem [88] : 
                        (N80)? \nz.mem [138] : 
                        (N82)? \nz.mem [188] : 
                        (N84)? \nz.mem [238] : 
                        (N86)? \nz.mem [288] : 
                        (N88)? \nz.mem [338] : 
                        (N90)? \nz.mem [388] : 
                        (N92)? \nz.mem [438] : 
                        (N94)? \nz.mem [488] : 
                        (N96)? \nz.mem [538] : 
                        (N98)? \nz.mem [588] : 
                        (N100)? \nz.mem [638] : 
                        (N102)? \nz.mem [688] : 
                        (N104)? \nz.mem [738] : 
                        (N106)? \nz.mem [788] : 
                        (N108)? \nz.mem [838] : 
                        (N110)? \nz.mem [888] : 
                        (N112)? \nz.mem [938] : 
                        (N114)? \nz.mem [988] : 
                        (N116)? \nz.mem [1038] : 
                        (N118)? \nz.mem [1088] : 
                        (N120)? \nz.mem [1138] : 
                        (N122)? \nz.mem [1188] : 
                        (N124)? \nz.mem [1238] : 
                        (N126)? \nz.mem [1288] : 
                        (N128)? \nz.mem [1338] : 
                        (N130)? \nz.mem [1388] : 
                        (N132)? \nz.mem [1438] : 
                        (N134)? \nz.mem [1488] : 
                        (N136)? \nz.mem [1538] : 
                        (N138)? \nz.mem [1588] : 
                        (N77)? \nz.mem [1638] : 
                        (N79)? \nz.mem [1688] : 
                        (N81)? \nz.mem [1738] : 
                        (N83)? \nz.mem [1788] : 
                        (N85)? \nz.mem [1838] : 
                        (N87)? \nz.mem [1888] : 
                        (N89)? \nz.mem [1938] : 
                        (N91)? \nz.mem [1988] : 
                        (N93)? \nz.mem [2038] : 
                        (N95)? \nz.mem [2088] : 
                        (N97)? \nz.mem [2138] : 
                        (N99)? \nz.mem [2188] : 
                        (N101)? \nz.mem [2238] : 
                        (N103)? \nz.mem [2288] : 
                        (N105)? \nz.mem [2338] : 
                        (N107)? \nz.mem [2388] : 
                        (N109)? \nz.mem [2438] : 
                        (N111)? \nz.mem [2488] : 
                        (N113)? \nz.mem [2538] : 
                        (N115)? \nz.mem [2588] : 
                        (N117)? \nz.mem [2638] : 
                        (N119)? \nz.mem [2688] : 
                        (N121)? \nz.mem [2738] : 
                        (N123)? \nz.mem [2788] : 
                        (N125)? \nz.mem [2838] : 
                        (N127)? \nz.mem [2888] : 
                        (N129)? \nz.mem [2938] : 
                        (N131)? \nz.mem [2988] : 
                        (N133)? \nz.mem [3038] : 
                        (N135)? \nz.mem [3088] : 
                        (N137)? \nz.mem [3138] : 
                        (N139)? \nz.mem [3188] : 1'b0;
  assign r_data_o[37] = (N76)? \nz.mem [37] : 
                        (N78)? \nz.mem [87] : 
                        (N80)? \nz.mem [137] : 
                        (N82)? \nz.mem [187] : 
                        (N84)? \nz.mem [237] : 
                        (N86)? \nz.mem [287] : 
                        (N88)? \nz.mem [337] : 
                        (N90)? \nz.mem [387] : 
                        (N92)? \nz.mem [437] : 
                        (N94)? \nz.mem [487] : 
                        (N96)? \nz.mem [537] : 
                        (N98)? \nz.mem [587] : 
                        (N100)? \nz.mem [637] : 
                        (N102)? \nz.mem [687] : 
                        (N104)? \nz.mem [737] : 
                        (N106)? \nz.mem [787] : 
                        (N108)? \nz.mem [837] : 
                        (N110)? \nz.mem [887] : 
                        (N112)? \nz.mem [937] : 
                        (N114)? \nz.mem [987] : 
                        (N116)? \nz.mem [1037] : 
                        (N118)? \nz.mem [1087] : 
                        (N120)? \nz.mem [1137] : 
                        (N122)? \nz.mem [1187] : 
                        (N124)? \nz.mem [1237] : 
                        (N126)? \nz.mem [1287] : 
                        (N128)? \nz.mem [1337] : 
                        (N130)? \nz.mem [1387] : 
                        (N132)? \nz.mem [1437] : 
                        (N134)? \nz.mem [1487] : 
                        (N136)? \nz.mem [1537] : 
                        (N138)? \nz.mem [1587] : 
                        (N77)? \nz.mem [1637] : 
                        (N79)? \nz.mem [1687] : 
                        (N81)? \nz.mem [1737] : 
                        (N83)? \nz.mem [1787] : 
                        (N85)? \nz.mem [1837] : 
                        (N87)? \nz.mem [1887] : 
                        (N89)? \nz.mem [1937] : 
                        (N91)? \nz.mem [1987] : 
                        (N93)? \nz.mem [2037] : 
                        (N95)? \nz.mem [2087] : 
                        (N97)? \nz.mem [2137] : 
                        (N99)? \nz.mem [2187] : 
                        (N101)? \nz.mem [2237] : 
                        (N103)? \nz.mem [2287] : 
                        (N105)? \nz.mem [2337] : 
                        (N107)? \nz.mem [2387] : 
                        (N109)? \nz.mem [2437] : 
                        (N111)? \nz.mem [2487] : 
                        (N113)? \nz.mem [2537] : 
                        (N115)? \nz.mem [2587] : 
                        (N117)? \nz.mem [2637] : 
                        (N119)? \nz.mem [2687] : 
                        (N121)? \nz.mem [2737] : 
                        (N123)? \nz.mem [2787] : 
                        (N125)? \nz.mem [2837] : 
                        (N127)? \nz.mem [2887] : 
                        (N129)? \nz.mem [2937] : 
                        (N131)? \nz.mem [2987] : 
                        (N133)? \nz.mem [3037] : 
                        (N135)? \nz.mem [3087] : 
                        (N137)? \nz.mem [3137] : 
                        (N139)? \nz.mem [3187] : 1'b0;
  assign r_data_o[36] = (N76)? \nz.mem [36] : 
                        (N78)? \nz.mem [86] : 
                        (N80)? \nz.mem [136] : 
                        (N82)? \nz.mem [186] : 
                        (N84)? \nz.mem [236] : 
                        (N86)? \nz.mem [286] : 
                        (N88)? \nz.mem [336] : 
                        (N90)? \nz.mem [386] : 
                        (N92)? \nz.mem [436] : 
                        (N94)? \nz.mem [486] : 
                        (N96)? \nz.mem [536] : 
                        (N98)? \nz.mem [586] : 
                        (N100)? \nz.mem [636] : 
                        (N102)? \nz.mem [686] : 
                        (N104)? \nz.mem [736] : 
                        (N106)? \nz.mem [786] : 
                        (N108)? \nz.mem [836] : 
                        (N110)? \nz.mem [886] : 
                        (N112)? \nz.mem [936] : 
                        (N114)? \nz.mem [986] : 
                        (N116)? \nz.mem [1036] : 
                        (N118)? \nz.mem [1086] : 
                        (N120)? \nz.mem [1136] : 
                        (N122)? \nz.mem [1186] : 
                        (N124)? \nz.mem [1236] : 
                        (N126)? \nz.mem [1286] : 
                        (N128)? \nz.mem [1336] : 
                        (N130)? \nz.mem [1386] : 
                        (N132)? \nz.mem [1436] : 
                        (N134)? \nz.mem [1486] : 
                        (N136)? \nz.mem [1536] : 
                        (N138)? \nz.mem [1586] : 
                        (N77)? \nz.mem [1636] : 
                        (N79)? \nz.mem [1686] : 
                        (N81)? \nz.mem [1736] : 
                        (N83)? \nz.mem [1786] : 
                        (N85)? \nz.mem [1836] : 
                        (N87)? \nz.mem [1886] : 
                        (N89)? \nz.mem [1936] : 
                        (N91)? \nz.mem [1986] : 
                        (N93)? \nz.mem [2036] : 
                        (N95)? \nz.mem [2086] : 
                        (N97)? \nz.mem [2136] : 
                        (N99)? \nz.mem [2186] : 
                        (N101)? \nz.mem [2236] : 
                        (N103)? \nz.mem [2286] : 
                        (N105)? \nz.mem [2336] : 
                        (N107)? \nz.mem [2386] : 
                        (N109)? \nz.mem [2436] : 
                        (N111)? \nz.mem [2486] : 
                        (N113)? \nz.mem [2536] : 
                        (N115)? \nz.mem [2586] : 
                        (N117)? \nz.mem [2636] : 
                        (N119)? \nz.mem [2686] : 
                        (N121)? \nz.mem [2736] : 
                        (N123)? \nz.mem [2786] : 
                        (N125)? \nz.mem [2836] : 
                        (N127)? \nz.mem [2886] : 
                        (N129)? \nz.mem [2936] : 
                        (N131)? \nz.mem [2986] : 
                        (N133)? \nz.mem [3036] : 
                        (N135)? \nz.mem [3086] : 
                        (N137)? \nz.mem [3136] : 
                        (N139)? \nz.mem [3186] : 1'b0;
  assign r_data_o[35] = (N76)? \nz.mem [35] : 
                        (N78)? \nz.mem [85] : 
                        (N80)? \nz.mem [135] : 
                        (N82)? \nz.mem [185] : 
                        (N84)? \nz.mem [235] : 
                        (N86)? \nz.mem [285] : 
                        (N88)? \nz.mem [335] : 
                        (N90)? \nz.mem [385] : 
                        (N92)? \nz.mem [435] : 
                        (N94)? \nz.mem [485] : 
                        (N96)? \nz.mem [535] : 
                        (N98)? \nz.mem [585] : 
                        (N100)? \nz.mem [635] : 
                        (N102)? \nz.mem [685] : 
                        (N104)? \nz.mem [735] : 
                        (N106)? \nz.mem [785] : 
                        (N108)? \nz.mem [835] : 
                        (N110)? \nz.mem [885] : 
                        (N112)? \nz.mem [935] : 
                        (N114)? \nz.mem [985] : 
                        (N116)? \nz.mem [1035] : 
                        (N118)? \nz.mem [1085] : 
                        (N120)? \nz.mem [1135] : 
                        (N122)? \nz.mem [1185] : 
                        (N124)? \nz.mem [1235] : 
                        (N126)? \nz.mem [1285] : 
                        (N128)? \nz.mem [1335] : 
                        (N130)? \nz.mem [1385] : 
                        (N132)? \nz.mem [1435] : 
                        (N134)? \nz.mem [1485] : 
                        (N136)? \nz.mem [1535] : 
                        (N138)? \nz.mem [1585] : 
                        (N77)? \nz.mem [1635] : 
                        (N79)? \nz.mem [1685] : 
                        (N81)? \nz.mem [1735] : 
                        (N83)? \nz.mem [1785] : 
                        (N85)? \nz.mem [1835] : 
                        (N87)? \nz.mem [1885] : 
                        (N89)? \nz.mem [1935] : 
                        (N91)? \nz.mem [1985] : 
                        (N93)? \nz.mem [2035] : 
                        (N95)? \nz.mem [2085] : 
                        (N97)? \nz.mem [2135] : 
                        (N99)? \nz.mem [2185] : 
                        (N101)? \nz.mem [2235] : 
                        (N103)? \nz.mem [2285] : 
                        (N105)? \nz.mem [2335] : 
                        (N107)? \nz.mem [2385] : 
                        (N109)? \nz.mem [2435] : 
                        (N111)? \nz.mem [2485] : 
                        (N113)? \nz.mem [2535] : 
                        (N115)? \nz.mem [2585] : 
                        (N117)? \nz.mem [2635] : 
                        (N119)? \nz.mem [2685] : 
                        (N121)? \nz.mem [2735] : 
                        (N123)? \nz.mem [2785] : 
                        (N125)? \nz.mem [2835] : 
                        (N127)? \nz.mem [2885] : 
                        (N129)? \nz.mem [2935] : 
                        (N131)? \nz.mem [2985] : 
                        (N133)? \nz.mem [3035] : 
                        (N135)? \nz.mem [3085] : 
                        (N137)? \nz.mem [3135] : 
                        (N139)? \nz.mem [3185] : 1'b0;
  assign r_data_o[34] = (N76)? \nz.mem [34] : 
                        (N78)? \nz.mem [84] : 
                        (N80)? \nz.mem [134] : 
                        (N82)? \nz.mem [184] : 
                        (N84)? \nz.mem [234] : 
                        (N86)? \nz.mem [284] : 
                        (N88)? \nz.mem [334] : 
                        (N90)? \nz.mem [384] : 
                        (N92)? \nz.mem [434] : 
                        (N94)? \nz.mem [484] : 
                        (N96)? \nz.mem [534] : 
                        (N98)? \nz.mem [584] : 
                        (N100)? \nz.mem [634] : 
                        (N102)? \nz.mem [684] : 
                        (N104)? \nz.mem [734] : 
                        (N106)? \nz.mem [784] : 
                        (N108)? \nz.mem [834] : 
                        (N110)? \nz.mem [884] : 
                        (N112)? \nz.mem [934] : 
                        (N114)? \nz.mem [984] : 
                        (N116)? \nz.mem [1034] : 
                        (N118)? \nz.mem [1084] : 
                        (N120)? \nz.mem [1134] : 
                        (N122)? \nz.mem [1184] : 
                        (N124)? \nz.mem [1234] : 
                        (N126)? \nz.mem [1284] : 
                        (N128)? \nz.mem [1334] : 
                        (N130)? \nz.mem [1384] : 
                        (N132)? \nz.mem [1434] : 
                        (N134)? \nz.mem [1484] : 
                        (N136)? \nz.mem [1534] : 
                        (N138)? \nz.mem [1584] : 
                        (N77)? \nz.mem [1634] : 
                        (N79)? \nz.mem [1684] : 
                        (N81)? \nz.mem [1734] : 
                        (N83)? \nz.mem [1784] : 
                        (N85)? \nz.mem [1834] : 
                        (N87)? \nz.mem [1884] : 
                        (N89)? \nz.mem [1934] : 
                        (N91)? \nz.mem [1984] : 
                        (N93)? \nz.mem [2034] : 
                        (N95)? \nz.mem [2084] : 
                        (N97)? \nz.mem [2134] : 
                        (N99)? \nz.mem [2184] : 
                        (N101)? \nz.mem [2234] : 
                        (N103)? \nz.mem [2284] : 
                        (N105)? \nz.mem [2334] : 
                        (N107)? \nz.mem [2384] : 
                        (N109)? \nz.mem [2434] : 
                        (N111)? \nz.mem [2484] : 
                        (N113)? \nz.mem [2534] : 
                        (N115)? \nz.mem [2584] : 
                        (N117)? \nz.mem [2634] : 
                        (N119)? \nz.mem [2684] : 
                        (N121)? \nz.mem [2734] : 
                        (N123)? \nz.mem [2784] : 
                        (N125)? \nz.mem [2834] : 
                        (N127)? \nz.mem [2884] : 
                        (N129)? \nz.mem [2934] : 
                        (N131)? \nz.mem [2984] : 
                        (N133)? \nz.mem [3034] : 
                        (N135)? \nz.mem [3084] : 
                        (N137)? \nz.mem [3134] : 
                        (N139)? \nz.mem [3184] : 1'b0;
  assign r_data_o[33] = (N76)? \nz.mem [33] : 
                        (N78)? \nz.mem [83] : 
                        (N80)? \nz.mem [133] : 
                        (N82)? \nz.mem [183] : 
                        (N84)? \nz.mem [233] : 
                        (N86)? \nz.mem [283] : 
                        (N88)? \nz.mem [333] : 
                        (N90)? \nz.mem [383] : 
                        (N92)? \nz.mem [433] : 
                        (N94)? \nz.mem [483] : 
                        (N96)? \nz.mem [533] : 
                        (N98)? \nz.mem [583] : 
                        (N100)? \nz.mem [633] : 
                        (N102)? \nz.mem [683] : 
                        (N104)? \nz.mem [733] : 
                        (N106)? \nz.mem [783] : 
                        (N108)? \nz.mem [833] : 
                        (N110)? \nz.mem [883] : 
                        (N112)? \nz.mem [933] : 
                        (N114)? \nz.mem [983] : 
                        (N116)? \nz.mem [1033] : 
                        (N118)? \nz.mem [1083] : 
                        (N120)? \nz.mem [1133] : 
                        (N122)? \nz.mem [1183] : 
                        (N124)? \nz.mem [1233] : 
                        (N126)? \nz.mem [1283] : 
                        (N128)? \nz.mem [1333] : 
                        (N130)? \nz.mem [1383] : 
                        (N132)? \nz.mem [1433] : 
                        (N134)? \nz.mem [1483] : 
                        (N136)? \nz.mem [1533] : 
                        (N138)? \nz.mem [1583] : 
                        (N77)? \nz.mem [1633] : 
                        (N79)? \nz.mem [1683] : 
                        (N81)? \nz.mem [1733] : 
                        (N83)? \nz.mem [1783] : 
                        (N85)? \nz.mem [1833] : 
                        (N87)? \nz.mem [1883] : 
                        (N89)? \nz.mem [1933] : 
                        (N91)? \nz.mem [1983] : 
                        (N93)? \nz.mem [2033] : 
                        (N95)? \nz.mem [2083] : 
                        (N97)? \nz.mem [2133] : 
                        (N99)? \nz.mem [2183] : 
                        (N101)? \nz.mem [2233] : 
                        (N103)? \nz.mem [2283] : 
                        (N105)? \nz.mem [2333] : 
                        (N107)? \nz.mem [2383] : 
                        (N109)? \nz.mem [2433] : 
                        (N111)? \nz.mem [2483] : 
                        (N113)? \nz.mem [2533] : 
                        (N115)? \nz.mem [2583] : 
                        (N117)? \nz.mem [2633] : 
                        (N119)? \nz.mem [2683] : 
                        (N121)? \nz.mem [2733] : 
                        (N123)? \nz.mem [2783] : 
                        (N125)? \nz.mem [2833] : 
                        (N127)? \nz.mem [2883] : 
                        (N129)? \nz.mem [2933] : 
                        (N131)? \nz.mem [2983] : 
                        (N133)? \nz.mem [3033] : 
                        (N135)? \nz.mem [3083] : 
                        (N137)? \nz.mem [3133] : 
                        (N139)? \nz.mem [3183] : 1'b0;
  assign r_data_o[32] = (N76)? \nz.mem [32] : 
                        (N78)? \nz.mem [82] : 
                        (N80)? \nz.mem [132] : 
                        (N82)? \nz.mem [182] : 
                        (N84)? \nz.mem [232] : 
                        (N86)? \nz.mem [282] : 
                        (N88)? \nz.mem [332] : 
                        (N90)? \nz.mem [382] : 
                        (N92)? \nz.mem [432] : 
                        (N94)? \nz.mem [482] : 
                        (N96)? \nz.mem [532] : 
                        (N98)? \nz.mem [582] : 
                        (N100)? \nz.mem [632] : 
                        (N102)? \nz.mem [682] : 
                        (N104)? \nz.mem [732] : 
                        (N106)? \nz.mem [782] : 
                        (N108)? \nz.mem [832] : 
                        (N110)? \nz.mem [882] : 
                        (N112)? \nz.mem [932] : 
                        (N114)? \nz.mem [982] : 
                        (N116)? \nz.mem [1032] : 
                        (N118)? \nz.mem [1082] : 
                        (N120)? \nz.mem [1132] : 
                        (N122)? \nz.mem [1182] : 
                        (N124)? \nz.mem [1232] : 
                        (N126)? \nz.mem [1282] : 
                        (N128)? \nz.mem [1332] : 
                        (N130)? \nz.mem [1382] : 
                        (N132)? \nz.mem [1432] : 
                        (N134)? \nz.mem [1482] : 
                        (N136)? \nz.mem [1532] : 
                        (N138)? \nz.mem [1582] : 
                        (N77)? \nz.mem [1632] : 
                        (N79)? \nz.mem [1682] : 
                        (N81)? \nz.mem [1732] : 
                        (N83)? \nz.mem [1782] : 
                        (N85)? \nz.mem [1832] : 
                        (N87)? \nz.mem [1882] : 
                        (N89)? \nz.mem [1932] : 
                        (N91)? \nz.mem [1982] : 
                        (N93)? \nz.mem [2032] : 
                        (N95)? \nz.mem [2082] : 
                        (N97)? \nz.mem [2132] : 
                        (N99)? \nz.mem [2182] : 
                        (N101)? \nz.mem [2232] : 
                        (N103)? \nz.mem [2282] : 
                        (N105)? \nz.mem [2332] : 
                        (N107)? \nz.mem [2382] : 
                        (N109)? \nz.mem [2432] : 
                        (N111)? \nz.mem [2482] : 
                        (N113)? \nz.mem [2532] : 
                        (N115)? \nz.mem [2582] : 
                        (N117)? \nz.mem [2632] : 
                        (N119)? \nz.mem [2682] : 
                        (N121)? \nz.mem [2732] : 
                        (N123)? \nz.mem [2782] : 
                        (N125)? \nz.mem [2832] : 
                        (N127)? \nz.mem [2882] : 
                        (N129)? \nz.mem [2932] : 
                        (N131)? \nz.mem [2982] : 
                        (N133)? \nz.mem [3032] : 
                        (N135)? \nz.mem [3082] : 
                        (N137)? \nz.mem [3132] : 
                        (N139)? \nz.mem [3182] : 1'b0;
  assign r_data_o[31] = (N76)? \nz.mem [31] : 
                        (N78)? \nz.mem [81] : 
                        (N80)? \nz.mem [131] : 
                        (N82)? \nz.mem [181] : 
                        (N84)? \nz.mem [231] : 
                        (N86)? \nz.mem [281] : 
                        (N88)? \nz.mem [331] : 
                        (N90)? \nz.mem [381] : 
                        (N92)? \nz.mem [431] : 
                        (N94)? \nz.mem [481] : 
                        (N96)? \nz.mem [531] : 
                        (N98)? \nz.mem [581] : 
                        (N100)? \nz.mem [631] : 
                        (N102)? \nz.mem [681] : 
                        (N104)? \nz.mem [731] : 
                        (N106)? \nz.mem [781] : 
                        (N108)? \nz.mem [831] : 
                        (N110)? \nz.mem [881] : 
                        (N112)? \nz.mem [931] : 
                        (N114)? \nz.mem [981] : 
                        (N116)? \nz.mem [1031] : 
                        (N118)? \nz.mem [1081] : 
                        (N120)? \nz.mem [1131] : 
                        (N122)? \nz.mem [1181] : 
                        (N124)? \nz.mem [1231] : 
                        (N126)? \nz.mem [1281] : 
                        (N128)? \nz.mem [1331] : 
                        (N130)? \nz.mem [1381] : 
                        (N132)? \nz.mem [1431] : 
                        (N134)? \nz.mem [1481] : 
                        (N136)? \nz.mem [1531] : 
                        (N138)? \nz.mem [1581] : 
                        (N77)? \nz.mem [1631] : 
                        (N79)? \nz.mem [1681] : 
                        (N81)? \nz.mem [1731] : 
                        (N83)? \nz.mem [1781] : 
                        (N85)? \nz.mem [1831] : 
                        (N87)? \nz.mem [1881] : 
                        (N89)? \nz.mem [1931] : 
                        (N91)? \nz.mem [1981] : 
                        (N93)? \nz.mem [2031] : 
                        (N95)? \nz.mem [2081] : 
                        (N97)? \nz.mem [2131] : 
                        (N99)? \nz.mem [2181] : 
                        (N101)? \nz.mem [2231] : 
                        (N103)? \nz.mem [2281] : 
                        (N105)? \nz.mem [2331] : 
                        (N107)? \nz.mem [2381] : 
                        (N109)? \nz.mem [2431] : 
                        (N111)? \nz.mem [2481] : 
                        (N113)? \nz.mem [2531] : 
                        (N115)? \nz.mem [2581] : 
                        (N117)? \nz.mem [2631] : 
                        (N119)? \nz.mem [2681] : 
                        (N121)? \nz.mem [2731] : 
                        (N123)? \nz.mem [2781] : 
                        (N125)? \nz.mem [2831] : 
                        (N127)? \nz.mem [2881] : 
                        (N129)? \nz.mem [2931] : 
                        (N131)? \nz.mem [2981] : 
                        (N133)? \nz.mem [3031] : 
                        (N135)? \nz.mem [3081] : 
                        (N137)? \nz.mem [3131] : 
                        (N139)? \nz.mem [3181] : 1'b0;
  assign r_data_o[30] = (N76)? \nz.mem [30] : 
                        (N78)? \nz.mem [80] : 
                        (N80)? \nz.mem [130] : 
                        (N82)? \nz.mem [180] : 
                        (N84)? \nz.mem [230] : 
                        (N86)? \nz.mem [280] : 
                        (N88)? \nz.mem [330] : 
                        (N90)? \nz.mem [380] : 
                        (N92)? \nz.mem [430] : 
                        (N94)? \nz.mem [480] : 
                        (N96)? \nz.mem [530] : 
                        (N98)? \nz.mem [580] : 
                        (N100)? \nz.mem [630] : 
                        (N102)? \nz.mem [680] : 
                        (N104)? \nz.mem [730] : 
                        (N106)? \nz.mem [780] : 
                        (N108)? \nz.mem [830] : 
                        (N110)? \nz.mem [880] : 
                        (N112)? \nz.mem [930] : 
                        (N114)? \nz.mem [980] : 
                        (N116)? \nz.mem [1030] : 
                        (N118)? \nz.mem [1080] : 
                        (N120)? \nz.mem [1130] : 
                        (N122)? \nz.mem [1180] : 
                        (N124)? \nz.mem [1230] : 
                        (N126)? \nz.mem [1280] : 
                        (N128)? \nz.mem [1330] : 
                        (N130)? \nz.mem [1380] : 
                        (N132)? \nz.mem [1430] : 
                        (N134)? \nz.mem [1480] : 
                        (N136)? \nz.mem [1530] : 
                        (N138)? \nz.mem [1580] : 
                        (N77)? \nz.mem [1630] : 
                        (N79)? \nz.mem [1680] : 
                        (N81)? \nz.mem [1730] : 
                        (N83)? \nz.mem [1780] : 
                        (N85)? \nz.mem [1830] : 
                        (N87)? \nz.mem [1880] : 
                        (N89)? \nz.mem [1930] : 
                        (N91)? \nz.mem [1980] : 
                        (N93)? \nz.mem [2030] : 
                        (N95)? \nz.mem [2080] : 
                        (N97)? \nz.mem [2130] : 
                        (N99)? \nz.mem [2180] : 
                        (N101)? \nz.mem [2230] : 
                        (N103)? \nz.mem [2280] : 
                        (N105)? \nz.mem [2330] : 
                        (N107)? \nz.mem [2380] : 
                        (N109)? \nz.mem [2430] : 
                        (N111)? \nz.mem [2480] : 
                        (N113)? \nz.mem [2530] : 
                        (N115)? \nz.mem [2580] : 
                        (N117)? \nz.mem [2630] : 
                        (N119)? \nz.mem [2680] : 
                        (N121)? \nz.mem [2730] : 
                        (N123)? \nz.mem [2780] : 
                        (N125)? \nz.mem [2830] : 
                        (N127)? \nz.mem [2880] : 
                        (N129)? \nz.mem [2930] : 
                        (N131)? \nz.mem [2980] : 
                        (N133)? \nz.mem [3030] : 
                        (N135)? \nz.mem [3080] : 
                        (N137)? \nz.mem [3130] : 
                        (N139)? \nz.mem [3180] : 1'b0;
  assign r_data_o[29] = (N76)? \nz.mem [29] : 
                        (N78)? \nz.mem [79] : 
                        (N80)? \nz.mem [129] : 
                        (N82)? \nz.mem [179] : 
                        (N84)? \nz.mem [229] : 
                        (N86)? \nz.mem [279] : 
                        (N88)? \nz.mem [329] : 
                        (N90)? \nz.mem [379] : 
                        (N92)? \nz.mem [429] : 
                        (N94)? \nz.mem [479] : 
                        (N96)? \nz.mem [529] : 
                        (N98)? \nz.mem [579] : 
                        (N100)? \nz.mem [629] : 
                        (N102)? \nz.mem [679] : 
                        (N104)? \nz.mem [729] : 
                        (N106)? \nz.mem [779] : 
                        (N108)? \nz.mem [829] : 
                        (N110)? \nz.mem [879] : 
                        (N112)? \nz.mem [929] : 
                        (N114)? \nz.mem [979] : 
                        (N116)? \nz.mem [1029] : 
                        (N118)? \nz.mem [1079] : 
                        (N120)? \nz.mem [1129] : 
                        (N122)? \nz.mem [1179] : 
                        (N124)? \nz.mem [1229] : 
                        (N126)? \nz.mem [1279] : 
                        (N128)? \nz.mem [1329] : 
                        (N130)? \nz.mem [1379] : 
                        (N132)? \nz.mem [1429] : 
                        (N134)? \nz.mem [1479] : 
                        (N136)? \nz.mem [1529] : 
                        (N138)? \nz.mem [1579] : 
                        (N77)? \nz.mem [1629] : 
                        (N79)? \nz.mem [1679] : 
                        (N81)? \nz.mem [1729] : 
                        (N83)? \nz.mem [1779] : 
                        (N85)? \nz.mem [1829] : 
                        (N87)? \nz.mem [1879] : 
                        (N89)? \nz.mem [1929] : 
                        (N91)? \nz.mem [1979] : 
                        (N93)? \nz.mem [2029] : 
                        (N95)? \nz.mem [2079] : 
                        (N97)? \nz.mem [2129] : 
                        (N99)? \nz.mem [2179] : 
                        (N101)? \nz.mem [2229] : 
                        (N103)? \nz.mem [2279] : 
                        (N105)? \nz.mem [2329] : 
                        (N107)? \nz.mem [2379] : 
                        (N109)? \nz.mem [2429] : 
                        (N111)? \nz.mem [2479] : 
                        (N113)? \nz.mem [2529] : 
                        (N115)? \nz.mem [2579] : 
                        (N117)? \nz.mem [2629] : 
                        (N119)? \nz.mem [2679] : 
                        (N121)? \nz.mem [2729] : 
                        (N123)? \nz.mem [2779] : 
                        (N125)? \nz.mem [2829] : 
                        (N127)? \nz.mem [2879] : 
                        (N129)? \nz.mem [2929] : 
                        (N131)? \nz.mem [2979] : 
                        (N133)? \nz.mem [3029] : 
                        (N135)? \nz.mem [3079] : 
                        (N137)? \nz.mem [3129] : 
                        (N139)? \nz.mem [3179] : 1'b0;
  assign r_data_o[28] = (N76)? \nz.mem [28] : 
                        (N78)? \nz.mem [78] : 
                        (N80)? \nz.mem [128] : 
                        (N82)? \nz.mem [178] : 
                        (N84)? \nz.mem [228] : 
                        (N86)? \nz.mem [278] : 
                        (N88)? \nz.mem [328] : 
                        (N90)? \nz.mem [378] : 
                        (N92)? \nz.mem [428] : 
                        (N94)? \nz.mem [478] : 
                        (N96)? \nz.mem [528] : 
                        (N98)? \nz.mem [578] : 
                        (N100)? \nz.mem [628] : 
                        (N102)? \nz.mem [678] : 
                        (N104)? \nz.mem [728] : 
                        (N106)? \nz.mem [778] : 
                        (N108)? \nz.mem [828] : 
                        (N110)? \nz.mem [878] : 
                        (N112)? \nz.mem [928] : 
                        (N114)? \nz.mem [978] : 
                        (N116)? \nz.mem [1028] : 
                        (N118)? \nz.mem [1078] : 
                        (N120)? \nz.mem [1128] : 
                        (N122)? \nz.mem [1178] : 
                        (N124)? \nz.mem [1228] : 
                        (N126)? \nz.mem [1278] : 
                        (N128)? \nz.mem [1328] : 
                        (N130)? \nz.mem [1378] : 
                        (N132)? \nz.mem [1428] : 
                        (N134)? \nz.mem [1478] : 
                        (N136)? \nz.mem [1528] : 
                        (N138)? \nz.mem [1578] : 
                        (N77)? \nz.mem [1628] : 
                        (N79)? \nz.mem [1678] : 
                        (N81)? \nz.mem [1728] : 
                        (N83)? \nz.mem [1778] : 
                        (N85)? \nz.mem [1828] : 
                        (N87)? \nz.mem [1878] : 
                        (N89)? \nz.mem [1928] : 
                        (N91)? \nz.mem [1978] : 
                        (N93)? \nz.mem [2028] : 
                        (N95)? \nz.mem [2078] : 
                        (N97)? \nz.mem [2128] : 
                        (N99)? \nz.mem [2178] : 
                        (N101)? \nz.mem [2228] : 
                        (N103)? \nz.mem [2278] : 
                        (N105)? \nz.mem [2328] : 
                        (N107)? \nz.mem [2378] : 
                        (N109)? \nz.mem [2428] : 
                        (N111)? \nz.mem [2478] : 
                        (N113)? \nz.mem [2528] : 
                        (N115)? \nz.mem [2578] : 
                        (N117)? \nz.mem [2628] : 
                        (N119)? \nz.mem [2678] : 
                        (N121)? \nz.mem [2728] : 
                        (N123)? \nz.mem [2778] : 
                        (N125)? \nz.mem [2828] : 
                        (N127)? \nz.mem [2878] : 
                        (N129)? \nz.mem [2928] : 
                        (N131)? \nz.mem [2978] : 
                        (N133)? \nz.mem [3028] : 
                        (N135)? \nz.mem [3078] : 
                        (N137)? \nz.mem [3128] : 
                        (N139)? \nz.mem [3178] : 1'b0;
  assign r_data_o[27] = (N76)? \nz.mem [27] : 
                        (N78)? \nz.mem [77] : 
                        (N80)? \nz.mem [127] : 
                        (N82)? \nz.mem [177] : 
                        (N84)? \nz.mem [227] : 
                        (N86)? \nz.mem [277] : 
                        (N88)? \nz.mem [327] : 
                        (N90)? \nz.mem [377] : 
                        (N92)? \nz.mem [427] : 
                        (N94)? \nz.mem [477] : 
                        (N96)? \nz.mem [527] : 
                        (N98)? \nz.mem [577] : 
                        (N100)? \nz.mem [627] : 
                        (N102)? \nz.mem [677] : 
                        (N104)? \nz.mem [727] : 
                        (N106)? \nz.mem [777] : 
                        (N108)? \nz.mem [827] : 
                        (N110)? \nz.mem [877] : 
                        (N112)? \nz.mem [927] : 
                        (N114)? \nz.mem [977] : 
                        (N116)? \nz.mem [1027] : 
                        (N118)? \nz.mem [1077] : 
                        (N120)? \nz.mem [1127] : 
                        (N122)? \nz.mem [1177] : 
                        (N124)? \nz.mem [1227] : 
                        (N126)? \nz.mem [1277] : 
                        (N128)? \nz.mem [1327] : 
                        (N130)? \nz.mem [1377] : 
                        (N132)? \nz.mem [1427] : 
                        (N134)? \nz.mem [1477] : 
                        (N136)? \nz.mem [1527] : 
                        (N138)? \nz.mem [1577] : 
                        (N77)? \nz.mem [1627] : 
                        (N79)? \nz.mem [1677] : 
                        (N81)? \nz.mem [1727] : 
                        (N83)? \nz.mem [1777] : 
                        (N85)? \nz.mem [1827] : 
                        (N87)? \nz.mem [1877] : 
                        (N89)? \nz.mem [1927] : 
                        (N91)? \nz.mem [1977] : 
                        (N93)? \nz.mem [2027] : 
                        (N95)? \nz.mem [2077] : 
                        (N97)? \nz.mem [2127] : 
                        (N99)? \nz.mem [2177] : 
                        (N101)? \nz.mem [2227] : 
                        (N103)? \nz.mem [2277] : 
                        (N105)? \nz.mem [2327] : 
                        (N107)? \nz.mem [2377] : 
                        (N109)? \nz.mem [2427] : 
                        (N111)? \nz.mem [2477] : 
                        (N113)? \nz.mem [2527] : 
                        (N115)? \nz.mem [2577] : 
                        (N117)? \nz.mem [2627] : 
                        (N119)? \nz.mem [2677] : 
                        (N121)? \nz.mem [2727] : 
                        (N123)? \nz.mem [2777] : 
                        (N125)? \nz.mem [2827] : 
                        (N127)? \nz.mem [2877] : 
                        (N129)? \nz.mem [2927] : 
                        (N131)? \nz.mem [2977] : 
                        (N133)? \nz.mem [3027] : 
                        (N135)? \nz.mem [3077] : 
                        (N137)? \nz.mem [3127] : 
                        (N139)? \nz.mem [3177] : 1'b0;
  assign r_data_o[26] = (N76)? \nz.mem [26] : 
                        (N78)? \nz.mem [76] : 
                        (N80)? \nz.mem [126] : 
                        (N82)? \nz.mem [176] : 
                        (N84)? \nz.mem [226] : 
                        (N86)? \nz.mem [276] : 
                        (N88)? \nz.mem [326] : 
                        (N90)? \nz.mem [376] : 
                        (N92)? \nz.mem [426] : 
                        (N94)? \nz.mem [476] : 
                        (N96)? \nz.mem [526] : 
                        (N98)? \nz.mem [576] : 
                        (N100)? \nz.mem [626] : 
                        (N102)? \nz.mem [676] : 
                        (N104)? \nz.mem [726] : 
                        (N106)? \nz.mem [776] : 
                        (N108)? \nz.mem [826] : 
                        (N110)? \nz.mem [876] : 
                        (N112)? \nz.mem [926] : 
                        (N114)? \nz.mem [976] : 
                        (N116)? \nz.mem [1026] : 
                        (N118)? \nz.mem [1076] : 
                        (N120)? \nz.mem [1126] : 
                        (N122)? \nz.mem [1176] : 
                        (N124)? \nz.mem [1226] : 
                        (N126)? \nz.mem [1276] : 
                        (N128)? \nz.mem [1326] : 
                        (N130)? \nz.mem [1376] : 
                        (N132)? \nz.mem [1426] : 
                        (N134)? \nz.mem [1476] : 
                        (N136)? \nz.mem [1526] : 
                        (N138)? \nz.mem [1576] : 
                        (N77)? \nz.mem [1626] : 
                        (N79)? \nz.mem [1676] : 
                        (N81)? \nz.mem [1726] : 
                        (N83)? \nz.mem [1776] : 
                        (N85)? \nz.mem [1826] : 
                        (N87)? \nz.mem [1876] : 
                        (N89)? \nz.mem [1926] : 
                        (N91)? \nz.mem [1976] : 
                        (N93)? \nz.mem [2026] : 
                        (N95)? \nz.mem [2076] : 
                        (N97)? \nz.mem [2126] : 
                        (N99)? \nz.mem [2176] : 
                        (N101)? \nz.mem [2226] : 
                        (N103)? \nz.mem [2276] : 
                        (N105)? \nz.mem [2326] : 
                        (N107)? \nz.mem [2376] : 
                        (N109)? \nz.mem [2426] : 
                        (N111)? \nz.mem [2476] : 
                        (N113)? \nz.mem [2526] : 
                        (N115)? \nz.mem [2576] : 
                        (N117)? \nz.mem [2626] : 
                        (N119)? \nz.mem [2676] : 
                        (N121)? \nz.mem [2726] : 
                        (N123)? \nz.mem [2776] : 
                        (N125)? \nz.mem [2826] : 
                        (N127)? \nz.mem [2876] : 
                        (N129)? \nz.mem [2926] : 
                        (N131)? \nz.mem [2976] : 
                        (N133)? \nz.mem [3026] : 
                        (N135)? \nz.mem [3076] : 
                        (N137)? \nz.mem [3126] : 
                        (N139)? \nz.mem [3176] : 1'b0;
  assign r_data_o[25] = (N76)? \nz.mem [25] : 
                        (N78)? \nz.mem [75] : 
                        (N80)? \nz.mem [125] : 
                        (N82)? \nz.mem [175] : 
                        (N84)? \nz.mem [225] : 
                        (N86)? \nz.mem [275] : 
                        (N88)? \nz.mem [325] : 
                        (N90)? \nz.mem [375] : 
                        (N92)? \nz.mem [425] : 
                        (N94)? \nz.mem [475] : 
                        (N96)? \nz.mem [525] : 
                        (N98)? \nz.mem [575] : 
                        (N100)? \nz.mem [625] : 
                        (N102)? \nz.mem [675] : 
                        (N104)? \nz.mem [725] : 
                        (N106)? \nz.mem [775] : 
                        (N108)? \nz.mem [825] : 
                        (N110)? \nz.mem [875] : 
                        (N112)? \nz.mem [925] : 
                        (N114)? \nz.mem [975] : 
                        (N116)? \nz.mem [1025] : 
                        (N118)? \nz.mem [1075] : 
                        (N120)? \nz.mem [1125] : 
                        (N122)? \nz.mem [1175] : 
                        (N124)? \nz.mem [1225] : 
                        (N126)? \nz.mem [1275] : 
                        (N128)? \nz.mem [1325] : 
                        (N130)? \nz.mem [1375] : 
                        (N132)? \nz.mem [1425] : 
                        (N134)? \nz.mem [1475] : 
                        (N136)? \nz.mem [1525] : 
                        (N138)? \nz.mem [1575] : 
                        (N77)? \nz.mem [1625] : 
                        (N79)? \nz.mem [1675] : 
                        (N81)? \nz.mem [1725] : 
                        (N83)? \nz.mem [1775] : 
                        (N85)? \nz.mem [1825] : 
                        (N87)? \nz.mem [1875] : 
                        (N89)? \nz.mem [1925] : 
                        (N91)? \nz.mem [1975] : 
                        (N93)? \nz.mem [2025] : 
                        (N95)? \nz.mem [2075] : 
                        (N97)? \nz.mem [2125] : 
                        (N99)? \nz.mem [2175] : 
                        (N101)? \nz.mem [2225] : 
                        (N103)? \nz.mem [2275] : 
                        (N105)? \nz.mem [2325] : 
                        (N107)? \nz.mem [2375] : 
                        (N109)? \nz.mem [2425] : 
                        (N111)? \nz.mem [2475] : 
                        (N113)? \nz.mem [2525] : 
                        (N115)? \nz.mem [2575] : 
                        (N117)? \nz.mem [2625] : 
                        (N119)? \nz.mem [2675] : 
                        (N121)? \nz.mem [2725] : 
                        (N123)? \nz.mem [2775] : 
                        (N125)? \nz.mem [2825] : 
                        (N127)? \nz.mem [2875] : 
                        (N129)? \nz.mem [2925] : 
                        (N131)? \nz.mem [2975] : 
                        (N133)? \nz.mem [3025] : 
                        (N135)? \nz.mem [3075] : 
                        (N137)? \nz.mem [3125] : 
                        (N139)? \nz.mem [3175] : 1'b0;
  assign r_data_o[24] = (N76)? \nz.mem [24] : 
                        (N78)? \nz.mem [74] : 
                        (N80)? \nz.mem [124] : 
                        (N82)? \nz.mem [174] : 
                        (N84)? \nz.mem [224] : 
                        (N86)? \nz.mem [274] : 
                        (N88)? \nz.mem [324] : 
                        (N90)? \nz.mem [374] : 
                        (N92)? \nz.mem [424] : 
                        (N94)? \nz.mem [474] : 
                        (N96)? \nz.mem [524] : 
                        (N98)? \nz.mem [574] : 
                        (N100)? \nz.mem [624] : 
                        (N102)? \nz.mem [674] : 
                        (N104)? \nz.mem [724] : 
                        (N106)? \nz.mem [774] : 
                        (N108)? \nz.mem [824] : 
                        (N110)? \nz.mem [874] : 
                        (N112)? \nz.mem [924] : 
                        (N114)? \nz.mem [974] : 
                        (N116)? \nz.mem [1024] : 
                        (N118)? \nz.mem [1074] : 
                        (N120)? \nz.mem [1124] : 
                        (N122)? \nz.mem [1174] : 
                        (N124)? \nz.mem [1224] : 
                        (N126)? \nz.mem [1274] : 
                        (N128)? \nz.mem [1324] : 
                        (N130)? \nz.mem [1374] : 
                        (N132)? \nz.mem [1424] : 
                        (N134)? \nz.mem [1474] : 
                        (N136)? \nz.mem [1524] : 
                        (N138)? \nz.mem [1574] : 
                        (N77)? \nz.mem [1624] : 
                        (N79)? \nz.mem [1674] : 
                        (N81)? \nz.mem [1724] : 
                        (N83)? \nz.mem [1774] : 
                        (N85)? \nz.mem [1824] : 
                        (N87)? \nz.mem [1874] : 
                        (N89)? \nz.mem [1924] : 
                        (N91)? \nz.mem [1974] : 
                        (N93)? \nz.mem [2024] : 
                        (N95)? \nz.mem [2074] : 
                        (N97)? \nz.mem [2124] : 
                        (N99)? \nz.mem [2174] : 
                        (N101)? \nz.mem [2224] : 
                        (N103)? \nz.mem [2274] : 
                        (N105)? \nz.mem [2324] : 
                        (N107)? \nz.mem [2374] : 
                        (N109)? \nz.mem [2424] : 
                        (N111)? \nz.mem [2474] : 
                        (N113)? \nz.mem [2524] : 
                        (N115)? \nz.mem [2574] : 
                        (N117)? \nz.mem [2624] : 
                        (N119)? \nz.mem [2674] : 
                        (N121)? \nz.mem [2724] : 
                        (N123)? \nz.mem [2774] : 
                        (N125)? \nz.mem [2824] : 
                        (N127)? \nz.mem [2874] : 
                        (N129)? \nz.mem [2924] : 
                        (N131)? \nz.mem [2974] : 
                        (N133)? \nz.mem [3024] : 
                        (N135)? \nz.mem [3074] : 
                        (N137)? \nz.mem [3124] : 
                        (N139)? \nz.mem [3174] : 1'b0;
  assign r_data_o[23] = (N76)? \nz.mem [23] : 
                        (N78)? \nz.mem [73] : 
                        (N80)? \nz.mem [123] : 
                        (N82)? \nz.mem [173] : 
                        (N84)? \nz.mem [223] : 
                        (N86)? \nz.mem [273] : 
                        (N88)? \nz.mem [323] : 
                        (N90)? \nz.mem [373] : 
                        (N92)? \nz.mem [423] : 
                        (N94)? \nz.mem [473] : 
                        (N96)? \nz.mem [523] : 
                        (N98)? \nz.mem [573] : 
                        (N100)? \nz.mem [623] : 
                        (N102)? \nz.mem [673] : 
                        (N104)? \nz.mem [723] : 
                        (N106)? \nz.mem [773] : 
                        (N108)? \nz.mem [823] : 
                        (N110)? \nz.mem [873] : 
                        (N112)? \nz.mem [923] : 
                        (N114)? \nz.mem [973] : 
                        (N116)? \nz.mem [1023] : 
                        (N118)? \nz.mem [1073] : 
                        (N120)? \nz.mem [1123] : 
                        (N122)? \nz.mem [1173] : 
                        (N124)? \nz.mem [1223] : 
                        (N126)? \nz.mem [1273] : 
                        (N128)? \nz.mem [1323] : 
                        (N130)? \nz.mem [1373] : 
                        (N132)? \nz.mem [1423] : 
                        (N134)? \nz.mem [1473] : 
                        (N136)? \nz.mem [1523] : 
                        (N138)? \nz.mem [1573] : 
                        (N77)? \nz.mem [1623] : 
                        (N79)? \nz.mem [1673] : 
                        (N81)? \nz.mem [1723] : 
                        (N83)? \nz.mem [1773] : 
                        (N85)? \nz.mem [1823] : 
                        (N87)? \nz.mem [1873] : 
                        (N89)? \nz.mem [1923] : 
                        (N91)? \nz.mem [1973] : 
                        (N93)? \nz.mem [2023] : 
                        (N95)? \nz.mem [2073] : 
                        (N97)? \nz.mem [2123] : 
                        (N99)? \nz.mem [2173] : 
                        (N101)? \nz.mem [2223] : 
                        (N103)? \nz.mem [2273] : 
                        (N105)? \nz.mem [2323] : 
                        (N107)? \nz.mem [2373] : 
                        (N109)? \nz.mem [2423] : 
                        (N111)? \nz.mem [2473] : 
                        (N113)? \nz.mem [2523] : 
                        (N115)? \nz.mem [2573] : 
                        (N117)? \nz.mem [2623] : 
                        (N119)? \nz.mem [2673] : 
                        (N121)? \nz.mem [2723] : 
                        (N123)? \nz.mem [2773] : 
                        (N125)? \nz.mem [2823] : 
                        (N127)? \nz.mem [2873] : 
                        (N129)? \nz.mem [2923] : 
                        (N131)? \nz.mem [2973] : 
                        (N133)? \nz.mem [3023] : 
                        (N135)? \nz.mem [3073] : 
                        (N137)? \nz.mem [3123] : 
                        (N139)? \nz.mem [3173] : 1'b0;
  assign r_data_o[22] = (N76)? \nz.mem [22] : 
                        (N78)? \nz.mem [72] : 
                        (N80)? \nz.mem [122] : 
                        (N82)? \nz.mem [172] : 
                        (N84)? \nz.mem [222] : 
                        (N86)? \nz.mem [272] : 
                        (N88)? \nz.mem [322] : 
                        (N90)? \nz.mem [372] : 
                        (N92)? \nz.mem [422] : 
                        (N94)? \nz.mem [472] : 
                        (N96)? \nz.mem [522] : 
                        (N98)? \nz.mem [572] : 
                        (N100)? \nz.mem [622] : 
                        (N102)? \nz.mem [672] : 
                        (N104)? \nz.mem [722] : 
                        (N106)? \nz.mem [772] : 
                        (N108)? \nz.mem [822] : 
                        (N110)? \nz.mem [872] : 
                        (N112)? \nz.mem [922] : 
                        (N114)? \nz.mem [972] : 
                        (N116)? \nz.mem [1022] : 
                        (N118)? \nz.mem [1072] : 
                        (N120)? \nz.mem [1122] : 
                        (N122)? \nz.mem [1172] : 
                        (N124)? \nz.mem [1222] : 
                        (N126)? \nz.mem [1272] : 
                        (N128)? \nz.mem [1322] : 
                        (N130)? \nz.mem [1372] : 
                        (N132)? \nz.mem [1422] : 
                        (N134)? \nz.mem [1472] : 
                        (N136)? \nz.mem [1522] : 
                        (N138)? \nz.mem [1572] : 
                        (N77)? \nz.mem [1622] : 
                        (N79)? \nz.mem [1672] : 
                        (N81)? \nz.mem [1722] : 
                        (N83)? \nz.mem [1772] : 
                        (N85)? \nz.mem [1822] : 
                        (N87)? \nz.mem [1872] : 
                        (N89)? \nz.mem [1922] : 
                        (N91)? \nz.mem [1972] : 
                        (N93)? \nz.mem [2022] : 
                        (N95)? \nz.mem [2072] : 
                        (N97)? \nz.mem [2122] : 
                        (N99)? \nz.mem [2172] : 
                        (N101)? \nz.mem [2222] : 
                        (N103)? \nz.mem [2272] : 
                        (N105)? \nz.mem [2322] : 
                        (N107)? \nz.mem [2372] : 
                        (N109)? \nz.mem [2422] : 
                        (N111)? \nz.mem [2472] : 
                        (N113)? \nz.mem [2522] : 
                        (N115)? \nz.mem [2572] : 
                        (N117)? \nz.mem [2622] : 
                        (N119)? \nz.mem [2672] : 
                        (N121)? \nz.mem [2722] : 
                        (N123)? \nz.mem [2772] : 
                        (N125)? \nz.mem [2822] : 
                        (N127)? \nz.mem [2872] : 
                        (N129)? \nz.mem [2922] : 
                        (N131)? \nz.mem [2972] : 
                        (N133)? \nz.mem [3022] : 
                        (N135)? \nz.mem [3072] : 
                        (N137)? \nz.mem [3122] : 
                        (N139)? \nz.mem [3172] : 1'b0;
  assign r_data_o[21] = (N76)? \nz.mem [21] : 
                        (N78)? \nz.mem [71] : 
                        (N80)? \nz.mem [121] : 
                        (N82)? \nz.mem [171] : 
                        (N84)? \nz.mem [221] : 
                        (N86)? \nz.mem [271] : 
                        (N88)? \nz.mem [321] : 
                        (N90)? \nz.mem [371] : 
                        (N92)? \nz.mem [421] : 
                        (N94)? \nz.mem [471] : 
                        (N96)? \nz.mem [521] : 
                        (N98)? \nz.mem [571] : 
                        (N100)? \nz.mem [621] : 
                        (N102)? \nz.mem [671] : 
                        (N104)? \nz.mem [721] : 
                        (N106)? \nz.mem [771] : 
                        (N108)? \nz.mem [821] : 
                        (N110)? \nz.mem [871] : 
                        (N112)? \nz.mem [921] : 
                        (N114)? \nz.mem [971] : 
                        (N116)? \nz.mem [1021] : 
                        (N118)? \nz.mem [1071] : 
                        (N120)? \nz.mem [1121] : 
                        (N122)? \nz.mem [1171] : 
                        (N124)? \nz.mem [1221] : 
                        (N126)? \nz.mem [1271] : 
                        (N128)? \nz.mem [1321] : 
                        (N130)? \nz.mem [1371] : 
                        (N132)? \nz.mem [1421] : 
                        (N134)? \nz.mem [1471] : 
                        (N136)? \nz.mem [1521] : 
                        (N138)? \nz.mem [1571] : 
                        (N77)? \nz.mem [1621] : 
                        (N79)? \nz.mem [1671] : 
                        (N81)? \nz.mem [1721] : 
                        (N83)? \nz.mem [1771] : 
                        (N85)? \nz.mem [1821] : 
                        (N87)? \nz.mem [1871] : 
                        (N89)? \nz.mem [1921] : 
                        (N91)? \nz.mem [1971] : 
                        (N93)? \nz.mem [2021] : 
                        (N95)? \nz.mem [2071] : 
                        (N97)? \nz.mem [2121] : 
                        (N99)? \nz.mem [2171] : 
                        (N101)? \nz.mem [2221] : 
                        (N103)? \nz.mem [2271] : 
                        (N105)? \nz.mem [2321] : 
                        (N107)? \nz.mem [2371] : 
                        (N109)? \nz.mem [2421] : 
                        (N111)? \nz.mem [2471] : 
                        (N113)? \nz.mem [2521] : 
                        (N115)? \nz.mem [2571] : 
                        (N117)? \nz.mem [2621] : 
                        (N119)? \nz.mem [2671] : 
                        (N121)? \nz.mem [2721] : 
                        (N123)? \nz.mem [2771] : 
                        (N125)? \nz.mem [2821] : 
                        (N127)? \nz.mem [2871] : 
                        (N129)? \nz.mem [2921] : 
                        (N131)? \nz.mem [2971] : 
                        (N133)? \nz.mem [3021] : 
                        (N135)? \nz.mem [3071] : 
                        (N137)? \nz.mem [3121] : 
                        (N139)? \nz.mem [3171] : 1'b0;
  assign r_data_o[20] = (N76)? \nz.mem [20] : 
                        (N78)? \nz.mem [70] : 
                        (N80)? \nz.mem [120] : 
                        (N82)? \nz.mem [170] : 
                        (N84)? \nz.mem [220] : 
                        (N86)? \nz.mem [270] : 
                        (N88)? \nz.mem [320] : 
                        (N90)? \nz.mem [370] : 
                        (N92)? \nz.mem [420] : 
                        (N94)? \nz.mem [470] : 
                        (N96)? \nz.mem [520] : 
                        (N98)? \nz.mem [570] : 
                        (N100)? \nz.mem [620] : 
                        (N102)? \nz.mem [670] : 
                        (N104)? \nz.mem [720] : 
                        (N106)? \nz.mem [770] : 
                        (N108)? \nz.mem [820] : 
                        (N110)? \nz.mem [870] : 
                        (N112)? \nz.mem [920] : 
                        (N114)? \nz.mem [970] : 
                        (N116)? \nz.mem [1020] : 
                        (N118)? \nz.mem [1070] : 
                        (N120)? \nz.mem [1120] : 
                        (N122)? \nz.mem [1170] : 
                        (N124)? \nz.mem [1220] : 
                        (N126)? \nz.mem [1270] : 
                        (N128)? \nz.mem [1320] : 
                        (N130)? \nz.mem [1370] : 
                        (N132)? \nz.mem [1420] : 
                        (N134)? \nz.mem [1470] : 
                        (N136)? \nz.mem [1520] : 
                        (N138)? \nz.mem [1570] : 
                        (N77)? \nz.mem [1620] : 
                        (N79)? \nz.mem [1670] : 
                        (N81)? \nz.mem [1720] : 
                        (N83)? \nz.mem [1770] : 
                        (N85)? \nz.mem [1820] : 
                        (N87)? \nz.mem [1870] : 
                        (N89)? \nz.mem [1920] : 
                        (N91)? \nz.mem [1970] : 
                        (N93)? \nz.mem [2020] : 
                        (N95)? \nz.mem [2070] : 
                        (N97)? \nz.mem [2120] : 
                        (N99)? \nz.mem [2170] : 
                        (N101)? \nz.mem [2220] : 
                        (N103)? \nz.mem [2270] : 
                        (N105)? \nz.mem [2320] : 
                        (N107)? \nz.mem [2370] : 
                        (N109)? \nz.mem [2420] : 
                        (N111)? \nz.mem [2470] : 
                        (N113)? \nz.mem [2520] : 
                        (N115)? \nz.mem [2570] : 
                        (N117)? \nz.mem [2620] : 
                        (N119)? \nz.mem [2670] : 
                        (N121)? \nz.mem [2720] : 
                        (N123)? \nz.mem [2770] : 
                        (N125)? \nz.mem [2820] : 
                        (N127)? \nz.mem [2870] : 
                        (N129)? \nz.mem [2920] : 
                        (N131)? \nz.mem [2970] : 
                        (N133)? \nz.mem [3020] : 
                        (N135)? \nz.mem [3070] : 
                        (N137)? \nz.mem [3120] : 
                        (N139)? \nz.mem [3170] : 1'b0;
  assign r_data_o[19] = (N76)? \nz.mem [19] : 
                        (N78)? \nz.mem [69] : 
                        (N80)? \nz.mem [119] : 
                        (N82)? \nz.mem [169] : 
                        (N84)? \nz.mem [219] : 
                        (N86)? \nz.mem [269] : 
                        (N88)? \nz.mem [319] : 
                        (N90)? \nz.mem [369] : 
                        (N92)? \nz.mem [419] : 
                        (N94)? \nz.mem [469] : 
                        (N96)? \nz.mem [519] : 
                        (N98)? \nz.mem [569] : 
                        (N100)? \nz.mem [619] : 
                        (N102)? \nz.mem [669] : 
                        (N104)? \nz.mem [719] : 
                        (N106)? \nz.mem [769] : 
                        (N108)? \nz.mem [819] : 
                        (N110)? \nz.mem [869] : 
                        (N112)? \nz.mem [919] : 
                        (N114)? \nz.mem [969] : 
                        (N116)? \nz.mem [1019] : 
                        (N118)? \nz.mem [1069] : 
                        (N120)? \nz.mem [1119] : 
                        (N122)? \nz.mem [1169] : 
                        (N124)? \nz.mem [1219] : 
                        (N126)? \nz.mem [1269] : 
                        (N128)? \nz.mem [1319] : 
                        (N130)? \nz.mem [1369] : 
                        (N132)? \nz.mem [1419] : 
                        (N134)? \nz.mem [1469] : 
                        (N136)? \nz.mem [1519] : 
                        (N138)? \nz.mem [1569] : 
                        (N77)? \nz.mem [1619] : 
                        (N79)? \nz.mem [1669] : 
                        (N81)? \nz.mem [1719] : 
                        (N83)? \nz.mem [1769] : 
                        (N85)? \nz.mem [1819] : 
                        (N87)? \nz.mem [1869] : 
                        (N89)? \nz.mem [1919] : 
                        (N91)? \nz.mem [1969] : 
                        (N93)? \nz.mem [2019] : 
                        (N95)? \nz.mem [2069] : 
                        (N97)? \nz.mem [2119] : 
                        (N99)? \nz.mem [2169] : 
                        (N101)? \nz.mem [2219] : 
                        (N103)? \nz.mem [2269] : 
                        (N105)? \nz.mem [2319] : 
                        (N107)? \nz.mem [2369] : 
                        (N109)? \nz.mem [2419] : 
                        (N111)? \nz.mem [2469] : 
                        (N113)? \nz.mem [2519] : 
                        (N115)? \nz.mem [2569] : 
                        (N117)? \nz.mem [2619] : 
                        (N119)? \nz.mem [2669] : 
                        (N121)? \nz.mem [2719] : 
                        (N123)? \nz.mem [2769] : 
                        (N125)? \nz.mem [2819] : 
                        (N127)? \nz.mem [2869] : 
                        (N129)? \nz.mem [2919] : 
                        (N131)? \nz.mem [2969] : 
                        (N133)? \nz.mem [3019] : 
                        (N135)? \nz.mem [3069] : 
                        (N137)? \nz.mem [3119] : 
                        (N139)? \nz.mem [3169] : 1'b0;
  assign r_data_o[18] = (N76)? \nz.mem [18] : 
                        (N78)? \nz.mem [68] : 
                        (N80)? \nz.mem [118] : 
                        (N82)? \nz.mem [168] : 
                        (N84)? \nz.mem [218] : 
                        (N86)? \nz.mem [268] : 
                        (N88)? \nz.mem [318] : 
                        (N90)? \nz.mem [368] : 
                        (N92)? \nz.mem [418] : 
                        (N94)? \nz.mem [468] : 
                        (N96)? \nz.mem [518] : 
                        (N98)? \nz.mem [568] : 
                        (N100)? \nz.mem [618] : 
                        (N102)? \nz.mem [668] : 
                        (N104)? \nz.mem [718] : 
                        (N106)? \nz.mem [768] : 
                        (N108)? \nz.mem [818] : 
                        (N110)? \nz.mem [868] : 
                        (N112)? \nz.mem [918] : 
                        (N114)? \nz.mem [968] : 
                        (N116)? \nz.mem [1018] : 
                        (N118)? \nz.mem [1068] : 
                        (N120)? \nz.mem [1118] : 
                        (N122)? \nz.mem [1168] : 
                        (N124)? \nz.mem [1218] : 
                        (N126)? \nz.mem [1268] : 
                        (N128)? \nz.mem [1318] : 
                        (N130)? \nz.mem [1368] : 
                        (N132)? \nz.mem [1418] : 
                        (N134)? \nz.mem [1468] : 
                        (N136)? \nz.mem [1518] : 
                        (N138)? \nz.mem [1568] : 
                        (N77)? \nz.mem [1618] : 
                        (N79)? \nz.mem [1668] : 
                        (N81)? \nz.mem [1718] : 
                        (N83)? \nz.mem [1768] : 
                        (N85)? \nz.mem [1818] : 
                        (N87)? \nz.mem [1868] : 
                        (N89)? \nz.mem [1918] : 
                        (N91)? \nz.mem [1968] : 
                        (N93)? \nz.mem [2018] : 
                        (N95)? \nz.mem [2068] : 
                        (N97)? \nz.mem [2118] : 
                        (N99)? \nz.mem [2168] : 
                        (N101)? \nz.mem [2218] : 
                        (N103)? \nz.mem [2268] : 
                        (N105)? \nz.mem [2318] : 
                        (N107)? \nz.mem [2368] : 
                        (N109)? \nz.mem [2418] : 
                        (N111)? \nz.mem [2468] : 
                        (N113)? \nz.mem [2518] : 
                        (N115)? \nz.mem [2568] : 
                        (N117)? \nz.mem [2618] : 
                        (N119)? \nz.mem [2668] : 
                        (N121)? \nz.mem [2718] : 
                        (N123)? \nz.mem [2768] : 
                        (N125)? \nz.mem [2818] : 
                        (N127)? \nz.mem [2868] : 
                        (N129)? \nz.mem [2918] : 
                        (N131)? \nz.mem [2968] : 
                        (N133)? \nz.mem [3018] : 
                        (N135)? \nz.mem [3068] : 
                        (N137)? \nz.mem [3118] : 
                        (N139)? \nz.mem [3168] : 1'b0;
  assign r_data_o[17] = (N76)? \nz.mem [17] : 
                        (N78)? \nz.mem [67] : 
                        (N80)? \nz.mem [117] : 
                        (N82)? \nz.mem [167] : 
                        (N84)? \nz.mem [217] : 
                        (N86)? \nz.mem [267] : 
                        (N88)? \nz.mem [317] : 
                        (N90)? \nz.mem [367] : 
                        (N92)? \nz.mem [417] : 
                        (N94)? \nz.mem [467] : 
                        (N96)? \nz.mem [517] : 
                        (N98)? \nz.mem [567] : 
                        (N100)? \nz.mem [617] : 
                        (N102)? \nz.mem [667] : 
                        (N104)? \nz.mem [717] : 
                        (N106)? \nz.mem [767] : 
                        (N108)? \nz.mem [817] : 
                        (N110)? \nz.mem [867] : 
                        (N112)? \nz.mem [917] : 
                        (N114)? \nz.mem [967] : 
                        (N116)? \nz.mem [1017] : 
                        (N118)? \nz.mem [1067] : 
                        (N120)? \nz.mem [1117] : 
                        (N122)? \nz.mem [1167] : 
                        (N124)? \nz.mem [1217] : 
                        (N126)? \nz.mem [1267] : 
                        (N128)? \nz.mem [1317] : 
                        (N130)? \nz.mem [1367] : 
                        (N132)? \nz.mem [1417] : 
                        (N134)? \nz.mem [1467] : 
                        (N136)? \nz.mem [1517] : 
                        (N138)? \nz.mem [1567] : 
                        (N77)? \nz.mem [1617] : 
                        (N79)? \nz.mem [1667] : 
                        (N81)? \nz.mem [1717] : 
                        (N83)? \nz.mem [1767] : 
                        (N85)? \nz.mem [1817] : 
                        (N87)? \nz.mem [1867] : 
                        (N89)? \nz.mem [1917] : 
                        (N91)? \nz.mem [1967] : 
                        (N93)? \nz.mem [2017] : 
                        (N95)? \nz.mem [2067] : 
                        (N97)? \nz.mem [2117] : 
                        (N99)? \nz.mem [2167] : 
                        (N101)? \nz.mem [2217] : 
                        (N103)? \nz.mem [2267] : 
                        (N105)? \nz.mem [2317] : 
                        (N107)? \nz.mem [2367] : 
                        (N109)? \nz.mem [2417] : 
                        (N111)? \nz.mem [2467] : 
                        (N113)? \nz.mem [2517] : 
                        (N115)? \nz.mem [2567] : 
                        (N117)? \nz.mem [2617] : 
                        (N119)? \nz.mem [2667] : 
                        (N121)? \nz.mem [2717] : 
                        (N123)? \nz.mem [2767] : 
                        (N125)? \nz.mem [2817] : 
                        (N127)? \nz.mem [2867] : 
                        (N129)? \nz.mem [2917] : 
                        (N131)? \nz.mem [2967] : 
                        (N133)? \nz.mem [3017] : 
                        (N135)? \nz.mem [3067] : 
                        (N137)? \nz.mem [3117] : 
                        (N139)? \nz.mem [3167] : 1'b0;
  assign r_data_o[16] = (N76)? \nz.mem [16] : 
                        (N78)? \nz.mem [66] : 
                        (N80)? \nz.mem [116] : 
                        (N82)? \nz.mem [166] : 
                        (N84)? \nz.mem [216] : 
                        (N86)? \nz.mem [266] : 
                        (N88)? \nz.mem [316] : 
                        (N90)? \nz.mem [366] : 
                        (N92)? \nz.mem [416] : 
                        (N94)? \nz.mem [466] : 
                        (N96)? \nz.mem [516] : 
                        (N98)? \nz.mem [566] : 
                        (N100)? \nz.mem [616] : 
                        (N102)? \nz.mem [666] : 
                        (N104)? \nz.mem [716] : 
                        (N106)? \nz.mem [766] : 
                        (N108)? \nz.mem [816] : 
                        (N110)? \nz.mem [866] : 
                        (N112)? \nz.mem [916] : 
                        (N114)? \nz.mem [966] : 
                        (N116)? \nz.mem [1016] : 
                        (N118)? \nz.mem [1066] : 
                        (N120)? \nz.mem [1116] : 
                        (N122)? \nz.mem [1166] : 
                        (N124)? \nz.mem [1216] : 
                        (N126)? \nz.mem [1266] : 
                        (N128)? \nz.mem [1316] : 
                        (N130)? \nz.mem [1366] : 
                        (N132)? \nz.mem [1416] : 
                        (N134)? \nz.mem [1466] : 
                        (N136)? \nz.mem [1516] : 
                        (N138)? \nz.mem [1566] : 
                        (N77)? \nz.mem [1616] : 
                        (N79)? \nz.mem [1666] : 
                        (N81)? \nz.mem [1716] : 
                        (N83)? \nz.mem [1766] : 
                        (N85)? \nz.mem [1816] : 
                        (N87)? \nz.mem [1866] : 
                        (N89)? \nz.mem [1916] : 
                        (N91)? \nz.mem [1966] : 
                        (N93)? \nz.mem [2016] : 
                        (N95)? \nz.mem [2066] : 
                        (N97)? \nz.mem [2116] : 
                        (N99)? \nz.mem [2166] : 
                        (N101)? \nz.mem [2216] : 
                        (N103)? \nz.mem [2266] : 
                        (N105)? \nz.mem [2316] : 
                        (N107)? \nz.mem [2366] : 
                        (N109)? \nz.mem [2416] : 
                        (N111)? \nz.mem [2466] : 
                        (N113)? \nz.mem [2516] : 
                        (N115)? \nz.mem [2566] : 
                        (N117)? \nz.mem [2616] : 
                        (N119)? \nz.mem [2666] : 
                        (N121)? \nz.mem [2716] : 
                        (N123)? \nz.mem [2766] : 
                        (N125)? \nz.mem [2816] : 
                        (N127)? \nz.mem [2866] : 
                        (N129)? \nz.mem [2916] : 
                        (N131)? \nz.mem [2966] : 
                        (N133)? \nz.mem [3016] : 
                        (N135)? \nz.mem [3066] : 
                        (N137)? \nz.mem [3116] : 
                        (N139)? \nz.mem [3166] : 1'b0;
  assign r_data_o[15] = (N76)? \nz.mem [15] : 
                        (N78)? \nz.mem [65] : 
                        (N80)? \nz.mem [115] : 
                        (N82)? \nz.mem [165] : 
                        (N84)? \nz.mem [215] : 
                        (N86)? \nz.mem [265] : 
                        (N88)? \nz.mem [315] : 
                        (N90)? \nz.mem [365] : 
                        (N92)? \nz.mem [415] : 
                        (N94)? \nz.mem [465] : 
                        (N96)? \nz.mem [515] : 
                        (N98)? \nz.mem [565] : 
                        (N100)? \nz.mem [615] : 
                        (N102)? \nz.mem [665] : 
                        (N104)? \nz.mem [715] : 
                        (N106)? \nz.mem [765] : 
                        (N108)? \nz.mem [815] : 
                        (N110)? \nz.mem [865] : 
                        (N112)? \nz.mem [915] : 
                        (N114)? \nz.mem [965] : 
                        (N116)? \nz.mem [1015] : 
                        (N118)? \nz.mem [1065] : 
                        (N120)? \nz.mem [1115] : 
                        (N122)? \nz.mem [1165] : 
                        (N124)? \nz.mem [1215] : 
                        (N126)? \nz.mem [1265] : 
                        (N128)? \nz.mem [1315] : 
                        (N130)? \nz.mem [1365] : 
                        (N132)? \nz.mem [1415] : 
                        (N134)? \nz.mem [1465] : 
                        (N136)? \nz.mem [1515] : 
                        (N138)? \nz.mem [1565] : 
                        (N77)? \nz.mem [1615] : 
                        (N79)? \nz.mem [1665] : 
                        (N81)? \nz.mem [1715] : 
                        (N83)? \nz.mem [1765] : 
                        (N85)? \nz.mem [1815] : 
                        (N87)? \nz.mem [1865] : 
                        (N89)? \nz.mem [1915] : 
                        (N91)? \nz.mem [1965] : 
                        (N93)? \nz.mem [2015] : 
                        (N95)? \nz.mem [2065] : 
                        (N97)? \nz.mem [2115] : 
                        (N99)? \nz.mem [2165] : 
                        (N101)? \nz.mem [2215] : 
                        (N103)? \nz.mem [2265] : 
                        (N105)? \nz.mem [2315] : 
                        (N107)? \nz.mem [2365] : 
                        (N109)? \nz.mem [2415] : 
                        (N111)? \nz.mem [2465] : 
                        (N113)? \nz.mem [2515] : 
                        (N115)? \nz.mem [2565] : 
                        (N117)? \nz.mem [2615] : 
                        (N119)? \nz.mem [2665] : 
                        (N121)? \nz.mem [2715] : 
                        (N123)? \nz.mem [2765] : 
                        (N125)? \nz.mem [2815] : 
                        (N127)? \nz.mem [2865] : 
                        (N129)? \nz.mem [2915] : 
                        (N131)? \nz.mem [2965] : 
                        (N133)? \nz.mem [3015] : 
                        (N135)? \nz.mem [3065] : 
                        (N137)? \nz.mem [3115] : 
                        (N139)? \nz.mem [3165] : 1'b0;
  assign r_data_o[14] = (N76)? \nz.mem [14] : 
                        (N78)? \nz.mem [64] : 
                        (N80)? \nz.mem [114] : 
                        (N82)? \nz.mem [164] : 
                        (N84)? \nz.mem [214] : 
                        (N86)? \nz.mem [264] : 
                        (N88)? \nz.mem [314] : 
                        (N90)? \nz.mem [364] : 
                        (N92)? \nz.mem [414] : 
                        (N94)? \nz.mem [464] : 
                        (N96)? \nz.mem [514] : 
                        (N98)? \nz.mem [564] : 
                        (N100)? \nz.mem [614] : 
                        (N102)? \nz.mem [664] : 
                        (N104)? \nz.mem [714] : 
                        (N106)? \nz.mem [764] : 
                        (N108)? \nz.mem [814] : 
                        (N110)? \nz.mem [864] : 
                        (N112)? \nz.mem [914] : 
                        (N114)? \nz.mem [964] : 
                        (N116)? \nz.mem [1014] : 
                        (N118)? \nz.mem [1064] : 
                        (N120)? \nz.mem [1114] : 
                        (N122)? \nz.mem [1164] : 
                        (N124)? \nz.mem [1214] : 
                        (N126)? \nz.mem [1264] : 
                        (N128)? \nz.mem [1314] : 
                        (N130)? \nz.mem [1364] : 
                        (N132)? \nz.mem [1414] : 
                        (N134)? \nz.mem [1464] : 
                        (N136)? \nz.mem [1514] : 
                        (N138)? \nz.mem [1564] : 
                        (N77)? \nz.mem [1614] : 
                        (N79)? \nz.mem [1664] : 
                        (N81)? \nz.mem [1714] : 
                        (N83)? \nz.mem [1764] : 
                        (N85)? \nz.mem [1814] : 
                        (N87)? \nz.mem [1864] : 
                        (N89)? \nz.mem [1914] : 
                        (N91)? \nz.mem [1964] : 
                        (N93)? \nz.mem [2014] : 
                        (N95)? \nz.mem [2064] : 
                        (N97)? \nz.mem [2114] : 
                        (N99)? \nz.mem [2164] : 
                        (N101)? \nz.mem [2214] : 
                        (N103)? \nz.mem [2264] : 
                        (N105)? \nz.mem [2314] : 
                        (N107)? \nz.mem [2364] : 
                        (N109)? \nz.mem [2414] : 
                        (N111)? \nz.mem [2464] : 
                        (N113)? \nz.mem [2514] : 
                        (N115)? \nz.mem [2564] : 
                        (N117)? \nz.mem [2614] : 
                        (N119)? \nz.mem [2664] : 
                        (N121)? \nz.mem [2714] : 
                        (N123)? \nz.mem [2764] : 
                        (N125)? \nz.mem [2814] : 
                        (N127)? \nz.mem [2864] : 
                        (N129)? \nz.mem [2914] : 
                        (N131)? \nz.mem [2964] : 
                        (N133)? \nz.mem [3014] : 
                        (N135)? \nz.mem [3064] : 
                        (N137)? \nz.mem [3114] : 
                        (N139)? \nz.mem [3164] : 1'b0;
  assign r_data_o[13] = (N76)? \nz.mem [13] : 
                        (N78)? \nz.mem [63] : 
                        (N80)? \nz.mem [113] : 
                        (N82)? \nz.mem [163] : 
                        (N84)? \nz.mem [213] : 
                        (N86)? \nz.mem [263] : 
                        (N88)? \nz.mem [313] : 
                        (N90)? \nz.mem [363] : 
                        (N92)? \nz.mem [413] : 
                        (N94)? \nz.mem [463] : 
                        (N96)? \nz.mem [513] : 
                        (N98)? \nz.mem [563] : 
                        (N100)? \nz.mem [613] : 
                        (N102)? \nz.mem [663] : 
                        (N104)? \nz.mem [713] : 
                        (N106)? \nz.mem [763] : 
                        (N108)? \nz.mem [813] : 
                        (N110)? \nz.mem [863] : 
                        (N112)? \nz.mem [913] : 
                        (N114)? \nz.mem [963] : 
                        (N116)? \nz.mem [1013] : 
                        (N118)? \nz.mem [1063] : 
                        (N120)? \nz.mem [1113] : 
                        (N122)? \nz.mem [1163] : 
                        (N124)? \nz.mem [1213] : 
                        (N126)? \nz.mem [1263] : 
                        (N128)? \nz.mem [1313] : 
                        (N130)? \nz.mem [1363] : 
                        (N132)? \nz.mem [1413] : 
                        (N134)? \nz.mem [1463] : 
                        (N136)? \nz.mem [1513] : 
                        (N138)? \nz.mem [1563] : 
                        (N77)? \nz.mem [1613] : 
                        (N79)? \nz.mem [1663] : 
                        (N81)? \nz.mem [1713] : 
                        (N83)? \nz.mem [1763] : 
                        (N85)? \nz.mem [1813] : 
                        (N87)? \nz.mem [1863] : 
                        (N89)? \nz.mem [1913] : 
                        (N91)? \nz.mem [1963] : 
                        (N93)? \nz.mem [2013] : 
                        (N95)? \nz.mem [2063] : 
                        (N97)? \nz.mem [2113] : 
                        (N99)? \nz.mem [2163] : 
                        (N101)? \nz.mem [2213] : 
                        (N103)? \nz.mem [2263] : 
                        (N105)? \nz.mem [2313] : 
                        (N107)? \nz.mem [2363] : 
                        (N109)? \nz.mem [2413] : 
                        (N111)? \nz.mem [2463] : 
                        (N113)? \nz.mem [2513] : 
                        (N115)? \nz.mem [2563] : 
                        (N117)? \nz.mem [2613] : 
                        (N119)? \nz.mem [2663] : 
                        (N121)? \nz.mem [2713] : 
                        (N123)? \nz.mem [2763] : 
                        (N125)? \nz.mem [2813] : 
                        (N127)? \nz.mem [2863] : 
                        (N129)? \nz.mem [2913] : 
                        (N131)? \nz.mem [2963] : 
                        (N133)? \nz.mem [3013] : 
                        (N135)? \nz.mem [3063] : 
                        (N137)? \nz.mem [3113] : 
                        (N139)? \nz.mem [3163] : 1'b0;
  assign r_data_o[12] = (N76)? \nz.mem [12] : 
                        (N78)? \nz.mem [62] : 
                        (N80)? \nz.mem [112] : 
                        (N82)? \nz.mem [162] : 
                        (N84)? \nz.mem [212] : 
                        (N86)? \nz.mem [262] : 
                        (N88)? \nz.mem [312] : 
                        (N90)? \nz.mem [362] : 
                        (N92)? \nz.mem [412] : 
                        (N94)? \nz.mem [462] : 
                        (N96)? \nz.mem [512] : 
                        (N98)? \nz.mem [562] : 
                        (N100)? \nz.mem [612] : 
                        (N102)? \nz.mem [662] : 
                        (N104)? \nz.mem [712] : 
                        (N106)? \nz.mem [762] : 
                        (N108)? \nz.mem [812] : 
                        (N110)? \nz.mem [862] : 
                        (N112)? \nz.mem [912] : 
                        (N114)? \nz.mem [962] : 
                        (N116)? \nz.mem [1012] : 
                        (N118)? \nz.mem [1062] : 
                        (N120)? \nz.mem [1112] : 
                        (N122)? \nz.mem [1162] : 
                        (N124)? \nz.mem [1212] : 
                        (N126)? \nz.mem [1262] : 
                        (N128)? \nz.mem [1312] : 
                        (N130)? \nz.mem [1362] : 
                        (N132)? \nz.mem [1412] : 
                        (N134)? \nz.mem [1462] : 
                        (N136)? \nz.mem [1512] : 
                        (N138)? \nz.mem [1562] : 
                        (N77)? \nz.mem [1612] : 
                        (N79)? \nz.mem [1662] : 
                        (N81)? \nz.mem [1712] : 
                        (N83)? \nz.mem [1762] : 
                        (N85)? \nz.mem [1812] : 
                        (N87)? \nz.mem [1862] : 
                        (N89)? \nz.mem [1912] : 
                        (N91)? \nz.mem [1962] : 
                        (N93)? \nz.mem [2012] : 
                        (N95)? \nz.mem [2062] : 
                        (N97)? \nz.mem [2112] : 
                        (N99)? \nz.mem [2162] : 
                        (N101)? \nz.mem [2212] : 
                        (N103)? \nz.mem [2262] : 
                        (N105)? \nz.mem [2312] : 
                        (N107)? \nz.mem [2362] : 
                        (N109)? \nz.mem [2412] : 
                        (N111)? \nz.mem [2462] : 
                        (N113)? \nz.mem [2512] : 
                        (N115)? \nz.mem [2562] : 
                        (N117)? \nz.mem [2612] : 
                        (N119)? \nz.mem [2662] : 
                        (N121)? \nz.mem [2712] : 
                        (N123)? \nz.mem [2762] : 
                        (N125)? \nz.mem [2812] : 
                        (N127)? \nz.mem [2862] : 
                        (N129)? \nz.mem [2912] : 
                        (N131)? \nz.mem [2962] : 
                        (N133)? \nz.mem [3012] : 
                        (N135)? \nz.mem [3062] : 
                        (N137)? \nz.mem [3112] : 
                        (N139)? \nz.mem [3162] : 1'b0;
  assign r_data_o[11] = (N76)? \nz.mem [11] : 
                        (N78)? \nz.mem [61] : 
                        (N80)? \nz.mem [111] : 
                        (N82)? \nz.mem [161] : 
                        (N84)? \nz.mem [211] : 
                        (N86)? \nz.mem [261] : 
                        (N88)? \nz.mem [311] : 
                        (N90)? \nz.mem [361] : 
                        (N92)? \nz.mem [411] : 
                        (N94)? \nz.mem [461] : 
                        (N96)? \nz.mem [511] : 
                        (N98)? \nz.mem [561] : 
                        (N100)? \nz.mem [611] : 
                        (N102)? \nz.mem [661] : 
                        (N104)? \nz.mem [711] : 
                        (N106)? \nz.mem [761] : 
                        (N108)? \nz.mem [811] : 
                        (N110)? \nz.mem [861] : 
                        (N112)? \nz.mem [911] : 
                        (N114)? \nz.mem [961] : 
                        (N116)? \nz.mem [1011] : 
                        (N118)? \nz.mem [1061] : 
                        (N120)? \nz.mem [1111] : 
                        (N122)? \nz.mem [1161] : 
                        (N124)? \nz.mem [1211] : 
                        (N126)? \nz.mem [1261] : 
                        (N128)? \nz.mem [1311] : 
                        (N130)? \nz.mem [1361] : 
                        (N132)? \nz.mem [1411] : 
                        (N134)? \nz.mem [1461] : 
                        (N136)? \nz.mem [1511] : 
                        (N138)? \nz.mem [1561] : 
                        (N77)? \nz.mem [1611] : 
                        (N79)? \nz.mem [1661] : 
                        (N81)? \nz.mem [1711] : 
                        (N83)? \nz.mem [1761] : 
                        (N85)? \nz.mem [1811] : 
                        (N87)? \nz.mem [1861] : 
                        (N89)? \nz.mem [1911] : 
                        (N91)? \nz.mem [1961] : 
                        (N93)? \nz.mem [2011] : 
                        (N95)? \nz.mem [2061] : 
                        (N97)? \nz.mem [2111] : 
                        (N99)? \nz.mem [2161] : 
                        (N101)? \nz.mem [2211] : 
                        (N103)? \nz.mem [2261] : 
                        (N105)? \nz.mem [2311] : 
                        (N107)? \nz.mem [2361] : 
                        (N109)? \nz.mem [2411] : 
                        (N111)? \nz.mem [2461] : 
                        (N113)? \nz.mem [2511] : 
                        (N115)? \nz.mem [2561] : 
                        (N117)? \nz.mem [2611] : 
                        (N119)? \nz.mem [2661] : 
                        (N121)? \nz.mem [2711] : 
                        (N123)? \nz.mem [2761] : 
                        (N125)? \nz.mem [2811] : 
                        (N127)? \nz.mem [2861] : 
                        (N129)? \nz.mem [2911] : 
                        (N131)? \nz.mem [2961] : 
                        (N133)? \nz.mem [3011] : 
                        (N135)? \nz.mem [3061] : 
                        (N137)? \nz.mem [3111] : 
                        (N139)? \nz.mem [3161] : 1'b0;
  assign r_data_o[10] = (N76)? \nz.mem [10] : 
                        (N78)? \nz.mem [60] : 
                        (N80)? \nz.mem [110] : 
                        (N82)? \nz.mem [160] : 
                        (N84)? \nz.mem [210] : 
                        (N86)? \nz.mem [260] : 
                        (N88)? \nz.mem [310] : 
                        (N90)? \nz.mem [360] : 
                        (N92)? \nz.mem [410] : 
                        (N94)? \nz.mem [460] : 
                        (N96)? \nz.mem [510] : 
                        (N98)? \nz.mem [560] : 
                        (N100)? \nz.mem [610] : 
                        (N102)? \nz.mem [660] : 
                        (N104)? \nz.mem [710] : 
                        (N106)? \nz.mem [760] : 
                        (N108)? \nz.mem [810] : 
                        (N110)? \nz.mem [860] : 
                        (N112)? \nz.mem [910] : 
                        (N114)? \nz.mem [960] : 
                        (N116)? \nz.mem [1010] : 
                        (N118)? \nz.mem [1060] : 
                        (N120)? \nz.mem [1110] : 
                        (N122)? \nz.mem [1160] : 
                        (N124)? \nz.mem [1210] : 
                        (N126)? \nz.mem [1260] : 
                        (N128)? \nz.mem [1310] : 
                        (N130)? \nz.mem [1360] : 
                        (N132)? \nz.mem [1410] : 
                        (N134)? \nz.mem [1460] : 
                        (N136)? \nz.mem [1510] : 
                        (N138)? \nz.mem [1560] : 
                        (N77)? \nz.mem [1610] : 
                        (N79)? \nz.mem [1660] : 
                        (N81)? \nz.mem [1710] : 
                        (N83)? \nz.mem [1760] : 
                        (N85)? \nz.mem [1810] : 
                        (N87)? \nz.mem [1860] : 
                        (N89)? \nz.mem [1910] : 
                        (N91)? \nz.mem [1960] : 
                        (N93)? \nz.mem [2010] : 
                        (N95)? \nz.mem [2060] : 
                        (N97)? \nz.mem [2110] : 
                        (N99)? \nz.mem [2160] : 
                        (N101)? \nz.mem [2210] : 
                        (N103)? \nz.mem [2260] : 
                        (N105)? \nz.mem [2310] : 
                        (N107)? \nz.mem [2360] : 
                        (N109)? \nz.mem [2410] : 
                        (N111)? \nz.mem [2460] : 
                        (N113)? \nz.mem [2510] : 
                        (N115)? \nz.mem [2560] : 
                        (N117)? \nz.mem [2610] : 
                        (N119)? \nz.mem [2660] : 
                        (N121)? \nz.mem [2710] : 
                        (N123)? \nz.mem [2760] : 
                        (N125)? \nz.mem [2810] : 
                        (N127)? \nz.mem [2860] : 
                        (N129)? \nz.mem [2910] : 
                        (N131)? \nz.mem [2960] : 
                        (N133)? \nz.mem [3010] : 
                        (N135)? \nz.mem [3060] : 
                        (N137)? \nz.mem [3110] : 
                        (N139)? \nz.mem [3160] : 1'b0;
  assign r_data_o[9] = (N76)? \nz.mem [9] : 
                       (N78)? \nz.mem [59] : 
                       (N80)? \nz.mem [109] : 
                       (N82)? \nz.mem [159] : 
                       (N84)? \nz.mem [209] : 
                       (N86)? \nz.mem [259] : 
                       (N88)? \nz.mem [309] : 
                       (N90)? \nz.mem [359] : 
                       (N92)? \nz.mem [409] : 
                       (N94)? \nz.mem [459] : 
                       (N96)? \nz.mem [509] : 
                       (N98)? \nz.mem [559] : 
                       (N100)? \nz.mem [609] : 
                       (N102)? \nz.mem [659] : 
                       (N104)? \nz.mem [709] : 
                       (N106)? \nz.mem [759] : 
                       (N108)? \nz.mem [809] : 
                       (N110)? \nz.mem [859] : 
                       (N112)? \nz.mem [909] : 
                       (N114)? \nz.mem [959] : 
                       (N116)? \nz.mem [1009] : 
                       (N118)? \nz.mem [1059] : 
                       (N120)? \nz.mem [1109] : 
                       (N122)? \nz.mem [1159] : 
                       (N124)? \nz.mem [1209] : 
                       (N126)? \nz.mem [1259] : 
                       (N128)? \nz.mem [1309] : 
                       (N130)? \nz.mem [1359] : 
                       (N132)? \nz.mem [1409] : 
                       (N134)? \nz.mem [1459] : 
                       (N136)? \nz.mem [1509] : 
                       (N138)? \nz.mem [1559] : 
                       (N77)? \nz.mem [1609] : 
                       (N79)? \nz.mem [1659] : 
                       (N81)? \nz.mem [1709] : 
                       (N83)? \nz.mem [1759] : 
                       (N85)? \nz.mem [1809] : 
                       (N87)? \nz.mem [1859] : 
                       (N89)? \nz.mem [1909] : 
                       (N91)? \nz.mem [1959] : 
                       (N93)? \nz.mem [2009] : 
                       (N95)? \nz.mem [2059] : 
                       (N97)? \nz.mem [2109] : 
                       (N99)? \nz.mem [2159] : 
                       (N101)? \nz.mem [2209] : 
                       (N103)? \nz.mem [2259] : 
                       (N105)? \nz.mem [2309] : 
                       (N107)? \nz.mem [2359] : 
                       (N109)? \nz.mem [2409] : 
                       (N111)? \nz.mem [2459] : 
                       (N113)? \nz.mem [2509] : 
                       (N115)? \nz.mem [2559] : 
                       (N117)? \nz.mem [2609] : 
                       (N119)? \nz.mem [2659] : 
                       (N121)? \nz.mem [2709] : 
                       (N123)? \nz.mem [2759] : 
                       (N125)? \nz.mem [2809] : 
                       (N127)? \nz.mem [2859] : 
                       (N129)? \nz.mem [2909] : 
                       (N131)? \nz.mem [2959] : 
                       (N133)? \nz.mem [3009] : 
                       (N135)? \nz.mem [3059] : 
                       (N137)? \nz.mem [3109] : 
                       (N139)? \nz.mem [3159] : 1'b0;
  assign r_data_o[8] = (N76)? \nz.mem [8] : 
                       (N78)? \nz.mem [58] : 
                       (N80)? \nz.mem [108] : 
                       (N82)? \nz.mem [158] : 
                       (N84)? \nz.mem [208] : 
                       (N86)? \nz.mem [258] : 
                       (N88)? \nz.mem [308] : 
                       (N90)? \nz.mem [358] : 
                       (N92)? \nz.mem [408] : 
                       (N94)? \nz.mem [458] : 
                       (N96)? \nz.mem [508] : 
                       (N98)? \nz.mem [558] : 
                       (N100)? \nz.mem [608] : 
                       (N102)? \nz.mem [658] : 
                       (N104)? \nz.mem [708] : 
                       (N106)? \nz.mem [758] : 
                       (N108)? \nz.mem [808] : 
                       (N110)? \nz.mem [858] : 
                       (N112)? \nz.mem [908] : 
                       (N114)? \nz.mem [958] : 
                       (N116)? \nz.mem [1008] : 
                       (N118)? \nz.mem [1058] : 
                       (N120)? \nz.mem [1108] : 
                       (N122)? \nz.mem [1158] : 
                       (N124)? \nz.mem [1208] : 
                       (N126)? \nz.mem [1258] : 
                       (N128)? \nz.mem [1308] : 
                       (N130)? \nz.mem [1358] : 
                       (N132)? \nz.mem [1408] : 
                       (N134)? \nz.mem [1458] : 
                       (N136)? \nz.mem [1508] : 
                       (N138)? \nz.mem [1558] : 
                       (N77)? \nz.mem [1608] : 
                       (N79)? \nz.mem [1658] : 
                       (N81)? \nz.mem [1708] : 
                       (N83)? \nz.mem [1758] : 
                       (N85)? \nz.mem [1808] : 
                       (N87)? \nz.mem [1858] : 
                       (N89)? \nz.mem [1908] : 
                       (N91)? \nz.mem [1958] : 
                       (N93)? \nz.mem [2008] : 
                       (N95)? \nz.mem [2058] : 
                       (N97)? \nz.mem [2108] : 
                       (N99)? \nz.mem [2158] : 
                       (N101)? \nz.mem [2208] : 
                       (N103)? \nz.mem [2258] : 
                       (N105)? \nz.mem [2308] : 
                       (N107)? \nz.mem [2358] : 
                       (N109)? \nz.mem [2408] : 
                       (N111)? \nz.mem [2458] : 
                       (N113)? \nz.mem [2508] : 
                       (N115)? \nz.mem [2558] : 
                       (N117)? \nz.mem [2608] : 
                       (N119)? \nz.mem [2658] : 
                       (N121)? \nz.mem [2708] : 
                       (N123)? \nz.mem [2758] : 
                       (N125)? \nz.mem [2808] : 
                       (N127)? \nz.mem [2858] : 
                       (N129)? \nz.mem [2908] : 
                       (N131)? \nz.mem [2958] : 
                       (N133)? \nz.mem [3008] : 
                       (N135)? \nz.mem [3058] : 
                       (N137)? \nz.mem [3108] : 
                       (N139)? \nz.mem [3158] : 1'b0;
  assign r_data_o[7] = (N76)? \nz.mem [7] : 
                       (N78)? \nz.mem [57] : 
                       (N80)? \nz.mem [107] : 
                       (N82)? \nz.mem [157] : 
                       (N84)? \nz.mem [207] : 
                       (N86)? \nz.mem [257] : 
                       (N88)? \nz.mem [307] : 
                       (N90)? \nz.mem [357] : 
                       (N92)? \nz.mem [407] : 
                       (N94)? \nz.mem [457] : 
                       (N96)? \nz.mem [507] : 
                       (N98)? \nz.mem [557] : 
                       (N100)? \nz.mem [607] : 
                       (N102)? \nz.mem [657] : 
                       (N104)? \nz.mem [707] : 
                       (N106)? \nz.mem [757] : 
                       (N108)? \nz.mem [807] : 
                       (N110)? \nz.mem [857] : 
                       (N112)? \nz.mem [907] : 
                       (N114)? \nz.mem [957] : 
                       (N116)? \nz.mem [1007] : 
                       (N118)? \nz.mem [1057] : 
                       (N120)? \nz.mem [1107] : 
                       (N122)? \nz.mem [1157] : 
                       (N124)? \nz.mem [1207] : 
                       (N126)? \nz.mem [1257] : 
                       (N128)? \nz.mem [1307] : 
                       (N130)? \nz.mem [1357] : 
                       (N132)? \nz.mem [1407] : 
                       (N134)? \nz.mem [1457] : 
                       (N136)? \nz.mem [1507] : 
                       (N138)? \nz.mem [1557] : 
                       (N77)? \nz.mem [1607] : 
                       (N79)? \nz.mem [1657] : 
                       (N81)? \nz.mem [1707] : 
                       (N83)? \nz.mem [1757] : 
                       (N85)? \nz.mem [1807] : 
                       (N87)? \nz.mem [1857] : 
                       (N89)? \nz.mem [1907] : 
                       (N91)? \nz.mem [1957] : 
                       (N93)? \nz.mem [2007] : 
                       (N95)? \nz.mem [2057] : 
                       (N97)? \nz.mem [2107] : 
                       (N99)? \nz.mem [2157] : 
                       (N101)? \nz.mem [2207] : 
                       (N103)? \nz.mem [2257] : 
                       (N105)? \nz.mem [2307] : 
                       (N107)? \nz.mem [2357] : 
                       (N109)? \nz.mem [2407] : 
                       (N111)? \nz.mem [2457] : 
                       (N113)? \nz.mem [2507] : 
                       (N115)? \nz.mem [2557] : 
                       (N117)? \nz.mem [2607] : 
                       (N119)? \nz.mem [2657] : 
                       (N121)? \nz.mem [2707] : 
                       (N123)? \nz.mem [2757] : 
                       (N125)? \nz.mem [2807] : 
                       (N127)? \nz.mem [2857] : 
                       (N129)? \nz.mem [2907] : 
                       (N131)? \nz.mem [2957] : 
                       (N133)? \nz.mem [3007] : 
                       (N135)? \nz.mem [3057] : 
                       (N137)? \nz.mem [3107] : 
                       (N139)? \nz.mem [3157] : 1'b0;
  assign r_data_o[6] = (N76)? \nz.mem [6] : 
                       (N78)? \nz.mem [56] : 
                       (N80)? \nz.mem [106] : 
                       (N82)? \nz.mem [156] : 
                       (N84)? \nz.mem [206] : 
                       (N86)? \nz.mem [256] : 
                       (N88)? \nz.mem [306] : 
                       (N90)? \nz.mem [356] : 
                       (N92)? \nz.mem [406] : 
                       (N94)? \nz.mem [456] : 
                       (N96)? \nz.mem [506] : 
                       (N98)? \nz.mem [556] : 
                       (N100)? \nz.mem [606] : 
                       (N102)? \nz.mem [656] : 
                       (N104)? \nz.mem [706] : 
                       (N106)? \nz.mem [756] : 
                       (N108)? \nz.mem [806] : 
                       (N110)? \nz.mem [856] : 
                       (N112)? \nz.mem [906] : 
                       (N114)? \nz.mem [956] : 
                       (N116)? \nz.mem [1006] : 
                       (N118)? \nz.mem [1056] : 
                       (N120)? \nz.mem [1106] : 
                       (N122)? \nz.mem [1156] : 
                       (N124)? \nz.mem [1206] : 
                       (N126)? \nz.mem [1256] : 
                       (N128)? \nz.mem [1306] : 
                       (N130)? \nz.mem [1356] : 
                       (N132)? \nz.mem [1406] : 
                       (N134)? \nz.mem [1456] : 
                       (N136)? \nz.mem [1506] : 
                       (N138)? \nz.mem [1556] : 
                       (N77)? \nz.mem [1606] : 
                       (N79)? \nz.mem [1656] : 
                       (N81)? \nz.mem [1706] : 
                       (N83)? \nz.mem [1756] : 
                       (N85)? \nz.mem [1806] : 
                       (N87)? \nz.mem [1856] : 
                       (N89)? \nz.mem [1906] : 
                       (N91)? \nz.mem [1956] : 
                       (N93)? \nz.mem [2006] : 
                       (N95)? \nz.mem [2056] : 
                       (N97)? \nz.mem [2106] : 
                       (N99)? \nz.mem [2156] : 
                       (N101)? \nz.mem [2206] : 
                       (N103)? \nz.mem [2256] : 
                       (N105)? \nz.mem [2306] : 
                       (N107)? \nz.mem [2356] : 
                       (N109)? \nz.mem [2406] : 
                       (N111)? \nz.mem [2456] : 
                       (N113)? \nz.mem [2506] : 
                       (N115)? \nz.mem [2556] : 
                       (N117)? \nz.mem [2606] : 
                       (N119)? \nz.mem [2656] : 
                       (N121)? \nz.mem [2706] : 
                       (N123)? \nz.mem [2756] : 
                       (N125)? \nz.mem [2806] : 
                       (N127)? \nz.mem [2856] : 
                       (N129)? \nz.mem [2906] : 
                       (N131)? \nz.mem [2956] : 
                       (N133)? \nz.mem [3006] : 
                       (N135)? \nz.mem [3056] : 
                       (N137)? \nz.mem [3106] : 
                       (N139)? \nz.mem [3156] : 1'b0;
  assign r_data_o[5] = (N76)? \nz.mem [5] : 
                       (N78)? \nz.mem [55] : 
                       (N80)? \nz.mem [105] : 
                       (N82)? \nz.mem [155] : 
                       (N84)? \nz.mem [205] : 
                       (N86)? \nz.mem [255] : 
                       (N88)? \nz.mem [305] : 
                       (N90)? \nz.mem [355] : 
                       (N92)? \nz.mem [405] : 
                       (N94)? \nz.mem [455] : 
                       (N96)? \nz.mem [505] : 
                       (N98)? \nz.mem [555] : 
                       (N100)? \nz.mem [605] : 
                       (N102)? \nz.mem [655] : 
                       (N104)? \nz.mem [705] : 
                       (N106)? \nz.mem [755] : 
                       (N108)? \nz.mem [805] : 
                       (N110)? \nz.mem [855] : 
                       (N112)? \nz.mem [905] : 
                       (N114)? \nz.mem [955] : 
                       (N116)? \nz.mem [1005] : 
                       (N118)? \nz.mem [1055] : 
                       (N120)? \nz.mem [1105] : 
                       (N122)? \nz.mem [1155] : 
                       (N124)? \nz.mem [1205] : 
                       (N126)? \nz.mem [1255] : 
                       (N128)? \nz.mem [1305] : 
                       (N130)? \nz.mem [1355] : 
                       (N132)? \nz.mem [1405] : 
                       (N134)? \nz.mem [1455] : 
                       (N136)? \nz.mem [1505] : 
                       (N138)? \nz.mem [1555] : 
                       (N77)? \nz.mem [1605] : 
                       (N79)? \nz.mem [1655] : 
                       (N81)? \nz.mem [1705] : 
                       (N83)? \nz.mem [1755] : 
                       (N85)? \nz.mem [1805] : 
                       (N87)? \nz.mem [1855] : 
                       (N89)? \nz.mem [1905] : 
                       (N91)? \nz.mem [1955] : 
                       (N93)? \nz.mem [2005] : 
                       (N95)? \nz.mem [2055] : 
                       (N97)? \nz.mem [2105] : 
                       (N99)? \nz.mem [2155] : 
                       (N101)? \nz.mem [2205] : 
                       (N103)? \nz.mem [2255] : 
                       (N105)? \nz.mem [2305] : 
                       (N107)? \nz.mem [2355] : 
                       (N109)? \nz.mem [2405] : 
                       (N111)? \nz.mem [2455] : 
                       (N113)? \nz.mem [2505] : 
                       (N115)? \nz.mem [2555] : 
                       (N117)? \nz.mem [2605] : 
                       (N119)? \nz.mem [2655] : 
                       (N121)? \nz.mem [2705] : 
                       (N123)? \nz.mem [2755] : 
                       (N125)? \nz.mem [2805] : 
                       (N127)? \nz.mem [2855] : 
                       (N129)? \nz.mem [2905] : 
                       (N131)? \nz.mem [2955] : 
                       (N133)? \nz.mem [3005] : 
                       (N135)? \nz.mem [3055] : 
                       (N137)? \nz.mem [3105] : 
                       (N139)? \nz.mem [3155] : 1'b0;
  assign r_data_o[4] = (N76)? \nz.mem [4] : 
                       (N78)? \nz.mem [54] : 
                       (N80)? \nz.mem [104] : 
                       (N82)? \nz.mem [154] : 
                       (N84)? \nz.mem [204] : 
                       (N86)? \nz.mem [254] : 
                       (N88)? \nz.mem [304] : 
                       (N90)? \nz.mem [354] : 
                       (N92)? \nz.mem [404] : 
                       (N94)? \nz.mem [454] : 
                       (N96)? \nz.mem [504] : 
                       (N98)? \nz.mem [554] : 
                       (N100)? \nz.mem [604] : 
                       (N102)? \nz.mem [654] : 
                       (N104)? \nz.mem [704] : 
                       (N106)? \nz.mem [754] : 
                       (N108)? \nz.mem [804] : 
                       (N110)? \nz.mem [854] : 
                       (N112)? \nz.mem [904] : 
                       (N114)? \nz.mem [954] : 
                       (N116)? \nz.mem [1004] : 
                       (N118)? \nz.mem [1054] : 
                       (N120)? \nz.mem [1104] : 
                       (N122)? \nz.mem [1154] : 
                       (N124)? \nz.mem [1204] : 
                       (N126)? \nz.mem [1254] : 
                       (N128)? \nz.mem [1304] : 
                       (N130)? \nz.mem [1354] : 
                       (N132)? \nz.mem [1404] : 
                       (N134)? \nz.mem [1454] : 
                       (N136)? \nz.mem [1504] : 
                       (N138)? \nz.mem [1554] : 
                       (N77)? \nz.mem [1604] : 
                       (N79)? \nz.mem [1654] : 
                       (N81)? \nz.mem [1704] : 
                       (N83)? \nz.mem [1754] : 
                       (N85)? \nz.mem [1804] : 
                       (N87)? \nz.mem [1854] : 
                       (N89)? \nz.mem [1904] : 
                       (N91)? \nz.mem [1954] : 
                       (N93)? \nz.mem [2004] : 
                       (N95)? \nz.mem [2054] : 
                       (N97)? \nz.mem [2104] : 
                       (N99)? \nz.mem [2154] : 
                       (N101)? \nz.mem [2204] : 
                       (N103)? \nz.mem [2254] : 
                       (N105)? \nz.mem [2304] : 
                       (N107)? \nz.mem [2354] : 
                       (N109)? \nz.mem [2404] : 
                       (N111)? \nz.mem [2454] : 
                       (N113)? \nz.mem [2504] : 
                       (N115)? \nz.mem [2554] : 
                       (N117)? \nz.mem [2604] : 
                       (N119)? \nz.mem [2654] : 
                       (N121)? \nz.mem [2704] : 
                       (N123)? \nz.mem [2754] : 
                       (N125)? \nz.mem [2804] : 
                       (N127)? \nz.mem [2854] : 
                       (N129)? \nz.mem [2904] : 
                       (N131)? \nz.mem [2954] : 
                       (N133)? \nz.mem [3004] : 
                       (N135)? \nz.mem [3054] : 
                       (N137)? \nz.mem [3104] : 
                       (N139)? \nz.mem [3154] : 1'b0;
  assign r_data_o[3] = (N76)? \nz.mem [3] : 
                       (N78)? \nz.mem [53] : 
                       (N80)? \nz.mem [103] : 
                       (N82)? \nz.mem [153] : 
                       (N84)? \nz.mem [203] : 
                       (N86)? \nz.mem [253] : 
                       (N88)? \nz.mem [303] : 
                       (N90)? \nz.mem [353] : 
                       (N92)? \nz.mem [403] : 
                       (N94)? \nz.mem [453] : 
                       (N96)? \nz.mem [503] : 
                       (N98)? \nz.mem [553] : 
                       (N100)? \nz.mem [603] : 
                       (N102)? \nz.mem [653] : 
                       (N104)? \nz.mem [703] : 
                       (N106)? \nz.mem [753] : 
                       (N108)? \nz.mem [803] : 
                       (N110)? \nz.mem [853] : 
                       (N112)? \nz.mem [903] : 
                       (N114)? \nz.mem [953] : 
                       (N116)? \nz.mem [1003] : 
                       (N118)? \nz.mem [1053] : 
                       (N120)? \nz.mem [1103] : 
                       (N122)? \nz.mem [1153] : 
                       (N124)? \nz.mem [1203] : 
                       (N126)? \nz.mem [1253] : 
                       (N128)? \nz.mem [1303] : 
                       (N130)? \nz.mem [1353] : 
                       (N132)? \nz.mem [1403] : 
                       (N134)? \nz.mem [1453] : 
                       (N136)? \nz.mem [1503] : 
                       (N138)? \nz.mem [1553] : 
                       (N77)? \nz.mem [1603] : 
                       (N79)? \nz.mem [1653] : 
                       (N81)? \nz.mem [1703] : 
                       (N83)? \nz.mem [1753] : 
                       (N85)? \nz.mem [1803] : 
                       (N87)? \nz.mem [1853] : 
                       (N89)? \nz.mem [1903] : 
                       (N91)? \nz.mem [1953] : 
                       (N93)? \nz.mem [2003] : 
                       (N95)? \nz.mem [2053] : 
                       (N97)? \nz.mem [2103] : 
                       (N99)? \nz.mem [2153] : 
                       (N101)? \nz.mem [2203] : 
                       (N103)? \nz.mem [2253] : 
                       (N105)? \nz.mem [2303] : 
                       (N107)? \nz.mem [2353] : 
                       (N109)? \nz.mem [2403] : 
                       (N111)? \nz.mem [2453] : 
                       (N113)? \nz.mem [2503] : 
                       (N115)? \nz.mem [2553] : 
                       (N117)? \nz.mem [2603] : 
                       (N119)? \nz.mem [2653] : 
                       (N121)? \nz.mem [2703] : 
                       (N123)? \nz.mem [2753] : 
                       (N125)? \nz.mem [2803] : 
                       (N127)? \nz.mem [2853] : 
                       (N129)? \nz.mem [2903] : 
                       (N131)? \nz.mem [2953] : 
                       (N133)? \nz.mem [3003] : 
                       (N135)? \nz.mem [3053] : 
                       (N137)? \nz.mem [3103] : 
                       (N139)? \nz.mem [3153] : 1'b0;
  assign r_data_o[2] = (N76)? \nz.mem [2] : 
                       (N78)? \nz.mem [52] : 
                       (N80)? \nz.mem [102] : 
                       (N82)? \nz.mem [152] : 
                       (N84)? \nz.mem [202] : 
                       (N86)? \nz.mem [252] : 
                       (N88)? \nz.mem [302] : 
                       (N90)? \nz.mem [352] : 
                       (N92)? \nz.mem [402] : 
                       (N94)? \nz.mem [452] : 
                       (N96)? \nz.mem [502] : 
                       (N98)? \nz.mem [552] : 
                       (N100)? \nz.mem [602] : 
                       (N102)? \nz.mem [652] : 
                       (N104)? \nz.mem [702] : 
                       (N106)? \nz.mem [752] : 
                       (N108)? \nz.mem [802] : 
                       (N110)? \nz.mem [852] : 
                       (N112)? \nz.mem [902] : 
                       (N114)? \nz.mem [952] : 
                       (N116)? \nz.mem [1002] : 
                       (N118)? \nz.mem [1052] : 
                       (N120)? \nz.mem [1102] : 
                       (N122)? \nz.mem [1152] : 
                       (N124)? \nz.mem [1202] : 
                       (N126)? \nz.mem [1252] : 
                       (N128)? \nz.mem [1302] : 
                       (N130)? \nz.mem [1352] : 
                       (N132)? \nz.mem [1402] : 
                       (N134)? \nz.mem [1452] : 
                       (N136)? \nz.mem [1502] : 
                       (N138)? \nz.mem [1552] : 
                       (N77)? \nz.mem [1602] : 
                       (N79)? \nz.mem [1652] : 
                       (N81)? \nz.mem [1702] : 
                       (N83)? \nz.mem [1752] : 
                       (N85)? \nz.mem [1802] : 
                       (N87)? \nz.mem [1852] : 
                       (N89)? \nz.mem [1902] : 
                       (N91)? \nz.mem [1952] : 
                       (N93)? \nz.mem [2002] : 
                       (N95)? \nz.mem [2052] : 
                       (N97)? \nz.mem [2102] : 
                       (N99)? \nz.mem [2152] : 
                       (N101)? \nz.mem [2202] : 
                       (N103)? \nz.mem [2252] : 
                       (N105)? \nz.mem [2302] : 
                       (N107)? \nz.mem [2352] : 
                       (N109)? \nz.mem [2402] : 
                       (N111)? \nz.mem [2452] : 
                       (N113)? \nz.mem [2502] : 
                       (N115)? \nz.mem [2552] : 
                       (N117)? \nz.mem [2602] : 
                       (N119)? \nz.mem [2652] : 
                       (N121)? \nz.mem [2702] : 
                       (N123)? \nz.mem [2752] : 
                       (N125)? \nz.mem [2802] : 
                       (N127)? \nz.mem [2852] : 
                       (N129)? \nz.mem [2902] : 
                       (N131)? \nz.mem [2952] : 
                       (N133)? \nz.mem [3002] : 
                       (N135)? \nz.mem [3052] : 
                       (N137)? \nz.mem [3102] : 
                       (N139)? \nz.mem [3152] : 1'b0;
  assign r_data_o[1] = (N76)? \nz.mem [1] : 
                       (N78)? \nz.mem [51] : 
                       (N80)? \nz.mem [101] : 
                       (N82)? \nz.mem [151] : 
                       (N84)? \nz.mem [201] : 
                       (N86)? \nz.mem [251] : 
                       (N88)? \nz.mem [301] : 
                       (N90)? \nz.mem [351] : 
                       (N92)? \nz.mem [401] : 
                       (N94)? \nz.mem [451] : 
                       (N96)? \nz.mem [501] : 
                       (N98)? \nz.mem [551] : 
                       (N100)? \nz.mem [601] : 
                       (N102)? \nz.mem [651] : 
                       (N104)? \nz.mem [701] : 
                       (N106)? \nz.mem [751] : 
                       (N108)? \nz.mem [801] : 
                       (N110)? \nz.mem [851] : 
                       (N112)? \nz.mem [901] : 
                       (N114)? \nz.mem [951] : 
                       (N116)? \nz.mem [1001] : 
                       (N118)? \nz.mem [1051] : 
                       (N120)? \nz.mem [1101] : 
                       (N122)? \nz.mem [1151] : 
                       (N124)? \nz.mem [1201] : 
                       (N126)? \nz.mem [1251] : 
                       (N128)? \nz.mem [1301] : 
                       (N130)? \nz.mem [1351] : 
                       (N132)? \nz.mem [1401] : 
                       (N134)? \nz.mem [1451] : 
                       (N136)? \nz.mem [1501] : 
                       (N138)? \nz.mem [1551] : 
                       (N77)? \nz.mem [1601] : 
                       (N79)? \nz.mem [1651] : 
                       (N81)? \nz.mem [1701] : 
                       (N83)? \nz.mem [1751] : 
                       (N85)? \nz.mem [1801] : 
                       (N87)? \nz.mem [1851] : 
                       (N89)? \nz.mem [1901] : 
                       (N91)? \nz.mem [1951] : 
                       (N93)? \nz.mem [2001] : 
                       (N95)? \nz.mem [2051] : 
                       (N97)? \nz.mem [2101] : 
                       (N99)? \nz.mem [2151] : 
                       (N101)? \nz.mem [2201] : 
                       (N103)? \nz.mem [2251] : 
                       (N105)? \nz.mem [2301] : 
                       (N107)? \nz.mem [2351] : 
                       (N109)? \nz.mem [2401] : 
                       (N111)? \nz.mem [2451] : 
                       (N113)? \nz.mem [2501] : 
                       (N115)? \nz.mem [2551] : 
                       (N117)? \nz.mem [2601] : 
                       (N119)? \nz.mem [2651] : 
                       (N121)? \nz.mem [2701] : 
                       (N123)? \nz.mem [2751] : 
                       (N125)? \nz.mem [2801] : 
                       (N127)? \nz.mem [2851] : 
                       (N129)? \nz.mem [2901] : 
                       (N131)? \nz.mem [2951] : 
                       (N133)? \nz.mem [3001] : 
                       (N135)? \nz.mem [3051] : 
                       (N137)? \nz.mem [3101] : 
                       (N139)? \nz.mem [3151] : 1'b0;
  assign r_data_o[0] = (N76)? \nz.mem [0] : 
                       (N78)? \nz.mem [50] : 
                       (N80)? \nz.mem [100] : 
                       (N82)? \nz.mem [150] : 
                       (N84)? \nz.mem [200] : 
                       (N86)? \nz.mem [250] : 
                       (N88)? \nz.mem [300] : 
                       (N90)? \nz.mem [350] : 
                       (N92)? \nz.mem [400] : 
                       (N94)? \nz.mem [450] : 
                       (N96)? \nz.mem [500] : 
                       (N98)? \nz.mem [550] : 
                       (N100)? \nz.mem [600] : 
                       (N102)? \nz.mem [650] : 
                       (N104)? \nz.mem [700] : 
                       (N106)? \nz.mem [750] : 
                       (N108)? \nz.mem [800] : 
                       (N110)? \nz.mem [850] : 
                       (N112)? \nz.mem [900] : 
                       (N114)? \nz.mem [950] : 
                       (N116)? \nz.mem [1000] : 
                       (N118)? \nz.mem [1050] : 
                       (N120)? \nz.mem [1100] : 
                       (N122)? \nz.mem [1150] : 
                       (N124)? \nz.mem [1200] : 
                       (N126)? \nz.mem [1250] : 
                       (N128)? \nz.mem [1300] : 
                       (N130)? \nz.mem [1350] : 
                       (N132)? \nz.mem [1400] : 
                       (N134)? \nz.mem [1450] : 
                       (N136)? \nz.mem [1500] : 
                       (N138)? \nz.mem [1550] : 
                       (N77)? \nz.mem [1600] : 
                       (N79)? \nz.mem [1650] : 
                       (N81)? \nz.mem [1700] : 
                       (N83)? \nz.mem [1750] : 
                       (N85)? \nz.mem [1800] : 
                       (N87)? \nz.mem [1850] : 
                       (N89)? \nz.mem [1900] : 
                       (N91)? \nz.mem [1950] : 
                       (N93)? \nz.mem [2000] : 
                       (N95)? \nz.mem [2050] : 
                       (N97)? \nz.mem [2100] : 
                       (N99)? \nz.mem [2150] : 
                       (N101)? \nz.mem [2200] : 
                       (N103)? \nz.mem [2250] : 
                       (N105)? \nz.mem [2300] : 
                       (N107)? \nz.mem [2350] : 
                       (N109)? \nz.mem [2400] : 
                       (N111)? \nz.mem [2450] : 
                       (N113)? \nz.mem [2500] : 
                       (N115)? \nz.mem [2550] : 
                       (N117)? \nz.mem [2600] : 
                       (N119)? \nz.mem [2650] : 
                       (N121)? \nz.mem [2700] : 
                       (N123)? \nz.mem [2750] : 
                       (N125)? \nz.mem [2800] : 
                       (N127)? \nz.mem [2850] : 
                       (N129)? \nz.mem [2900] : 
                       (N131)? \nz.mem [2950] : 
                       (N133)? \nz.mem [3000] : 
                       (N135)? \nz.mem [3050] : 
                       (N137)? \nz.mem [3100] : 
                       (N139)? \nz.mem [3150] : 1'b0;
  assign N269 = ~w_addr_i[5];
  assign N270 = w_addr_i[3] & w_addr_i[4];
  assign N271 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N272 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N273 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N274 = w_addr_i[5] & N270;
  assign N275 = w_addr_i[5] & N271;
  assign N276 = w_addr_i[5] & N272;
  assign N277 = w_addr_i[5] & N273;
  assign N278 = N269 & N270;
  assign N279 = N269 & N271;
  assign N280 = N269 & N272;
  assign N281 = N269 & N273;
  assign N282 = ~w_addr_i[2];
  assign N283 = w_addr_i[0] & w_addr_i[1];
  assign N284 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N285 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N286 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N287 = w_addr_i[2] & N283;
  assign N288 = w_addr_i[2] & N284;
  assign N289 = w_addr_i[2] & N285;
  assign N290 = w_addr_i[2] & N286;
  assign N291 = N282 & N283;
  assign N292 = N282 & N284;
  assign N293 = N282 & N285;
  assign N294 = N282 & N286;
  assign N204 = N274 & N287;
  assign N203 = N274 & N288;
  assign N202 = N274 & N289;
  assign N201 = N274 & N290;
  assign N200 = N274 & N291;
  assign N199 = N274 & N292;
  assign N198 = N274 & N293;
  assign N197 = N274 & N294;
  assign N196 = N275 & N287;
  assign N195 = N275 & N288;
  assign N194 = N275 & N289;
  assign N193 = N275 & N290;
  assign N192 = N275 & N291;
  assign N191 = N275 & N292;
  assign N190 = N275 & N293;
  assign N189 = N275 & N294;
  assign N188 = N276 & N287;
  assign N187 = N276 & N288;
  assign N186 = N276 & N289;
  assign N185 = N276 & N290;
  assign N184 = N276 & N291;
  assign N183 = N276 & N292;
  assign N182 = N276 & N293;
  assign N181 = N276 & N294;
  assign N180 = N277 & N287;
  assign N179 = N277 & N288;
  assign N178 = N277 & N289;
  assign N177 = N277 & N290;
  assign N176 = N277 & N291;
  assign N175 = N277 & N292;
  assign N174 = N277 & N293;
  assign N173 = N277 & N294;
  assign N172 = N278 & N287;
  assign N171 = N278 & N288;
  assign N170 = N278 & N289;
  assign N169 = N278 & N290;
  assign N168 = N278 & N291;
  assign N167 = N278 & N292;
  assign N166 = N278 & N293;
  assign N165 = N278 & N294;
  assign N164 = N279 & N287;
  assign N163 = N279 & N288;
  assign N162 = N279 & N289;
  assign N161 = N279 & N290;
  assign N160 = N279 & N291;
  assign N159 = N279 & N292;
  assign N158 = N279 & N293;
  assign N157 = N279 & N294;
  assign N156 = N280 & N287;
  assign N155 = N280 & N288;
  assign N154 = N280 & N289;
  assign N153 = N280 & N290;
  assign N152 = N280 & N291;
  assign N151 = N280 & N292;
  assign N150 = N280 & N293;
  assign N149 = N280 & N294;
  assign N148 = N281 & N287;
  assign N147 = N281 & N288;
  assign N146 = N281 & N289;
  assign N145 = N281 & N290;
  assign N144 = N281 & N291;
  assign N143 = N281 & N292;
  assign N142 = N281 & N293;
  assign N141 = N281 & N294;
  assign { N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205 } = (N8)? { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~r_addr_i[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r_addr_i[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r_addr_i[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r_addr_i[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r_addr_i[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r_addr_i[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r_addr_i[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r_addr_i[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r_addr_i[3];
  assign N42 = ~r_addr_i[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r_addr_i[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r_addr_i[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r_addr_i[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r_addr_i[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r_addr_i[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r_addr_i[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r_addr_i[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r_addr_i[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r_addr_i[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r_addr_i[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r_addr_i[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r_addr_i[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r_addr_i[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r_addr_i[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r_addr_i[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r_addr_i[4];
  assign N75 = ~r_addr_i[5];
  assign N76 = N43 & N75;
  assign N77 = N43 & r_addr_i[5];
  assign N78 = N45 & N75;
  assign N79 = N45 & r_addr_i[5];
  assign N80 = N47 & N75;
  assign N81 = N47 & r_addr_i[5];
  assign N82 = N49 & N75;
  assign N83 = N49 & r_addr_i[5];
  assign N84 = N51 & N75;
  assign N85 = N51 & r_addr_i[5];
  assign N86 = N53 & N75;
  assign N87 = N53 & r_addr_i[5];
  assign N88 = N55 & N75;
  assign N89 = N55 & r_addr_i[5];
  assign N90 = N57 & N75;
  assign N91 = N57 & r_addr_i[5];
  assign N92 = N59 & N75;
  assign N93 = N59 & r_addr_i[5];
  assign N94 = N61 & N75;
  assign N95 = N61 & r_addr_i[5];
  assign N96 = N63 & N75;
  assign N97 = N63 & r_addr_i[5];
  assign N98 = N65 & N75;
  assign N99 = N65 & r_addr_i[5];
  assign N100 = N67 & N75;
  assign N101 = N67 & r_addr_i[5];
  assign N102 = N69 & N75;
  assign N103 = N69 & r_addr_i[5];
  assign N104 = N71 & N75;
  assign N105 = N71 & r_addr_i[5];
  assign N106 = N73 & N75;
  assign N107 = N73 & r_addr_i[5];
  assign N108 = N44 & N75;
  assign N109 = N44 & r_addr_i[5];
  assign N110 = N46 & N75;
  assign N111 = N46 & r_addr_i[5];
  assign N112 = N48 & N75;
  assign N113 = N48 & r_addr_i[5];
  assign N114 = N50 & N75;
  assign N115 = N50 & r_addr_i[5];
  assign N116 = N52 & N75;
  assign N117 = N52 & r_addr_i[5];
  assign N118 = N54 & N75;
  assign N119 = N54 & r_addr_i[5];
  assign N120 = N56 & N75;
  assign N121 = N56 & r_addr_i[5];
  assign N122 = N58 & N75;
  assign N123 = N58 & r_addr_i[5];
  assign N124 = N60 & N75;
  assign N125 = N60 & r_addr_i[5];
  assign N126 = N62 & N75;
  assign N127 = N62 & r_addr_i[5];
  assign N128 = N64 & N75;
  assign N129 = N64 & r_addr_i[5];
  assign N130 = N66 & N75;
  assign N131 = N66 & r_addr_i[5];
  assign N132 = N68 & N75;
  assign N133 = N68 & r_addr_i[5];
  assign N134 = N70 & N75;
  assign N135 = N70 & r_addr_i[5];
  assign N136 = N72 & N75;
  assign N137 = N72 & r_addr_i[5];
  assign N138 = N74 & N75;
  assign N139 = N74 & r_addr_i[5];
  assign N140 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N268) begin
      \nz.mem_3199_sv2v_reg  <= w_data_i[49];
      \nz.mem_3198_sv2v_reg  <= w_data_i[48];
      \nz.mem_3197_sv2v_reg  <= w_data_i[47];
      \nz.mem_3196_sv2v_reg  <= w_data_i[46];
      \nz.mem_3195_sv2v_reg  <= w_data_i[45];
      \nz.mem_3194_sv2v_reg  <= w_data_i[44];
      \nz.mem_3193_sv2v_reg  <= w_data_i[43];
      \nz.mem_3192_sv2v_reg  <= w_data_i[42];
      \nz.mem_3191_sv2v_reg  <= w_data_i[41];
      \nz.mem_3190_sv2v_reg  <= w_data_i[40];
      \nz.mem_3189_sv2v_reg  <= w_data_i[39];
      \nz.mem_3188_sv2v_reg  <= w_data_i[38];
      \nz.mem_3187_sv2v_reg  <= w_data_i[37];
      \nz.mem_3186_sv2v_reg  <= w_data_i[36];
      \nz.mem_3185_sv2v_reg  <= w_data_i[35];
      \nz.mem_3184_sv2v_reg  <= w_data_i[34];
      \nz.mem_3183_sv2v_reg  <= w_data_i[33];
      \nz.mem_3182_sv2v_reg  <= w_data_i[32];
      \nz.mem_3181_sv2v_reg  <= w_data_i[31];
      \nz.mem_3180_sv2v_reg  <= w_data_i[30];
      \nz.mem_3179_sv2v_reg  <= w_data_i[29];
      \nz.mem_3178_sv2v_reg  <= w_data_i[28];
      \nz.mem_3177_sv2v_reg  <= w_data_i[27];
      \nz.mem_3176_sv2v_reg  <= w_data_i[26];
      \nz.mem_3175_sv2v_reg  <= w_data_i[25];
      \nz.mem_3174_sv2v_reg  <= w_data_i[24];
      \nz.mem_3173_sv2v_reg  <= w_data_i[23];
      \nz.mem_3172_sv2v_reg  <= w_data_i[22];
      \nz.mem_3171_sv2v_reg  <= w_data_i[21];
      \nz.mem_3170_sv2v_reg  <= w_data_i[20];
      \nz.mem_3169_sv2v_reg  <= w_data_i[19];
      \nz.mem_3168_sv2v_reg  <= w_data_i[18];
      \nz.mem_3167_sv2v_reg  <= w_data_i[17];
      \nz.mem_3166_sv2v_reg  <= w_data_i[16];
      \nz.mem_3165_sv2v_reg  <= w_data_i[15];
      \nz.mem_3164_sv2v_reg  <= w_data_i[14];
      \nz.mem_3163_sv2v_reg  <= w_data_i[13];
      \nz.mem_3162_sv2v_reg  <= w_data_i[12];
      \nz.mem_3161_sv2v_reg  <= w_data_i[11];
      \nz.mem_3160_sv2v_reg  <= w_data_i[10];
      \nz.mem_3159_sv2v_reg  <= w_data_i[9];
      \nz.mem_3158_sv2v_reg  <= w_data_i[8];
      \nz.mem_3157_sv2v_reg  <= w_data_i[7];
      \nz.mem_3156_sv2v_reg  <= w_data_i[6];
      \nz.mem_3155_sv2v_reg  <= w_data_i[5];
      \nz.mem_3154_sv2v_reg  <= w_data_i[4];
      \nz.mem_3153_sv2v_reg  <= w_data_i[3];
      \nz.mem_3152_sv2v_reg  <= w_data_i[2];
      \nz.mem_3151_sv2v_reg  <= w_data_i[1];
      \nz.mem_3150_sv2v_reg  <= w_data_i[0];
    end 
    if(N267) begin
      \nz.mem_3149_sv2v_reg  <= w_data_i[49];
      \nz.mem_3148_sv2v_reg  <= w_data_i[48];
      \nz.mem_3147_sv2v_reg  <= w_data_i[47];
      \nz.mem_3146_sv2v_reg  <= w_data_i[46];
      \nz.mem_3145_sv2v_reg  <= w_data_i[45];
      \nz.mem_3144_sv2v_reg  <= w_data_i[44];
      \nz.mem_3143_sv2v_reg  <= w_data_i[43];
      \nz.mem_3142_sv2v_reg  <= w_data_i[42];
      \nz.mem_3141_sv2v_reg  <= w_data_i[41];
      \nz.mem_3140_sv2v_reg  <= w_data_i[40];
      \nz.mem_3139_sv2v_reg  <= w_data_i[39];
      \nz.mem_3138_sv2v_reg  <= w_data_i[38];
      \nz.mem_3137_sv2v_reg  <= w_data_i[37];
      \nz.mem_3136_sv2v_reg  <= w_data_i[36];
      \nz.mem_3135_sv2v_reg  <= w_data_i[35];
      \nz.mem_3134_sv2v_reg  <= w_data_i[34];
      \nz.mem_3133_sv2v_reg  <= w_data_i[33];
      \nz.mem_3132_sv2v_reg  <= w_data_i[32];
      \nz.mem_3131_sv2v_reg  <= w_data_i[31];
      \nz.mem_3130_sv2v_reg  <= w_data_i[30];
      \nz.mem_3129_sv2v_reg  <= w_data_i[29];
      \nz.mem_3128_sv2v_reg  <= w_data_i[28];
      \nz.mem_3127_sv2v_reg  <= w_data_i[27];
      \nz.mem_3126_sv2v_reg  <= w_data_i[26];
      \nz.mem_3125_sv2v_reg  <= w_data_i[25];
      \nz.mem_3124_sv2v_reg  <= w_data_i[24];
      \nz.mem_3123_sv2v_reg  <= w_data_i[23];
      \nz.mem_3122_sv2v_reg  <= w_data_i[22];
      \nz.mem_3121_sv2v_reg  <= w_data_i[21];
      \nz.mem_3120_sv2v_reg  <= w_data_i[20];
      \nz.mem_3119_sv2v_reg  <= w_data_i[19];
      \nz.mem_3118_sv2v_reg  <= w_data_i[18];
      \nz.mem_3117_sv2v_reg  <= w_data_i[17];
      \nz.mem_3116_sv2v_reg  <= w_data_i[16];
      \nz.mem_3115_sv2v_reg  <= w_data_i[15];
      \nz.mem_3114_sv2v_reg  <= w_data_i[14];
      \nz.mem_3113_sv2v_reg  <= w_data_i[13];
      \nz.mem_3112_sv2v_reg  <= w_data_i[12];
      \nz.mem_3111_sv2v_reg  <= w_data_i[11];
      \nz.mem_3110_sv2v_reg  <= w_data_i[10];
      \nz.mem_3109_sv2v_reg  <= w_data_i[9];
      \nz.mem_3108_sv2v_reg  <= w_data_i[8];
      \nz.mem_3107_sv2v_reg  <= w_data_i[7];
      \nz.mem_3106_sv2v_reg  <= w_data_i[6];
      \nz.mem_3105_sv2v_reg  <= w_data_i[5];
      \nz.mem_3104_sv2v_reg  <= w_data_i[4];
      \nz.mem_3103_sv2v_reg  <= w_data_i[3];
      \nz.mem_3102_sv2v_reg  <= w_data_i[2];
      \nz.mem_3101_sv2v_reg  <= w_data_i[1];
      \nz.mem_3100_sv2v_reg  <= w_data_i[0];
    end 
    if(N266) begin
      \nz.mem_3099_sv2v_reg  <= w_data_i[49];
      \nz.mem_3098_sv2v_reg  <= w_data_i[48];
      \nz.mem_3097_sv2v_reg  <= w_data_i[47];
      \nz.mem_3096_sv2v_reg  <= w_data_i[46];
      \nz.mem_3095_sv2v_reg  <= w_data_i[45];
      \nz.mem_3094_sv2v_reg  <= w_data_i[44];
      \nz.mem_3093_sv2v_reg  <= w_data_i[43];
      \nz.mem_3092_sv2v_reg  <= w_data_i[42];
      \nz.mem_3091_sv2v_reg  <= w_data_i[41];
      \nz.mem_3090_sv2v_reg  <= w_data_i[40];
      \nz.mem_3089_sv2v_reg  <= w_data_i[39];
      \nz.mem_3088_sv2v_reg  <= w_data_i[38];
      \nz.mem_3087_sv2v_reg  <= w_data_i[37];
      \nz.mem_3086_sv2v_reg  <= w_data_i[36];
      \nz.mem_3085_sv2v_reg  <= w_data_i[35];
      \nz.mem_3084_sv2v_reg  <= w_data_i[34];
      \nz.mem_3083_sv2v_reg  <= w_data_i[33];
      \nz.mem_3082_sv2v_reg  <= w_data_i[32];
      \nz.mem_3081_sv2v_reg  <= w_data_i[31];
      \nz.mem_3080_sv2v_reg  <= w_data_i[30];
      \nz.mem_3079_sv2v_reg  <= w_data_i[29];
      \nz.mem_3078_sv2v_reg  <= w_data_i[28];
      \nz.mem_3077_sv2v_reg  <= w_data_i[27];
      \nz.mem_3076_sv2v_reg  <= w_data_i[26];
      \nz.mem_3075_sv2v_reg  <= w_data_i[25];
      \nz.mem_3074_sv2v_reg  <= w_data_i[24];
      \nz.mem_3073_sv2v_reg  <= w_data_i[23];
      \nz.mem_3072_sv2v_reg  <= w_data_i[22];
      \nz.mem_3071_sv2v_reg  <= w_data_i[21];
      \nz.mem_3070_sv2v_reg  <= w_data_i[20];
      \nz.mem_3069_sv2v_reg  <= w_data_i[19];
      \nz.mem_3068_sv2v_reg  <= w_data_i[18];
      \nz.mem_3067_sv2v_reg  <= w_data_i[17];
      \nz.mem_3066_sv2v_reg  <= w_data_i[16];
      \nz.mem_3065_sv2v_reg  <= w_data_i[15];
      \nz.mem_3064_sv2v_reg  <= w_data_i[14];
      \nz.mem_3063_sv2v_reg  <= w_data_i[13];
      \nz.mem_3062_sv2v_reg  <= w_data_i[12];
      \nz.mem_3061_sv2v_reg  <= w_data_i[11];
      \nz.mem_3060_sv2v_reg  <= w_data_i[10];
      \nz.mem_3059_sv2v_reg  <= w_data_i[9];
      \nz.mem_3058_sv2v_reg  <= w_data_i[8];
      \nz.mem_3057_sv2v_reg  <= w_data_i[7];
      \nz.mem_3056_sv2v_reg  <= w_data_i[6];
      \nz.mem_3055_sv2v_reg  <= w_data_i[5];
      \nz.mem_3054_sv2v_reg  <= w_data_i[4];
      \nz.mem_3053_sv2v_reg  <= w_data_i[3];
      \nz.mem_3052_sv2v_reg  <= w_data_i[2];
      \nz.mem_3051_sv2v_reg  <= w_data_i[1];
      \nz.mem_3050_sv2v_reg  <= w_data_i[0];
    end 
    if(N265) begin
      \nz.mem_3049_sv2v_reg  <= w_data_i[49];
      \nz.mem_3048_sv2v_reg  <= w_data_i[48];
      \nz.mem_3047_sv2v_reg  <= w_data_i[47];
      \nz.mem_3046_sv2v_reg  <= w_data_i[46];
      \nz.mem_3045_sv2v_reg  <= w_data_i[45];
      \nz.mem_3044_sv2v_reg  <= w_data_i[44];
      \nz.mem_3043_sv2v_reg  <= w_data_i[43];
      \nz.mem_3042_sv2v_reg  <= w_data_i[42];
      \nz.mem_3041_sv2v_reg  <= w_data_i[41];
      \nz.mem_3040_sv2v_reg  <= w_data_i[40];
      \nz.mem_3039_sv2v_reg  <= w_data_i[39];
      \nz.mem_3038_sv2v_reg  <= w_data_i[38];
      \nz.mem_3037_sv2v_reg  <= w_data_i[37];
      \nz.mem_3036_sv2v_reg  <= w_data_i[36];
      \nz.mem_3035_sv2v_reg  <= w_data_i[35];
      \nz.mem_3034_sv2v_reg  <= w_data_i[34];
      \nz.mem_3033_sv2v_reg  <= w_data_i[33];
      \nz.mem_3032_sv2v_reg  <= w_data_i[32];
      \nz.mem_3031_sv2v_reg  <= w_data_i[31];
      \nz.mem_3030_sv2v_reg  <= w_data_i[30];
      \nz.mem_3029_sv2v_reg  <= w_data_i[29];
      \nz.mem_3028_sv2v_reg  <= w_data_i[28];
      \nz.mem_3027_sv2v_reg  <= w_data_i[27];
      \nz.mem_3026_sv2v_reg  <= w_data_i[26];
      \nz.mem_3025_sv2v_reg  <= w_data_i[25];
      \nz.mem_3024_sv2v_reg  <= w_data_i[24];
      \nz.mem_3023_sv2v_reg  <= w_data_i[23];
      \nz.mem_3022_sv2v_reg  <= w_data_i[22];
      \nz.mem_3021_sv2v_reg  <= w_data_i[21];
      \nz.mem_3020_sv2v_reg  <= w_data_i[20];
      \nz.mem_3019_sv2v_reg  <= w_data_i[19];
      \nz.mem_3018_sv2v_reg  <= w_data_i[18];
      \nz.mem_3017_sv2v_reg  <= w_data_i[17];
      \nz.mem_3016_sv2v_reg  <= w_data_i[16];
      \nz.mem_3015_sv2v_reg  <= w_data_i[15];
      \nz.mem_3014_sv2v_reg  <= w_data_i[14];
      \nz.mem_3013_sv2v_reg  <= w_data_i[13];
      \nz.mem_3012_sv2v_reg  <= w_data_i[12];
      \nz.mem_3011_sv2v_reg  <= w_data_i[11];
      \nz.mem_3010_sv2v_reg  <= w_data_i[10];
      \nz.mem_3009_sv2v_reg  <= w_data_i[9];
      \nz.mem_3008_sv2v_reg  <= w_data_i[8];
      \nz.mem_3007_sv2v_reg  <= w_data_i[7];
      \nz.mem_3006_sv2v_reg  <= w_data_i[6];
      \nz.mem_3005_sv2v_reg  <= w_data_i[5];
      \nz.mem_3004_sv2v_reg  <= w_data_i[4];
      \nz.mem_3003_sv2v_reg  <= w_data_i[3];
      \nz.mem_3002_sv2v_reg  <= w_data_i[2];
      \nz.mem_3001_sv2v_reg  <= w_data_i[1];
      \nz.mem_3000_sv2v_reg  <= w_data_i[0];
    end 
    if(N264) begin
      \nz.mem_2999_sv2v_reg  <= w_data_i[49];
      \nz.mem_2998_sv2v_reg  <= w_data_i[48];
      \nz.mem_2997_sv2v_reg  <= w_data_i[47];
      \nz.mem_2996_sv2v_reg  <= w_data_i[46];
      \nz.mem_2995_sv2v_reg  <= w_data_i[45];
      \nz.mem_2994_sv2v_reg  <= w_data_i[44];
      \nz.mem_2993_sv2v_reg  <= w_data_i[43];
      \nz.mem_2992_sv2v_reg  <= w_data_i[42];
      \nz.mem_2991_sv2v_reg  <= w_data_i[41];
      \nz.mem_2990_sv2v_reg  <= w_data_i[40];
      \nz.mem_2989_sv2v_reg  <= w_data_i[39];
      \nz.mem_2988_sv2v_reg  <= w_data_i[38];
      \nz.mem_2987_sv2v_reg  <= w_data_i[37];
      \nz.mem_2986_sv2v_reg  <= w_data_i[36];
      \nz.mem_2985_sv2v_reg  <= w_data_i[35];
      \nz.mem_2984_sv2v_reg  <= w_data_i[34];
      \nz.mem_2983_sv2v_reg  <= w_data_i[33];
      \nz.mem_2982_sv2v_reg  <= w_data_i[32];
      \nz.mem_2981_sv2v_reg  <= w_data_i[31];
      \nz.mem_2980_sv2v_reg  <= w_data_i[30];
      \nz.mem_2979_sv2v_reg  <= w_data_i[29];
      \nz.mem_2978_sv2v_reg  <= w_data_i[28];
      \nz.mem_2977_sv2v_reg  <= w_data_i[27];
      \nz.mem_2976_sv2v_reg  <= w_data_i[26];
      \nz.mem_2975_sv2v_reg  <= w_data_i[25];
      \nz.mem_2974_sv2v_reg  <= w_data_i[24];
      \nz.mem_2973_sv2v_reg  <= w_data_i[23];
      \nz.mem_2972_sv2v_reg  <= w_data_i[22];
      \nz.mem_2971_sv2v_reg  <= w_data_i[21];
      \nz.mem_2970_sv2v_reg  <= w_data_i[20];
      \nz.mem_2969_sv2v_reg  <= w_data_i[19];
      \nz.mem_2968_sv2v_reg  <= w_data_i[18];
      \nz.mem_2967_sv2v_reg  <= w_data_i[17];
      \nz.mem_2966_sv2v_reg  <= w_data_i[16];
      \nz.mem_2965_sv2v_reg  <= w_data_i[15];
      \nz.mem_2964_sv2v_reg  <= w_data_i[14];
      \nz.mem_2963_sv2v_reg  <= w_data_i[13];
      \nz.mem_2962_sv2v_reg  <= w_data_i[12];
      \nz.mem_2961_sv2v_reg  <= w_data_i[11];
      \nz.mem_2960_sv2v_reg  <= w_data_i[10];
      \nz.mem_2959_sv2v_reg  <= w_data_i[9];
      \nz.mem_2958_sv2v_reg  <= w_data_i[8];
      \nz.mem_2957_sv2v_reg  <= w_data_i[7];
      \nz.mem_2956_sv2v_reg  <= w_data_i[6];
      \nz.mem_2955_sv2v_reg  <= w_data_i[5];
      \nz.mem_2954_sv2v_reg  <= w_data_i[4];
      \nz.mem_2953_sv2v_reg  <= w_data_i[3];
      \nz.mem_2952_sv2v_reg  <= w_data_i[2];
      \nz.mem_2951_sv2v_reg  <= w_data_i[1];
      \nz.mem_2950_sv2v_reg  <= w_data_i[0];
    end 
    if(N263) begin
      \nz.mem_2949_sv2v_reg  <= w_data_i[49];
      \nz.mem_2948_sv2v_reg  <= w_data_i[48];
      \nz.mem_2947_sv2v_reg  <= w_data_i[47];
      \nz.mem_2946_sv2v_reg  <= w_data_i[46];
      \nz.mem_2945_sv2v_reg  <= w_data_i[45];
      \nz.mem_2944_sv2v_reg  <= w_data_i[44];
      \nz.mem_2943_sv2v_reg  <= w_data_i[43];
      \nz.mem_2942_sv2v_reg  <= w_data_i[42];
      \nz.mem_2941_sv2v_reg  <= w_data_i[41];
      \nz.mem_2940_sv2v_reg  <= w_data_i[40];
      \nz.mem_2939_sv2v_reg  <= w_data_i[39];
      \nz.mem_2938_sv2v_reg  <= w_data_i[38];
      \nz.mem_2937_sv2v_reg  <= w_data_i[37];
      \nz.mem_2936_sv2v_reg  <= w_data_i[36];
      \nz.mem_2935_sv2v_reg  <= w_data_i[35];
      \nz.mem_2934_sv2v_reg  <= w_data_i[34];
      \nz.mem_2933_sv2v_reg  <= w_data_i[33];
      \nz.mem_2932_sv2v_reg  <= w_data_i[32];
      \nz.mem_2931_sv2v_reg  <= w_data_i[31];
      \nz.mem_2930_sv2v_reg  <= w_data_i[30];
      \nz.mem_2929_sv2v_reg  <= w_data_i[29];
      \nz.mem_2928_sv2v_reg  <= w_data_i[28];
      \nz.mem_2927_sv2v_reg  <= w_data_i[27];
      \nz.mem_2926_sv2v_reg  <= w_data_i[26];
      \nz.mem_2925_sv2v_reg  <= w_data_i[25];
      \nz.mem_2924_sv2v_reg  <= w_data_i[24];
      \nz.mem_2923_sv2v_reg  <= w_data_i[23];
      \nz.mem_2922_sv2v_reg  <= w_data_i[22];
      \nz.mem_2921_sv2v_reg  <= w_data_i[21];
      \nz.mem_2920_sv2v_reg  <= w_data_i[20];
      \nz.mem_2919_sv2v_reg  <= w_data_i[19];
      \nz.mem_2918_sv2v_reg  <= w_data_i[18];
      \nz.mem_2917_sv2v_reg  <= w_data_i[17];
      \nz.mem_2916_sv2v_reg  <= w_data_i[16];
      \nz.mem_2915_sv2v_reg  <= w_data_i[15];
      \nz.mem_2914_sv2v_reg  <= w_data_i[14];
      \nz.mem_2913_sv2v_reg  <= w_data_i[13];
      \nz.mem_2912_sv2v_reg  <= w_data_i[12];
      \nz.mem_2911_sv2v_reg  <= w_data_i[11];
      \nz.mem_2910_sv2v_reg  <= w_data_i[10];
      \nz.mem_2909_sv2v_reg  <= w_data_i[9];
      \nz.mem_2908_sv2v_reg  <= w_data_i[8];
      \nz.mem_2907_sv2v_reg  <= w_data_i[7];
      \nz.mem_2906_sv2v_reg  <= w_data_i[6];
      \nz.mem_2905_sv2v_reg  <= w_data_i[5];
      \nz.mem_2904_sv2v_reg  <= w_data_i[4];
      \nz.mem_2903_sv2v_reg  <= w_data_i[3];
      \nz.mem_2902_sv2v_reg  <= w_data_i[2];
      \nz.mem_2901_sv2v_reg  <= w_data_i[1];
      \nz.mem_2900_sv2v_reg  <= w_data_i[0];
    end 
    if(N262) begin
      \nz.mem_2899_sv2v_reg  <= w_data_i[49];
      \nz.mem_2898_sv2v_reg  <= w_data_i[48];
      \nz.mem_2897_sv2v_reg  <= w_data_i[47];
      \nz.mem_2896_sv2v_reg  <= w_data_i[46];
      \nz.mem_2895_sv2v_reg  <= w_data_i[45];
      \nz.mem_2894_sv2v_reg  <= w_data_i[44];
      \nz.mem_2893_sv2v_reg  <= w_data_i[43];
      \nz.mem_2892_sv2v_reg  <= w_data_i[42];
      \nz.mem_2891_sv2v_reg  <= w_data_i[41];
      \nz.mem_2890_sv2v_reg  <= w_data_i[40];
      \nz.mem_2889_sv2v_reg  <= w_data_i[39];
      \nz.mem_2888_sv2v_reg  <= w_data_i[38];
      \nz.mem_2887_sv2v_reg  <= w_data_i[37];
      \nz.mem_2886_sv2v_reg  <= w_data_i[36];
      \nz.mem_2885_sv2v_reg  <= w_data_i[35];
      \nz.mem_2884_sv2v_reg  <= w_data_i[34];
      \nz.mem_2883_sv2v_reg  <= w_data_i[33];
      \nz.mem_2882_sv2v_reg  <= w_data_i[32];
      \nz.mem_2881_sv2v_reg  <= w_data_i[31];
      \nz.mem_2880_sv2v_reg  <= w_data_i[30];
      \nz.mem_2879_sv2v_reg  <= w_data_i[29];
      \nz.mem_2878_sv2v_reg  <= w_data_i[28];
      \nz.mem_2877_sv2v_reg  <= w_data_i[27];
      \nz.mem_2876_sv2v_reg  <= w_data_i[26];
      \nz.mem_2875_sv2v_reg  <= w_data_i[25];
      \nz.mem_2874_sv2v_reg  <= w_data_i[24];
      \nz.mem_2873_sv2v_reg  <= w_data_i[23];
      \nz.mem_2872_sv2v_reg  <= w_data_i[22];
      \nz.mem_2871_sv2v_reg  <= w_data_i[21];
      \nz.mem_2870_sv2v_reg  <= w_data_i[20];
      \nz.mem_2869_sv2v_reg  <= w_data_i[19];
      \nz.mem_2868_sv2v_reg  <= w_data_i[18];
      \nz.mem_2867_sv2v_reg  <= w_data_i[17];
      \nz.mem_2866_sv2v_reg  <= w_data_i[16];
      \nz.mem_2865_sv2v_reg  <= w_data_i[15];
      \nz.mem_2864_sv2v_reg  <= w_data_i[14];
      \nz.mem_2863_sv2v_reg  <= w_data_i[13];
      \nz.mem_2862_sv2v_reg  <= w_data_i[12];
      \nz.mem_2861_sv2v_reg  <= w_data_i[11];
      \nz.mem_2860_sv2v_reg  <= w_data_i[10];
      \nz.mem_2859_sv2v_reg  <= w_data_i[9];
      \nz.mem_2858_sv2v_reg  <= w_data_i[8];
      \nz.mem_2857_sv2v_reg  <= w_data_i[7];
      \nz.mem_2856_sv2v_reg  <= w_data_i[6];
      \nz.mem_2855_sv2v_reg  <= w_data_i[5];
      \nz.mem_2854_sv2v_reg  <= w_data_i[4];
      \nz.mem_2853_sv2v_reg  <= w_data_i[3];
      \nz.mem_2852_sv2v_reg  <= w_data_i[2];
      \nz.mem_2851_sv2v_reg  <= w_data_i[1];
      \nz.mem_2850_sv2v_reg  <= w_data_i[0];
    end 
    if(N261) begin
      \nz.mem_2849_sv2v_reg  <= w_data_i[49];
      \nz.mem_2848_sv2v_reg  <= w_data_i[48];
      \nz.mem_2847_sv2v_reg  <= w_data_i[47];
      \nz.mem_2846_sv2v_reg  <= w_data_i[46];
      \nz.mem_2845_sv2v_reg  <= w_data_i[45];
      \nz.mem_2844_sv2v_reg  <= w_data_i[44];
      \nz.mem_2843_sv2v_reg  <= w_data_i[43];
      \nz.mem_2842_sv2v_reg  <= w_data_i[42];
      \nz.mem_2841_sv2v_reg  <= w_data_i[41];
      \nz.mem_2840_sv2v_reg  <= w_data_i[40];
      \nz.mem_2839_sv2v_reg  <= w_data_i[39];
      \nz.mem_2838_sv2v_reg  <= w_data_i[38];
      \nz.mem_2837_sv2v_reg  <= w_data_i[37];
      \nz.mem_2836_sv2v_reg  <= w_data_i[36];
      \nz.mem_2835_sv2v_reg  <= w_data_i[35];
      \nz.mem_2834_sv2v_reg  <= w_data_i[34];
      \nz.mem_2833_sv2v_reg  <= w_data_i[33];
      \nz.mem_2832_sv2v_reg  <= w_data_i[32];
      \nz.mem_2831_sv2v_reg  <= w_data_i[31];
      \nz.mem_2830_sv2v_reg  <= w_data_i[30];
      \nz.mem_2829_sv2v_reg  <= w_data_i[29];
      \nz.mem_2828_sv2v_reg  <= w_data_i[28];
      \nz.mem_2827_sv2v_reg  <= w_data_i[27];
      \nz.mem_2826_sv2v_reg  <= w_data_i[26];
      \nz.mem_2825_sv2v_reg  <= w_data_i[25];
      \nz.mem_2824_sv2v_reg  <= w_data_i[24];
      \nz.mem_2823_sv2v_reg  <= w_data_i[23];
      \nz.mem_2822_sv2v_reg  <= w_data_i[22];
      \nz.mem_2821_sv2v_reg  <= w_data_i[21];
      \nz.mem_2820_sv2v_reg  <= w_data_i[20];
      \nz.mem_2819_sv2v_reg  <= w_data_i[19];
      \nz.mem_2818_sv2v_reg  <= w_data_i[18];
      \nz.mem_2817_sv2v_reg  <= w_data_i[17];
      \nz.mem_2816_sv2v_reg  <= w_data_i[16];
      \nz.mem_2815_sv2v_reg  <= w_data_i[15];
      \nz.mem_2814_sv2v_reg  <= w_data_i[14];
      \nz.mem_2813_sv2v_reg  <= w_data_i[13];
      \nz.mem_2812_sv2v_reg  <= w_data_i[12];
      \nz.mem_2811_sv2v_reg  <= w_data_i[11];
      \nz.mem_2810_sv2v_reg  <= w_data_i[10];
      \nz.mem_2809_sv2v_reg  <= w_data_i[9];
      \nz.mem_2808_sv2v_reg  <= w_data_i[8];
      \nz.mem_2807_sv2v_reg  <= w_data_i[7];
      \nz.mem_2806_sv2v_reg  <= w_data_i[6];
      \nz.mem_2805_sv2v_reg  <= w_data_i[5];
      \nz.mem_2804_sv2v_reg  <= w_data_i[4];
      \nz.mem_2803_sv2v_reg  <= w_data_i[3];
      \nz.mem_2802_sv2v_reg  <= w_data_i[2];
      \nz.mem_2801_sv2v_reg  <= w_data_i[1];
      \nz.mem_2800_sv2v_reg  <= w_data_i[0];
    end 
    if(N260) begin
      \nz.mem_2799_sv2v_reg  <= w_data_i[49];
      \nz.mem_2798_sv2v_reg  <= w_data_i[48];
      \nz.mem_2797_sv2v_reg  <= w_data_i[47];
      \nz.mem_2796_sv2v_reg  <= w_data_i[46];
      \nz.mem_2795_sv2v_reg  <= w_data_i[45];
      \nz.mem_2794_sv2v_reg  <= w_data_i[44];
      \nz.mem_2793_sv2v_reg  <= w_data_i[43];
      \nz.mem_2792_sv2v_reg  <= w_data_i[42];
      \nz.mem_2791_sv2v_reg  <= w_data_i[41];
      \nz.mem_2790_sv2v_reg  <= w_data_i[40];
      \nz.mem_2789_sv2v_reg  <= w_data_i[39];
      \nz.mem_2788_sv2v_reg  <= w_data_i[38];
      \nz.mem_2787_sv2v_reg  <= w_data_i[37];
      \nz.mem_2786_sv2v_reg  <= w_data_i[36];
      \nz.mem_2785_sv2v_reg  <= w_data_i[35];
      \nz.mem_2784_sv2v_reg  <= w_data_i[34];
      \nz.mem_2783_sv2v_reg  <= w_data_i[33];
      \nz.mem_2782_sv2v_reg  <= w_data_i[32];
      \nz.mem_2781_sv2v_reg  <= w_data_i[31];
      \nz.mem_2780_sv2v_reg  <= w_data_i[30];
      \nz.mem_2779_sv2v_reg  <= w_data_i[29];
      \nz.mem_2778_sv2v_reg  <= w_data_i[28];
      \nz.mem_2777_sv2v_reg  <= w_data_i[27];
      \nz.mem_2776_sv2v_reg  <= w_data_i[26];
      \nz.mem_2775_sv2v_reg  <= w_data_i[25];
      \nz.mem_2774_sv2v_reg  <= w_data_i[24];
      \nz.mem_2773_sv2v_reg  <= w_data_i[23];
      \nz.mem_2772_sv2v_reg  <= w_data_i[22];
      \nz.mem_2771_sv2v_reg  <= w_data_i[21];
      \nz.mem_2770_sv2v_reg  <= w_data_i[20];
      \nz.mem_2769_sv2v_reg  <= w_data_i[19];
      \nz.mem_2768_sv2v_reg  <= w_data_i[18];
      \nz.mem_2767_sv2v_reg  <= w_data_i[17];
      \nz.mem_2766_sv2v_reg  <= w_data_i[16];
      \nz.mem_2765_sv2v_reg  <= w_data_i[15];
      \nz.mem_2764_sv2v_reg  <= w_data_i[14];
      \nz.mem_2763_sv2v_reg  <= w_data_i[13];
      \nz.mem_2762_sv2v_reg  <= w_data_i[12];
      \nz.mem_2761_sv2v_reg  <= w_data_i[11];
      \nz.mem_2760_sv2v_reg  <= w_data_i[10];
      \nz.mem_2759_sv2v_reg  <= w_data_i[9];
      \nz.mem_2758_sv2v_reg  <= w_data_i[8];
      \nz.mem_2757_sv2v_reg  <= w_data_i[7];
      \nz.mem_2756_sv2v_reg  <= w_data_i[6];
      \nz.mem_2755_sv2v_reg  <= w_data_i[5];
      \nz.mem_2754_sv2v_reg  <= w_data_i[4];
      \nz.mem_2753_sv2v_reg  <= w_data_i[3];
      \nz.mem_2752_sv2v_reg  <= w_data_i[2];
      \nz.mem_2751_sv2v_reg  <= w_data_i[1];
      \nz.mem_2750_sv2v_reg  <= w_data_i[0];
    end 
    if(N259) begin
      \nz.mem_2749_sv2v_reg  <= w_data_i[49];
      \nz.mem_2748_sv2v_reg  <= w_data_i[48];
      \nz.mem_2747_sv2v_reg  <= w_data_i[47];
      \nz.mem_2746_sv2v_reg  <= w_data_i[46];
      \nz.mem_2745_sv2v_reg  <= w_data_i[45];
      \nz.mem_2744_sv2v_reg  <= w_data_i[44];
      \nz.mem_2743_sv2v_reg  <= w_data_i[43];
      \nz.mem_2742_sv2v_reg  <= w_data_i[42];
      \nz.mem_2741_sv2v_reg  <= w_data_i[41];
      \nz.mem_2740_sv2v_reg  <= w_data_i[40];
      \nz.mem_2739_sv2v_reg  <= w_data_i[39];
      \nz.mem_2738_sv2v_reg  <= w_data_i[38];
      \nz.mem_2737_sv2v_reg  <= w_data_i[37];
      \nz.mem_2736_sv2v_reg  <= w_data_i[36];
      \nz.mem_2735_sv2v_reg  <= w_data_i[35];
      \nz.mem_2734_sv2v_reg  <= w_data_i[34];
      \nz.mem_2733_sv2v_reg  <= w_data_i[33];
      \nz.mem_2732_sv2v_reg  <= w_data_i[32];
      \nz.mem_2731_sv2v_reg  <= w_data_i[31];
      \nz.mem_2730_sv2v_reg  <= w_data_i[30];
      \nz.mem_2729_sv2v_reg  <= w_data_i[29];
      \nz.mem_2728_sv2v_reg  <= w_data_i[28];
      \nz.mem_2727_sv2v_reg  <= w_data_i[27];
      \nz.mem_2726_sv2v_reg  <= w_data_i[26];
      \nz.mem_2725_sv2v_reg  <= w_data_i[25];
      \nz.mem_2724_sv2v_reg  <= w_data_i[24];
      \nz.mem_2723_sv2v_reg  <= w_data_i[23];
      \nz.mem_2722_sv2v_reg  <= w_data_i[22];
      \nz.mem_2721_sv2v_reg  <= w_data_i[21];
      \nz.mem_2720_sv2v_reg  <= w_data_i[20];
      \nz.mem_2719_sv2v_reg  <= w_data_i[19];
      \nz.mem_2718_sv2v_reg  <= w_data_i[18];
      \nz.mem_2717_sv2v_reg  <= w_data_i[17];
      \nz.mem_2716_sv2v_reg  <= w_data_i[16];
      \nz.mem_2715_sv2v_reg  <= w_data_i[15];
      \nz.mem_2714_sv2v_reg  <= w_data_i[14];
      \nz.mem_2713_sv2v_reg  <= w_data_i[13];
      \nz.mem_2712_sv2v_reg  <= w_data_i[12];
      \nz.mem_2711_sv2v_reg  <= w_data_i[11];
      \nz.mem_2710_sv2v_reg  <= w_data_i[10];
      \nz.mem_2709_sv2v_reg  <= w_data_i[9];
      \nz.mem_2708_sv2v_reg  <= w_data_i[8];
      \nz.mem_2707_sv2v_reg  <= w_data_i[7];
      \nz.mem_2706_sv2v_reg  <= w_data_i[6];
      \nz.mem_2705_sv2v_reg  <= w_data_i[5];
      \nz.mem_2704_sv2v_reg  <= w_data_i[4];
      \nz.mem_2703_sv2v_reg  <= w_data_i[3];
      \nz.mem_2702_sv2v_reg  <= w_data_i[2];
      \nz.mem_2701_sv2v_reg  <= w_data_i[1];
      \nz.mem_2700_sv2v_reg  <= w_data_i[0];
    end 
    if(N258) begin
      \nz.mem_2699_sv2v_reg  <= w_data_i[49];
      \nz.mem_2698_sv2v_reg  <= w_data_i[48];
      \nz.mem_2697_sv2v_reg  <= w_data_i[47];
      \nz.mem_2696_sv2v_reg  <= w_data_i[46];
      \nz.mem_2695_sv2v_reg  <= w_data_i[45];
      \nz.mem_2694_sv2v_reg  <= w_data_i[44];
      \nz.mem_2693_sv2v_reg  <= w_data_i[43];
      \nz.mem_2692_sv2v_reg  <= w_data_i[42];
      \nz.mem_2691_sv2v_reg  <= w_data_i[41];
      \nz.mem_2690_sv2v_reg  <= w_data_i[40];
      \nz.mem_2689_sv2v_reg  <= w_data_i[39];
      \nz.mem_2688_sv2v_reg  <= w_data_i[38];
      \nz.mem_2687_sv2v_reg  <= w_data_i[37];
      \nz.mem_2686_sv2v_reg  <= w_data_i[36];
      \nz.mem_2685_sv2v_reg  <= w_data_i[35];
      \nz.mem_2684_sv2v_reg  <= w_data_i[34];
      \nz.mem_2683_sv2v_reg  <= w_data_i[33];
      \nz.mem_2682_sv2v_reg  <= w_data_i[32];
      \nz.mem_2681_sv2v_reg  <= w_data_i[31];
      \nz.mem_2680_sv2v_reg  <= w_data_i[30];
      \nz.mem_2679_sv2v_reg  <= w_data_i[29];
      \nz.mem_2678_sv2v_reg  <= w_data_i[28];
      \nz.mem_2677_sv2v_reg  <= w_data_i[27];
      \nz.mem_2676_sv2v_reg  <= w_data_i[26];
      \nz.mem_2675_sv2v_reg  <= w_data_i[25];
      \nz.mem_2674_sv2v_reg  <= w_data_i[24];
      \nz.mem_2673_sv2v_reg  <= w_data_i[23];
      \nz.mem_2672_sv2v_reg  <= w_data_i[22];
      \nz.mem_2671_sv2v_reg  <= w_data_i[21];
      \nz.mem_2670_sv2v_reg  <= w_data_i[20];
      \nz.mem_2669_sv2v_reg  <= w_data_i[19];
      \nz.mem_2668_sv2v_reg  <= w_data_i[18];
      \nz.mem_2667_sv2v_reg  <= w_data_i[17];
      \nz.mem_2666_sv2v_reg  <= w_data_i[16];
      \nz.mem_2665_sv2v_reg  <= w_data_i[15];
      \nz.mem_2664_sv2v_reg  <= w_data_i[14];
      \nz.mem_2663_sv2v_reg  <= w_data_i[13];
      \nz.mem_2662_sv2v_reg  <= w_data_i[12];
      \nz.mem_2661_sv2v_reg  <= w_data_i[11];
      \nz.mem_2660_sv2v_reg  <= w_data_i[10];
      \nz.mem_2659_sv2v_reg  <= w_data_i[9];
      \nz.mem_2658_sv2v_reg  <= w_data_i[8];
      \nz.mem_2657_sv2v_reg  <= w_data_i[7];
      \nz.mem_2656_sv2v_reg  <= w_data_i[6];
      \nz.mem_2655_sv2v_reg  <= w_data_i[5];
      \nz.mem_2654_sv2v_reg  <= w_data_i[4];
      \nz.mem_2653_sv2v_reg  <= w_data_i[3];
      \nz.mem_2652_sv2v_reg  <= w_data_i[2];
      \nz.mem_2651_sv2v_reg  <= w_data_i[1];
      \nz.mem_2650_sv2v_reg  <= w_data_i[0];
    end 
    if(N257) begin
      \nz.mem_2649_sv2v_reg  <= w_data_i[49];
      \nz.mem_2648_sv2v_reg  <= w_data_i[48];
      \nz.mem_2647_sv2v_reg  <= w_data_i[47];
      \nz.mem_2646_sv2v_reg  <= w_data_i[46];
      \nz.mem_2645_sv2v_reg  <= w_data_i[45];
      \nz.mem_2644_sv2v_reg  <= w_data_i[44];
      \nz.mem_2643_sv2v_reg  <= w_data_i[43];
      \nz.mem_2642_sv2v_reg  <= w_data_i[42];
      \nz.mem_2641_sv2v_reg  <= w_data_i[41];
      \nz.mem_2640_sv2v_reg  <= w_data_i[40];
      \nz.mem_2639_sv2v_reg  <= w_data_i[39];
      \nz.mem_2638_sv2v_reg  <= w_data_i[38];
      \nz.mem_2637_sv2v_reg  <= w_data_i[37];
      \nz.mem_2636_sv2v_reg  <= w_data_i[36];
      \nz.mem_2635_sv2v_reg  <= w_data_i[35];
      \nz.mem_2634_sv2v_reg  <= w_data_i[34];
      \nz.mem_2633_sv2v_reg  <= w_data_i[33];
      \nz.mem_2632_sv2v_reg  <= w_data_i[32];
      \nz.mem_2631_sv2v_reg  <= w_data_i[31];
      \nz.mem_2630_sv2v_reg  <= w_data_i[30];
      \nz.mem_2629_sv2v_reg  <= w_data_i[29];
      \nz.mem_2628_sv2v_reg  <= w_data_i[28];
      \nz.mem_2627_sv2v_reg  <= w_data_i[27];
      \nz.mem_2626_sv2v_reg  <= w_data_i[26];
      \nz.mem_2625_sv2v_reg  <= w_data_i[25];
      \nz.mem_2624_sv2v_reg  <= w_data_i[24];
      \nz.mem_2623_sv2v_reg  <= w_data_i[23];
      \nz.mem_2622_sv2v_reg  <= w_data_i[22];
      \nz.mem_2621_sv2v_reg  <= w_data_i[21];
      \nz.mem_2620_sv2v_reg  <= w_data_i[20];
      \nz.mem_2619_sv2v_reg  <= w_data_i[19];
      \nz.mem_2618_sv2v_reg  <= w_data_i[18];
      \nz.mem_2617_sv2v_reg  <= w_data_i[17];
      \nz.mem_2616_sv2v_reg  <= w_data_i[16];
      \nz.mem_2615_sv2v_reg  <= w_data_i[15];
      \nz.mem_2614_sv2v_reg  <= w_data_i[14];
      \nz.mem_2613_sv2v_reg  <= w_data_i[13];
      \nz.mem_2612_sv2v_reg  <= w_data_i[12];
      \nz.mem_2611_sv2v_reg  <= w_data_i[11];
      \nz.mem_2610_sv2v_reg  <= w_data_i[10];
      \nz.mem_2609_sv2v_reg  <= w_data_i[9];
      \nz.mem_2608_sv2v_reg  <= w_data_i[8];
      \nz.mem_2607_sv2v_reg  <= w_data_i[7];
      \nz.mem_2606_sv2v_reg  <= w_data_i[6];
      \nz.mem_2605_sv2v_reg  <= w_data_i[5];
      \nz.mem_2604_sv2v_reg  <= w_data_i[4];
      \nz.mem_2603_sv2v_reg  <= w_data_i[3];
      \nz.mem_2602_sv2v_reg  <= w_data_i[2];
      \nz.mem_2601_sv2v_reg  <= w_data_i[1];
      \nz.mem_2600_sv2v_reg  <= w_data_i[0];
    end 
    if(N256) begin
      \nz.mem_2599_sv2v_reg  <= w_data_i[49];
      \nz.mem_2598_sv2v_reg  <= w_data_i[48];
      \nz.mem_2597_sv2v_reg  <= w_data_i[47];
      \nz.mem_2596_sv2v_reg  <= w_data_i[46];
      \nz.mem_2595_sv2v_reg  <= w_data_i[45];
      \nz.mem_2594_sv2v_reg  <= w_data_i[44];
      \nz.mem_2593_sv2v_reg  <= w_data_i[43];
      \nz.mem_2592_sv2v_reg  <= w_data_i[42];
      \nz.mem_2591_sv2v_reg  <= w_data_i[41];
      \nz.mem_2590_sv2v_reg  <= w_data_i[40];
      \nz.mem_2589_sv2v_reg  <= w_data_i[39];
      \nz.mem_2588_sv2v_reg  <= w_data_i[38];
      \nz.mem_2587_sv2v_reg  <= w_data_i[37];
      \nz.mem_2586_sv2v_reg  <= w_data_i[36];
      \nz.mem_2585_sv2v_reg  <= w_data_i[35];
      \nz.mem_2584_sv2v_reg  <= w_data_i[34];
      \nz.mem_2583_sv2v_reg  <= w_data_i[33];
      \nz.mem_2582_sv2v_reg  <= w_data_i[32];
      \nz.mem_2581_sv2v_reg  <= w_data_i[31];
      \nz.mem_2580_sv2v_reg  <= w_data_i[30];
      \nz.mem_2579_sv2v_reg  <= w_data_i[29];
      \nz.mem_2578_sv2v_reg  <= w_data_i[28];
      \nz.mem_2577_sv2v_reg  <= w_data_i[27];
      \nz.mem_2576_sv2v_reg  <= w_data_i[26];
      \nz.mem_2575_sv2v_reg  <= w_data_i[25];
      \nz.mem_2574_sv2v_reg  <= w_data_i[24];
      \nz.mem_2573_sv2v_reg  <= w_data_i[23];
      \nz.mem_2572_sv2v_reg  <= w_data_i[22];
      \nz.mem_2571_sv2v_reg  <= w_data_i[21];
      \nz.mem_2570_sv2v_reg  <= w_data_i[20];
      \nz.mem_2569_sv2v_reg  <= w_data_i[19];
      \nz.mem_2568_sv2v_reg  <= w_data_i[18];
      \nz.mem_2567_sv2v_reg  <= w_data_i[17];
      \nz.mem_2566_sv2v_reg  <= w_data_i[16];
      \nz.mem_2565_sv2v_reg  <= w_data_i[15];
      \nz.mem_2564_sv2v_reg  <= w_data_i[14];
      \nz.mem_2563_sv2v_reg  <= w_data_i[13];
      \nz.mem_2562_sv2v_reg  <= w_data_i[12];
      \nz.mem_2561_sv2v_reg  <= w_data_i[11];
      \nz.mem_2560_sv2v_reg  <= w_data_i[10];
      \nz.mem_2559_sv2v_reg  <= w_data_i[9];
      \nz.mem_2558_sv2v_reg  <= w_data_i[8];
      \nz.mem_2557_sv2v_reg  <= w_data_i[7];
      \nz.mem_2556_sv2v_reg  <= w_data_i[6];
      \nz.mem_2555_sv2v_reg  <= w_data_i[5];
      \nz.mem_2554_sv2v_reg  <= w_data_i[4];
      \nz.mem_2553_sv2v_reg  <= w_data_i[3];
      \nz.mem_2552_sv2v_reg  <= w_data_i[2];
      \nz.mem_2551_sv2v_reg  <= w_data_i[1];
      \nz.mem_2550_sv2v_reg  <= w_data_i[0];
    end 
    if(N255) begin
      \nz.mem_2549_sv2v_reg  <= w_data_i[49];
      \nz.mem_2548_sv2v_reg  <= w_data_i[48];
      \nz.mem_2547_sv2v_reg  <= w_data_i[47];
      \nz.mem_2546_sv2v_reg  <= w_data_i[46];
      \nz.mem_2545_sv2v_reg  <= w_data_i[45];
      \nz.mem_2544_sv2v_reg  <= w_data_i[44];
      \nz.mem_2543_sv2v_reg  <= w_data_i[43];
      \nz.mem_2542_sv2v_reg  <= w_data_i[42];
      \nz.mem_2541_sv2v_reg  <= w_data_i[41];
      \nz.mem_2540_sv2v_reg  <= w_data_i[40];
      \nz.mem_2539_sv2v_reg  <= w_data_i[39];
      \nz.mem_2538_sv2v_reg  <= w_data_i[38];
      \nz.mem_2537_sv2v_reg  <= w_data_i[37];
      \nz.mem_2536_sv2v_reg  <= w_data_i[36];
      \nz.mem_2535_sv2v_reg  <= w_data_i[35];
      \nz.mem_2534_sv2v_reg  <= w_data_i[34];
      \nz.mem_2533_sv2v_reg  <= w_data_i[33];
      \nz.mem_2532_sv2v_reg  <= w_data_i[32];
      \nz.mem_2531_sv2v_reg  <= w_data_i[31];
      \nz.mem_2530_sv2v_reg  <= w_data_i[30];
      \nz.mem_2529_sv2v_reg  <= w_data_i[29];
      \nz.mem_2528_sv2v_reg  <= w_data_i[28];
      \nz.mem_2527_sv2v_reg  <= w_data_i[27];
      \nz.mem_2526_sv2v_reg  <= w_data_i[26];
      \nz.mem_2525_sv2v_reg  <= w_data_i[25];
      \nz.mem_2524_sv2v_reg  <= w_data_i[24];
      \nz.mem_2523_sv2v_reg  <= w_data_i[23];
      \nz.mem_2522_sv2v_reg  <= w_data_i[22];
      \nz.mem_2521_sv2v_reg  <= w_data_i[21];
      \nz.mem_2520_sv2v_reg  <= w_data_i[20];
      \nz.mem_2519_sv2v_reg  <= w_data_i[19];
      \nz.mem_2518_sv2v_reg  <= w_data_i[18];
      \nz.mem_2517_sv2v_reg  <= w_data_i[17];
      \nz.mem_2516_sv2v_reg  <= w_data_i[16];
      \nz.mem_2515_sv2v_reg  <= w_data_i[15];
      \nz.mem_2514_sv2v_reg  <= w_data_i[14];
      \nz.mem_2513_sv2v_reg  <= w_data_i[13];
      \nz.mem_2512_sv2v_reg  <= w_data_i[12];
      \nz.mem_2511_sv2v_reg  <= w_data_i[11];
      \nz.mem_2510_sv2v_reg  <= w_data_i[10];
      \nz.mem_2509_sv2v_reg  <= w_data_i[9];
      \nz.mem_2508_sv2v_reg  <= w_data_i[8];
      \nz.mem_2507_sv2v_reg  <= w_data_i[7];
      \nz.mem_2506_sv2v_reg  <= w_data_i[6];
      \nz.mem_2505_sv2v_reg  <= w_data_i[5];
      \nz.mem_2504_sv2v_reg  <= w_data_i[4];
      \nz.mem_2503_sv2v_reg  <= w_data_i[3];
      \nz.mem_2502_sv2v_reg  <= w_data_i[2];
      \nz.mem_2501_sv2v_reg  <= w_data_i[1];
      \nz.mem_2500_sv2v_reg  <= w_data_i[0];
    end 
    if(N254) begin
      \nz.mem_2499_sv2v_reg  <= w_data_i[49];
      \nz.mem_2498_sv2v_reg  <= w_data_i[48];
      \nz.mem_2497_sv2v_reg  <= w_data_i[47];
      \nz.mem_2496_sv2v_reg  <= w_data_i[46];
      \nz.mem_2495_sv2v_reg  <= w_data_i[45];
      \nz.mem_2494_sv2v_reg  <= w_data_i[44];
      \nz.mem_2493_sv2v_reg  <= w_data_i[43];
      \nz.mem_2492_sv2v_reg  <= w_data_i[42];
      \nz.mem_2491_sv2v_reg  <= w_data_i[41];
      \nz.mem_2490_sv2v_reg  <= w_data_i[40];
      \nz.mem_2489_sv2v_reg  <= w_data_i[39];
      \nz.mem_2488_sv2v_reg  <= w_data_i[38];
      \nz.mem_2487_sv2v_reg  <= w_data_i[37];
      \nz.mem_2486_sv2v_reg  <= w_data_i[36];
      \nz.mem_2485_sv2v_reg  <= w_data_i[35];
      \nz.mem_2484_sv2v_reg  <= w_data_i[34];
      \nz.mem_2483_sv2v_reg  <= w_data_i[33];
      \nz.mem_2482_sv2v_reg  <= w_data_i[32];
      \nz.mem_2481_sv2v_reg  <= w_data_i[31];
      \nz.mem_2480_sv2v_reg  <= w_data_i[30];
      \nz.mem_2479_sv2v_reg  <= w_data_i[29];
      \nz.mem_2478_sv2v_reg  <= w_data_i[28];
      \nz.mem_2477_sv2v_reg  <= w_data_i[27];
      \nz.mem_2476_sv2v_reg  <= w_data_i[26];
      \nz.mem_2475_sv2v_reg  <= w_data_i[25];
      \nz.mem_2474_sv2v_reg  <= w_data_i[24];
      \nz.mem_2473_sv2v_reg  <= w_data_i[23];
      \nz.mem_2472_sv2v_reg  <= w_data_i[22];
      \nz.mem_2471_sv2v_reg  <= w_data_i[21];
      \nz.mem_2470_sv2v_reg  <= w_data_i[20];
      \nz.mem_2469_sv2v_reg  <= w_data_i[19];
      \nz.mem_2468_sv2v_reg  <= w_data_i[18];
      \nz.mem_2467_sv2v_reg  <= w_data_i[17];
      \nz.mem_2466_sv2v_reg  <= w_data_i[16];
      \nz.mem_2465_sv2v_reg  <= w_data_i[15];
      \nz.mem_2464_sv2v_reg  <= w_data_i[14];
      \nz.mem_2463_sv2v_reg  <= w_data_i[13];
      \nz.mem_2462_sv2v_reg  <= w_data_i[12];
      \nz.mem_2461_sv2v_reg  <= w_data_i[11];
      \nz.mem_2460_sv2v_reg  <= w_data_i[10];
      \nz.mem_2459_sv2v_reg  <= w_data_i[9];
      \nz.mem_2458_sv2v_reg  <= w_data_i[8];
      \nz.mem_2457_sv2v_reg  <= w_data_i[7];
      \nz.mem_2456_sv2v_reg  <= w_data_i[6];
      \nz.mem_2455_sv2v_reg  <= w_data_i[5];
      \nz.mem_2454_sv2v_reg  <= w_data_i[4];
      \nz.mem_2453_sv2v_reg  <= w_data_i[3];
      \nz.mem_2452_sv2v_reg  <= w_data_i[2];
      \nz.mem_2451_sv2v_reg  <= w_data_i[1];
      \nz.mem_2450_sv2v_reg  <= w_data_i[0];
    end 
    if(N253) begin
      \nz.mem_2449_sv2v_reg  <= w_data_i[49];
      \nz.mem_2448_sv2v_reg  <= w_data_i[48];
      \nz.mem_2447_sv2v_reg  <= w_data_i[47];
      \nz.mem_2446_sv2v_reg  <= w_data_i[46];
      \nz.mem_2445_sv2v_reg  <= w_data_i[45];
      \nz.mem_2444_sv2v_reg  <= w_data_i[44];
      \nz.mem_2443_sv2v_reg  <= w_data_i[43];
      \nz.mem_2442_sv2v_reg  <= w_data_i[42];
      \nz.mem_2441_sv2v_reg  <= w_data_i[41];
      \nz.mem_2440_sv2v_reg  <= w_data_i[40];
      \nz.mem_2439_sv2v_reg  <= w_data_i[39];
      \nz.mem_2438_sv2v_reg  <= w_data_i[38];
      \nz.mem_2437_sv2v_reg  <= w_data_i[37];
      \nz.mem_2436_sv2v_reg  <= w_data_i[36];
      \nz.mem_2435_sv2v_reg  <= w_data_i[35];
      \nz.mem_2434_sv2v_reg  <= w_data_i[34];
      \nz.mem_2433_sv2v_reg  <= w_data_i[33];
      \nz.mem_2432_sv2v_reg  <= w_data_i[32];
      \nz.mem_2431_sv2v_reg  <= w_data_i[31];
      \nz.mem_2430_sv2v_reg  <= w_data_i[30];
      \nz.mem_2429_sv2v_reg  <= w_data_i[29];
      \nz.mem_2428_sv2v_reg  <= w_data_i[28];
      \nz.mem_2427_sv2v_reg  <= w_data_i[27];
      \nz.mem_2426_sv2v_reg  <= w_data_i[26];
      \nz.mem_2425_sv2v_reg  <= w_data_i[25];
      \nz.mem_2424_sv2v_reg  <= w_data_i[24];
      \nz.mem_2423_sv2v_reg  <= w_data_i[23];
      \nz.mem_2422_sv2v_reg  <= w_data_i[22];
      \nz.mem_2421_sv2v_reg  <= w_data_i[21];
      \nz.mem_2420_sv2v_reg  <= w_data_i[20];
      \nz.mem_2419_sv2v_reg  <= w_data_i[19];
      \nz.mem_2418_sv2v_reg  <= w_data_i[18];
      \nz.mem_2417_sv2v_reg  <= w_data_i[17];
      \nz.mem_2416_sv2v_reg  <= w_data_i[16];
      \nz.mem_2415_sv2v_reg  <= w_data_i[15];
      \nz.mem_2414_sv2v_reg  <= w_data_i[14];
      \nz.mem_2413_sv2v_reg  <= w_data_i[13];
      \nz.mem_2412_sv2v_reg  <= w_data_i[12];
      \nz.mem_2411_sv2v_reg  <= w_data_i[11];
      \nz.mem_2410_sv2v_reg  <= w_data_i[10];
      \nz.mem_2409_sv2v_reg  <= w_data_i[9];
      \nz.mem_2408_sv2v_reg  <= w_data_i[8];
      \nz.mem_2407_sv2v_reg  <= w_data_i[7];
      \nz.mem_2406_sv2v_reg  <= w_data_i[6];
      \nz.mem_2405_sv2v_reg  <= w_data_i[5];
      \nz.mem_2404_sv2v_reg  <= w_data_i[4];
      \nz.mem_2403_sv2v_reg  <= w_data_i[3];
      \nz.mem_2402_sv2v_reg  <= w_data_i[2];
      \nz.mem_2401_sv2v_reg  <= w_data_i[1];
      \nz.mem_2400_sv2v_reg  <= w_data_i[0];
    end 
    if(N252) begin
      \nz.mem_2399_sv2v_reg  <= w_data_i[49];
      \nz.mem_2398_sv2v_reg  <= w_data_i[48];
      \nz.mem_2397_sv2v_reg  <= w_data_i[47];
      \nz.mem_2396_sv2v_reg  <= w_data_i[46];
      \nz.mem_2395_sv2v_reg  <= w_data_i[45];
      \nz.mem_2394_sv2v_reg  <= w_data_i[44];
      \nz.mem_2393_sv2v_reg  <= w_data_i[43];
      \nz.mem_2392_sv2v_reg  <= w_data_i[42];
      \nz.mem_2391_sv2v_reg  <= w_data_i[41];
      \nz.mem_2390_sv2v_reg  <= w_data_i[40];
      \nz.mem_2389_sv2v_reg  <= w_data_i[39];
      \nz.mem_2388_sv2v_reg  <= w_data_i[38];
      \nz.mem_2387_sv2v_reg  <= w_data_i[37];
      \nz.mem_2386_sv2v_reg  <= w_data_i[36];
      \nz.mem_2385_sv2v_reg  <= w_data_i[35];
      \nz.mem_2384_sv2v_reg  <= w_data_i[34];
      \nz.mem_2383_sv2v_reg  <= w_data_i[33];
      \nz.mem_2382_sv2v_reg  <= w_data_i[32];
      \nz.mem_2381_sv2v_reg  <= w_data_i[31];
      \nz.mem_2380_sv2v_reg  <= w_data_i[30];
      \nz.mem_2379_sv2v_reg  <= w_data_i[29];
      \nz.mem_2378_sv2v_reg  <= w_data_i[28];
      \nz.mem_2377_sv2v_reg  <= w_data_i[27];
      \nz.mem_2376_sv2v_reg  <= w_data_i[26];
      \nz.mem_2375_sv2v_reg  <= w_data_i[25];
      \nz.mem_2374_sv2v_reg  <= w_data_i[24];
      \nz.mem_2373_sv2v_reg  <= w_data_i[23];
      \nz.mem_2372_sv2v_reg  <= w_data_i[22];
      \nz.mem_2371_sv2v_reg  <= w_data_i[21];
      \nz.mem_2370_sv2v_reg  <= w_data_i[20];
      \nz.mem_2369_sv2v_reg  <= w_data_i[19];
      \nz.mem_2368_sv2v_reg  <= w_data_i[18];
      \nz.mem_2367_sv2v_reg  <= w_data_i[17];
      \nz.mem_2366_sv2v_reg  <= w_data_i[16];
      \nz.mem_2365_sv2v_reg  <= w_data_i[15];
      \nz.mem_2364_sv2v_reg  <= w_data_i[14];
      \nz.mem_2363_sv2v_reg  <= w_data_i[13];
      \nz.mem_2362_sv2v_reg  <= w_data_i[12];
      \nz.mem_2361_sv2v_reg  <= w_data_i[11];
      \nz.mem_2360_sv2v_reg  <= w_data_i[10];
      \nz.mem_2359_sv2v_reg  <= w_data_i[9];
      \nz.mem_2358_sv2v_reg  <= w_data_i[8];
      \nz.mem_2357_sv2v_reg  <= w_data_i[7];
      \nz.mem_2356_sv2v_reg  <= w_data_i[6];
      \nz.mem_2355_sv2v_reg  <= w_data_i[5];
      \nz.mem_2354_sv2v_reg  <= w_data_i[4];
      \nz.mem_2353_sv2v_reg  <= w_data_i[3];
      \nz.mem_2352_sv2v_reg  <= w_data_i[2];
      \nz.mem_2351_sv2v_reg  <= w_data_i[1];
      \nz.mem_2350_sv2v_reg  <= w_data_i[0];
    end 
    if(N251) begin
      \nz.mem_2349_sv2v_reg  <= w_data_i[49];
      \nz.mem_2348_sv2v_reg  <= w_data_i[48];
      \nz.mem_2347_sv2v_reg  <= w_data_i[47];
      \nz.mem_2346_sv2v_reg  <= w_data_i[46];
      \nz.mem_2345_sv2v_reg  <= w_data_i[45];
      \nz.mem_2344_sv2v_reg  <= w_data_i[44];
      \nz.mem_2343_sv2v_reg  <= w_data_i[43];
      \nz.mem_2342_sv2v_reg  <= w_data_i[42];
      \nz.mem_2341_sv2v_reg  <= w_data_i[41];
      \nz.mem_2340_sv2v_reg  <= w_data_i[40];
      \nz.mem_2339_sv2v_reg  <= w_data_i[39];
      \nz.mem_2338_sv2v_reg  <= w_data_i[38];
      \nz.mem_2337_sv2v_reg  <= w_data_i[37];
      \nz.mem_2336_sv2v_reg  <= w_data_i[36];
      \nz.mem_2335_sv2v_reg  <= w_data_i[35];
      \nz.mem_2334_sv2v_reg  <= w_data_i[34];
      \nz.mem_2333_sv2v_reg  <= w_data_i[33];
      \nz.mem_2332_sv2v_reg  <= w_data_i[32];
      \nz.mem_2331_sv2v_reg  <= w_data_i[31];
      \nz.mem_2330_sv2v_reg  <= w_data_i[30];
      \nz.mem_2329_sv2v_reg  <= w_data_i[29];
      \nz.mem_2328_sv2v_reg  <= w_data_i[28];
      \nz.mem_2327_sv2v_reg  <= w_data_i[27];
      \nz.mem_2326_sv2v_reg  <= w_data_i[26];
      \nz.mem_2325_sv2v_reg  <= w_data_i[25];
      \nz.mem_2324_sv2v_reg  <= w_data_i[24];
      \nz.mem_2323_sv2v_reg  <= w_data_i[23];
      \nz.mem_2322_sv2v_reg  <= w_data_i[22];
      \nz.mem_2321_sv2v_reg  <= w_data_i[21];
      \nz.mem_2320_sv2v_reg  <= w_data_i[20];
      \nz.mem_2319_sv2v_reg  <= w_data_i[19];
      \nz.mem_2318_sv2v_reg  <= w_data_i[18];
      \nz.mem_2317_sv2v_reg  <= w_data_i[17];
      \nz.mem_2316_sv2v_reg  <= w_data_i[16];
      \nz.mem_2315_sv2v_reg  <= w_data_i[15];
      \nz.mem_2314_sv2v_reg  <= w_data_i[14];
      \nz.mem_2313_sv2v_reg  <= w_data_i[13];
      \nz.mem_2312_sv2v_reg  <= w_data_i[12];
      \nz.mem_2311_sv2v_reg  <= w_data_i[11];
      \nz.mem_2310_sv2v_reg  <= w_data_i[10];
      \nz.mem_2309_sv2v_reg  <= w_data_i[9];
      \nz.mem_2308_sv2v_reg  <= w_data_i[8];
      \nz.mem_2307_sv2v_reg  <= w_data_i[7];
      \nz.mem_2306_sv2v_reg  <= w_data_i[6];
      \nz.mem_2305_sv2v_reg  <= w_data_i[5];
      \nz.mem_2304_sv2v_reg  <= w_data_i[4];
      \nz.mem_2303_sv2v_reg  <= w_data_i[3];
      \nz.mem_2302_sv2v_reg  <= w_data_i[2];
      \nz.mem_2301_sv2v_reg  <= w_data_i[1];
      \nz.mem_2300_sv2v_reg  <= w_data_i[0];
    end 
    if(N250) begin
      \nz.mem_2299_sv2v_reg  <= w_data_i[49];
      \nz.mem_2298_sv2v_reg  <= w_data_i[48];
      \nz.mem_2297_sv2v_reg  <= w_data_i[47];
      \nz.mem_2296_sv2v_reg  <= w_data_i[46];
      \nz.mem_2295_sv2v_reg  <= w_data_i[45];
      \nz.mem_2294_sv2v_reg  <= w_data_i[44];
      \nz.mem_2293_sv2v_reg  <= w_data_i[43];
      \nz.mem_2292_sv2v_reg  <= w_data_i[42];
      \nz.mem_2291_sv2v_reg  <= w_data_i[41];
      \nz.mem_2290_sv2v_reg  <= w_data_i[40];
      \nz.mem_2289_sv2v_reg  <= w_data_i[39];
      \nz.mem_2288_sv2v_reg  <= w_data_i[38];
      \nz.mem_2287_sv2v_reg  <= w_data_i[37];
      \nz.mem_2286_sv2v_reg  <= w_data_i[36];
      \nz.mem_2285_sv2v_reg  <= w_data_i[35];
      \nz.mem_2284_sv2v_reg  <= w_data_i[34];
      \nz.mem_2283_sv2v_reg  <= w_data_i[33];
      \nz.mem_2282_sv2v_reg  <= w_data_i[32];
      \nz.mem_2281_sv2v_reg  <= w_data_i[31];
      \nz.mem_2280_sv2v_reg  <= w_data_i[30];
      \nz.mem_2279_sv2v_reg  <= w_data_i[29];
      \nz.mem_2278_sv2v_reg  <= w_data_i[28];
      \nz.mem_2277_sv2v_reg  <= w_data_i[27];
      \nz.mem_2276_sv2v_reg  <= w_data_i[26];
      \nz.mem_2275_sv2v_reg  <= w_data_i[25];
      \nz.mem_2274_sv2v_reg  <= w_data_i[24];
      \nz.mem_2273_sv2v_reg  <= w_data_i[23];
      \nz.mem_2272_sv2v_reg  <= w_data_i[22];
      \nz.mem_2271_sv2v_reg  <= w_data_i[21];
      \nz.mem_2270_sv2v_reg  <= w_data_i[20];
      \nz.mem_2269_sv2v_reg  <= w_data_i[19];
      \nz.mem_2268_sv2v_reg  <= w_data_i[18];
      \nz.mem_2267_sv2v_reg  <= w_data_i[17];
      \nz.mem_2266_sv2v_reg  <= w_data_i[16];
      \nz.mem_2265_sv2v_reg  <= w_data_i[15];
      \nz.mem_2264_sv2v_reg  <= w_data_i[14];
      \nz.mem_2263_sv2v_reg  <= w_data_i[13];
      \nz.mem_2262_sv2v_reg  <= w_data_i[12];
      \nz.mem_2261_sv2v_reg  <= w_data_i[11];
      \nz.mem_2260_sv2v_reg  <= w_data_i[10];
      \nz.mem_2259_sv2v_reg  <= w_data_i[9];
      \nz.mem_2258_sv2v_reg  <= w_data_i[8];
      \nz.mem_2257_sv2v_reg  <= w_data_i[7];
      \nz.mem_2256_sv2v_reg  <= w_data_i[6];
      \nz.mem_2255_sv2v_reg  <= w_data_i[5];
      \nz.mem_2254_sv2v_reg  <= w_data_i[4];
      \nz.mem_2253_sv2v_reg  <= w_data_i[3];
      \nz.mem_2252_sv2v_reg  <= w_data_i[2];
      \nz.mem_2251_sv2v_reg  <= w_data_i[1];
      \nz.mem_2250_sv2v_reg  <= w_data_i[0];
    end 
    if(N249) begin
      \nz.mem_2249_sv2v_reg  <= w_data_i[49];
      \nz.mem_2248_sv2v_reg  <= w_data_i[48];
      \nz.mem_2247_sv2v_reg  <= w_data_i[47];
      \nz.mem_2246_sv2v_reg  <= w_data_i[46];
      \nz.mem_2245_sv2v_reg  <= w_data_i[45];
      \nz.mem_2244_sv2v_reg  <= w_data_i[44];
      \nz.mem_2243_sv2v_reg  <= w_data_i[43];
      \nz.mem_2242_sv2v_reg  <= w_data_i[42];
      \nz.mem_2241_sv2v_reg  <= w_data_i[41];
      \nz.mem_2240_sv2v_reg  <= w_data_i[40];
      \nz.mem_2239_sv2v_reg  <= w_data_i[39];
      \nz.mem_2238_sv2v_reg  <= w_data_i[38];
      \nz.mem_2237_sv2v_reg  <= w_data_i[37];
      \nz.mem_2236_sv2v_reg  <= w_data_i[36];
      \nz.mem_2235_sv2v_reg  <= w_data_i[35];
      \nz.mem_2234_sv2v_reg  <= w_data_i[34];
      \nz.mem_2233_sv2v_reg  <= w_data_i[33];
      \nz.mem_2232_sv2v_reg  <= w_data_i[32];
      \nz.mem_2231_sv2v_reg  <= w_data_i[31];
      \nz.mem_2230_sv2v_reg  <= w_data_i[30];
      \nz.mem_2229_sv2v_reg  <= w_data_i[29];
      \nz.mem_2228_sv2v_reg  <= w_data_i[28];
      \nz.mem_2227_sv2v_reg  <= w_data_i[27];
      \nz.mem_2226_sv2v_reg  <= w_data_i[26];
      \nz.mem_2225_sv2v_reg  <= w_data_i[25];
      \nz.mem_2224_sv2v_reg  <= w_data_i[24];
      \nz.mem_2223_sv2v_reg  <= w_data_i[23];
      \nz.mem_2222_sv2v_reg  <= w_data_i[22];
      \nz.mem_2221_sv2v_reg  <= w_data_i[21];
      \nz.mem_2220_sv2v_reg  <= w_data_i[20];
      \nz.mem_2219_sv2v_reg  <= w_data_i[19];
      \nz.mem_2218_sv2v_reg  <= w_data_i[18];
      \nz.mem_2217_sv2v_reg  <= w_data_i[17];
      \nz.mem_2216_sv2v_reg  <= w_data_i[16];
      \nz.mem_2215_sv2v_reg  <= w_data_i[15];
      \nz.mem_2214_sv2v_reg  <= w_data_i[14];
      \nz.mem_2213_sv2v_reg  <= w_data_i[13];
      \nz.mem_2212_sv2v_reg  <= w_data_i[12];
      \nz.mem_2211_sv2v_reg  <= w_data_i[11];
      \nz.mem_2210_sv2v_reg  <= w_data_i[10];
      \nz.mem_2209_sv2v_reg  <= w_data_i[9];
      \nz.mem_2208_sv2v_reg  <= w_data_i[8];
      \nz.mem_2207_sv2v_reg  <= w_data_i[7];
      \nz.mem_2206_sv2v_reg  <= w_data_i[6];
      \nz.mem_2205_sv2v_reg  <= w_data_i[5];
      \nz.mem_2204_sv2v_reg  <= w_data_i[4];
      \nz.mem_2203_sv2v_reg  <= w_data_i[3];
      \nz.mem_2202_sv2v_reg  <= w_data_i[2];
      \nz.mem_2201_sv2v_reg  <= w_data_i[1];
      \nz.mem_2200_sv2v_reg  <= w_data_i[0];
    end 
    if(N248) begin
      \nz.mem_2199_sv2v_reg  <= w_data_i[49];
      \nz.mem_2198_sv2v_reg  <= w_data_i[48];
      \nz.mem_2197_sv2v_reg  <= w_data_i[47];
      \nz.mem_2196_sv2v_reg  <= w_data_i[46];
      \nz.mem_2195_sv2v_reg  <= w_data_i[45];
      \nz.mem_2194_sv2v_reg  <= w_data_i[44];
      \nz.mem_2193_sv2v_reg  <= w_data_i[43];
      \nz.mem_2192_sv2v_reg  <= w_data_i[42];
      \nz.mem_2191_sv2v_reg  <= w_data_i[41];
      \nz.mem_2190_sv2v_reg  <= w_data_i[40];
      \nz.mem_2189_sv2v_reg  <= w_data_i[39];
      \nz.mem_2188_sv2v_reg  <= w_data_i[38];
      \nz.mem_2187_sv2v_reg  <= w_data_i[37];
      \nz.mem_2186_sv2v_reg  <= w_data_i[36];
      \nz.mem_2185_sv2v_reg  <= w_data_i[35];
      \nz.mem_2184_sv2v_reg  <= w_data_i[34];
      \nz.mem_2183_sv2v_reg  <= w_data_i[33];
      \nz.mem_2182_sv2v_reg  <= w_data_i[32];
      \nz.mem_2181_sv2v_reg  <= w_data_i[31];
      \nz.mem_2180_sv2v_reg  <= w_data_i[30];
      \nz.mem_2179_sv2v_reg  <= w_data_i[29];
      \nz.mem_2178_sv2v_reg  <= w_data_i[28];
      \nz.mem_2177_sv2v_reg  <= w_data_i[27];
      \nz.mem_2176_sv2v_reg  <= w_data_i[26];
      \nz.mem_2175_sv2v_reg  <= w_data_i[25];
      \nz.mem_2174_sv2v_reg  <= w_data_i[24];
      \nz.mem_2173_sv2v_reg  <= w_data_i[23];
      \nz.mem_2172_sv2v_reg  <= w_data_i[22];
      \nz.mem_2171_sv2v_reg  <= w_data_i[21];
      \nz.mem_2170_sv2v_reg  <= w_data_i[20];
      \nz.mem_2169_sv2v_reg  <= w_data_i[19];
      \nz.mem_2168_sv2v_reg  <= w_data_i[18];
      \nz.mem_2167_sv2v_reg  <= w_data_i[17];
      \nz.mem_2166_sv2v_reg  <= w_data_i[16];
      \nz.mem_2165_sv2v_reg  <= w_data_i[15];
      \nz.mem_2164_sv2v_reg  <= w_data_i[14];
      \nz.mem_2163_sv2v_reg  <= w_data_i[13];
      \nz.mem_2162_sv2v_reg  <= w_data_i[12];
      \nz.mem_2161_sv2v_reg  <= w_data_i[11];
      \nz.mem_2160_sv2v_reg  <= w_data_i[10];
      \nz.mem_2159_sv2v_reg  <= w_data_i[9];
      \nz.mem_2158_sv2v_reg  <= w_data_i[8];
      \nz.mem_2157_sv2v_reg  <= w_data_i[7];
      \nz.mem_2156_sv2v_reg  <= w_data_i[6];
      \nz.mem_2155_sv2v_reg  <= w_data_i[5];
      \nz.mem_2154_sv2v_reg  <= w_data_i[4];
      \nz.mem_2153_sv2v_reg  <= w_data_i[3];
      \nz.mem_2152_sv2v_reg  <= w_data_i[2];
      \nz.mem_2151_sv2v_reg  <= w_data_i[1];
      \nz.mem_2150_sv2v_reg  <= w_data_i[0];
    end 
    if(N247) begin
      \nz.mem_2149_sv2v_reg  <= w_data_i[49];
      \nz.mem_2148_sv2v_reg  <= w_data_i[48];
      \nz.mem_2147_sv2v_reg  <= w_data_i[47];
      \nz.mem_2146_sv2v_reg  <= w_data_i[46];
      \nz.mem_2145_sv2v_reg  <= w_data_i[45];
      \nz.mem_2144_sv2v_reg  <= w_data_i[44];
      \nz.mem_2143_sv2v_reg  <= w_data_i[43];
      \nz.mem_2142_sv2v_reg  <= w_data_i[42];
      \nz.mem_2141_sv2v_reg  <= w_data_i[41];
      \nz.mem_2140_sv2v_reg  <= w_data_i[40];
      \nz.mem_2139_sv2v_reg  <= w_data_i[39];
      \nz.mem_2138_sv2v_reg  <= w_data_i[38];
      \nz.mem_2137_sv2v_reg  <= w_data_i[37];
      \nz.mem_2136_sv2v_reg  <= w_data_i[36];
      \nz.mem_2135_sv2v_reg  <= w_data_i[35];
      \nz.mem_2134_sv2v_reg  <= w_data_i[34];
      \nz.mem_2133_sv2v_reg  <= w_data_i[33];
      \nz.mem_2132_sv2v_reg  <= w_data_i[32];
      \nz.mem_2131_sv2v_reg  <= w_data_i[31];
      \nz.mem_2130_sv2v_reg  <= w_data_i[30];
      \nz.mem_2129_sv2v_reg  <= w_data_i[29];
      \nz.mem_2128_sv2v_reg  <= w_data_i[28];
      \nz.mem_2127_sv2v_reg  <= w_data_i[27];
      \nz.mem_2126_sv2v_reg  <= w_data_i[26];
      \nz.mem_2125_sv2v_reg  <= w_data_i[25];
      \nz.mem_2124_sv2v_reg  <= w_data_i[24];
      \nz.mem_2123_sv2v_reg  <= w_data_i[23];
      \nz.mem_2122_sv2v_reg  <= w_data_i[22];
      \nz.mem_2121_sv2v_reg  <= w_data_i[21];
      \nz.mem_2120_sv2v_reg  <= w_data_i[20];
      \nz.mem_2119_sv2v_reg  <= w_data_i[19];
      \nz.mem_2118_sv2v_reg  <= w_data_i[18];
      \nz.mem_2117_sv2v_reg  <= w_data_i[17];
      \nz.mem_2116_sv2v_reg  <= w_data_i[16];
      \nz.mem_2115_sv2v_reg  <= w_data_i[15];
      \nz.mem_2114_sv2v_reg  <= w_data_i[14];
      \nz.mem_2113_sv2v_reg  <= w_data_i[13];
      \nz.mem_2112_sv2v_reg  <= w_data_i[12];
      \nz.mem_2111_sv2v_reg  <= w_data_i[11];
      \nz.mem_2110_sv2v_reg  <= w_data_i[10];
      \nz.mem_2109_sv2v_reg  <= w_data_i[9];
      \nz.mem_2108_sv2v_reg  <= w_data_i[8];
      \nz.mem_2107_sv2v_reg  <= w_data_i[7];
      \nz.mem_2106_sv2v_reg  <= w_data_i[6];
      \nz.mem_2105_sv2v_reg  <= w_data_i[5];
      \nz.mem_2104_sv2v_reg  <= w_data_i[4];
      \nz.mem_2103_sv2v_reg  <= w_data_i[3];
      \nz.mem_2102_sv2v_reg  <= w_data_i[2];
      \nz.mem_2101_sv2v_reg  <= w_data_i[1];
      \nz.mem_2100_sv2v_reg  <= w_data_i[0];
    end 
    if(N246) begin
      \nz.mem_2099_sv2v_reg  <= w_data_i[49];
      \nz.mem_2098_sv2v_reg  <= w_data_i[48];
      \nz.mem_2097_sv2v_reg  <= w_data_i[47];
      \nz.mem_2096_sv2v_reg  <= w_data_i[46];
      \nz.mem_2095_sv2v_reg  <= w_data_i[45];
      \nz.mem_2094_sv2v_reg  <= w_data_i[44];
      \nz.mem_2093_sv2v_reg  <= w_data_i[43];
      \nz.mem_2092_sv2v_reg  <= w_data_i[42];
      \nz.mem_2091_sv2v_reg  <= w_data_i[41];
      \nz.mem_2090_sv2v_reg  <= w_data_i[40];
      \nz.mem_2089_sv2v_reg  <= w_data_i[39];
      \nz.mem_2088_sv2v_reg  <= w_data_i[38];
      \nz.mem_2087_sv2v_reg  <= w_data_i[37];
      \nz.mem_2086_sv2v_reg  <= w_data_i[36];
      \nz.mem_2085_sv2v_reg  <= w_data_i[35];
      \nz.mem_2084_sv2v_reg  <= w_data_i[34];
      \nz.mem_2083_sv2v_reg  <= w_data_i[33];
      \nz.mem_2082_sv2v_reg  <= w_data_i[32];
      \nz.mem_2081_sv2v_reg  <= w_data_i[31];
      \nz.mem_2080_sv2v_reg  <= w_data_i[30];
      \nz.mem_2079_sv2v_reg  <= w_data_i[29];
      \nz.mem_2078_sv2v_reg  <= w_data_i[28];
      \nz.mem_2077_sv2v_reg  <= w_data_i[27];
      \nz.mem_2076_sv2v_reg  <= w_data_i[26];
      \nz.mem_2075_sv2v_reg  <= w_data_i[25];
      \nz.mem_2074_sv2v_reg  <= w_data_i[24];
      \nz.mem_2073_sv2v_reg  <= w_data_i[23];
      \nz.mem_2072_sv2v_reg  <= w_data_i[22];
      \nz.mem_2071_sv2v_reg  <= w_data_i[21];
      \nz.mem_2070_sv2v_reg  <= w_data_i[20];
      \nz.mem_2069_sv2v_reg  <= w_data_i[19];
      \nz.mem_2068_sv2v_reg  <= w_data_i[18];
      \nz.mem_2067_sv2v_reg  <= w_data_i[17];
      \nz.mem_2066_sv2v_reg  <= w_data_i[16];
      \nz.mem_2065_sv2v_reg  <= w_data_i[15];
      \nz.mem_2064_sv2v_reg  <= w_data_i[14];
      \nz.mem_2063_sv2v_reg  <= w_data_i[13];
      \nz.mem_2062_sv2v_reg  <= w_data_i[12];
      \nz.mem_2061_sv2v_reg  <= w_data_i[11];
      \nz.mem_2060_sv2v_reg  <= w_data_i[10];
      \nz.mem_2059_sv2v_reg  <= w_data_i[9];
      \nz.mem_2058_sv2v_reg  <= w_data_i[8];
      \nz.mem_2057_sv2v_reg  <= w_data_i[7];
      \nz.mem_2056_sv2v_reg  <= w_data_i[6];
      \nz.mem_2055_sv2v_reg  <= w_data_i[5];
      \nz.mem_2054_sv2v_reg  <= w_data_i[4];
      \nz.mem_2053_sv2v_reg  <= w_data_i[3];
      \nz.mem_2052_sv2v_reg  <= w_data_i[2];
      \nz.mem_2051_sv2v_reg  <= w_data_i[1];
      \nz.mem_2050_sv2v_reg  <= w_data_i[0];
    end 
    if(N245) begin
      \nz.mem_2049_sv2v_reg  <= w_data_i[49];
      \nz.mem_2048_sv2v_reg  <= w_data_i[48];
      \nz.mem_2047_sv2v_reg  <= w_data_i[47];
      \nz.mem_2046_sv2v_reg  <= w_data_i[46];
      \nz.mem_2045_sv2v_reg  <= w_data_i[45];
      \nz.mem_2044_sv2v_reg  <= w_data_i[44];
      \nz.mem_2043_sv2v_reg  <= w_data_i[43];
      \nz.mem_2042_sv2v_reg  <= w_data_i[42];
      \nz.mem_2041_sv2v_reg  <= w_data_i[41];
      \nz.mem_2040_sv2v_reg  <= w_data_i[40];
      \nz.mem_2039_sv2v_reg  <= w_data_i[39];
      \nz.mem_2038_sv2v_reg  <= w_data_i[38];
      \nz.mem_2037_sv2v_reg  <= w_data_i[37];
      \nz.mem_2036_sv2v_reg  <= w_data_i[36];
      \nz.mem_2035_sv2v_reg  <= w_data_i[35];
      \nz.mem_2034_sv2v_reg  <= w_data_i[34];
      \nz.mem_2033_sv2v_reg  <= w_data_i[33];
      \nz.mem_2032_sv2v_reg  <= w_data_i[32];
      \nz.mem_2031_sv2v_reg  <= w_data_i[31];
      \nz.mem_2030_sv2v_reg  <= w_data_i[30];
      \nz.mem_2029_sv2v_reg  <= w_data_i[29];
      \nz.mem_2028_sv2v_reg  <= w_data_i[28];
      \nz.mem_2027_sv2v_reg  <= w_data_i[27];
      \nz.mem_2026_sv2v_reg  <= w_data_i[26];
      \nz.mem_2025_sv2v_reg  <= w_data_i[25];
      \nz.mem_2024_sv2v_reg  <= w_data_i[24];
      \nz.mem_2023_sv2v_reg  <= w_data_i[23];
      \nz.mem_2022_sv2v_reg  <= w_data_i[22];
      \nz.mem_2021_sv2v_reg  <= w_data_i[21];
      \nz.mem_2020_sv2v_reg  <= w_data_i[20];
      \nz.mem_2019_sv2v_reg  <= w_data_i[19];
      \nz.mem_2018_sv2v_reg  <= w_data_i[18];
      \nz.mem_2017_sv2v_reg  <= w_data_i[17];
      \nz.mem_2016_sv2v_reg  <= w_data_i[16];
      \nz.mem_2015_sv2v_reg  <= w_data_i[15];
      \nz.mem_2014_sv2v_reg  <= w_data_i[14];
      \nz.mem_2013_sv2v_reg  <= w_data_i[13];
      \nz.mem_2012_sv2v_reg  <= w_data_i[12];
      \nz.mem_2011_sv2v_reg  <= w_data_i[11];
      \nz.mem_2010_sv2v_reg  <= w_data_i[10];
      \nz.mem_2009_sv2v_reg  <= w_data_i[9];
      \nz.mem_2008_sv2v_reg  <= w_data_i[8];
      \nz.mem_2007_sv2v_reg  <= w_data_i[7];
      \nz.mem_2006_sv2v_reg  <= w_data_i[6];
      \nz.mem_2005_sv2v_reg  <= w_data_i[5];
      \nz.mem_2004_sv2v_reg  <= w_data_i[4];
      \nz.mem_2003_sv2v_reg  <= w_data_i[3];
      \nz.mem_2002_sv2v_reg  <= w_data_i[2];
      \nz.mem_2001_sv2v_reg  <= w_data_i[1];
      \nz.mem_2000_sv2v_reg  <= w_data_i[0];
    end 
    if(N244) begin
      \nz.mem_1999_sv2v_reg  <= w_data_i[49];
      \nz.mem_1998_sv2v_reg  <= w_data_i[48];
      \nz.mem_1997_sv2v_reg  <= w_data_i[47];
      \nz.mem_1996_sv2v_reg  <= w_data_i[46];
      \nz.mem_1995_sv2v_reg  <= w_data_i[45];
      \nz.mem_1994_sv2v_reg  <= w_data_i[44];
      \nz.mem_1993_sv2v_reg  <= w_data_i[43];
      \nz.mem_1992_sv2v_reg  <= w_data_i[42];
      \nz.mem_1991_sv2v_reg  <= w_data_i[41];
      \nz.mem_1990_sv2v_reg  <= w_data_i[40];
      \nz.mem_1989_sv2v_reg  <= w_data_i[39];
      \nz.mem_1988_sv2v_reg  <= w_data_i[38];
      \nz.mem_1987_sv2v_reg  <= w_data_i[37];
      \nz.mem_1986_sv2v_reg  <= w_data_i[36];
      \nz.mem_1985_sv2v_reg  <= w_data_i[35];
      \nz.mem_1984_sv2v_reg  <= w_data_i[34];
      \nz.mem_1983_sv2v_reg  <= w_data_i[33];
      \nz.mem_1982_sv2v_reg  <= w_data_i[32];
      \nz.mem_1981_sv2v_reg  <= w_data_i[31];
      \nz.mem_1980_sv2v_reg  <= w_data_i[30];
      \nz.mem_1979_sv2v_reg  <= w_data_i[29];
      \nz.mem_1978_sv2v_reg  <= w_data_i[28];
      \nz.mem_1977_sv2v_reg  <= w_data_i[27];
      \nz.mem_1976_sv2v_reg  <= w_data_i[26];
      \nz.mem_1975_sv2v_reg  <= w_data_i[25];
      \nz.mem_1974_sv2v_reg  <= w_data_i[24];
      \nz.mem_1973_sv2v_reg  <= w_data_i[23];
      \nz.mem_1972_sv2v_reg  <= w_data_i[22];
      \nz.mem_1971_sv2v_reg  <= w_data_i[21];
      \nz.mem_1970_sv2v_reg  <= w_data_i[20];
      \nz.mem_1969_sv2v_reg  <= w_data_i[19];
      \nz.mem_1968_sv2v_reg  <= w_data_i[18];
      \nz.mem_1967_sv2v_reg  <= w_data_i[17];
      \nz.mem_1966_sv2v_reg  <= w_data_i[16];
      \nz.mem_1965_sv2v_reg  <= w_data_i[15];
      \nz.mem_1964_sv2v_reg  <= w_data_i[14];
      \nz.mem_1963_sv2v_reg  <= w_data_i[13];
      \nz.mem_1962_sv2v_reg  <= w_data_i[12];
      \nz.mem_1961_sv2v_reg  <= w_data_i[11];
      \nz.mem_1960_sv2v_reg  <= w_data_i[10];
      \nz.mem_1959_sv2v_reg  <= w_data_i[9];
      \nz.mem_1958_sv2v_reg  <= w_data_i[8];
      \nz.mem_1957_sv2v_reg  <= w_data_i[7];
      \nz.mem_1956_sv2v_reg  <= w_data_i[6];
      \nz.mem_1955_sv2v_reg  <= w_data_i[5];
      \nz.mem_1954_sv2v_reg  <= w_data_i[4];
      \nz.mem_1953_sv2v_reg  <= w_data_i[3];
      \nz.mem_1952_sv2v_reg  <= w_data_i[2];
      \nz.mem_1951_sv2v_reg  <= w_data_i[1];
      \nz.mem_1950_sv2v_reg  <= w_data_i[0];
    end 
    if(N243) begin
      \nz.mem_1949_sv2v_reg  <= w_data_i[49];
      \nz.mem_1948_sv2v_reg  <= w_data_i[48];
      \nz.mem_1947_sv2v_reg  <= w_data_i[47];
      \nz.mem_1946_sv2v_reg  <= w_data_i[46];
      \nz.mem_1945_sv2v_reg  <= w_data_i[45];
      \nz.mem_1944_sv2v_reg  <= w_data_i[44];
      \nz.mem_1943_sv2v_reg  <= w_data_i[43];
      \nz.mem_1942_sv2v_reg  <= w_data_i[42];
      \nz.mem_1941_sv2v_reg  <= w_data_i[41];
      \nz.mem_1940_sv2v_reg  <= w_data_i[40];
      \nz.mem_1939_sv2v_reg  <= w_data_i[39];
      \nz.mem_1938_sv2v_reg  <= w_data_i[38];
      \nz.mem_1937_sv2v_reg  <= w_data_i[37];
      \nz.mem_1936_sv2v_reg  <= w_data_i[36];
      \nz.mem_1935_sv2v_reg  <= w_data_i[35];
      \nz.mem_1934_sv2v_reg  <= w_data_i[34];
      \nz.mem_1933_sv2v_reg  <= w_data_i[33];
      \nz.mem_1932_sv2v_reg  <= w_data_i[32];
      \nz.mem_1931_sv2v_reg  <= w_data_i[31];
      \nz.mem_1930_sv2v_reg  <= w_data_i[30];
      \nz.mem_1929_sv2v_reg  <= w_data_i[29];
      \nz.mem_1928_sv2v_reg  <= w_data_i[28];
      \nz.mem_1927_sv2v_reg  <= w_data_i[27];
      \nz.mem_1926_sv2v_reg  <= w_data_i[26];
      \nz.mem_1925_sv2v_reg  <= w_data_i[25];
      \nz.mem_1924_sv2v_reg  <= w_data_i[24];
      \nz.mem_1923_sv2v_reg  <= w_data_i[23];
      \nz.mem_1922_sv2v_reg  <= w_data_i[22];
      \nz.mem_1921_sv2v_reg  <= w_data_i[21];
      \nz.mem_1920_sv2v_reg  <= w_data_i[20];
      \nz.mem_1919_sv2v_reg  <= w_data_i[19];
      \nz.mem_1918_sv2v_reg  <= w_data_i[18];
      \nz.mem_1917_sv2v_reg  <= w_data_i[17];
      \nz.mem_1916_sv2v_reg  <= w_data_i[16];
      \nz.mem_1915_sv2v_reg  <= w_data_i[15];
      \nz.mem_1914_sv2v_reg  <= w_data_i[14];
      \nz.mem_1913_sv2v_reg  <= w_data_i[13];
      \nz.mem_1912_sv2v_reg  <= w_data_i[12];
      \nz.mem_1911_sv2v_reg  <= w_data_i[11];
      \nz.mem_1910_sv2v_reg  <= w_data_i[10];
      \nz.mem_1909_sv2v_reg  <= w_data_i[9];
      \nz.mem_1908_sv2v_reg  <= w_data_i[8];
      \nz.mem_1907_sv2v_reg  <= w_data_i[7];
      \nz.mem_1906_sv2v_reg  <= w_data_i[6];
      \nz.mem_1905_sv2v_reg  <= w_data_i[5];
      \nz.mem_1904_sv2v_reg  <= w_data_i[4];
      \nz.mem_1903_sv2v_reg  <= w_data_i[3];
      \nz.mem_1902_sv2v_reg  <= w_data_i[2];
      \nz.mem_1901_sv2v_reg  <= w_data_i[1];
      \nz.mem_1900_sv2v_reg  <= w_data_i[0];
    end 
    if(N242) begin
      \nz.mem_1899_sv2v_reg  <= w_data_i[49];
      \nz.mem_1898_sv2v_reg  <= w_data_i[48];
      \nz.mem_1897_sv2v_reg  <= w_data_i[47];
      \nz.mem_1896_sv2v_reg  <= w_data_i[46];
      \nz.mem_1895_sv2v_reg  <= w_data_i[45];
      \nz.mem_1894_sv2v_reg  <= w_data_i[44];
      \nz.mem_1893_sv2v_reg  <= w_data_i[43];
      \nz.mem_1892_sv2v_reg  <= w_data_i[42];
      \nz.mem_1891_sv2v_reg  <= w_data_i[41];
      \nz.mem_1890_sv2v_reg  <= w_data_i[40];
      \nz.mem_1889_sv2v_reg  <= w_data_i[39];
      \nz.mem_1888_sv2v_reg  <= w_data_i[38];
      \nz.mem_1887_sv2v_reg  <= w_data_i[37];
      \nz.mem_1886_sv2v_reg  <= w_data_i[36];
      \nz.mem_1885_sv2v_reg  <= w_data_i[35];
      \nz.mem_1884_sv2v_reg  <= w_data_i[34];
      \nz.mem_1883_sv2v_reg  <= w_data_i[33];
      \nz.mem_1882_sv2v_reg  <= w_data_i[32];
      \nz.mem_1881_sv2v_reg  <= w_data_i[31];
      \nz.mem_1880_sv2v_reg  <= w_data_i[30];
      \nz.mem_1879_sv2v_reg  <= w_data_i[29];
      \nz.mem_1878_sv2v_reg  <= w_data_i[28];
      \nz.mem_1877_sv2v_reg  <= w_data_i[27];
      \nz.mem_1876_sv2v_reg  <= w_data_i[26];
      \nz.mem_1875_sv2v_reg  <= w_data_i[25];
      \nz.mem_1874_sv2v_reg  <= w_data_i[24];
      \nz.mem_1873_sv2v_reg  <= w_data_i[23];
      \nz.mem_1872_sv2v_reg  <= w_data_i[22];
      \nz.mem_1871_sv2v_reg  <= w_data_i[21];
      \nz.mem_1870_sv2v_reg  <= w_data_i[20];
      \nz.mem_1869_sv2v_reg  <= w_data_i[19];
      \nz.mem_1868_sv2v_reg  <= w_data_i[18];
      \nz.mem_1867_sv2v_reg  <= w_data_i[17];
      \nz.mem_1866_sv2v_reg  <= w_data_i[16];
      \nz.mem_1865_sv2v_reg  <= w_data_i[15];
      \nz.mem_1864_sv2v_reg  <= w_data_i[14];
      \nz.mem_1863_sv2v_reg  <= w_data_i[13];
      \nz.mem_1862_sv2v_reg  <= w_data_i[12];
      \nz.mem_1861_sv2v_reg  <= w_data_i[11];
      \nz.mem_1860_sv2v_reg  <= w_data_i[10];
      \nz.mem_1859_sv2v_reg  <= w_data_i[9];
      \nz.mem_1858_sv2v_reg  <= w_data_i[8];
      \nz.mem_1857_sv2v_reg  <= w_data_i[7];
      \nz.mem_1856_sv2v_reg  <= w_data_i[6];
      \nz.mem_1855_sv2v_reg  <= w_data_i[5];
      \nz.mem_1854_sv2v_reg  <= w_data_i[4];
      \nz.mem_1853_sv2v_reg  <= w_data_i[3];
      \nz.mem_1852_sv2v_reg  <= w_data_i[2];
      \nz.mem_1851_sv2v_reg  <= w_data_i[1];
      \nz.mem_1850_sv2v_reg  <= w_data_i[0];
    end 
    if(N241) begin
      \nz.mem_1849_sv2v_reg  <= w_data_i[49];
      \nz.mem_1848_sv2v_reg  <= w_data_i[48];
      \nz.mem_1847_sv2v_reg  <= w_data_i[47];
      \nz.mem_1846_sv2v_reg  <= w_data_i[46];
      \nz.mem_1845_sv2v_reg  <= w_data_i[45];
      \nz.mem_1844_sv2v_reg  <= w_data_i[44];
      \nz.mem_1843_sv2v_reg  <= w_data_i[43];
      \nz.mem_1842_sv2v_reg  <= w_data_i[42];
      \nz.mem_1841_sv2v_reg  <= w_data_i[41];
      \nz.mem_1840_sv2v_reg  <= w_data_i[40];
      \nz.mem_1839_sv2v_reg  <= w_data_i[39];
      \nz.mem_1838_sv2v_reg  <= w_data_i[38];
      \nz.mem_1837_sv2v_reg  <= w_data_i[37];
      \nz.mem_1836_sv2v_reg  <= w_data_i[36];
      \nz.mem_1835_sv2v_reg  <= w_data_i[35];
      \nz.mem_1834_sv2v_reg  <= w_data_i[34];
      \nz.mem_1833_sv2v_reg  <= w_data_i[33];
      \nz.mem_1832_sv2v_reg  <= w_data_i[32];
      \nz.mem_1831_sv2v_reg  <= w_data_i[31];
      \nz.mem_1830_sv2v_reg  <= w_data_i[30];
      \nz.mem_1829_sv2v_reg  <= w_data_i[29];
      \nz.mem_1828_sv2v_reg  <= w_data_i[28];
      \nz.mem_1827_sv2v_reg  <= w_data_i[27];
      \nz.mem_1826_sv2v_reg  <= w_data_i[26];
      \nz.mem_1825_sv2v_reg  <= w_data_i[25];
      \nz.mem_1824_sv2v_reg  <= w_data_i[24];
      \nz.mem_1823_sv2v_reg  <= w_data_i[23];
      \nz.mem_1822_sv2v_reg  <= w_data_i[22];
      \nz.mem_1821_sv2v_reg  <= w_data_i[21];
      \nz.mem_1820_sv2v_reg  <= w_data_i[20];
      \nz.mem_1819_sv2v_reg  <= w_data_i[19];
      \nz.mem_1818_sv2v_reg  <= w_data_i[18];
      \nz.mem_1817_sv2v_reg  <= w_data_i[17];
      \nz.mem_1816_sv2v_reg  <= w_data_i[16];
      \nz.mem_1815_sv2v_reg  <= w_data_i[15];
      \nz.mem_1814_sv2v_reg  <= w_data_i[14];
      \nz.mem_1813_sv2v_reg  <= w_data_i[13];
      \nz.mem_1812_sv2v_reg  <= w_data_i[12];
      \nz.mem_1811_sv2v_reg  <= w_data_i[11];
      \nz.mem_1810_sv2v_reg  <= w_data_i[10];
      \nz.mem_1809_sv2v_reg  <= w_data_i[9];
      \nz.mem_1808_sv2v_reg  <= w_data_i[8];
      \nz.mem_1807_sv2v_reg  <= w_data_i[7];
      \nz.mem_1806_sv2v_reg  <= w_data_i[6];
      \nz.mem_1805_sv2v_reg  <= w_data_i[5];
      \nz.mem_1804_sv2v_reg  <= w_data_i[4];
      \nz.mem_1803_sv2v_reg  <= w_data_i[3];
      \nz.mem_1802_sv2v_reg  <= w_data_i[2];
      \nz.mem_1801_sv2v_reg  <= w_data_i[1];
      \nz.mem_1800_sv2v_reg  <= w_data_i[0];
    end 
    if(N240) begin
      \nz.mem_1799_sv2v_reg  <= w_data_i[49];
      \nz.mem_1798_sv2v_reg  <= w_data_i[48];
      \nz.mem_1797_sv2v_reg  <= w_data_i[47];
      \nz.mem_1796_sv2v_reg  <= w_data_i[46];
      \nz.mem_1795_sv2v_reg  <= w_data_i[45];
      \nz.mem_1794_sv2v_reg  <= w_data_i[44];
      \nz.mem_1793_sv2v_reg  <= w_data_i[43];
      \nz.mem_1792_sv2v_reg  <= w_data_i[42];
      \nz.mem_1791_sv2v_reg  <= w_data_i[41];
      \nz.mem_1790_sv2v_reg  <= w_data_i[40];
      \nz.mem_1789_sv2v_reg  <= w_data_i[39];
      \nz.mem_1788_sv2v_reg  <= w_data_i[38];
      \nz.mem_1787_sv2v_reg  <= w_data_i[37];
      \nz.mem_1786_sv2v_reg  <= w_data_i[36];
      \nz.mem_1785_sv2v_reg  <= w_data_i[35];
      \nz.mem_1784_sv2v_reg  <= w_data_i[34];
      \nz.mem_1783_sv2v_reg  <= w_data_i[33];
      \nz.mem_1782_sv2v_reg  <= w_data_i[32];
      \nz.mem_1781_sv2v_reg  <= w_data_i[31];
      \nz.mem_1780_sv2v_reg  <= w_data_i[30];
      \nz.mem_1779_sv2v_reg  <= w_data_i[29];
      \nz.mem_1778_sv2v_reg  <= w_data_i[28];
      \nz.mem_1777_sv2v_reg  <= w_data_i[27];
      \nz.mem_1776_sv2v_reg  <= w_data_i[26];
      \nz.mem_1775_sv2v_reg  <= w_data_i[25];
      \nz.mem_1774_sv2v_reg  <= w_data_i[24];
      \nz.mem_1773_sv2v_reg  <= w_data_i[23];
      \nz.mem_1772_sv2v_reg  <= w_data_i[22];
      \nz.mem_1771_sv2v_reg  <= w_data_i[21];
      \nz.mem_1770_sv2v_reg  <= w_data_i[20];
      \nz.mem_1769_sv2v_reg  <= w_data_i[19];
      \nz.mem_1768_sv2v_reg  <= w_data_i[18];
      \nz.mem_1767_sv2v_reg  <= w_data_i[17];
      \nz.mem_1766_sv2v_reg  <= w_data_i[16];
      \nz.mem_1765_sv2v_reg  <= w_data_i[15];
      \nz.mem_1764_sv2v_reg  <= w_data_i[14];
      \nz.mem_1763_sv2v_reg  <= w_data_i[13];
      \nz.mem_1762_sv2v_reg  <= w_data_i[12];
      \nz.mem_1761_sv2v_reg  <= w_data_i[11];
      \nz.mem_1760_sv2v_reg  <= w_data_i[10];
      \nz.mem_1759_sv2v_reg  <= w_data_i[9];
      \nz.mem_1758_sv2v_reg  <= w_data_i[8];
      \nz.mem_1757_sv2v_reg  <= w_data_i[7];
      \nz.mem_1756_sv2v_reg  <= w_data_i[6];
      \nz.mem_1755_sv2v_reg  <= w_data_i[5];
      \nz.mem_1754_sv2v_reg  <= w_data_i[4];
      \nz.mem_1753_sv2v_reg  <= w_data_i[3];
      \nz.mem_1752_sv2v_reg  <= w_data_i[2];
      \nz.mem_1751_sv2v_reg  <= w_data_i[1];
      \nz.mem_1750_sv2v_reg  <= w_data_i[0];
    end 
    if(N239) begin
      \nz.mem_1749_sv2v_reg  <= w_data_i[49];
      \nz.mem_1748_sv2v_reg  <= w_data_i[48];
      \nz.mem_1747_sv2v_reg  <= w_data_i[47];
      \nz.mem_1746_sv2v_reg  <= w_data_i[46];
      \nz.mem_1745_sv2v_reg  <= w_data_i[45];
      \nz.mem_1744_sv2v_reg  <= w_data_i[44];
      \nz.mem_1743_sv2v_reg  <= w_data_i[43];
      \nz.mem_1742_sv2v_reg  <= w_data_i[42];
      \nz.mem_1741_sv2v_reg  <= w_data_i[41];
      \nz.mem_1740_sv2v_reg  <= w_data_i[40];
      \nz.mem_1739_sv2v_reg  <= w_data_i[39];
      \nz.mem_1738_sv2v_reg  <= w_data_i[38];
      \nz.mem_1737_sv2v_reg  <= w_data_i[37];
      \nz.mem_1736_sv2v_reg  <= w_data_i[36];
      \nz.mem_1735_sv2v_reg  <= w_data_i[35];
      \nz.mem_1734_sv2v_reg  <= w_data_i[34];
      \nz.mem_1733_sv2v_reg  <= w_data_i[33];
      \nz.mem_1732_sv2v_reg  <= w_data_i[32];
      \nz.mem_1731_sv2v_reg  <= w_data_i[31];
      \nz.mem_1730_sv2v_reg  <= w_data_i[30];
      \nz.mem_1729_sv2v_reg  <= w_data_i[29];
      \nz.mem_1728_sv2v_reg  <= w_data_i[28];
      \nz.mem_1727_sv2v_reg  <= w_data_i[27];
      \nz.mem_1726_sv2v_reg  <= w_data_i[26];
      \nz.mem_1725_sv2v_reg  <= w_data_i[25];
      \nz.mem_1724_sv2v_reg  <= w_data_i[24];
      \nz.mem_1723_sv2v_reg  <= w_data_i[23];
      \nz.mem_1722_sv2v_reg  <= w_data_i[22];
      \nz.mem_1721_sv2v_reg  <= w_data_i[21];
      \nz.mem_1720_sv2v_reg  <= w_data_i[20];
      \nz.mem_1719_sv2v_reg  <= w_data_i[19];
      \nz.mem_1718_sv2v_reg  <= w_data_i[18];
      \nz.mem_1717_sv2v_reg  <= w_data_i[17];
      \nz.mem_1716_sv2v_reg  <= w_data_i[16];
      \nz.mem_1715_sv2v_reg  <= w_data_i[15];
      \nz.mem_1714_sv2v_reg  <= w_data_i[14];
      \nz.mem_1713_sv2v_reg  <= w_data_i[13];
      \nz.mem_1712_sv2v_reg  <= w_data_i[12];
      \nz.mem_1711_sv2v_reg  <= w_data_i[11];
      \nz.mem_1710_sv2v_reg  <= w_data_i[10];
      \nz.mem_1709_sv2v_reg  <= w_data_i[9];
      \nz.mem_1708_sv2v_reg  <= w_data_i[8];
      \nz.mem_1707_sv2v_reg  <= w_data_i[7];
      \nz.mem_1706_sv2v_reg  <= w_data_i[6];
      \nz.mem_1705_sv2v_reg  <= w_data_i[5];
      \nz.mem_1704_sv2v_reg  <= w_data_i[4];
      \nz.mem_1703_sv2v_reg  <= w_data_i[3];
      \nz.mem_1702_sv2v_reg  <= w_data_i[2];
      \nz.mem_1701_sv2v_reg  <= w_data_i[1];
      \nz.mem_1700_sv2v_reg  <= w_data_i[0];
    end 
    if(N238) begin
      \nz.mem_1699_sv2v_reg  <= w_data_i[49];
      \nz.mem_1698_sv2v_reg  <= w_data_i[48];
      \nz.mem_1697_sv2v_reg  <= w_data_i[47];
      \nz.mem_1696_sv2v_reg  <= w_data_i[46];
      \nz.mem_1695_sv2v_reg  <= w_data_i[45];
      \nz.mem_1694_sv2v_reg  <= w_data_i[44];
      \nz.mem_1693_sv2v_reg  <= w_data_i[43];
      \nz.mem_1692_sv2v_reg  <= w_data_i[42];
      \nz.mem_1691_sv2v_reg  <= w_data_i[41];
      \nz.mem_1690_sv2v_reg  <= w_data_i[40];
      \nz.mem_1689_sv2v_reg  <= w_data_i[39];
      \nz.mem_1688_sv2v_reg  <= w_data_i[38];
      \nz.mem_1687_sv2v_reg  <= w_data_i[37];
      \nz.mem_1686_sv2v_reg  <= w_data_i[36];
      \nz.mem_1685_sv2v_reg  <= w_data_i[35];
      \nz.mem_1684_sv2v_reg  <= w_data_i[34];
      \nz.mem_1683_sv2v_reg  <= w_data_i[33];
      \nz.mem_1682_sv2v_reg  <= w_data_i[32];
      \nz.mem_1681_sv2v_reg  <= w_data_i[31];
      \nz.mem_1680_sv2v_reg  <= w_data_i[30];
      \nz.mem_1679_sv2v_reg  <= w_data_i[29];
      \nz.mem_1678_sv2v_reg  <= w_data_i[28];
      \nz.mem_1677_sv2v_reg  <= w_data_i[27];
      \nz.mem_1676_sv2v_reg  <= w_data_i[26];
      \nz.mem_1675_sv2v_reg  <= w_data_i[25];
      \nz.mem_1674_sv2v_reg  <= w_data_i[24];
      \nz.mem_1673_sv2v_reg  <= w_data_i[23];
      \nz.mem_1672_sv2v_reg  <= w_data_i[22];
      \nz.mem_1671_sv2v_reg  <= w_data_i[21];
      \nz.mem_1670_sv2v_reg  <= w_data_i[20];
      \nz.mem_1669_sv2v_reg  <= w_data_i[19];
      \nz.mem_1668_sv2v_reg  <= w_data_i[18];
      \nz.mem_1667_sv2v_reg  <= w_data_i[17];
      \nz.mem_1666_sv2v_reg  <= w_data_i[16];
      \nz.mem_1665_sv2v_reg  <= w_data_i[15];
      \nz.mem_1664_sv2v_reg  <= w_data_i[14];
      \nz.mem_1663_sv2v_reg  <= w_data_i[13];
      \nz.mem_1662_sv2v_reg  <= w_data_i[12];
      \nz.mem_1661_sv2v_reg  <= w_data_i[11];
      \nz.mem_1660_sv2v_reg  <= w_data_i[10];
      \nz.mem_1659_sv2v_reg  <= w_data_i[9];
      \nz.mem_1658_sv2v_reg  <= w_data_i[8];
      \nz.mem_1657_sv2v_reg  <= w_data_i[7];
      \nz.mem_1656_sv2v_reg  <= w_data_i[6];
      \nz.mem_1655_sv2v_reg  <= w_data_i[5];
      \nz.mem_1654_sv2v_reg  <= w_data_i[4];
      \nz.mem_1653_sv2v_reg  <= w_data_i[3];
      \nz.mem_1652_sv2v_reg  <= w_data_i[2];
      \nz.mem_1651_sv2v_reg  <= w_data_i[1];
      \nz.mem_1650_sv2v_reg  <= w_data_i[0];
    end 
    if(N237) begin
      \nz.mem_1649_sv2v_reg  <= w_data_i[49];
      \nz.mem_1648_sv2v_reg  <= w_data_i[48];
      \nz.mem_1647_sv2v_reg  <= w_data_i[47];
      \nz.mem_1646_sv2v_reg  <= w_data_i[46];
      \nz.mem_1645_sv2v_reg  <= w_data_i[45];
      \nz.mem_1644_sv2v_reg  <= w_data_i[44];
      \nz.mem_1643_sv2v_reg  <= w_data_i[43];
      \nz.mem_1642_sv2v_reg  <= w_data_i[42];
      \nz.mem_1641_sv2v_reg  <= w_data_i[41];
      \nz.mem_1640_sv2v_reg  <= w_data_i[40];
      \nz.mem_1639_sv2v_reg  <= w_data_i[39];
      \nz.mem_1638_sv2v_reg  <= w_data_i[38];
      \nz.mem_1637_sv2v_reg  <= w_data_i[37];
      \nz.mem_1636_sv2v_reg  <= w_data_i[36];
      \nz.mem_1635_sv2v_reg  <= w_data_i[35];
      \nz.mem_1634_sv2v_reg  <= w_data_i[34];
      \nz.mem_1633_sv2v_reg  <= w_data_i[33];
      \nz.mem_1632_sv2v_reg  <= w_data_i[32];
      \nz.mem_1631_sv2v_reg  <= w_data_i[31];
      \nz.mem_1630_sv2v_reg  <= w_data_i[30];
      \nz.mem_1629_sv2v_reg  <= w_data_i[29];
      \nz.mem_1628_sv2v_reg  <= w_data_i[28];
      \nz.mem_1627_sv2v_reg  <= w_data_i[27];
      \nz.mem_1626_sv2v_reg  <= w_data_i[26];
      \nz.mem_1625_sv2v_reg  <= w_data_i[25];
      \nz.mem_1624_sv2v_reg  <= w_data_i[24];
      \nz.mem_1623_sv2v_reg  <= w_data_i[23];
      \nz.mem_1622_sv2v_reg  <= w_data_i[22];
      \nz.mem_1621_sv2v_reg  <= w_data_i[21];
      \nz.mem_1620_sv2v_reg  <= w_data_i[20];
      \nz.mem_1619_sv2v_reg  <= w_data_i[19];
      \nz.mem_1618_sv2v_reg  <= w_data_i[18];
      \nz.mem_1617_sv2v_reg  <= w_data_i[17];
      \nz.mem_1616_sv2v_reg  <= w_data_i[16];
      \nz.mem_1615_sv2v_reg  <= w_data_i[15];
      \nz.mem_1614_sv2v_reg  <= w_data_i[14];
      \nz.mem_1613_sv2v_reg  <= w_data_i[13];
      \nz.mem_1612_sv2v_reg  <= w_data_i[12];
      \nz.mem_1611_sv2v_reg  <= w_data_i[11];
      \nz.mem_1610_sv2v_reg  <= w_data_i[10];
      \nz.mem_1609_sv2v_reg  <= w_data_i[9];
      \nz.mem_1608_sv2v_reg  <= w_data_i[8];
      \nz.mem_1607_sv2v_reg  <= w_data_i[7];
      \nz.mem_1606_sv2v_reg  <= w_data_i[6];
      \nz.mem_1605_sv2v_reg  <= w_data_i[5];
      \nz.mem_1604_sv2v_reg  <= w_data_i[4];
      \nz.mem_1603_sv2v_reg  <= w_data_i[3];
      \nz.mem_1602_sv2v_reg  <= w_data_i[2];
      \nz.mem_1601_sv2v_reg  <= w_data_i[1];
      \nz.mem_1600_sv2v_reg  <= w_data_i[0];
    end 
    if(N236) begin
      \nz.mem_1599_sv2v_reg  <= w_data_i[49];
      \nz.mem_1598_sv2v_reg  <= w_data_i[48];
      \nz.mem_1597_sv2v_reg  <= w_data_i[47];
      \nz.mem_1596_sv2v_reg  <= w_data_i[46];
      \nz.mem_1595_sv2v_reg  <= w_data_i[45];
      \nz.mem_1594_sv2v_reg  <= w_data_i[44];
      \nz.mem_1593_sv2v_reg  <= w_data_i[43];
      \nz.mem_1592_sv2v_reg  <= w_data_i[42];
      \nz.mem_1591_sv2v_reg  <= w_data_i[41];
      \nz.mem_1590_sv2v_reg  <= w_data_i[40];
      \nz.mem_1589_sv2v_reg  <= w_data_i[39];
      \nz.mem_1588_sv2v_reg  <= w_data_i[38];
      \nz.mem_1587_sv2v_reg  <= w_data_i[37];
      \nz.mem_1586_sv2v_reg  <= w_data_i[36];
      \nz.mem_1585_sv2v_reg  <= w_data_i[35];
      \nz.mem_1584_sv2v_reg  <= w_data_i[34];
      \nz.mem_1583_sv2v_reg  <= w_data_i[33];
      \nz.mem_1582_sv2v_reg  <= w_data_i[32];
      \nz.mem_1581_sv2v_reg  <= w_data_i[31];
      \nz.mem_1580_sv2v_reg  <= w_data_i[30];
      \nz.mem_1579_sv2v_reg  <= w_data_i[29];
      \nz.mem_1578_sv2v_reg  <= w_data_i[28];
      \nz.mem_1577_sv2v_reg  <= w_data_i[27];
      \nz.mem_1576_sv2v_reg  <= w_data_i[26];
      \nz.mem_1575_sv2v_reg  <= w_data_i[25];
      \nz.mem_1574_sv2v_reg  <= w_data_i[24];
      \nz.mem_1573_sv2v_reg  <= w_data_i[23];
      \nz.mem_1572_sv2v_reg  <= w_data_i[22];
      \nz.mem_1571_sv2v_reg  <= w_data_i[21];
      \nz.mem_1570_sv2v_reg  <= w_data_i[20];
      \nz.mem_1569_sv2v_reg  <= w_data_i[19];
      \nz.mem_1568_sv2v_reg  <= w_data_i[18];
      \nz.mem_1567_sv2v_reg  <= w_data_i[17];
      \nz.mem_1566_sv2v_reg  <= w_data_i[16];
      \nz.mem_1565_sv2v_reg  <= w_data_i[15];
      \nz.mem_1564_sv2v_reg  <= w_data_i[14];
      \nz.mem_1563_sv2v_reg  <= w_data_i[13];
      \nz.mem_1562_sv2v_reg  <= w_data_i[12];
      \nz.mem_1561_sv2v_reg  <= w_data_i[11];
      \nz.mem_1560_sv2v_reg  <= w_data_i[10];
      \nz.mem_1559_sv2v_reg  <= w_data_i[9];
      \nz.mem_1558_sv2v_reg  <= w_data_i[8];
      \nz.mem_1557_sv2v_reg  <= w_data_i[7];
      \nz.mem_1556_sv2v_reg  <= w_data_i[6];
      \nz.mem_1555_sv2v_reg  <= w_data_i[5];
      \nz.mem_1554_sv2v_reg  <= w_data_i[4];
      \nz.mem_1553_sv2v_reg  <= w_data_i[3];
      \nz.mem_1552_sv2v_reg  <= w_data_i[2];
      \nz.mem_1551_sv2v_reg  <= w_data_i[1];
      \nz.mem_1550_sv2v_reg  <= w_data_i[0];
    end 
    if(N235) begin
      \nz.mem_1549_sv2v_reg  <= w_data_i[49];
      \nz.mem_1548_sv2v_reg  <= w_data_i[48];
      \nz.mem_1547_sv2v_reg  <= w_data_i[47];
      \nz.mem_1546_sv2v_reg  <= w_data_i[46];
      \nz.mem_1545_sv2v_reg  <= w_data_i[45];
      \nz.mem_1544_sv2v_reg  <= w_data_i[44];
      \nz.mem_1543_sv2v_reg  <= w_data_i[43];
      \nz.mem_1542_sv2v_reg  <= w_data_i[42];
      \nz.mem_1541_sv2v_reg  <= w_data_i[41];
      \nz.mem_1540_sv2v_reg  <= w_data_i[40];
      \nz.mem_1539_sv2v_reg  <= w_data_i[39];
      \nz.mem_1538_sv2v_reg  <= w_data_i[38];
      \nz.mem_1537_sv2v_reg  <= w_data_i[37];
      \nz.mem_1536_sv2v_reg  <= w_data_i[36];
      \nz.mem_1535_sv2v_reg  <= w_data_i[35];
      \nz.mem_1534_sv2v_reg  <= w_data_i[34];
      \nz.mem_1533_sv2v_reg  <= w_data_i[33];
      \nz.mem_1532_sv2v_reg  <= w_data_i[32];
      \nz.mem_1531_sv2v_reg  <= w_data_i[31];
      \nz.mem_1530_sv2v_reg  <= w_data_i[30];
      \nz.mem_1529_sv2v_reg  <= w_data_i[29];
      \nz.mem_1528_sv2v_reg  <= w_data_i[28];
      \nz.mem_1527_sv2v_reg  <= w_data_i[27];
      \nz.mem_1526_sv2v_reg  <= w_data_i[26];
      \nz.mem_1525_sv2v_reg  <= w_data_i[25];
      \nz.mem_1524_sv2v_reg  <= w_data_i[24];
      \nz.mem_1523_sv2v_reg  <= w_data_i[23];
      \nz.mem_1522_sv2v_reg  <= w_data_i[22];
      \nz.mem_1521_sv2v_reg  <= w_data_i[21];
      \nz.mem_1520_sv2v_reg  <= w_data_i[20];
      \nz.mem_1519_sv2v_reg  <= w_data_i[19];
      \nz.mem_1518_sv2v_reg  <= w_data_i[18];
      \nz.mem_1517_sv2v_reg  <= w_data_i[17];
      \nz.mem_1516_sv2v_reg  <= w_data_i[16];
      \nz.mem_1515_sv2v_reg  <= w_data_i[15];
      \nz.mem_1514_sv2v_reg  <= w_data_i[14];
      \nz.mem_1513_sv2v_reg  <= w_data_i[13];
      \nz.mem_1512_sv2v_reg  <= w_data_i[12];
      \nz.mem_1511_sv2v_reg  <= w_data_i[11];
      \nz.mem_1510_sv2v_reg  <= w_data_i[10];
      \nz.mem_1509_sv2v_reg  <= w_data_i[9];
      \nz.mem_1508_sv2v_reg  <= w_data_i[8];
      \nz.mem_1507_sv2v_reg  <= w_data_i[7];
      \nz.mem_1506_sv2v_reg  <= w_data_i[6];
      \nz.mem_1505_sv2v_reg  <= w_data_i[5];
      \nz.mem_1504_sv2v_reg  <= w_data_i[4];
      \nz.mem_1503_sv2v_reg  <= w_data_i[3];
      \nz.mem_1502_sv2v_reg  <= w_data_i[2];
      \nz.mem_1501_sv2v_reg  <= w_data_i[1];
      \nz.mem_1500_sv2v_reg  <= w_data_i[0];
    end 
    if(N234) begin
      \nz.mem_1499_sv2v_reg  <= w_data_i[49];
      \nz.mem_1498_sv2v_reg  <= w_data_i[48];
      \nz.mem_1497_sv2v_reg  <= w_data_i[47];
      \nz.mem_1496_sv2v_reg  <= w_data_i[46];
      \nz.mem_1495_sv2v_reg  <= w_data_i[45];
      \nz.mem_1494_sv2v_reg  <= w_data_i[44];
      \nz.mem_1493_sv2v_reg  <= w_data_i[43];
      \nz.mem_1492_sv2v_reg  <= w_data_i[42];
      \nz.mem_1491_sv2v_reg  <= w_data_i[41];
      \nz.mem_1490_sv2v_reg  <= w_data_i[40];
      \nz.mem_1489_sv2v_reg  <= w_data_i[39];
      \nz.mem_1488_sv2v_reg  <= w_data_i[38];
      \nz.mem_1487_sv2v_reg  <= w_data_i[37];
      \nz.mem_1486_sv2v_reg  <= w_data_i[36];
      \nz.mem_1485_sv2v_reg  <= w_data_i[35];
      \nz.mem_1484_sv2v_reg  <= w_data_i[34];
      \nz.mem_1483_sv2v_reg  <= w_data_i[33];
      \nz.mem_1482_sv2v_reg  <= w_data_i[32];
      \nz.mem_1481_sv2v_reg  <= w_data_i[31];
      \nz.mem_1480_sv2v_reg  <= w_data_i[30];
      \nz.mem_1479_sv2v_reg  <= w_data_i[29];
      \nz.mem_1478_sv2v_reg  <= w_data_i[28];
      \nz.mem_1477_sv2v_reg  <= w_data_i[27];
      \nz.mem_1476_sv2v_reg  <= w_data_i[26];
      \nz.mem_1475_sv2v_reg  <= w_data_i[25];
      \nz.mem_1474_sv2v_reg  <= w_data_i[24];
      \nz.mem_1473_sv2v_reg  <= w_data_i[23];
      \nz.mem_1472_sv2v_reg  <= w_data_i[22];
      \nz.mem_1471_sv2v_reg  <= w_data_i[21];
      \nz.mem_1470_sv2v_reg  <= w_data_i[20];
      \nz.mem_1469_sv2v_reg  <= w_data_i[19];
      \nz.mem_1468_sv2v_reg  <= w_data_i[18];
      \nz.mem_1467_sv2v_reg  <= w_data_i[17];
      \nz.mem_1466_sv2v_reg  <= w_data_i[16];
      \nz.mem_1465_sv2v_reg  <= w_data_i[15];
      \nz.mem_1464_sv2v_reg  <= w_data_i[14];
      \nz.mem_1463_sv2v_reg  <= w_data_i[13];
      \nz.mem_1462_sv2v_reg  <= w_data_i[12];
      \nz.mem_1461_sv2v_reg  <= w_data_i[11];
      \nz.mem_1460_sv2v_reg  <= w_data_i[10];
      \nz.mem_1459_sv2v_reg  <= w_data_i[9];
      \nz.mem_1458_sv2v_reg  <= w_data_i[8];
      \nz.mem_1457_sv2v_reg  <= w_data_i[7];
      \nz.mem_1456_sv2v_reg  <= w_data_i[6];
      \nz.mem_1455_sv2v_reg  <= w_data_i[5];
      \nz.mem_1454_sv2v_reg  <= w_data_i[4];
      \nz.mem_1453_sv2v_reg  <= w_data_i[3];
      \nz.mem_1452_sv2v_reg  <= w_data_i[2];
      \nz.mem_1451_sv2v_reg  <= w_data_i[1];
      \nz.mem_1450_sv2v_reg  <= w_data_i[0];
    end 
    if(N233) begin
      \nz.mem_1449_sv2v_reg  <= w_data_i[49];
      \nz.mem_1448_sv2v_reg  <= w_data_i[48];
      \nz.mem_1447_sv2v_reg  <= w_data_i[47];
      \nz.mem_1446_sv2v_reg  <= w_data_i[46];
      \nz.mem_1445_sv2v_reg  <= w_data_i[45];
      \nz.mem_1444_sv2v_reg  <= w_data_i[44];
      \nz.mem_1443_sv2v_reg  <= w_data_i[43];
      \nz.mem_1442_sv2v_reg  <= w_data_i[42];
      \nz.mem_1441_sv2v_reg  <= w_data_i[41];
      \nz.mem_1440_sv2v_reg  <= w_data_i[40];
      \nz.mem_1439_sv2v_reg  <= w_data_i[39];
      \nz.mem_1438_sv2v_reg  <= w_data_i[38];
      \nz.mem_1437_sv2v_reg  <= w_data_i[37];
      \nz.mem_1436_sv2v_reg  <= w_data_i[36];
      \nz.mem_1435_sv2v_reg  <= w_data_i[35];
      \nz.mem_1434_sv2v_reg  <= w_data_i[34];
      \nz.mem_1433_sv2v_reg  <= w_data_i[33];
      \nz.mem_1432_sv2v_reg  <= w_data_i[32];
      \nz.mem_1431_sv2v_reg  <= w_data_i[31];
      \nz.mem_1430_sv2v_reg  <= w_data_i[30];
      \nz.mem_1429_sv2v_reg  <= w_data_i[29];
      \nz.mem_1428_sv2v_reg  <= w_data_i[28];
      \nz.mem_1427_sv2v_reg  <= w_data_i[27];
      \nz.mem_1426_sv2v_reg  <= w_data_i[26];
      \nz.mem_1425_sv2v_reg  <= w_data_i[25];
      \nz.mem_1424_sv2v_reg  <= w_data_i[24];
      \nz.mem_1423_sv2v_reg  <= w_data_i[23];
      \nz.mem_1422_sv2v_reg  <= w_data_i[22];
      \nz.mem_1421_sv2v_reg  <= w_data_i[21];
      \nz.mem_1420_sv2v_reg  <= w_data_i[20];
      \nz.mem_1419_sv2v_reg  <= w_data_i[19];
      \nz.mem_1418_sv2v_reg  <= w_data_i[18];
      \nz.mem_1417_sv2v_reg  <= w_data_i[17];
      \nz.mem_1416_sv2v_reg  <= w_data_i[16];
      \nz.mem_1415_sv2v_reg  <= w_data_i[15];
      \nz.mem_1414_sv2v_reg  <= w_data_i[14];
      \nz.mem_1413_sv2v_reg  <= w_data_i[13];
      \nz.mem_1412_sv2v_reg  <= w_data_i[12];
      \nz.mem_1411_sv2v_reg  <= w_data_i[11];
      \nz.mem_1410_sv2v_reg  <= w_data_i[10];
      \nz.mem_1409_sv2v_reg  <= w_data_i[9];
      \nz.mem_1408_sv2v_reg  <= w_data_i[8];
      \nz.mem_1407_sv2v_reg  <= w_data_i[7];
      \nz.mem_1406_sv2v_reg  <= w_data_i[6];
      \nz.mem_1405_sv2v_reg  <= w_data_i[5];
      \nz.mem_1404_sv2v_reg  <= w_data_i[4];
      \nz.mem_1403_sv2v_reg  <= w_data_i[3];
      \nz.mem_1402_sv2v_reg  <= w_data_i[2];
      \nz.mem_1401_sv2v_reg  <= w_data_i[1];
      \nz.mem_1400_sv2v_reg  <= w_data_i[0];
    end 
    if(N232) begin
      \nz.mem_1399_sv2v_reg  <= w_data_i[49];
      \nz.mem_1398_sv2v_reg  <= w_data_i[48];
      \nz.mem_1397_sv2v_reg  <= w_data_i[47];
      \nz.mem_1396_sv2v_reg  <= w_data_i[46];
      \nz.mem_1395_sv2v_reg  <= w_data_i[45];
      \nz.mem_1394_sv2v_reg  <= w_data_i[44];
      \nz.mem_1393_sv2v_reg  <= w_data_i[43];
      \nz.mem_1392_sv2v_reg  <= w_data_i[42];
      \nz.mem_1391_sv2v_reg  <= w_data_i[41];
      \nz.mem_1390_sv2v_reg  <= w_data_i[40];
      \nz.mem_1389_sv2v_reg  <= w_data_i[39];
      \nz.mem_1388_sv2v_reg  <= w_data_i[38];
      \nz.mem_1387_sv2v_reg  <= w_data_i[37];
      \nz.mem_1386_sv2v_reg  <= w_data_i[36];
      \nz.mem_1385_sv2v_reg  <= w_data_i[35];
      \nz.mem_1384_sv2v_reg  <= w_data_i[34];
      \nz.mem_1383_sv2v_reg  <= w_data_i[33];
      \nz.mem_1382_sv2v_reg  <= w_data_i[32];
      \nz.mem_1381_sv2v_reg  <= w_data_i[31];
      \nz.mem_1380_sv2v_reg  <= w_data_i[30];
      \nz.mem_1379_sv2v_reg  <= w_data_i[29];
      \nz.mem_1378_sv2v_reg  <= w_data_i[28];
      \nz.mem_1377_sv2v_reg  <= w_data_i[27];
      \nz.mem_1376_sv2v_reg  <= w_data_i[26];
      \nz.mem_1375_sv2v_reg  <= w_data_i[25];
      \nz.mem_1374_sv2v_reg  <= w_data_i[24];
      \nz.mem_1373_sv2v_reg  <= w_data_i[23];
      \nz.mem_1372_sv2v_reg  <= w_data_i[22];
      \nz.mem_1371_sv2v_reg  <= w_data_i[21];
      \nz.mem_1370_sv2v_reg  <= w_data_i[20];
      \nz.mem_1369_sv2v_reg  <= w_data_i[19];
      \nz.mem_1368_sv2v_reg  <= w_data_i[18];
      \nz.mem_1367_sv2v_reg  <= w_data_i[17];
      \nz.mem_1366_sv2v_reg  <= w_data_i[16];
      \nz.mem_1365_sv2v_reg  <= w_data_i[15];
      \nz.mem_1364_sv2v_reg  <= w_data_i[14];
      \nz.mem_1363_sv2v_reg  <= w_data_i[13];
      \nz.mem_1362_sv2v_reg  <= w_data_i[12];
      \nz.mem_1361_sv2v_reg  <= w_data_i[11];
      \nz.mem_1360_sv2v_reg  <= w_data_i[10];
      \nz.mem_1359_sv2v_reg  <= w_data_i[9];
      \nz.mem_1358_sv2v_reg  <= w_data_i[8];
      \nz.mem_1357_sv2v_reg  <= w_data_i[7];
      \nz.mem_1356_sv2v_reg  <= w_data_i[6];
      \nz.mem_1355_sv2v_reg  <= w_data_i[5];
      \nz.mem_1354_sv2v_reg  <= w_data_i[4];
      \nz.mem_1353_sv2v_reg  <= w_data_i[3];
      \nz.mem_1352_sv2v_reg  <= w_data_i[2];
      \nz.mem_1351_sv2v_reg  <= w_data_i[1];
      \nz.mem_1350_sv2v_reg  <= w_data_i[0];
    end 
    if(N231) begin
      \nz.mem_1349_sv2v_reg  <= w_data_i[49];
      \nz.mem_1348_sv2v_reg  <= w_data_i[48];
      \nz.mem_1347_sv2v_reg  <= w_data_i[47];
      \nz.mem_1346_sv2v_reg  <= w_data_i[46];
      \nz.mem_1345_sv2v_reg  <= w_data_i[45];
      \nz.mem_1344_sv2v_reg  <= w_data_i[44];
      \nz.mem_1343_sv2v_reg  <= w_data_i[43];
      \nz.mem_1342_sv2v_reg  <= w_data_i[42];
      \nz.mem_1341_sv2v_reg  <= w_data_i[41];
      \nz.mem_1340_sv2v_reg  <= w_data_i[40];
      \nz.mem_1339_sv2v_reg  <= w_data_i[39];
      \nz.mem_1338_sv2v_reg  <= w_data_i[38];
      \nz.mem_1337_sv2v_reg  <= w_data_i[37];
      \nz.mem_1336_sv2v_reg  <= w_data_i[36];
      \nz.mem_1335_sv2v_reg  <= w_data_i[35];
      \nz.mem_1334_sv2v_reg  <= w_data_i[34];
      \nz.mem_1333_sv2v_reg  <= w_data_i[33];
      \nz.mem_1332_sv2v_reg  <= w_data_i[32];
      \nz.mem_1331_sv2v_reg  <= w_data_i[31];
      \nz.mem_1330_sv2v_reg  <= w_data_i[30];
      \nz.mem_1329_sv2v_reg  <= w_data_i[29];
      \nz.mem_1328_sv2v_reg  <= w_data_i[28];
      \nz.mem_1327_sv2v_reg  <= w_data_i[27];
      \nz.mem_1326_sv2v_reg  <= w_data_i[26];
      \nz.mem_1325_sv2v_reg  <= w_data_i[25];
      \nz.mem_1324_sv2v_reg  <= w_data_i[24];
      \nz.mem_1323_sv2v_reg  <= w_data_i[23];
      \nz.mem_1322_sv2v_reg  <= w_data_i[22];
      \nz.mem_1321_sv2v_reg  <= w_data_i[21];
      \nz.mem_1320_sv2v_reg  <= w_data_i[20];
      \nz.mem_1319_sv2v_reg  <= w_data_i[19];
      \nz.mem_1318_sv2v_reg  <= w_data_i[18];
      \nz.mem_1317_sv2v_reg  <= w_data_i[17];
      \nz.mem_1316_sv2v_reg  <= w_data_i[16];
      \nz.mem_1315_sv2v_reg  <= w_data_i[15];
      \nz.mem_1314_sv2v_reg  <= w_data_i[14];
      \nz.mem_1313_sv2v_reg  <= w_data_i[13];
      \nz.mem_1312_sv2v_reg  <= w_data_i[12];
      \nz.mem_1311_sv2v_reg  <= w_data_i[11];
      \nz.mem_1310_sv2v_reg  <= w_data_i[10];
      \nz.mem_1309_sv2v_reg  <= w_data_i[9];
      \nz.mem_1308_sv2v_reg  <= w_data_i[8];
      \nz.mem_1307_sv2v_reg  <= w_data_i[7];
      \nz.mem_1306_sv2v_reg  <= w_data_i[6];
      \nz.mem_1305_sv2v_reg  <= w_data_i[5];
      \nz.mem_1304_sv2v_reg  <= w_data_i[4];
      \nz.mem_1303_sv2v_reg  <= w_data_i[3];
      \nz.mem_1302_sv2v_reg  <= w_data_i[2];
      \nz.mem_1301_sv2v_reg  <= w_data_i[1];
      \nz.mem_1300_sv2v_reg  <= w_data_i[0];
    end 
    if(N230) begin
      \nz.mem_1299_sv2v_reg  <= w_data_i[49];
      \nz.mem_1298_sv2v_reg  <= w_data_i[48];
      \nz.mem_1297_sv2v_reg  <= w_data_i[47];
      \nz.mem_1296_sv2v_reg  <= w_data_i[46];
      \nz.mem_1295_sv2v_reg  <= w_data_i[45];
      \nz.mem_1294_sv2v_reg  <= w_data_i[44];
      \nz.mem_1293_sv2v_reg  <= w_data_i[43];
      \nz.mem_1292_sv2v_reg  <= w_data_i[42];
      \nz.mem_1291_sv2v_reg  <= w_data_i[41];
      \nz.mem_1290_sv2v_reg  <= w_data_i[40];
      \nz.mem_1289_sv2v_reg  <= w_data_i[39];
      \nz.mem_1288_sv2v_reg  <= w_data_i[38];
      \nz.mem_1287_sv2v_reg  <= w_data_i[37];
      \nz.mem_1286_sv2v_reg  <= w_data_i[36];
      \nz.mem_1285_sv2v_reg  <= w_data_i[35];
      \nz.mem_1284_sv2v_reg  <= w_data_i[34];
      \nz.mem_1283_sv2v_reg  <= w_data_i[33];
      \nz.mem_1282_sv2v_reg  <= w_data_i[32];
      \nz.mem_1281_sv2v_reg  <= w_data_i[31];
      \nz.mem_1280_sv2v_reg  <= w_data_i[30];
      \nz.mem_1279_sv2v_reg  <= w_data_i[29];
      \nz.mem_1278_sv2v_reg  <= w_data_i[28];
      \nz.mem_1277_sv2v_reg  <= w_data_i[27];
      \nz.mem_1276_sv2v_reg  <= w_data_i[26];
      \nz.mem_1275_sv2v_reg  <= w_data_i[25];
      \nz.mem_1274_sv2v_reg  <= w_data_i[24];
      \nz.mem_1273_sv2v_reg  <= w_data_i[23];
      \nz.mem_1272_sv2v_reg  <= w_data_i[22];
      \nz.mem_1271_sv2v_reg  <= w_data_i[21];
      \nz.mem_1270_sv2v_reg  <= w_data_i[20];
      \nz.mem_1269_sv2v_reg  <= w_data_i[19];
      \nz.mem_1268_sv2v_reg  <= w_data_i[18];
      \nz.mem_1267_sv2v_reg  <= w_data_i[17];
      \nz.mem_1266_sv2v_reg  <= w_data_i[16];
      \nz.mem_1265_sv2v_reg  <= w_data_i[15];
      \nz.mem_1264_sv2v_reg  <= w_data_i[14];
      \nz.mem_1263_sv2v_reg  <= w_data_i[13];
      \nz.mem_1262_sv2v_reg  <= w_data_i[12];
      \nz.mem_1261_sv2v_reg  <= w_data_i[11];
      \nz.mem_1260_sv2v_reg  <= w_data_i[10];
      \nz.mem_1259_sv2v_reg  <= w_data_i[9];
      \nz.mem_1258_sv2v_reg  <= w_data_i[8];
      \nz.mem_1257_sv2v_reg  <= w_data_i[7];
      \nz.mem_1256_sv2v_reg  <= w_data_i[6];
      \nz.mem_1255_sv2v_reg  <= w_data_i[5];
      \nz.mem_1254_sv2v_reg  <= w_data_i[4];
      \nz.mem_1253_sv2v_reg  <= w_data_i[3];
      \nz.mem_1252_sv2v_reg  <= w_data_i[2];
      \nz.mem_1251_sv2v_reg  <= w_data_i[1];
      \nz.mem_1250_sv2v_reg  <= w_data_i[0];
    end 
    if(N229) begin
      \nz.mem_1249_sv2v_reg  <= w_data_i[49];
      \nz.mem_1248_sv2v_reg  <= w_data_i[48];
      \nz.mem_1247_sv2v_reg  <= w_data_i[47];
      \nz.mem_1246_sv2v_reg  <= w_data_i[46];
      \nz.mem_1245_sv2v_reg  <= w_data_i[45];
      \nz.mem_1244_sv2v_reg  <= w_data_i[44];
      \nz.mem_1243_sv2v_reg  <= w_data_i[43];
      \nz.mem_1242_sv2v_reg  <= w_data_i[42];
      \nz.mem_1241_sv2v_reg  <= w_data_i[41];
      \nz.mem_1240_sv2v_reg  <= w_data_i[40];
      \nz.mem_1239_sv2v_reg  <= w_data_i[39];
      \nz.mem_1238_sv2v_reg  <= w_data_i[38];
      \nz.mem_1237_sv2v_reg  <= w_data_i[37];
      \nz.mem_1236_sv2v_reg  <= w_data_i[36];
      \nz.mem_1235_sv2v_reg  <= w_data_i[35];
      \nz.mem_1234_sv2v_reg  <= w_data_i[34];
      \nz.mem_1233_sv2v_reg  <= w_data_i[33];
      \nz.mem_1232_sv2v_reg  <= w_data_i[32];
      \nz.mem_1231_sv2v_reg  <= w_data_i[31];
      \nz.mem_1230_sv2v_reg  <= w_data_i[30];
      \nz.mem_1229_sv2v_reg  <= w_data_i[29];
      \nz.mem_1228_sv2v_reg  <= w_data_i[28];
      \nz.mem_1227_sv2v_reg  <= w_data_i[27];
      \nz.mem_1226_sv2v_reg  <= w_data_i[26];
      \nz.mem_1225_sv2v_reg  <= w_data_i[25];
      \nz.mem_1224_sv2v_reg  <= w_data_i[24];
      \nz.mem_1223_sv2v_reg  <= w_data_i[23];
      \nz.mem_1222_sv2v_reg  <= w_data_i[22];
      \nz.mem_1221_sv2v_reg  <= w_data_i[21];
      \nz.mem_1220_sv2v_reg  <= w_data_i[20];
      \nz.mem_1219_sv2v_reg  <= w_data_i[19];
      \nz.mem_1218_sv2v_reg  <= w_data_i[18];
      \nz.mem_1217_sv2v_reg  <= w_data_i[17];
      \nz.mem_1216_sv2v_reg  <= w_data_i[16];
      \nz.mem_1215_sv2v_reg  <= w_data_i[15];
      \nz.mem_1214_sv2v_reg  <= w_data_i[14];
      \nz.mem_1213_sv2v_reg  <= w_data_i[13];
      \nz.mem_1212_sv2v_reg  <= w_data_i[12];
      \nz.mem_1211_sv2v_reg  <= w_data_i[11];
      \nz.mem_1210_sv2v_reg  <= w_data_i[10];
      \nz.mem_1209_sv2v_reg  <= w_data_i[9];
      \nz.mem_1208_sv2v_reg  <= w_data_i[8];
      \nz.mem_1207_sv2v_reg  <= w_data_i[7];
      \nz.mem_1206_sv2v_reg  <= w_data_i[6];
      \nz.mem_1205_sv2v_reg  <= w_data_i[5];
      \nz.mem_1204_sv2v_reg  <= w_data_i[4];
      \nz.mem_1203_sv2v_reg  <= w_data_i[3];
      \nz.mem_1202_sv2v_reg  <= w_data_i[2];
      \nz.mem_1201_sv2v_reg  <= w_data_i[1];
      \nz.mem_1200_sv2v_reg  <= w_data_i[0];
    end 
    if(N228) begin
      \nz.mem_1199_sv2v_reg  <= w_data_i[49];
      \nz.mem_1198_sv2v_reg  <= w_data_i[48];
      \nz.mem_1197_sv2v_reg  <= w_data_i[47];
      \nz.mem_1196_sv2v_reg  <= w_data_i[46];
      \nz.mem_1195_sv2v_reg  <= w_data_i[45];
      \nz.mem_1194_sv2v_reg  <= w_data_i[44];
      \nz.mem_1193_sv2v_reg  <= w_data_i[43];
      \nz.mem_1192_sv2v_reg  <= w_data_i[42];
      \nz.mem_1191_sv2v_reg  <= w_data_i[41];
      \nz.mem_1190_sv2v_reg  <= w_data_i[40];
      \nz.mem_1189_sv2v_reg  <= w_data_i[39];
      \nz.mem_1188_sv2v_reg  <= w_data_i[38];
      \nz.mem_1187_sv2v_reg  <= w_data_i[37];
      \nz.mem_1186_sv2v_reg  <= w_data_i[36];
      \nz.mem_1185_sv2v_reg  <= w_data_i[35];
      \nz.mem_1184_sv2v_reg  <= w_data_i[34];
      \nz.mem_1183_sv2v_reg  <= w_data_i[33];
      \nz.mem_1182_sv2v_reg  <= w_data_i[32];
      \nz.mem_1181_sv2v_reg  <= w_data_i[31];
      \nz.mem_1180_sv2v_reg  <= w_data_i[30];
      \nz.mem_1179_sv2v_reg  <= w_data_i[29];
      \nz.mem_1178_sv2v_reg  <= w_data_i[28];
      \nz.mem_1177_sv2v_reg  <= w_data_i[27];
      \nz.mem_1176_sv2v_reg  <= w_data_i[26];
      \nz.mem_1175_sv2v_reg  <= w_data_i[25];
      \nz.mem_1174_sv2v_reg  <= w_data_i[24];
      \nz.mem_1173_sv2v_reg  <= w_data_i[23];
      \nz.mem_1172_sv2v_reg  <= w_data_i[22];
      \nz.mem_1171_sv2v_reg  <= w_data_i[21];
      \nz.mem_1170_sv2v_reg  <= w_data_i[20];
      \nz.mem_1169_sv2v_reg  <= w_data_i[19];
      \nz.mem_1168_sv2v_reg  <= w_data_i[18];
      \nz.mem_1167_sv2v_reg  <= w_data_i[17];
      \nz.mem_1166_sv2v_reg  <= w_data_i[16];
      \nz.mem_1165_sv2v_reg  <= w_data_i[15];
      \nz.mem_1164_sv2v_reg  <= w_data_i[14];
      \nz.mem_1163_sv2v_reg  <= w_data_i[13];
      \nz.mem_1162_sv2v_reg  <= w_data_i[12];
      \nz.mem_1161_sv2v_reg  <= w_data_i[11];
      \nz.mem_1160_sv2v_reg  <= w_data_i[10];
      \nz.mem_1159_sv2v_reg  <= w_data_i[9];
      \nz.mem_1158_sv2v_reg  <= w_data_i[8];
      \nz.mem_1157_sv2v_reg  <= w_data_i[7];
      \nz.mem_1156_sv2v_reg  <= w_data_i[6];
      \nz.mem_1155_sv2v_reg  <= w_data_i[5];
      \nz.mem_1154_sv2v_reg  <= w_data_i[4];
      \nz.mem_1153_sv2v_reg  <= w_data_i[3];
      \nz.mem_1152_sv2v_reg  <= w_data_i[2];
      \nz.mem_1151_sv2v_reg  <= w_data_i[1];
      \nz.mem_1150_sv2v_reg  <= w_data_i[0];
    end 
    if(N227) begin
      \nz.mem_1149_sv2v_reg  <= w_data_i[49];
      \nz.mem_1148_sv2v_reg  <= w_data_i[48];
      \nz.mem_1147_sv2v_reg  <= w_data_i[47];
      \nz.mem_1146_sv2v_reg  <= w_data_i[46];
      \nz.mem_1145_sv2v_reg  <= w_data_i[45];
      \nz.mem_1144_sv2v_reg  <= w_data_i[44];
      \nz.mem_1143_sv2v_reg  <= w_data_i[43];
      \nz.mem_1142_sv2v_reg  <= w_data_i[42];
      \nz.mem_1141_sv2v_reg  <= w_data_i[41];
      \nz.mem_1140_sv2v_reg  <= w_data_i[40];
      \nz.mem_1139_sv2v_reg  <= w_data_i[39];
      \nz.mem_1138_sv2v_reg  <= w_data_i[38];
      \nz.mem_1137_sv2v_reg  <= w_data_i[37];
      \nz.mem_1136_sv2v_reg  <= w_data_i[36];
      \nz.mem_1135_sv2v_reg  <= w_data_i[35];
      \nz.mem_1134_sv2v_reg  <= w_data_i[34];
      \nz.mem_1133_sv2v_reg  <= w_data_i[33];
      \nz.mem_1132_sv2v_reg  <= w_data_i[32];
      \nz.mem_1131_sv2v_reg  <= w_data_i[31];
      \nz.mem_1130_sv2v_reg  <= w_data_i[30];
      \nz.mem_1129_sv2v_reg  <= w_data_i[29];
      \nz.mem_1128_sv2v_reg  <= w_data_i[28];
      \nz.mem_1127_sv2v_reg  <= w_data_i[27];
      \nz.mem_1126_sv2v_reg  <= w_data_i[26];
      \nz.mem_1125_sv2v_reg  <= w_data_i[25];
      \nz.mem_1124_sv2v_reg  <= w_data_i[24];
      \nz.mem_1123_sv2v_reg  <= w_data_i[23];
      \nz.mem_1122_sv2v_reg  <= w_data_i[22];
      \nz.mem_1121_sv2v_reg  <= w_data_i[21];
      \nz.mem_1120_sv2v_reg  <= w_data_i[20];
      \nz.mem_1119_sv2v_reg  <= w_data_i[19];
      \nz.mem_1118_sv2v_reg  <= w_data_i[18];
      \nz.mem_1117_sv2v_reg  <= w_data_i[17];
      \nz.mem_1116_sv2v_reg  <= w_data_i[16];
      \nz.mem_1115_sv2v_reg  <= w_data_i[15];
      \nz.mem_1114_sv2v_reg  <= w_data_i[14];
      \nz.mem_1113_sv2v_reg  <= w_data_i[13];
      \nz.mem_1112_sv2v_reg  <= w_data_i[12];
      \nz.mem_1111_sv2v_reg  <= w_data_i[11];
      \nz.mem_1110_sv2v_reg  <= w_data_i[10];
      \nz.mem_1109_sv2v_reg  <= w_data_i[9];
      \nz.mem_1108_sv2v_reg  <= w_data_i[8];
      \nz.mem_1107_sv2v_reg  <= w_data_i[7];
      \nz.mem_1106_sv2v_reg  <= w_data_i[6];
      \nz.mem_1105_sv2v_reg  <= w_data_i[5];
      \nz.mem_1104_sv2v_reg  <= w_data_i[4];
      \nz.mem_1103_sv2v_reg  <= w_data_i[3];
      \nz.mem_1102_sv2v_reg  <= w_data_i[2];
      \nz.mem_1101_sv2v_reg  <= w_data_i[1];
      \nz.mem_1100_sv2v_reg  <= w_data_i[0];
    end 
    if(N226) begin
      \nz.mem_1099_sv2v_reg  <= w_data_i[49];
      \nz.mem_1098_sv2v_reg  <= w_data_i[48];
      \nz.mem_1097_sv2v_reg  <= w_data_i[47];
      \nz.mem_1096_sv2v_reg  <= w_data_i[46];
      \nz.mem_1095_sv2v_reg  <= w_data_i[45];
      \nz.mem_1094_sv2v_reg  <= w_data_i[44];
      \nz.mem_1093_sv2v_reg  <= w_data_i[43];
      \nz.mem_1092_sv2v_reg  <= w_data_i[42];
      \nz.mem_1091_sv2v_reg  <= w_data_i[41];
      \nz.mem_1090_sv2v_reg  <= w_data_i[40];
      \nz.mem_1089_sv2v_reg  <= w_data_i[39];
      \nz.mem_1088_sv2v_reg  <= w_data_i[38];
      \nz.mem_1087_sv2v_reg  <= w_data_i[37];
      \nz.mem_1086_sv2v_reg  <= w_data_i[36];
      \nz.mem_1085_sv2v_reg  <= w_data_i[35];
      \nz.mem_1084_sv2v_reg  <= w_data_i[34];
      \nz.mem_1083_sv2v_reg  <= w_data_i[33];
      \nz.mem_1082_sv2v_reg  <= w_data_i[32];
      \nz.mem_1081_sv2v_reg  <= w_data_i[31];
      \nz.mem_1080_sv2v_reg  <= w_data_i[30];
      \nz.mem_1079_sv2v_reg  <= w_data_i[29];
      \nz.mem_1078_sv2v_reg  <= w_data_i[28];
      \nz.mem_1077_sv2v_reg  <= w_data_i[27];
      \nz.mem_1076_sv2v_reg  <= w_data_i[26];
      \nz.mem_1075_sv2v_reg  <= w_data_i[25];
      \nz.mem_1074_sv2v_reg  <= w_data_i[24];
      \nz.mem_1073_sv2v_reg  <= w_data_i[23];
      \nz.mem_1072_sv2v_reg  <= w_data_i[22];
      \nz.mem_1071_sv2v_reg  <= w_data_i[21];
      \nz.mem_1070_sv2v_reg  <= w_data_i[20];
      \nz.mem_1069_sv2v_reg  <= w_data_i[19];
      \nz.mem_1068_sv2v_reg  <= w_data_i[18];
      \nz.mem_1067_sv2v_reg  <= w_data_i[17];
      \nz.mem_1066_sv2v_reg  <= w_data_i[16];
      \nz.mem_1065_sv2v_reg  <= w_data_i[15];
      \nz.mem_1064_sv2v_reg  <= w_data_i[14];
      \nz.mem_1063_sv2v_reg  <= w_data_i[13];
      \nz.mem_1062_sv2v_reg  <= w_data_i[12];
      \nz.mem_1061_sv2v_reg  <= w_data_i[11];
      \nz.mem_1060_sv2v_reg  <= w_data_i[10];
      \nz.mem_1059_sv2v_reg  <= w_data_i[9];
      \nz.mem_1058_sv2v_reg  <= w_data_i[8];
      \nz.mem_1057_sv2v_reg  <= w_data_i[7];
      \nz.mem_1056_sv2v_reg  <= w_data_i[6];
      \nz.mem_1055_sv2v_reg  <= w_data_i[5];
      \nz.mem_1054_sv2v_reg  <= w_data_i[4];
      \nz.mem_1053_sv2v_reg  <= w_data_i[3];
      \nz.mem_1052_sv2v_reg  <= w_data_i[2];
      \nz.mem_1051_sv2v_reg  <= w_data_i[1];
      \nz.mem_1050_sv2v_reg  <= w_data_i[0];
    end 
    if(N225) begin
      \nz.mem_1049_sv2v_reg  <= w_data_i[49];
      \nz.mem_1048_sv2v_reg  <= w_data_i[48];
      \nz.mem_1047_sv2v_reg  <= w_data_i[47];
      \nz.mem_1046_sv2v_reg  <= w_data_i[46];
      \nz.mem_1045_sv2v_reg  <= w_data_i[45];
      \nz.mem_1044_sv2v_reg  <= w_data_i[44];
      \nz.mem_1043_sv2v_reg  <= w_data_i[43];
      \nz.mem_1042_sv2v_reg  <= w_data_i[42];
      \nz.mem_1041_sv2v_reg  <= w_data_i[41];
      \nz.mem_1040_sv2v_reg  <= w_data_i[40];
      \nz.mem_1039_sv2v_reg  <= w_data_i[39];
      \nz.mem_1038_sv2v_reg  <= w_data_i[38];
      \nz.mem_1037_sv2v_reg  <= w_data_i[37];
      \nz.mem_1036_sv2v_reg  <= w_data_i[36];
      \nz.mem_1035_sv2v_reg  <= w_data_i[35];
      \nz.mem_1034_sv2v_reg  <= w_data_i[34];
      \nz.mem_1033_sv2v_reg  <= w_data_i[33];
      \nz.mem_1032_sv2v_reg  <= w_data_i[32];
      \nz.mem_1031_sv2v_reg  <= w_data_i[31];
      \nz.mem_1030_sv2v_reg  <= w_data_i[30];
      \nz.mem_1029_sv2v_reg  <= w_data_i[29];
      \nz.mem_1028_sv2v_reg  <= w_data_i[28];
      \nz.mem_1027_sv2v_reg  <= w_data_i[27];
      \nz.mem_1026_sv2v_reg  <= w_data_i[26];
      \nz.mem_1025_sv2v_reg  <= w_data_i[25];
      \nz.mem_1024_sv2v_reg  <= w_data_i[24];
      \nz.mem_1023_sv2v_reg  <= w_data_i[23];
      \nz.mem_1022_sv2v_reg  <= w_data_i[22];
      \nz.mem_1021_sv2v_reg  <= w_data_i[21];
      \nz.mem_1020_sv2v_reg  <= w_data_i[20];
      \nz.mem_1019_sv2v_reg  <= w_data_i[19];
      \nz.mem_1018_sv2v_reg  <= w_data_i[18];
      \nz.mem_1017_sv2v_reg  <= w_data_i[17];
      \nz.mem_1016_sv2v_reg  <= w_data_i[16];
      \nz.mem_1015_sv2v_reg  <= w_data_i[15];
      \nz.mem_1014_sv2v_reg  <= w_data_i[14];
      \nz.mem_1013_sv2v_reg  <= w_data_i[13];
      \nz.mem_1012_sv2v_reg  <= w_data_i[12];
      \nz.mem_1011_sv2v_reg  <= w_data_i[11];
      \nz.mem_1010_sv2v_reg  <= w_data_i[10];
      \nz.mem_1009_sv2v_reg  <= w_data_i[9];
      \nz.mem_1008_sv2v_reg  <= w_data_i[8];
      \nz.mem_1007_sv2v_reg  <= w_data_i[7];
      \nz.mem_1006_sv2v_reg  <= w_data_i[6];
      \nz.mem_1005_sv2v_reg  <= w_data_i[5];
      \nz.mem_1004_sv2v_reg  <= w_data_i[4];
      \nz.mem_1003_sv2v_reg  <= w_data_i[3];
      \nz.mem_1002_sv2v_reg  <= w_data_i[2];
      \nz.mem_1001_sv2v_reg  <= w_data_i[1];
      \nz.mem_1000_sv2v_reg  <= w_data_i[0];
    end 
    if(N224) begin
      \nz.mem_999_sv2v_reg  <= w_data_i[49];
      \nz.mem_998_sv2v_reg  <= w_data_i[48];
      \nz.mem_997_sv2v_reg  <= w_data_i[47];
      \nz.mem_996_sv2v_reg  <= w_data_i[46];
      \nz.mem_995_sv2v_reg  <= w_data_i[45];
      \nz.mem_994_sv2v_reg  <= w_data_i[44];
      \nz.mem_993_sv2v_reg  <= w_data_i[43];
      \nz.mem_992_sv2v_reg  <= w_data_i[42];
      \nz.mem_991_sv2v_reg  <= w_data_i[41];
      \nz.mem_990_sv2v_reg  <= w_data_i[40];
      \nz.mem_989_sv2v_reg  <= w_data_i[39];
      \nz.mem_988_sv2v_reg  <= w_data_i[38];
      \nz.mem_987_sv2v_reg  <= w_data_i[37];
      \nz.mem_986_sv2v_reg  <= w_data_i[36];
      \nz.mem_985_sv2v_reg  <= w_data_i[35];
      \nz.mem_984_sv2v_reg  <= w_data_i[34];
      \nz.mem_983_sv2v_reg  <= w_data_i[33];
      \nz.mem_982_sv2v_reg  <= w_data_i[32];
      \nz.mem_981_sv2v_reg  <= w_data_i[31];
      \nz.mem_980_sv2v_reg  <= w_data_i[30];
      \nz.mem_979_sv2v_reg  <= w_data_i[29];
      \nz.mem_978_sv2v_reg  <= w_data_i[28];
      \nz.mem_977_sv2v_reg  <= w_data_i[27];
      \nz.mem_976_sv2v_reg  <= w_data_i[26];
      \nz.mem_975_sv2v_reg  <= w_data_i[25];
      \nz.mem_974_sv2v_reg  <= w_data_i[24];
      \nz.mem_973_sv2v_reg  <= w_data_i[23];
      \nz.mem_972_sv2v_reg  <= w_data_i[22];
      \nz.mem_971_sv2v_reg  <= w_data_i[21];
      \nz.mem_970_sv2v_reg  <= w_data_i[20];
      \nz.mem_969_sv2v_reg  <= w_data_i[19];
      \nz.mem_968_sv2v_reg  <= w_data_i[18];
      \nz.mem_967_sv2v_reg  <= w_data_i[17];
      \nz.mem_966_sv2v_reg  <= w_data_i[16];
      \nz.mem_965_sv2v_reg  <= w_data_i[15];
      \nz.mem_964_sv2v_reg  <= w_data_i[14];
      \nz.mem_963_sv2v_reg  <= w_data_i[13];
      \nz.mem_962_sv2v_reg  <= w_data_i[12];
      \nz.mem_961_sv2v_reg  <= w_data_i[11];
      \nz.mem_960_sv2v_reg  <= w_data_i[10];
      \nz.mem_959_sv2v_reg  <= w_data_i[9];
      \nz.mem_958_sv2v_reg  <= w_data_i[8];
      \nz.mem_957_sv2v_reg  <= w_data_i[7];
      \nz.mem_956_sv2v_reg  <= w_data_i[6];
      \nz.mem_955_sv2v_reg  <= w_data_i[5];
      \nz.mem_954_sv2v_reg  <= w_data_i[4];
      \nz.mem_953_sv2v_reg  <= w_data_i[3];
      \nz.mem_952_sv2v_reg  <= w_data_i[2];
      \nz.mem_951_sv2v_reg  <= w_data_i[1];
      \nz.mem_950_sv2v_reg  <= w_data_i[0];
    end 
    if(N223) begin
      \nz.mem_949_sv2v_reg  <= w_data_i[49];
      \nz.mem_948_sv2v_reg  <= w_data_i[48];
      \nz.mem_947_sv2v_reg  <= w_data_i[47];
      \nz.mem_946_sv2v_reg  <= w_data_i[46];
      \nz.mem_945_sv2v_reg  <= w_data_i[45];
      \nz.mem_944_sv2v_reg  <= w_data_i[44];
      \nz.mem_943_sv2v_reg  <= w_data_i[43];
      \nz.mem_942_sv2v_reg  <= w_data_i[42];
      \nz.mem_941_sv2v_reg  <= w_data_i[41];
      \nz.mem_940_sv2v_reg  <= w_data_i[40];
      \nz.mem_939_sv2v_reg  <= w_data_i[39];
      \nz.mem_938_sv2v_reg  <= w_data_i[38];
      \nz.mem_937_sv2v_reg  <= w_data_i[37];
      \nz.mem_936_sv2v_reg  <= w_data_i[36];
      \nz.mem_935_sv2v_reg  <= w_data_i[35];
      \nz.mem_934_sv2v_reg  <= w_data_i[34];
      \nz.mem_933_sv2v_reg  <= w_data_i[33];
      \nz.mem_932_sv2v_reg  <= w_data_i[32];
      \nz.mem_931_sv2v_reg  <= w_data_i[31];
      \nz.mem_930_sv2v_reg  <= w_data_i[30];
      \nz.mem_929_sv2v_reg  <= w_data_i[29];
      \nz.mem_928_sv2v_reg  <= w_data_i[28];
      \nz.mem_927_sv2v_reg  <= w_data_i[27];
      \nz.mem_926_sv2v_reg  <= w_data_i[26];
      \nz.mem_925_sv2v_reg  <= w_data_i[25];
      \nz.mem_924_sv2v_reg  <= w_data_i[24];
      \nz.mem_923_sv2v_reg  <= w_data_i[23];
      \nz.mem_922_sv2v_reg  <= w_data_i[22];
      \nz.mem_921_sv2v_reg  <= w_data_i[21];
      \nz.mem_920_sv2v_reg  <= w_data_i[20];
      \nz.mem_919_sv2v_reg  <= w_data_i[19];
      \nz.mem_918_sv2v_reg  <= w_data_i[18];
      \nz.mem_917_sv2v_reg  <= w_data_i[17];
      \nz.mem_916_sv2v_reg  <= w_data_i[16];
      \nz.mem_915_sv2v_reg  <= w_data_i[15];
      \nz.mem_914_sv2v_reg  <= w_data_i[14];
      \nz.mem_913_sv2v_reg  <= w_data_i[13];
      \nz.mem_912_sv2v_reg  <= w_data_i[12];
      \nz.mem_911_sv2v_reg  <= w_data_i[11];
      \nz.mem_910_sv2v_reg  <= w_data_i[10];
      \nz.mem_909_sv2v_reg  <= w_data_i[9];
      \nz.mem_908_sv2v_reg  <= w_data_i[8];
      \nz.mem_907_sv2v_reg  <= w_data_i[7];
      \nz.mem_906_sv2v_reg  <= w_data_i[6];
      \nz.mem_905_sv2v_reg  <= w_data_i[5];
      \nz.mem_904_sv2v_reg  <= w_data_i[4];
      \nz.mem_903_sv2v_reg  <= w_data_i[3];
      \nz.mem_902_sv2v_reg  <= w_data_i[2];
      \nz.mem_901_sv2v_reg  <= w_data_i[1];
      \nz.mem_900_sv2v_reg  <= w_data_i[0];
    end 
    if(N222) begin
      \nz.mem_899_sv2v_reg  <= w_data_i[49];
      \nz.mem_898_sv2v_reg  <= w_data_i[48];
      \nz.mem_897_sv2v_reg  <= w_data_i[47];
      \nz.mem_896_sv2v_reg  <= w_data_i[46];
      \nz.mem_895_sv2v_reg  <= w_data_i[45];
      \nz.mem_894_sv2v_reg  <= w_data_i[44];
      \nz.mem_893_sv2v_reg  <= w_data_i[43];
      \nz.mem_892_sv2v_reg  <= w_data_i[42];
      \nz.mem_891_sv2v_reg  <= w_data_i[41];
      \nz.mem_890_sv2v_reg  <= w_data_i[40];
      \nz.mem_889_sv2v_reg  <= w_data_i[39];
      \nz.mem_888_sv2v_reg  <= w_data_i[38];
      \nz.mem_887_sv2v_reg  <= w_data_i[37];
      \nz.mem_886_sv2v_reg  <= w_data_i[36];
      \nz.mem_885_sv2v_reg  <= w_data_i[35];
      \nz.mem_884_sv2v_reg  <= w_data_i[34];
      \nz.mem_883_sv2v_reg  <= w_data_i[33];
      \nz.mem_882_sv2v_reg  <= w_data_i[32];
      \nz.mem_881_sv2v_reg  <= w_data_i[31];
      \nz.mem_880_sv2v_reg  <= w_data_i[30];
      \nz.mem_879_sv2v_reg  <= w_data_i[29];
      \nz.mem_878_sv2v_reg  <= w_data_i[28];
      \nz.mem_877_sv2v_reg  <= w_data_i[27];
      \nz.mem_876_sv2v_reg  <= w_data_i[26];
      \nz.mem_875_sv2v_reg  <= w_data_i[25];
      \nz.mem_874_sv2v_reg  <= w_data_i[24];
      \nz.mem_873_sv2v_reg  <= w_data_i[23];
      \nz.mem_872_sv2v_reg  <= w_data_i[22];
      \nz.mem_871_sv2v_reg  <= w_data_i[21];
      \nz.mem_870_sv2v_reg  <= w_data_i[20];
      \nz.mem_869_sv2v_reg  <= w_data_i[19];
      \nz.mem_868_sv2v_reg  <= w_data_i[18];
      \nz.mem_867_sv2v_reg  <= w_data_i[17];
      \nz.mem_866_sv2v_reg  <= w_data_i[16];
      \nz.mem_865_sv2v_reg  <= w_data_i[15];
      \nz.mem_864_sv2v_reg  <= w_data_i[14];
      \nz.mem_863_sv2v_reg  <= w_data_i[13];
      \nz.mem_862_sv2v_reg  <= w_data_i[12];
      \nz.mem_861_sv2v_reg  <= w_data_i[11];
      \nz.mem_860_sv2v_reg  <= w_data_i[10];
      \nz.mem_859_sv2v_reg  <= w_data_i[9];
      \nz.mem_858_sv2v_reg  <= w_data_i[8];
      \nz.mem_857_sv2v_reg  <= w_data_i[7];
      \nz.mem_856_sv2v_reg  <= w_data_i[6];
      \nz.mem_855_sv2v_reg  <= w_data_i[5];
      \nz.mem_854_sv2v_reg  <= w_data_i[4];
      \nz.mem_853_sv2v_reg  <= w_data_i[3];
      \nz.mem_852_sv2v_reg  <= w_data_i[2];
      \nz.mem_851_sv2v_reg  <= w_data_i[1];
      \nz.mem_850_sv2v_reg  <= w_data_i[0];
    end 
    if(N221) begin
      \nz.mem_849_sv2v_reg  <= w_data_i[49];
      \nz.mem_848_sv2v_reg  <= w_data_i[48];
      \nz.mem_847_sv2v_reg  <= w_data_i[47];
      \nz.mem_846_sv2v_reg  <= w_data_i[46];
      \nz.mem_845_sv2v_reg  <= w_data_i[45];
      \nz.mem_844_sv2v_reg  <= w_data_i[44];
      \nz.mem_843_sv2v_reg  <= w_data_i[43];
      \nz.mem_842_sv2v_reg  <= w_data_i[42];
      \nz.mem_841_sv2v_reg  <= w_data_i[41];
      \nz.mem_840_sv2v_reg  <= w_data_i[40];
      \nz.mem_839_sv2v_reg  <= w_data_i[39];
      \nz.mem_838_sv2v_reg  <= w_data_i[38];
      \nz.mem_837_sv2v_reg  <= w_data_i[37];
      \nz.mem_836_sv2v_reg  <= w_data_i[36];
      \nz.mem_835_sv2v_reg  <= w_data_i[35];
      \nz.mem_834_sv2v_reg  <= w_data_i[34];
      \nz.mem_833_sv2v_reg  <= w_data_i[33];
      \nz.mem_832_sv2v_reg  <= w_data_i[32];
      \nz.mem_831_sv2v_reg  <= w_data_i[31];
      \nz.mem_830_sv2v_reg  <= w_data_i[30];
      \nz.mem_829_sv2v_reg  <= w_data_i[29];
      \nz.mem_828_sv2v_reg  <= w_data_i[28];
      \nz.mem_827_sv2v_reg  <= w_data_i[27];
      \nz.mem_826_sv2v_reg  <= w_data_i[26];
      \nz.mem_825_sv2v_reg  <= w_data_i[25];
      \nz.mem_824_sv2v_reg  <= w_data_i[24];
      \nz.mem_823_sv2v_reg  <= w_data_i[23];
      \nz.mem_822_sv2v_reg  <= w_data_i[22];
      \nz.mem_821_sv2v_reg  <= w_data_i[21];
      \nz.mem_820_sv2v_reg  <= w_data_i[20];
      \nz.mem_819_sv2v_reg  <= w_data_i[19];
      \nz.mem_818_sv2v_reg  <= w_data_i[18];
      \nz.mem_817_sv2v_reg  <= w_data_i[17];
      \nz.mem_816_sv2v_reg  <= w_data_i[16];
      \nz.mem_815_sv2v_reg  <= w_data_i[15];
      \nz.mem_814_sv2v_reg  <= w_data_i[14];
      \nz.mem_813_sv2v_reg  <= w_data_i[13];
      \nz.mem_812_sv2v_reg  <= w_data_i[12];
      \nz.mem_811_sv2v_reg  <= w_data_i[11];
      \nz.mem_810_sv2v_reg  <= w_data_i[10];
      \nz.mem_809_sv2v_reg  <= w_data_i[9];
      \nz.mem_808_sv2v_reg  <= w_data_i[8];
      \nz.mem_807_sv2v_reg  <= w_data_i[7];
      \nz.mem_806_sv2v_reg  <= w_data_i[6];
      \nz.mem_805_sv2v_reg  <= w_data_i[5];
      \nz.mem_804_sv2v_reg  <= w_data_i[4];
      \nz.mem_803_sv2v_reg  <= w_data_i[3];
      \nz.mem_802_sv2v_reg  <= w_data_i[2];
      \nz.mem_801_sv2v_reg  <= w_data_i[1];
      \nz.mem_800_sv2v_reg  <= w_data_i[0];
    end 
    if(N220) begin
      \nz.mem_799_sv2v_reg  <= w_data_i[49];
      \nz.mem_798_sv2v_reg  <= w_data_i[48];
      \nz.mem_797_sv2v_reg  <= w_data_i[47];
      \nz.mem_796_sv2v_reg  <= w_data_i[46];
      \nz.mem_795_sv2v_reg  <= w_data_i[45];
      \nz.mem_794_sv2v_reg  <= w_data_i[44];
      \nz.mem_793_sv2v_reg  <= w_data_i[43];
      \nz.mem_792_sv2v_reg  <= w_data_i[42];
      \nz.mem_791_sv2v_reg  <= w_data_i[41];
      \nz.mem_790_sv2v_reg  <= w_data_i[40];
      \nz.mem_789_sv2v_reg  <= w_data_i[39];
      \nz.mem_788_sv2v_reg  <= w_data_i[38];
      \nz.mem_787_sv2v_reg  <= w_data_i[37];
      \nz.mem_786_sv2v_reg  <= w_data_i[36];
      \nz.mem_785_sv2v_reg  <= w_data_i[35];
      \nz.mem_784_sv2v_reg  <= w_data_i[34];
      \nz.mem_783_sv2v_reg  <= w_data_i[33];
      \nz.mem_782_sv2v_reg  <= w_data_i[32];
      \nz.mem_781_sv2v_reg  <= w_data_i[31];
      \nz.mem_780_sv2v_reg  <= w_data_i[30];
      \nz.mem_779_sv2v_reg  <= w_data_i[29];
      \nz.mem_778_sv2v_reg  <= w_data_i[28];
      \nz.mem_777_sv2v_reg  <= w_data_i[27];
      \nz.mem_776_sv2v_reg  <= w_data_i[26];
      \nz.mem_775_sv2v_reg  <= w_data_i[25];
      \nz.mem_774_sv2v_reg  <= w_data_i[24];
      \nz.mem_773_sv2v_reg  <= w_data_i[23];
      \nz.mem_772_sv2v_reg  <= w_data_i[22];
      \nz.mem_771_sv2v_reg  <= w_data_i[21];
      \nz.mem_770_sv2v_reg  <= w_data_i[20];
      \nz.mem_769_sv2v_reg  <= w_data_i[19];
      \nz.mem_768_sv2v_reg  <= w_data_i[18];
      \nz.mem_767_sv2v_reg  <= w_data_i[17];
      \nz.mem_766_sv2v_reg  <= w_data_i[16];
      \nz.mem_765_sv2v_reg  <= w_data_i[15];
      \nz.mem_764_sv2v_reg  <= w_data_i[14];
      \nz.mem_763_sv2v_reg  <= w_data_i[13];
      \nz.mem_762_sv2v_reg  <= w_data_i[12];
      \nz.mem_761_sv2v_reg  <= w_data_i[11];
      \nz.mem_760_sv2v_reg  <= w_data_i[10];
      \nz.mem_759_sv2v_reg  <= w_data_i[9];
      \nz.mem_758_sv2v_reg  <= w_data_i[8];
      \nz.mem_757_sv2v_reg  <= w_data_i[7];
      \nz.mem_756_sv2v_reg  <= w_data_i[6];
      \nz.mem_755_sv2v_reg  <= w_data_i[5];
      \nz.mem_754_sv2v_reg  <= w_data_i[4];
      \nz.mem_753_sv2v_reg  <= w_data_i[3];
      \nz.mem_752_sv2v_reg  <= w_data_i[2];
      \nz.mem_751_sv2v_reg  <= w_data_i[1];
      \nz.mem_750_sv2v_reg  <= w_data_i[0];
    end 
    if(N219) begin
      \nz.mem_749_sv2v_reg  <= w_data_i[49];
      \nz.mem_748_sv2v_reg  <= w_data_i[48];
      \nz.mem_747_sv2v_reg  <= w_data_i[47];
      \nz.mem_746_sv2v_reg  <= w_data_i[46];
      \nz.mem_745_sv2v_reg  <= w_data_i[45];
      \nz.mem_744_sv2v_reg  <= w_data_i[44];
      \nz.mem_743_sv2v_reg  <= w_data_i[43];
      \nz.mem_742_sv2v_reg  <= w_data_i[42];
      \nz.mem_741_sv2v_reg  <= w_data_i[41];
      \nz.mem_740_sv2v_reg  <= w_data_i[40];
      \nz.mem_739_sv2v_reg  <= w_data_i[39];
      \nz.mem_738_sv2v_reg  <= w_data_i[38];
      \nz.mem_737_sv2v_reg  <= w_data_i[37];
      \nz.mem_736_sv2v_reg  <= w_data_i[36];
      \nz.mem_735_sv2v_reg  <= w_data_i[35];
      \nz.mem_734_sv2v_reg  <= w_data_i[34];
      \nz.mem_733_sv2v_reg  <= w_data_i[33];
      \nz.mem_732_sv2v_reg  <= w_data_i[32];
      \nz.mem_731_sv2v_reg  <= w_data_i[31];
      \nz.mem_730_sv2v_reg  <= w_data_i[30];
      \nz.mem_729_sv2v_reg  <= w_data_i[29];
      \nz.mem_728_sv2v_reg  <= w_data_i[28];
      \nz.mem_727_sv2v_reg  <= w_data_i[27];
      \nz.mem_726_sv2v_reg  <= w_data_i[26];
      \nz.mem_725_sv2v_reg  <= w_data_i[25];
      \nz.mem_724_sv2v_reg  <= w_data_i[24];
      \nz.mem_723_sv2v_reg  <= w_data_i[23];
      \nz.mem_722_sv2v_reg  <= w_data_i[22];
      \nz.mem_721_sv2v_reg  <= w_data_i[21];
      \nz.mem_720_sv2v_reg  <= w_data_i[20];
      \nz.mem_719_sv2v_reg  <= w_data_i[19];
      \nz.mem_718_sv2v_reg  <= w_data_i[18];
      \nz.mem_717_sv2v_reg  <= w_data_i[17];
      \nz.mem_716_sv2v_reg  <= w_data_i[16];
      \nz.mem_715_sv2v_reg  <= w_data_i[15];
      \nz.mem_714_sv2v_reg  <= w_data_i[14];
      \nz.mem_713_sv2v_reg  <= w_data_i[13];
      \nz.mem_712_sv2v_reg  <= w_data_i[12];
      \nz.mem_711_sv2v_reg  <= w_data_i[11];
      \nz.mem_710_sv2v_reg  <= w_data_i[10];
      \nz.mem_709_sv2v_reg  <= w_data_i[9];
      \nz.mem_708_sv2v_reg  <= w_data_i[8];
      \nz.mem_707_sv2v_reg  <= w_data_i[7];
      \nz.mem_706_sv2v_reg  <= w_data_i[6];
      \nz.mem_705_sv2v_reg  <= w_data_i[5];
      \nz.mem_704_sv2v_reg  <= w_data_i[4];
      \nz.mem_703_sv2v_reg  <= w_data_i[3];
      \nz.mem_702_sv2v_reg  <= w_data_i[2];
      \nz.mem_701_sv2v_reg  <= w_data_i[1];
      \nz.mem_700_sv2v_reg  <= w_data_i[0];
    end 
    if(N218) begin
      \nz.mem_699_sv2v_reg  <= w_data_i[49];
      \nz.mem_698_sv2v_reg  <= w_data_i[48];
      \nz.mem_697_sv2v_reg  <= w_data_i[47];
      \nz.mem_696_sv2v_reg  <= w_data_i[46];
      \nz.mem_695_sv2v_reg  <= w_data_i[45];
      \nz.mem_694_sv2v_reg  <= w_data_i[44];
      \nz.mem_693_sv2v_reg  <= w_data_i[43];
      \nz.mem_692_sv2v_reg  <= w_data_i[42];
      \nz.mem_691_sv2v_reg  <= w_data_i[41];
      \nz.mem_690_sv2v_reg  <= w_data_i[40];
      \nz.mem_689_sv2v_reg  <= w_data_i[39];
      \nz.mem_688_sv2v_reg  <= w_data_i[38];
      \nz.mem_687_sv2v_reg  <= w_data_i[37];
      \nz.mem_686_sv2v_reg  <= w_data_i[36];
      \nz.mem_685_sv2v_reg  <= w_data_i[35];
      \nz.mem_684_sv2v_reg  <= w_data_i[34];
      \nz.mem_683_sv2v_reg  <= w_data_i[33];
      \nz.mem_682_sv2v_reg  <= w_data_i[32];
      \nz.mem_681_sv2v_reg  <= w_data_i[31];
      \nz.mem_680_sv2v_reg  <= w_data_i[30];
      \nz.mem_679_sv2v_reg  <= w_data_i[29];
      \nz.mem_678_sv2v_reg  <= w_data_i[28];
      \nz.mem_677_sv2v_reg  <= w_data_i[27];
      \nz.mem_676_sv2v_reg  <= w_data_i[26];
      \nz.mem_675_sv2v_reg  <= w_data_i[25];
      \nz.mem_674_sv2v_reg  <= w_data_i[24];
      \nz.mem_673_sv2v_reg  <= w_data_i[23];
      \nz.mem_672_sv2v_reg  <= w_data_i[22];
      \nz.mem_671_sv2v_reg  <= w_data_i[21];
      \nz.mem_670_sv2v_reg  <= w_data_i[20];
      \nz.mem_669_sv2v_reg  <= w_data_i[19];
      \nz.mem_668_sv2v_reg  <= w_data_i[18];
      \nz.mem_667_sv2v_reg  <= w_data_i[17];
      \nz.mem_666_sv2v_reg  <= w_data_i[16];
      \nz.mem_665_sv2v_reg  <= w_data_i[15];
      \nz.mem_664_sv2v_reg  <= w_data_i[14];
      \nz.mem_663_sv2v_reg  <= w_data_i[13];
      \nz.mem_662_sv2v_reg  <= w_data_i[12];
      \nz.mem_661_sv2v_reg  <= w_data_i[11];
      \nz.mem_660_sv2v_reg  <= w_data_i[10];
      \nz.mem_659_sv2v_reg  <= w_data_i[9];
      \nz.mem_658_sv2v_reg  <= w_data_i[8];
      \nz.mem_657_sv2v_reg  <= w_data_i[7];
      \nz.mem_656_sv2v_reg  <= w_data_i[6];
      \nz.mem_655_sv2v_reg  <= w_data_i[5];
      \nz.mem_654_sv2v_reg  <= w_data_i[4];
      \nz.mem_653_sv2v_reg  <= w_data_i[3];
      \nz.mem_652_sv2v_reg  <= w_data_i[2];
      \nz.mem_651_sv2v_reg  <= w_data_i[1];
      \nz.mem_650_sv2v_reg  <= w_data_i[0];
    end 
    if(N217) begin
      \nz.mem_649_sv2v_reg  <= w_data_i[49];
      \nz.mem_648_sv2v_reg  <= w_data_i[48];
      \nz.mem_647_sv2v_reg  <= w_data_i[47];
      \nz.mem_646_sv2v_reg  <= w_data_i[46];
      \nz.mem_645_sv2v_reg  <= w_data_i[45];
      \nz.mem_644_sv2v_reg  <= w_data_i[44];
      \nz.mem_643_sv2v_reg  <= w_data_i[43];
      \nz.mem_642_sv2v_reg  <= w_data_i[42];
      \nz.mem_641_sv2v_reg  <= w_data_i[41];
      \nz.mem_640_sv2v_reg  <= w_data_i[40];
      \nz.mem_639_sv2v_reg  <= w_data_i[39];
      \nz.mem_638_sv2v_reg  <= w_data_i[38];
      \nz.mem_637_sv2v_reg  <= w_data_i[37];
      \nz.mem_636_sv2v_reg  <= w_data_i[36];
      \nz.mem_635_sv2v_reg  <= w_data_i[35];
      \nz.mem_634_sv2v_reg  <= w_data_i[34];
      \nz.mem_633_sv2v_reg  <= w_data_i[33];
      \nz.mem_632_sv2v_reg  <= w_data_i[32];
      \nz.mem_631_sv2v_reg  <= w_data_i[31];
      \nz.mem_630_sv2v_reg  <= w_data_i[30];
      \nz.mem_629_sv2v_reg  <= w_data_i[29];
      \nz.mem_628_sv2v_reg  <= w_data_i[28];
      \nz.mem_627_sv2v_reg  <= w_data_i[27];
      \nz.mem_626_sv2v_reg  <= w_data_i[26];
      \nz.mem_625_sv2v_reg  <= w_data_i[25];
      \nz.mem_624_sv2v_reg  <= w_data_i[24];
      \nz.mem_623_sv2v_reg  <= w_data_i[23];
      \nz.mem_622_sv2v_reg  <= w_data_i[22];
      \nz.mem_621_sv2v_reg  <= w_data_i[21];
      \nz.mem_620_sv2v_reg  <= w_data_i[20];
      \nz.mem_619_sv2v_reg  <= w_data_i[19];
      \nz.mem_618_sv2v_reg  <= w_data_i[18];
      \nz.mem_617_sv2v_reg  <= w_data_i[17];
      \nz.mem_616_sv2v_reg  <= w_data_i[16];
      \nz.mem_615_sv2v_reg  <= w_data_i[15];
      \nz.mem_614_sv2v_reg  <= w_data_i[14];
      \nz.mem_613_sv2v_reg  <= w_data_i[13];
      \nz.mem_612_sv2v_reg  <= w_data_i[12];
      \nz.mem_611_sv2v_reg  <= w_data_i[11];
      \nz.mem_610_sv2v_reg  <= w_data_i[10];
      \nz.mem_609_sv2v_reg  <= w_data_i[9];
      \nz.mem_608_sv2v_reg  <= w_data_i[8];
      \nz.mem_607_sv2v_reg  <= w_data_i[7];
      \nz.mem_606_sv2v_reg  <= w_data_i[6];
      \nz.mem_605_sv2v_reg  <= w_data_i[5];
      \nz.mem_604_sv2v_reg  <= w_data_i[4];
      \nz.mem_603_sv2v_reg  <= w_data_i[3];
      \nz.mem_602_sv2v_reg  <= w_data_i[2];
      \nz.mem_601_sv2v_reg  <= w_data_i[1];
      \nz.mem_600_sv2v_reg  <= w_data_i[0];
    end 
    if(N216) begin
      \nz.mem_599_sv2v_reg  <= w_data_i[49];
      \nz.mem_598_sv2v_reg  <= w_data_i[48];
      \nz.mem_597_sv2v_reg  <= w_data_i[47];
      \nz.mem_596_sv2v_reg  <= w_data_i[46];
      \nz.mem_595_sv2v_reg  <= w_data_i[45];
      \nz.mem_594_sv2v_reg  <= w_data_i[44];
      \nz.mem_593_sv2v_reg  <= w_data_i[43];
      \nz.mem_592_sv2v_reg  <= w_data_i[42];
      \nz.mem_591_sv2v_reg  <= w_data_i[41];
      \nz.mem_590_sv2v_reg  <= w_data_i[40];
      \nz.mem_589_sv2v_reg  <= w_data_i[39];
      \nz.mem_588_sv2v_reg  <= w_data_i[38];
      \nz.mem_587_sv2v_reg  <= w_data_i[37];
      \nz.mem_586_sv2v_reg  <= w_data_i[36];
      \nz.mem_585_sv2v_reg  <= w_data_i[35];
      \nz.mem_584_sv2v_reg  <= w_data_i[34];
      \nz.mem_583_sv2v_reg  <= w_data_i[33];
      \nz.mem_582_sv2v_reg  <= w_data_i[32];
      \nz.mem_581_sv2v_reg  <= w_data_i[31];
      \nz.mem_580_sv2v_reg  <= w_data_i[30];
      \nz.mem_579_sv2v_reg  <= w_data_i[29];
      \nz.mem_578_sv2v_reg  <= w_data_i[28];
      \nz.mem_577_sv2v_reg  <= w_data_i[27];
      \nz.mem_576_sv2v_reg  <= w_data_i[26];
      \nz.mem_575_sv2v_reg  <= w_data_i[25];
      \nz.mem_574_sv2v_reg  <= w_data_i[24];
      \nz.mem_573_sv2v_reg  <= w_data_i[23];
      \nz.mem_572_sv2v_reg  <= w_data_i[22];
      \nz.mem_571_sv2v_reg  <= w_data_i[21];
      \nz.mem_570_sv2v_reg  <= w_data_i[20];
      \nz.mem_569_sv2v_reg  <= w_data_i[19];
      \nz.mem_568_sv2v_reg  <= w_data_i[18];
      \nz.mem_567_sv2v_reg  <= w_data_i[17];
      \nz.mem_566_sv2v_reg  <= w_data_i[16];
      \nz.mem_565_sv2v_reg  <= w_data_i[15];
      \nz.mem_564_sv2v_reg  <= w_data_i[14];
      \nz.mem_563_sv2v_reg  <= w_data_i[13];
      \nz.mem_562_sv2v_reg  <= w_data_i[12];
      \nz.mem_561_sv2v_reg  <= w_data_i[11];
      \nz.mem_560_sv2v_reg  <= w_data_i[10];
      \nz.mem_559_sv2v_reg  <= w_data_i[9];
      \nz.mem_558_sv2v_reg  <= w_data_i[8];
      \nz.mem_557_sv2v_reg  <= w_data_i[7];
      \nz.mem_556_sv2v_reg  <= w_data_i[6];
      \nz.mem_555_sv2v_reg  <= w_data_i[5];
      \nz.mem_554_sv2v_reg  <= w_data_i[4];
      \nz.mem_553_sv2v_reg  <= w_data_i[3];
      \nz.mem_552_sv2v_reg  <= w_data_i[2];
      \nz.mem_551_sv2v_reg  <= w_data_i[1];
      \nz.mem_550_sv2v_reg  <= w_data_i[0];
    end 
    if(N215) begin
      \nz.mem_549_sv2v_reg  <= w_data_i[49];
      \nz.mem_548_sv2v_reg  <= w_data_i[48];
      \nz.mem_547_sv2v_reg  <= w_data_i[47];
      \nz.mem_546_sv2v_reg  <= w_data_i[46];
      \nz.mem_545_sv2v_reg  <= w_data_i[45];
      \nz.mem_544_sv2v_reg  <= w_data_i[44];
      \nz.mem_543_sv2v_reg  <= w_data_i[43];
      \nz.mem_542_sv2v_reg  <= w_data_i[42];
      \nz.mem_541_sv2v_reg  <= w_data_i[41];
      \nz.mem_540_sv2v_reg  <= w_data_i[40];
      \nz.mem_539_sv2v_reg  <= w_data_i[39];
      \nz.mem_538_sv2v_reg  <= w_data_i[38];
      \nz.mem_537_sv2v_reg  <= w_data_i[37];
      \nz.mem_536_sv2v_reg  <= w_data_i[36];
      \nz.mem_535_sv2v_reg  <= w_data_i[35];
      \nz.mem_534_sv2v_reg  <= w_data_i[34];
      \nz.mem_533_sv2v_reg  <= w_data_i[33];
      \nz.mem_532_sv2v_reg  <= w_data_i[32];
      \nz.mem_531_sv2v_reg  <= w_data_i[31];
      \nz.mem_530_sv2v_reg  <= w_data_i[30];
      \nz.mem_529_sv2v_reg  <= w_data_i[29];
      \nz.mem_528_sv2v_reg  <= w_data_i[28];
      \nz.mem_527_sv2v_reg  <= w_data_i[27];
      \nz.mem_526_sv2v_reg  <= w_data_i[26];
      \nz.mem_525_sv2v_reg  <= w_data_i[25];
      \nz.mem_524_sv2v_reg  <= w_data_i[24];
      \nz.mem_523_sv2v_reg  <= w_data_i[23];
      \nz.mem_522_sv2v_reg  <= w_data_i[22];
      \nz.mem_521_sv2v_reg  <= w_data_i[21];
      \nz.mem_520_sv2v_reg  <= w_data_i[20];
      \nz.mem_519_sv2v_reg  <= w_data_i[19];
      \nz.mem_518_sv2v_reg  <= w_data_i[18];
      \nz.mem_517_sv2v_reg  <= w_data_i[17];
      \nz.mem_516_sv2v_reg  <= w_data_i[16];
      \nz.mem_515_sv2v_reg  <= w_data_i[15];
      \nz.mem_514_sv2v_reg  <= w_data_i[14];
      \nz.mem_513_sv2v_reg  <= w_data_i[13];
      \nz.mem_512_sv2v_reg  <= w_data_i[12];
      \nz.mem_511_sv2v_reg  <= w_data_i[11];
      \nz.mem_510_sv2v_reg  <= w_data_i[10];
      \nz.mem_509_sv2v_reg  <= w_data_i[9];
      \nz.mem_508_sv2v_reg  <= w_data_i[8];
      \nz.mem_507_sv2v_reg  <= w_data_i[7];
      \nz.mem_506_sv2v_reg  <= w_data_i[6];
      \nz.mem_505_sv2v_reg  <= w_data_i[5];
      \nz.mem_504_sv2v_reg  <= w_data_i[4];
      \nz.mem_503_sv2v_reg  <= w_data_i[3];
      \nz.mem_502_sv2v_reg  <= w_data_i[2];
      \nz.mem_501_sv2v_reg  <= w_data_i[1];
      \nz.mem_500_sv2v_reg  <= w_data_i[0];
    end 
    if(N214) begin
      \nz.mem_499_sv2v_reg  <= w_data_i[49];
      \nz.mem_498_sv2v_reg  <= w_data_i[48];
      \nz.mem_497_sv2v_reg  <= w_data_i[47];
      \nz.mem_496_sv2v_reg  <= w_data_i[46];
      \nz.mem_495_sv2v_reg  <= w_data_i[45];
      \nz.mem_494_sv2v_reg  <= w_data_i[44];
      \nz.mem_493_sv2v_reg  <= w_data_i[43];
      \nz.mem_492_sv2v_reg  <= w_data_i[42];
      \nz.mem_491_sv2v_reg  <= w_data_i[41];
      \nz.mem_490_sv2v_reg  <= w_data_i[40];
      \nz.mem_489_sv2v_reg  <= w_data_i[39];
      \nz.mem_488_sv2v_reg  <= w_data_i[38];
      \nz.mem_487_sv2v_reg  <= w_data_i[37];
      \nz.mem_486_sv2v_reg  <= w_data_i[36];
      \nz.mem_485_sv2v_reg  <= w_data_i[35];
      \nz.mem_484_sv2v_reg  <= w_data_i[34];
      \nz.mem_483_sv2v_reg  <= w_data_i[33];
      \nz.mem_482_sv2v_reg  <= w_data_i[32];
      \nz.mem_481_sv2v_reg  <= w_data_i[31];
      \nz.mem_480_sv2v_reg  <= w_data_i[30];
      \nz.mem_479_sv2v_reg  <= w_data_i[29];
      \nz.mem_478_sv2v_reg  <= w_data_i[28];
      \nz.mem_477_sv2v_reg  <= w_data_i[27];
      \nz.mem_476_sv2v_reg  <= w_data_i[26];
      \nz.mem_475_sv2v_reg  <= w_data_i[25];
      \nz.mem_474_sv2v_reg  <= w_data_i[24];
      \nz.mem_473_sv2v_reg  <= w_data_i[23];
      \nz.mem_472_sv2v_reg  <= w_data_i[22];
      \nz.mem_471_sv2v_reg  <= w_data_i[21];
      \nz.mem_470_sv2v_reg  <= w_data_i[20];
      \nz.mem_469_sv2v_reg  <= w_data_i[19];
      \nz.mem_468_sv2v_reg  <= w_data_i[18];
      \nz.mem_467_sv2v_reg  <= w_data_i[17];
      \nz.mem_466_sv2v_reg  <= w_data_i[16];
      \nz.mem_465_sv2v_reg  <= w_data_i[15];
      \nz.mem_464_sv2v_reg  <= w_data_i[14];
      \nz.mem_463_sv2v_reg  <= w_data_i[13];
      \nz.mem_462_sv2v_reg  <= w_data_i[12];
      \nz.mem_461_sv2v_reg  <= w_data_i[11];
      \nz.mem_460_sv2v_reg  <= w_data_i[10];
      \nz.mem_459_sv2v_reg  <= w_data_i[9];
      \nz.mem_458_sv2v_reg  <= w_data_i[8];
      \nz.mem_457_sv2v_reg  <= w_data_i[7];
      \nz.mem_456_sv2v_reg  <= w_data_i[6];
      \nz.mem_455_sv2v_reg  <= w_data_i[5];
      \nz.mem_454_sv2v_reg  <= w_data_i[4];
      \nz.mem_453_sv2v_reg  <= w_data_i[3];
      \nz.mem_452_sv2v_reg  <= w_data_i[2];
      \nz.mem_451_sv2v_reg  <= w_data_i[1];
      \nz.mem_450_sv2v_reg  <= w_data_i[0];
    end 
    if(N213) begin
      \nz.mem_449_sv2v_reg  <= w_data_i[49];
      \nz.mem_448_sv2v_reg  <= w_data_i[48];
      \nz.mem_447_sv2v_reg  <= w_data_i[47];
      \nz.mem_446_sv2v_reg  <= w_data_i[46];
      \nz.mem_445_sv2v_reg  <= w_data_i[45];
      \nz.mem_444_sv2v_reg  <= w_data_i[44];
      \nz.mem_443_sv2v_reg  <= w_data_i[43];
      \nz.mem_442_sv2v_reg  <= w_data_i[42];
      \nz.mem_441_sv2v_reg  <= w_data_i[41];
      \nz.mem_440_sv2v_reg  <= w_data_i[40];
      \nz.mem_439_sv2v_reg  <= w_data_i[39];
      \nz.mem_438_sv2v_reg  <= w_data_i[38];
      \nz.mem_437_sv2v_reg  <= w_data_i[37];
      \nz.mem_436_sv2v_reg  <= w_data_i[36];
      \nz.mem_435_sv2v_reg  <= w_data_i[35];
      \nz.mem_434_sv2v_reg  <= w_data_i[34];
      \nz.mem_433_sv2v_reg  <= w_data_i[33];
      \nz.mem_432_sv2v_reg  <= w_data_i[32];
      \nz.mem_431_sv2v_reg  <= w_data_i[31];
      \nz.mem_430_sv2v_reg  <= w_data_i[30];
      \nz.mem_429_sv2v_reg  <= w_data_i[29];
      \nz.mem_428_sv2v_reg  <= w_data_i[28];
      \nz.mem_427_sv2v_reg  <= w_data_i[27];
      \nz.mem_426_sv2v_reg  <= w_data_i[26];
      \nz.mem_425_sv2v_reg  <= w_data_i[25];
      \nz.mem_424_sv2v_reg  <= w_data_i[24];
      \nz.mem_423_sv2v_reg  <= w_data_i[23];
      \nz.mem_422_sv2v_reg  <= w_data_i[22];
      \nz.mem_421_sv2v_reg  <= w_data_i[21];
      \nz.mem_420_sv2v_reg  <= w_data_i[20];
      \nz.mem_419_sv2v_reg  <= w_data_i[19];
      \nz.mem_418_sv2v_reg  <= w_data_i[18];
      \nz.mem_417_sv2v_reg  <= w_data_i[17];
      \nz.mem_416_sv2v_reg  <= w_data_i[16];
      \nz.mem_415_sv2v_reg  <= w_data_i[15];
      \nz.mem_414_sv2v_reg  <= w_data_i[14];
      \nz.mem_413_sv2v_reg  <= w_data_i[13];
      \nz.mem_412_sv2v_reg  <= w_data_i[12];
      \nz.mem_411_sv2v_reg  <= w_data_i[11];
      \nz.mem_410_sv2v_reg  <= w_data_i[10];
      \nz.mem_409_sv2v_reg  <= w_data_i[9];
      \nz.mem_408_sv2v_reg  <= w_data_i[8];
      \nz.mem_407_sv2v_reg  <= w_data_i[7];
      \nz.mem_406_sv2v_reg  <= w_data_i[6];
      \nz.mem_405_sv2v_reg  <= w_data_i[5];
      \nz.mem_404_sv2v_reg  <= w_data_i[4];
      \nz.mem_403_sv2v_reg  <= w_data_i[3];
      \nz.mem_402_sv2v_reg  <= w_data_i[2];
      \nz.mem_401_sv2v_reg  <= w_data_i[1];
      \nz.mem_400_sv2v_reg  <= w_data_i[0];
    end 
    if(N212) begin
      \nz.mem_399_sv2v_reg  <= w_data_i[49];
      \nz.mem_398_sv2v_reg  <= w_data_i[48];
      \nz.mem_397_sv2v_reg  <= w_data_i[47];
      \nz.mem_396_sv2v_reg  <= w_data_i[46];
      \nz.mem_395_sv2v_reg  <= w_data_i[45];
      \nz.mem_394_sv2v_reg  <= w_data_i[44];
      \nz.mem_393_sv2v_reg  <= w_data_i[43];
      \nz.mem_392_sv2v_reg  <= w_data_i[42];
      \nz.mem_391_sv2v_reg  <= w_data_i[41];
      \nz.mem_390_sv2v_reg  <= w_data_i[40];
      \nz.mem_389_sv2v_reg  <= w_data_i[39];
      \nz.mem_388_sv2v_reg  <= w_data_i[38];
      \nz.mem_387_sv2v_reg  <= w_data_i[37];
      \nz.mem_386_sv2v_reg  <= w_data_i[36];
      \nz.mem_385_sv2v_reg  <= w_data_i[35];
      \nz.mem_384_sv2v_reg  <= w_data_i[34];
      \nz.mem_383_sv2v_reg  <= w_data_i[33];
      \nz.mem_382_sv2v_reg  <= w_data_i[32];
      \nz.mem_381_sv2v_reg  <= w_data_i[31];
      \nz.mem_380_sv2v_reg  <= w_data_i[30];
      \nz.mem_379_sv2v_reg  <= w_data_i[29];
      \nz.mem_378_sv2v_reg  <= w_data_i[28];
      \nz.mem_377_sv2v_reg  <= w_data_i[27];
      \nz.mem_376_sv2v_reg  <= w_data_i[26];
      \nz.mem_375_sv2v_reg  <= w_data_i[25];
      \nz.mem_374_sv2v_reg  <= w_data_i[24];
      \nz.mem_373_sv2v_reg  <= w_data_i[23];
      \nz.mem_372_sv2v_reg  <= w_data_i[22];
      \nz.mem_371_sv2v_reg  <= w_data_i[21];
      \nz.mem_370_sv2v_reg  <= w_data_i[20];
      \nz.mem_369_sv2v_reg  <= w_data_i[19];
      \nz.mem_368_sv2v_reg  <= w_data_i[18];
      \nz.mem_367_sv2v_reg  <= w_data_i[17];
      \nz.mem_366_sv2v_reg  <= w_data_i[16];
      \nz.mem_365_sv2v_reg  <= w_data_i[15];
      \nz.mem_364_sv2v_reg  <= w_data_i[14];
      \nz.mem_363_sv2v_reg  <= w_data_i[13];
      \nz.mem_362_sv2v_reg  <= w_data_i[12];
      \nz.mem_361_sv2v_reg  <= w_data_i[11];
      \nz.mem_360_sv2v_reg  <= w_data_i[10];
      \nz.mem_359_sv2v_reg  <= w_data_i[9];
      \nz.mem_358_sv2v_reg  <= w_data_i[8];
      \nz.mem_357_sv2v_reg  <= w_data_i[7];
      \nz.mem_356_sv2v_reg  <= w_data_i[6];
      \nz.mem_355_sv2v_reg  <= w_data_i[5];
      \nz.mem_354_sv2v_reg  <= w_data_i[4];
      \nz.mem_353_sv2v_reg  <= w_data_i[3];
      \nz.mem_352_sv2v_reg  <= w_data_i[2];
      \nz.mem_351_sv2v_reg  <= w_data_i[1];
      \nz.mem_350_sv2v_reg  <= w_data_i[0];
    end 
    if(N211) begin
      \nz.mem_349_sv2v_reg  <= w_data_i[49];
      \nz.mem_348_sv2v_reg  <= w_data_i[48];
      \nz.mem_347_sv2v_reg  <= w_data_i[47];
      \nz.mem_346_sv2v_reg  <= w_data_i[46];
      \nz.mem_345_sv2v_reg  <= w_data_i[45];
      \nz.mem_344_sv2v_reg  <= w_data_i[44];
      \nz.mem_343_sv2v_reg  <= w_data_i[43];
      \nz.mem_342_sv2v_reg  <= w_data_i[42];
      \nz.mem_341_sv2v_reg  <= w_data_i[41];
      \nz.mem_340_sv2v_reg  <= w_data_i[40];
      \nz.mem_339_sv2v_reg  <= w_data_i[39];
      \nz.mem_338_sv2v_reg  <= w_data_i[38];
      \nz.mem_337_sv2v_reg  <= w_data_i[37];
      \nz.mem_336_sv2v_reg  <= w_data_i[36];
      \nz.mem_335_sv2v_reg  <= w_data_i[35];
      \nz.mem_334_sv2v_reg  <= w_data_i[34];
      \nz.mem_333_sv2v_reg  <= w_data_i[33];
      \nz.mem_332_sv2v_reg  <= w_data_i[32];
      \nz.mem_331_sv2v_reg  <= w_data_i[31];
      \nz.mem_330_sv2v_reg  <= w_data_i[30];
      \nz.mem_329_sv2v_reg  <= w_data_i[29];
      \nz.mem_328_sv2v_reg  <= w_data_i[28];
      \nz.mem_327_sv2v_reg  <= w_data_i[27];
      \nz.mem_326_sv2v_reg  <= w_data_i[26];
      \nz.mem_325_sv2v_reg  <= w_data_i[25];
      \nz.mem_324_sv2v_reg  <= w_data_i[24];
      \nz.mem_323_sv2v_reg  <= w_data_i[23];
      \nz.mem_322_sv2v_reg  <= w_data_i[22];
      \nz.mem_321_sv2v_reg  <= w_data_i[21];
      \nz.mem_320_sv2v_reg  <= w_data_i[20];
      \nz.mem_319_sv2v_reg  <= w_data_i[19];
      \nz.mem_318_sv2v_reg  <= w_data_i[18];
      \nz.mem_317_sv2v_reg  <= w_data_i[17];
      \nz.mem_316_sv2v_reg  <= w_data_i[16];
      \nz.mem_315_sv2v_reg  <= w_data_i[15];
      \nz.mem_314_sv2v_reg  <= w_data_i[14];
      \nz.mem_313_sv2v_reg  <= w_data_i[13];
      \nz.mem_312_sv2v_reg  <= w_data_i[12];
      \nz.mem_311_sv2v_reg  <= w_data_i[11];
      \nz.mem_310_sv2v_reg  <= w_data_i[10];
      \nz.mem_309_sv2v_reg  <= w_data_i[9];
      \nz.mem_308_sv2v_reg  <= w_data_i[8];
      \nz.mem_307_sv2v_reg  <= w_data_i[7];
      \nz.mem_306_sv2v_reg  <= w_data_i[6];
      \nz.mem_305_sv2v_reg  <= w_data_i[5];
      \nz.mem_304_sv2v_reg  <= w_data_i[4];
      \nz.mem_303_sv2v_reg  <= w_data_i[3];
      \nz.mem_302_sv2v_reg  <= w_data_i[2];
      \nz.mem_301_sv2v_reg  <= w_data_i[1];
      \nz.mem_300_sv2v_reg  <= w_data_i[0];
    end 
    if(N210) begin
      \nz.mem_299_sv2v_reg  <= w_data_i[49];
      \nz.mem_298_sv2v_reg  <= w_data_i[48];
      \nz.mem_297_sv2v_reg  <= w_data_i[47];
      \nz.mem_296_sv2v_reg  <= w_data_i[46];
      \nz.mem_295_sv2v_reg  <= w_data_i[45];
      \nz.mem_294_sv2v_reg  <= w_data_i[44];
      \nz.mem_293_sv2v_reg  <= w_data_i[43];
      \nz.mem_292_sv2v_reg  <= w_data_i[42];
      \nz.mem_291_sv2v_reg  <= w_data_i[41];
      \nz.mem_290_sv2v_reg  <= w_data_i[40];
      \nz.mem_289_sv2v_reg  <= w_data_i[39];
      \nz.mem_288_sv2v_reg  <= w_data_i[38];
      \nz.mem_287_sv2v_reg  <= w_data_i[37];
      \nz.mem_286_sv2v_reg  <= w_data_i[36];
      \nz.mem_285_sv2v_reg  <= w_data_i[35];
      \nz.mem_284_sv2v_reg  <= w_data_i[34];
      \nz.mem_283_sv2v_reg  <= w_data_i[33];
      \nz.mem_282_sv2v_reg  <= w_data_i[32];
      \nz.mem_281_sv2v_reg  <= w_data_i[31];
      \nz.mem_280_sv2v_reg  <= w_data_i[30];
      \nz.mem_279_sv2v_reg  <= w_data_i[29];
      \nz.mem_278_sv2v_reg  <= w_data_i[28];
      \nz.mem_277_sv2v_reg  <= w_data_i[27];
      \nz.mem_276_sv2v_reg  <= w_data_i[26];
      \nz.mem_275_sv2v_reg  <= w_data_i[25];
      \nz.mem_274_sv2v_reg  <= w_data_i[24];
      \nz.mem_273_sv2v_reg  <= w_data_i[23];
      \nz.mem_272_sv2v_reg  <= w_data_i[22];
      \nz.mem_271_sv2v_reg  <= w_data_i[21];
      \nz.mem_270_sv2v_reg  <= w_data_i[20];
      \nz.mem_269_sv2v_reg  <= w_data_i[19];
      \nz.mem_268_sv2v_reg  <= w_data_i[18];
      \nz.mem_267_sv2v_reg  <= w_data_i[17];
      \nz.mem_266_sv2v_reg  <= w_data_i[16];
      \nz.mem_265_sv2v_reg  <= w_data_i[15];
      \nz.mem_264_sv2v_reg  <= w_data_i[14];
      \nz.mem_263_sv2v_reg  <= w_data_i[13];
      \nz.mem_262_sv2v_reg  <= w_data_i[12];
      \nz.mem_261_sv2v_reg  <= w_data_i[11];
      \nz.mem_260_sv2v_reg  <= w_data_i[10];
      \nz.mem_259_sv2v_reg  <= w_data_i[9];
      \nz.mem_258_sv2v_reg  <= w_data_i[8];
      \nz.mem_257_sv2v_reg  <= w_data_i[7];
      \nz.mem_256_sv2v_reg  <= w_data_i[6];
      \nz.mem_255_sv2v_reg  <= w_data_i[5];
      \nz.mem_254_sv2v_reg  <= w_data_i[4];
      \nz.mem_253_sv2v_reg  <= w_data_i[3];
      \nz.mem_252_sv2v_reg  <= w_data_i[2];
      \nz.mem_251_sv2v_reg  <= w_data_i[1];
      \nz.mem_250_sv2v_reg  <= w_data_i[0];
    end 
    if(N209) begin
      \nz.mem_249_sv2v_reg  <= w_data_i[49];
      \nz.mem_248_sv2v_reg  <= w_data_i[48];
      \nz.mem_247_sv2v_reg  <= w_data_i[47];
      \nz.mem_246_sv2v_reg  <= w_data_i[46];
      \nz.mem_245_sv2v_reg  <= w_data_i[45];
      \nz.mem_244_sv2v_reg  <= w_data_i[44];
      \nz.mem_243_sv2v_reg  <= w_data_i[43];
      \nz.mem_242_sv2v_reg  <= w_data_i[42];
      \nz.mem_241_sv2v_reg  <= w_data_i[41];
      \nz.mem_240_sv2v_reg  <= w_data_i[40];
      \nz.mem_239_sv2v_reg  <= w_data_i[39];
      \nz.mem_238_sv2v_reg  <= w_data_i[38];
      \nz.mem_237_sv2v_reg  <= w_data_i[37];
      \nz.mem_236_sv2v_reg  <= w_data_i[36];
      \nz.mem_235_sv2v_reg  <= w_data_i[35];
      \nz.mem_234_sv2v_reg  <= w_data_i[34];
      \nz.mem_233_sv2v_reg  <= w_data_i[33];
      \nz.mem_232_sv2v_reg  <= w_data_i[32];
      \nz.mem_231_sv2v_reg  <= w_data_i[31];
      \nz.mem_230_sv2v_reg  <= w_data_i[30];
      \nz.mem_229_sv2v_reg  <= w_data_i[29];
      \nz.mem_228_sv2v_reg  <= w_data_i[28];
      \nz.mem_227_sv2v_reg  <= w_data_i[27];
      \nz.mem_226_sv2v_reg  <= w_data_i[26];
      \nz.mem_225_sv2v_reg  <= w_data_i[25];
      \nz.mem_224_sv2v_reg  <= w_data_i[24];
      \nz.mem_223_sv2v_reg  <= w_data_i[23];
      \nz.mem_222_sv2v_reg  <= w_data_i[22];
      \nz.mem_221_sv2v_reg  <= w_data_i[21];
      \nz.mem_220_sv2v_reg  <= w_data_i[20];
      \nz.mem_219_sv2v_reg  <= w_data_i[19];
      \nz.mem_218_sv2v_reg  <= w_data_i[18];
      \nz.mem_217_sv2v_reg  <= w_data_i[17];
      \nz.mem_216_sv2v_reg  <= w_data_i[16];
      \nz.mem_215_sv2v_reg  <= w_data_i[15];
      \nz.mem_214_sv2v_reg  <= w_data_i[14];
      \nz.mem_213_sv2v_reg  <= w_data_i[13];
      \nz.mem_212_sv2v_reg  <= w_data_i[12];
      \nz.mem_211_sv2v_reg  <= w_data_i[11];
      \nz.mem_210_sv2v_reg  <= w_data_i[10];
      \nz.mem_209_sv2v_reg  <= w_data_i[9];
      \nz.mem_208_sv2v_reg  <= w_data_i[8];
      \nz.mem_207_sv2v_reg  <= w_data_i[7];
      \nz.mem_206_sv2v_reg  <= w_data_i[6];
      \nz.mem_205_sv2v_reg  <= w_data_i[5];
      \nz.mem_204_sv2v_reg  <= w_data_i[4];
      \nz.mem_203_sv2v_reg  <= w_data_i[3];
      \nz.mem_202_sv2v_reg  <= w_data_i[2];
      \nz.mem_201_sv2v_reg  <= w_data_i[1];
      \nz.mem_200_sv2v_reg  <= w_data_i[0];
    end 
    if(N208) begin
      \nz.mem_199_sv2v_reg  <= w_data_i[49];
      \nz.mem_198_sv2v_reg  <= w_data_i[48];
      \nz.mem_197_sv2v_reg  <= w_data_i[47];
      \nz.mem_196_sv2v_reg  <= w_data_i[46];
      \nz.mem_195_sv2v_reg  <= w_data_i[45];
      \nz.mem_194_sv2v_reg  <= w_data_i[44];
      \nz.mem_193_sv2v_reg  <= w_data_i[43];
      \nz.mem_192_sv2v_reg  <= w_data_i[42];
      \nz.mem_191_sv2v_reg  <= w_data_i[41];
      \nz.mem_190_sv2v_reg  <= w_data_i[40];
      \nz.mem_189_sv2v_reg  <= w_data_i[39];
      \nz.mem_188_sv2v_reg  <= w_data_i[38];
      \nz.mem_187_sv2v_reg  <= w_data_i[37];
      \nz.mem_186_sv2v_reg  <= w_data_i[36];
      \nz.mem_185_sv2v_reg  <= w_data_i[35];
      \nz.mem_184_sv2v_reg  <= w_data_i[34];
      \nz.mem_183_sv2v_reg  <= w_data_i[33];
      \nz.mem_182_sv2v_reg  <= w_data_i[32];
      \nz.mem_181_sv2v_reg  <= w_data_i[31];
      \nz.mem_180_sv2v_reg  <= w_data_i[30];
      \nz.mem_179_sv2v_reg  <= w_data_i[29];
      \nz.mem_178_sv2v_reg  <= w_data_i[28];
      \nz.mem_177_sv2v_reg  <= w_data_i[27];
      \nz.mem_176_sv2v_reg  <= w_data_i[26];
      \nz.mem_175_sv2v_reg  <= w_data_i[25];
      \nz.mem_174_sv2v_reg  <= w_data_i[24];
      \nz.mem_173_sv2v_reg  <= w_data_i[23];
      \nz.mem_172_sv2v_reg  <= w_data_i[22];
      \nz.mem_171_sv2v_reg  <= w_data_i[21];
      \nz.mem_170_sv2v_reg  <= w_data_i[20];
      \nz.mem_169_sv2v_reg  <= w_data_i[19];
      \nz.mem_168_sv2v_reg  <= w_data_i[18];
      \nz.mem_167_sv2v_reg  <= w_data_i[17];
      \nz.mem_166_sv2v_reg  <= w_data_i[16];
      \nz.mem_165_sv2v_reg  <= w_data_i[15];
      \nz.mem_164_sv2v_reg  <= w_data_i[14];
      \nz.mem_163_sv2v_reg  <= w_data_i[13];
      \nz.mem_162_sv2v_reg  <= w_data_i[12];
      \nz.mem_161_sv2v_reg  <= w_data_i[11];
      \nz.mem_160_sv2v_reg  <= w_data_i[10];
      \nz.mem_159_sv2v_reg  <= w_data_i[9];
      \nz.mem_158_sv2v_reg  <= w_data_i[8];
      \nz.mem_157_sv2v_reg  <= w_data_i[7];
      \nz.mem_156_sv2v_reg  <= w_data_i[6];
      \nz.mem_155_sv2v_reg  <= w_data_i[5];
      \nz.mem_154_sv2v_reg  <= w_data_i[4];
      \nz.mem_153_sv2v_reg  <= w_data_i[3];
      \nz.mem_152_sv2v_reg  <= w_data_i[2];
      \nz.mem_151_sv2v_reg  <= w_data_i[1];
      \nz.mem_150_sv2v_reg  <= w_data_i[0];
    end 
    if(N207) begin
      \nz.mem_149_sv2v_reg  <= w_data_i[49];
      \nz.mem_148_sv2v_reg  <= w_data_i[48];
      \nz.mem_147_sv2v_reg  <= w_data_i[47];
      \nz.mem_146_sv2v_reg  <= w_data_i[46];
      \nz.mem_145_sv2v_reg  <= w_data_i[45];
      \nz.mem_144_sv2v_reg  <= w_data_i[44];
      \nz.mem_143_sv2v_reg  <= w_data_i[43];
      \nz.mem_142_sv2v_reg  <= w_data_i[42];
      \nz.mem_141_sv2v_reg  <= w_data_i[41];
      \nz.mem_140_sv2v_reg  <= w_data_i[40];
      \nz.mem_139_sv2v_reg  <= w_data_i[39];
      \nz.mem_138_sv2v_reg  <= w_data_i[38];
      \nz.mem_137_sv2v_reg  <= w_data_i[37];
      \nz.mem_136_sv2v_reg  <= w_data_i[36];
      \nz.mem_135_sv2v_reg  <= w_data_i[35];
      \nz.mem_134_sv2v_reg  <= w_data_i[34];
      \nz.mem_133_sv2v_reg  <= w_data_i[33];
      \nz.mem_132_sv2v_reg  <= w_data_i[32];
      \nz.mem_131_sv2v_reg  <= w_data_i[31];
      \nz.mem_130_sv2v_reg  <= w_data_i[30];
      \nz.mem_129_sv2v_reg  <= w_data_i[29];
      \nz.mem_128_sv2v_reg  <= w_data_i[28];
      \nz.mem_127_sv2v_reg  <= w_data_i[27];
      \nz.mem_126_sv2v_reg  <= w_data_i[26];
      \nz.mem_125_sv2v_reg  <= w_data_i[25];
      \nz.mem_124_sv2v_reg  <= w_data_i[24];
      \nz.mem_123_sv2v_reg  <= w_data_i[23];
      \nz.mem_122_sv2v_reg  <= w_data_i[22];
      \nz.mem_121_sv2v_reg  <= w_data_i[21];
      \nz.mem_120_sv2v_reg  <= w_data_i[20];
      \nz.mem_119_sv2v_reg  <= w_data_i[19];
      \nz.mem_118_sv2v_reg  <= w_data_i[18];
      \nz.mem_117_sv2v_reg  <= w_data_i[17];
      \nz.mem_116_sv2v_reg  <= w_data_i[16];
      \nz.mem_115_sv2v_reg  <= w_data_i[15];
      \nz.mem_114_sv2v_reg  <= w_data_i[14];
      \nz.mem_113_sv2v_reg  <= w_data_i[13];
      \nz.mem_112_sv2v_reg  <= w_data_i[12];
      \nz.mem_111_sv2v_reg  <= w_data_i[11];
      \nz.mem_110_sv2v_reg  <= w_data_i[10];
      \nz.mem_109_sv2v_reg  <= w_data_i[9];
      \nz.mem_108_sv2v_reg  <= w_data_i[8];
      \nz.mem_107_sv2v_reg  <= w_data_i[7];
      \nz.mem_106_sv2v_reg  <= w_data_i[6];
      \nz.mem_105_sv2v_reg  <= w_data_i[5];
      \nz.mem_104_sv2v_reg  <= w_data_i[4];
      \nz.mem_103_sv2v_reg  <= w_data_i[3];
      \nz.mem_102_sv2v_reg  <= w_data_i[2];
      \nz.mem_101_sv2v_reg  <= w_data_i[1];
      \nz.mem_100_sv2v_reg  <= w_data_i[0];
    end 
    if(N206) begin
      \nz.mem_99_sv2v_reg  <= w_data_i[49];
      \nz.mem_98_sv2v_reg  <= w_data_i[48];
      \nz.mem_97_sv2v_reg  <= w_data_i[47];
      \nz.mem_96_sv2v_reg  <= w_data_i[46];
      \nz.mem_95_sv2v_reg  <= w_data_i[45];
      \nz.mem_94_sv2v_reg  <= w_data_i[44];
      \nz.mem_93_sv2v_reg  <= w_data_i[43];
      \nz.mem_92_sv2v_reg  <= w_data_i[42];
      \nz.mem_91_sv2v_reg  <= w_data_i[41];
      \nz.mem_90_sv2v_reg  <= w_data_i[40];
      \nz.mem_89_sv2v_reg  <= w_data_i[39];
      \nz.mem_88_sv2v_reg  <= w_data_i[38];
      \nz.mem_87_sv2v_reg  <= w_data_i[37];
      \nz.mem_86_sv2v_reg  <= w_data_i[36];
      \nz.mem_85_sv2v_reg  <= w_data_i[35];
      \nz.mem_84_sv2v_reg  <= w_data_i[34];
      \nz.mem_83_sv2v_reg  <= w_data_i[33];
      \nz.mem_82_sv2v_reg  <= w_data_i[32];
      \nz.mem_81_sv2v_reg  <= w_data_i[31];
      \nz.mem_80_sv2v_reg  <= w_data_i[30];
      \nz.mem_79_sv2v_reg  <= w_data_i[29];
      \nz.mem_78_sv2v_reg  <= w_data_i[28];
      \nz.mem_77_sv2v_reg  <= w_data_i[27];
      \nz.mem_76_sv2v_reg  <= w_data_i[26];
      \nz.mem_75_sv2v_reg  <= w_data_i[25];
      \nz.mem_74_sv2v_reg  <= w_data_i[24];
      \nz.mem_73_sv2v_reg  <= w_data_i[23];
      \nz.mem_72_sv2v_reg  <= w_data_i[22];
      \nz.mem_71_sv2v_reg  <= w_data_i[21];
      \nz.mem_70_sv2v_reg  <= w_data_i[20];
      \nz.mem_69_sv2v_reg  <= w_data_i[19];
      \nz.mem_68_sv2v_reg  <= w_data_i[18];
      \nz.mem_67_sv2v_reg  <= w_data_i[17];
      \nz.mem_66_sv2v_reg  <= w_data_i[16];
      \nz.mem_65_sv2v_reg  <= w_data_i[15];
      \nz.mem_64_sv2v_reg  <= w_data_i[14];
      \nz.mem_63_sv2v_reg  <= w_data_i[13];
      \nz.mem_62_sv2v_reg  <= w_data_i[12];
      \nz.mem_61_sv2v_reg  <= w_data_i[11];
      \nz.mem_60_sv2v_reg  <= w_data_i[10];
      \nz.mem_59_sv2v_reg  <= w_data_i[9];
      \nz.mem_58_sv2v_reg  <= w_data_i[8];
      \nz.mem_57_sv2v_reg  <= w_data_i[7];
      \nz.mem_56_sv2v_reg  <= w_data_i[6];
      \nz.mem_55_sv2v_reg  <= w_data_i[5];
      \nz.mem_54_sv2v_reg  <= w_data_i[4];
      \nz.mem_53_sv2v_reg  <= w_data_i[3];
      \nz.mem_52_sv2v_reg  <= w_data_i[2];
      \nz.mem_51_sv2v_reg  <= w_data_i[1];
      \nz.mem_50_sv2v_reg  <= w_data_i[0];
    end 
    if(N205) begin
      \nz.mem_49_sv2v_reg  <= w_data_i[49];
      \nz.mem_48_sv2v_reg  <= w_data_i[48];
      \nz.mem_47_sv2v_reg  <= w_data_i[47];
      \nz.mem_46_sv2v_reg  <= w_data_i[46];
      \nz.mem_45_sv2v_reg  <= w_data_i[45];
      \nz.mem_44_sv2v_reg  <= w_data_i[44];
      \nz.mem_43_sv2v_reg  <= w_data_i[43];
      \nz.mem_42_sv2v_reg  <= w_data_i[42];
      \nz.mem_41_sv2v_reg  <= w_data_i[41];
      \nz.mem_40_sv2v_reg  <= w_data_i[40];
      \nz.mem_39_sv2v_reg  <= w_data_i[39];
      \nz.mem_38_sv2v_reg  <= w_data_i[38];
      \nz.mem_37_sv2v_reg  <= w_data_i[37];
      \nz.mem_36_sv2v_reg  <= w_data_i[36];
      \nz.mem_35_sv2v_reg  <= w_data_i[35];
      \nz.mem_34_sv2v_reg  <= w_data_i[34];
      \nz.mem_33_sv2v_reg  <= w_data_i[33];
      \nz.mem_32_sv2v_reg  <= w_data_i[32];
      \nz.mem_31_sv2v_reg  <= w_data_i[31];
      \nz.mem_30_sv2v_reg  <= w_data_i[30];
      \nz.mem_29_sv2v_reg  <= w_data_i[29];
      \nz.mem_28_sv2v_reg  <= w_data_i[28];
      \nz.mem_27_sv2v_reg  <= w_data_i[27];
      \nz.mem_26_sv2v_reg  <= w_data_i[26];
      \nz.mem_25_sv2v_reg  <= w_data_i[25];
      \nz.mem_24_sv2v_reg  <= w_data_i[24];
      \nz.mem_23_sv2v_reg  <= w_data_i[23];
      \nz.mem_22_sv2v_reg  <= w_data_i[22];
      \nz.mem_21_sv2v_reg  <= w_data_i[21];
      \nz.mem_20_sv2v_reg  <= w_data_i[20];
      \nz.mem_19_sv2v_reg  <= w_data_i[19];
      \nz.mem_18_sv2v_reg  <= w_data_i[18];
      \nz.mem_17_sv2v_reg  <= w_data_i[17];
      \nz.mem_16_sv2v_reg  <= w_data_i[16];
      \nz.mem_15_sv2v_reg  <= w_data_i[15];
      \nz.mem_14_sv2v_reg  <= w_data_i[14];
      \nz.mem_13_sv2v_reg  <= w_data_i[13];
      \nz.mem_12_sv2v_reg  <= w_data_i[12];
      \nz.mem_11_sv2v_reg  <= w_data_i[11];
      \nz.mem_10_sv2v_reg  <= w_data_i[10];
      \nz.mem_9_sv2v_reg  <= w_data_i[9];
      \nz.mem_8_sv2v_reg  <= w_data_i[8];
      \nz.mem_7_sv2v_reg  <= w_data_i[7];
      \nz.mem_6_sv2v_reg  <= w_data_i[6];
      \nz.mem_5_sv2v_reg  <= w_data_i[5];
      \nz.mem_4_sv2v_reg  <= w_data_i[4];
      \nz.mem_3_sv2v_reg  <= w_data_i[3];
      \nz.mem_2_sv2v_reg  <= w_data_i[2];
      \nz.mem_1_sv2v_reg  <= w_data_i[1];
      \nz.mem_0_sv2v_reg  <= w_data_i[0];
    end 
  end


endmodule



module bsg_mem_1r1w_width_p50_els_p64_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [5:0] w_addr_i;
  input [49:0] w_data_i;
  input [5:0] r_addr_i;
  output [49:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [49:0] r_data_o;

  bsg_mem_1r1w_synth_width_p50_els_p64_read_write_same_addr_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_launch_sync_sync_posedge_7_unit
(
  iclk_i,
  iclk_reset_i,
  oclk_i,
  iclk_data_i,
  iclk_data_o,
  oclk_data_o
);

  input [6:0] iclk_data_i;
  output [6:0] iclk_data_o;
  output [6:0] oclk_data_o;
  input iclk_i;
  input iclk_reset_i;
  input oclk_i;
  wire [6:0] iclk_data_o,oclk_data_o,bsg_SYNC_1_r;
  reg iclk_data_o_6_sv2v_reg,iclk_data_o_5_sv2v_reg,iclk_data_o_4_sv2v_reg,
  iclk_data_o_3_sv2v_reg,iclk_data_o_2_sv2v_reg,iclk_data_o_1_sv2v_reg,
  iclk_data_o_0_sv2v_reg,bsg_SYNC_1_r_6_sv2v_reg,bsg_SYNC_1_r_5_sv2v_reg,bsg_SYNC_1_r_4_sv2v_reg,
  bsg_SYNC_1_r_3_sv2v_reg,bsg_SYNC_1_r_2_sv2v_reg,bsg_SYNC_1_r_1_sv2v_reg,
  bsg_SYNC_1_r_0_sv2v_reg,oclk_data_o_6_sv2v_reg,oclk_data_o_5_sv2v_reg,oclk_data_o_4_sv2v_reg,
  oclk_data_o_3_sv2v_reg,oclk_data_o_2_sv2v_reg,oclk_data_o_1_sv2v_reg,
  oclk_data_o_0_sv2v_reg;
  assign iclk_data_o[6] = iclk_data_o_6_sv2v_reg;
  assign iclk_data_o[5] = iclk_data_o_5_sv2v_reg;
  assign iclk_data_o[4] = iclk_data_o_4_sv2v_reg;
  assign iclk_data_o[3] = iclk_data_o_3_sv2v_reg;
  assign iclk_data_o[2] = iclk_data_o_2_sv2v_reg;
  assign iclk_data_o[1] = iclk_data_o_1_sv2v_reg;
  assign iclk_data_o[0] = iclk_data_o_0_sv2v_reg;
  assign bsg_SYNC_1_r[6] = bsg_SYNC_1_r_6_sv2v_reg;
  assign bsg_SYNC_1_r[5] = bsg_SYNC_1_r_5_sv2v_reg;
  assign bsg_SYNC_1_r[4] = bsg_SYNC_1_r_4_sv2v_reg;
  assign bsg_SYNC_1_r[3] = bsg_SYNC_1_r_3_sv2v_reg;
  assign bsg_SYNC_1_r[2] = bsg_SYNC_1_r_2_sv2v_reg;
  assign bsg_SYNC_1_r[1] = bsg_SYNC_1_r_1_sv2v_reg;
  assign bsg_SYNC_1_r[0] = bsg_SYNC_1_r_0_sv2v_reg;
  assign oclk_data_o[6] = oclk_data_o_6_sv2v_reg;
  assign oclk_data_o[5] = oclk_data_o_5_sv2v_reg;
  assign oclk_data_o[4] = oclk_data_o_4_sv2v_reg;
  assign oclk_data_o[3] = oclk_data_o_3_sv2v_reg;
  assign oclk_data_o[2] = oclk_data_o_2_sv2v_reg;
  assign oclk_data_o[1] = oclk_data_o_1_sv2v_reg;
  assign oclk_data_o[0] = oclk_data_o_0_sv2v_reg;

  always @(posedge iclk_i) begin
    if(iclk_reset_i) begin
      iclk_data_o_6_sv2v_reg <= 1'b0;
      iclk_data_o_5_sv2v_reg <= 1'b0;
      iclk_data_o_4_sv2v_reg <= 1'b0;
      iclk_data_o_3_sv2v_reg <= 1'b0;
      iclk_data_o_2_sv2v_reg <= 1'b0;
      iclk_data_o_1_sv2v_reg <= 1'b0;
      iclk_data_o_0_sv2v_reg <= 1'b0;
    end else if(1'b1) begin
      iclk_data_o_6_sv2v_reg <= iclk_data_i[6];
      iclk_data_o_5_sv2v_reg <= iclk_data_i[5];
      iclk_data_o_4_sv2v_reg <= iclk_data_i[4];
      iclk_data_o_3_sv2v_reg <= iclk_data_i[3];
      iclk_data_o_2_sv2v_reg <= iclk_data_i[2];
      iclk_data_o_1_sv2v_reg <= iclk_data_i[1];
      iclk_data_o_0_sv2v_reg <= iclk_data_i[0];
    end 
  end


  always @(posedge oclk_i) begin
    if(1'b1) begin
      bsg_SYNC_1_r_6_sv2v_reg <= iclk_data_o[6];
      bsg_SYNC_1_r_5_sv2v_reg <= iclk_data_o[5];
      bsg_SYNC_1_r_4_sv2v_reg <= iclk_data_o[4];
      bsg_SYNC_1_r_3_sv2v_reg <= iclk_data_o[3];
      bsg_SYNC_1_r_2_sv2v_reg <= iclk_data_o[2];
      bsg_SYNC_1_r_1_sv2v_reg <= iclk_data_o[1];
      bsg_SYNC_1_r_0_sv2v_reg <= iclk_data_o[0];
      oclk_data_o_6_sv2v_reg <= bsg_SYNC_1_r[6];
      oclk_data_o_5_sv2v_reg <= bsg_SYNC_1_r[5];
      oclk_data_o_4_sv2v_reg <= bsg_SYNC_1_r[4];
      oclk_data_o_3_sv2v_reg <= bsg_SYNC_1_r[3];
      oclk_data_o_2_sv2v_reg <= bsg_SYNC_1_r[2];
      oclk_data_o_1_sv2v_reg <= bsg_SYNC_1_r[1];
      oclk_data_o_0_sv2v_reg <= bsg_SYNC_1_r[0];
    end 
  end


endmodule



module bsg_launch_sync_sync_width_p7_use_negedge_for_launch_p0_use_async_reset_p0
(
  iclk_i,
  iclk_reset_i,
  oclk_i,
  iclk_data_i,
  iclk_data_o,
  oclk_data_o
);

  input [6:0] iclk_data_i;
  output [6:0] iclk_data_o;
  output [6:0] oclk_data_o;
  input iclk_i;
  input iclk_reset_i;
  input oclk_i;
  wire [6:0] iclk_data_o,oclk_data_o;

  bsg_launch_sync_sync_posedge_7_unit
  \sync.p.z.blss 
  (
    .iclk_i(iclk_i),
    .iclk_reset_i(iclk_reset_i),
    .oclk_i(oclk_i),
    .iclk_data_i(iclk_data_i),
    .iclk_data_o(iclk_data_o),
    .oclk_data_o(oclk_data_o)
  );


endmodule



module bsg_async_ptr_gray_lg_size_p7
(
  w_clk_i,
  w_reset_i,
  w_inc_i,
  r_clk_i,
  w_ptr_binary_r_o,
  w_ptr_gray_r_o,
  w_ptr_gray_r_rsync_o
);

  output [6:0] w_ptr_binary_r_o;
  output [6:0] w_ptr_gray_r_o;
  output [6:0] w_ptr_gray_r_rsync_o;
  input w_clk_i;
  input w_reset_i;
  input w_inc_i;
  input r_clk_i;
  wire [6:0] w_ptr_binary_r_o,w_ptr_gray_r_o,w_ptr_gray_r_rsync_o,w_ptr_p1_r,w_ptr_p2,
  w_ptr_gray_n;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8;
  reg w_ptr_p1_r_6_sv2v_reg,w_ptr_p1_r_5_sv2v_reg,w_ptr_p1_r_4_sv2v_reg,
  w_ptr_p1_r_3_sv2v_reg,w_ptr_p1_r_2_sv2v_reg,w_ptr_p1_r_1_sv2v_reg,w_ptr_p1_r_0_sv2v_reg,
  w_ptr_binary_r_o_6_sv2v_reg,w_ptr_binary_r_o_5_sv2v_reg,w_ptr_binary_r_o_4_sv2v_reg,
  w_ptr_binary_r_o_3_sv2v_reg,w_ptr_binary_r_o_2_sv2v_reg,
  w_ptr_binary_r_o_1_sv2v_reg,w_ptr_binary_r_o_0_sv2v_reg;
  assign w_ptr_p1_r[6] = w_ptr_p1_r_6_sv2v_reg;
  assign w_ptr_p1_r[5] = w_ptr_p1_r_5_sv2v_reg;
  assign w_ptr_p1_r[4] = w_ptr_p1_r_4_sv2v_reg;
  assign w_ptr_p1_r[3] = w_ptr_p1_r_3_sv2v_reg;
  assign w_ptr_p1_r[2] = w_ptr_p1_r_2_sv2v_reg;
  assign w_ptr_p1_r[1] = w_ptr_p1_r_1_sv2v_reg;
  assign w_ptr_p1_r[0] = w_ptr_p1_r_0_sv2v_reg;
  assign w_ptr_binary_r_o[6] = w_ptr_binary_r_o_6_sv2v_reg;
  assign w_ptr_binary_r_o[5] = w_ptr_binary_r_o_5_sv2v_reg;
  assign w_ptr_binary_r_o[4] = w_ptr_binary_r_o_4_sv2v_reg;
  assign w_ptr_binary_r_o[3] = w_ptr_binary_r_o_3_sv2v_reg;
  assign w_ptr_binary_r_o[2] = w_ptr_binary_r_o_2_sv2v_reg;
  assign w_ptr_binary_r_o[1] = w_ptr_binary_r_o_1_sv2v_reg;
  assign w_ptr_binary_r_o[0] = w_ptr_binary_r_o_0_sv2v_reg;

  bsg_launch_sync_sync_width_p7_use_negedge_for_launch_p0_use_async_reset_p0
  ptr_sync
  (
    .iclk_i(w_clk_i),
    .iclk_reset_i(w_reset_i),
    .oclk_i(r_clk_i),
    .iclk_data_i(w_ptr_gray_n),
    .iclk_data_o(w_ptr_gray_r_o),
    .oclk_data_o(w_ptr_gray_r_rsync_o)
  );

  assign w_ptr_p2 = w_ptr_p1_r + 1'b1;
  assign w_ptr_gray_n = (N0)? { w_ptr_p1_r[6:6], N3, N4, N5, N6, N7, N8 } : 
                        (N1)? w_ptr_gray_r_o : 1'b0;
  assign N0 = w_inc_i;
  assign N1 = N2;
  assign N2 = ~w_inc_i;
  assign N3 = w_ptr_p1_r[6] ^ w_ptr_p1_r[5];
  assign N4 = w_ptr_p1_r[5] ^ w_ptr_p1_r[4];
  assign N5 = w_ptr_p1_r[4] ^ w_ptr_p1_r[3];
  assign N6 = w_ptr_p1_r[3] ^ w_ptr_p1_r[2];
  assign N7 = w_ptr_p1_r[2] ^ w_ptr_p1_r[1];
  assign N8 = w_ptr_p1_r[1] ^ w_ptr_p1_r[0];

  always @(posedge w_clk_i) begin
    if(w_reset_i) begin
      w_ptr_p1_r_6_sv2v_reg <= 1'b0;
      w_ptr_p1_r_5_sv2v_reg <= 1'b0;
      w_ptr_p1_r_4_sv2v_reg <= 1'b0;
      w_ptr_p1_r_3_sv2v_reg <= 1'b0;
      w_ptr_p1_r_2_sv2v_reg <= 1'b0;
      w_ptr_p1_r_1_sv2v_reg <= 1'b0;
      w_ptr_p1_r_0_sv2v_reg <= 1'b1;
      w_ptr_binary_r_o_6_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_5_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_4_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_3_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_2_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_1_sv2v_reg <= 1'b0;
      w_ptr_binary_r_o_0_sv2v_reg <= 1'b0;
    end else if(w_inc_i) begin
      w_ptr_p1_r_6_sv2v_reg <= w_ptr_p2[6];
      w_ptr_p1_r_5_sv2v_reg <= w_ptr_p2[5];
      w_ptr_p1_r_4_sv2v_reg <= w_ptr_p2[4];
      w_ptr_p1_r_3_sv2v_reg <= w_ptr_p2[3];
      w_ptr_p1_r_2_sv2v_reg <= w_ptr_p2[2];
      w_ptr_p1_r_1_sv2v_reg <= w_ptr_p2[1];
      w_ptr_p1_r_0_sv2v_reg <= w_ptr_p2[0];
      w_ptr_binary_r_o_6_sv2v_reg <= w_ptr_p1_r[6];
      w_ptr_binary_r_o_5_sv2v_reg <= w_ptr_p1_r[5];
      w_ptr_binary_r_o_4_sv2v_reg <= w_ptr_p1_r[4];
      w_ptr_binary_r_o_3_sv2v_reg <= w_ptr_p1_r[3];
      w_ptr_binary_r_o_2_sv2v_reg <= w_ptr_p1_r[2];
      w_ptr_binary_r_o_1_sv2v_reg <= w_ptr_p1_r[1];
      w_ptr_binary_r_o_0_sv2v_reg <= w_ptr_p1_r[0];
    end 
  end


endmodule



module bsg_async_fifo_lg_size_p6_width_p50
(
  w_clk_i,
  w_reset_i,
  w_enq_i,
  w_data_i,
  w_full_o,
  r_clk_i,
  r_reset_i,
  r_deq_i,
  r_data_o,
  r_valid_o
);

  input [49:0] w_data_i;
  output [49:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_enq_i;
  input r_clk_i;
  input r_reset_i;
  input r_deq_i;
  output w_full_o;
  output r_valid_o;
  wire [49:0] r_data_o;
  wire w_full_o,r_valid_o,N0,N1;
  wire [6:0] w_ptr_binary_r,r_ptr_binary_r,w_ptr_gray_r,w_ptr_gray_r_rsync,r_ptr_gray_r,
  r_ptr_gray_r_wsync;

  bsg_mem_1r1w_width_p50_els_p64_read_write_same_addr_p0
  MSYNC_1r1w
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_enq_i),
    .w_addr_i(w_ptr_binary_r[5:0]),
    .w_data_i(w_data_i),
    .r_v_i(r_valid_o),
    .r_addr_i(r_ptr_binary_r[5:0]),
    .r_data_o(r_data_o)
  );


  bsg_async_ptr_gray_lg_size_p7
  bapg_wr
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_inc_i(w_enq_i),
    .r_clk_i(r_clk_i),
    .w_ptr_binary_r_o(w_ptr_binary_r),
    .w_ptr_gray_r_o(w_ptr_gray_r),
    .w_ptr_gray_r_rsync_o(w_ptr_gray_r_rsync)
  );


  bsg_async_ptr_gray_lg_size_p7
  bapg_rd
  (
    .w_clk_i(r_clk_i),
    .w_reset_i(r_reset_i),
    .w_inc_i(r_deq_i),
    .r_clk_i(w_clk_i),
    .w_ptr_binary_r_o(r_ptr_binary_r),
    .w_ptr_gray_r_o(r_ptr_gray_r),
    .w_ptr_gray_r_rsync_o(r_ptr_gray_r_wsync)
  );

  assign r_valid_o = r_ptr_gray_r != w_ptr_gray_r_rsync;
  assign w_full_o = w_ptr_gray_r == { N0, N1, r_ptr_gray_r_wsync[4:0] };
  assign N0 = ~r_ptr_gray_r_wsync[6];
  assign N1 = ~r_ptr_gray_r_wsync[5];

endmodule



module bsg_sync_sync_1_unit
(
  oclk_i,
  iclk_data_i,
  oclk_data_o
);

  input [0:0] iclk_data_i;
  output [0:0] oclk_data_o;
  input oclk_i;
  wire [0:0] oclk_data_o,bsg_SYNC_1_r;
  reg bsg_SYNC_1_r_0_sv2v_reg,oclk_data_o_0_sv2v_reg;
  assign bsg_SYNC_1_r[0] = bsg_SYNC_1_r_0_sv2v_reg;
  assign oclk_data_o[0] = oclk_data_o_0_sv2v_reg;

  always @(posedge oclk_i) begin
    if(1'b1) begin
      bsg_SYNC_1_r_0_sv2v_reg <= iclk_data_i[0];
      oclk_data_o_0_sv2v_reg <= bsg_SYNC_1_r[0];
    end 
  end


endmodule



module bsg_sync_sync_width_p1
(
  oclk_i,
  iclk_data_i,
  oclk_data_o
);

  input [0:0] iclk_data_i;
  output [0:0] oclk_data_o;
  input oclk_i;
  wire [0:0] oclk_data_o;

  bsg_sync_sync_1_unit
  \z.bss 
  (
    .oclk_i(oclk_i),
    .iclk_data_i(iclk_data_i[0]),
    .oclk_data_o(oclk_data_o[0])
  );


endmodule



module bsg_fsb_node_async_buffer
(
  L_clk_i,
  L_reset_i,
  L_en_o,
  L_v_o,
  L_data_o,
  L_ready_i,
  L_v_i,
  L_data_i,
  L_yumi_o,
  R_clk_i,
  R_reset_i,
  R_en_i,
  R_v_i,
  R_data_i,
  R_ready_o,
  R_v_o,
  R_data_o,
  R_yumi_i
);

  output [49:0] L_data_o;
  input [49:0] L_data_i;
  input [49:0] R_data_i;
  output [49:0] R_data_o;
  input L_clk_i;
  input L_reset_i;
  input L_ready_i;
  input L_v_i;
  input R_clk_i;
  input R_reset_i;
  input R_en_i;
  input R_v_i;
  input R_yumi_i;
  output L_en_o;
  output L_v_o;
  output L_yumi_o;
  output R_ready_o;
  output R_v_o;
  wire [49:0] L_data_o,R_data_o;
  wire L_en_o,L_v_o,L_yumi_o,R_ready_o,R_v_o,R_w_full_lo,_0_net_,_1_net_,L_w_full_lo,
  N0,N1;

  bsg_async_fifo_lg_size_p6_width_p50
  r2l_fifo
  (
    .w_clk_i(R_clk_i),
    .w_reset_i(R_reset_i),
    .w_enq_i(_0_net_),
    .w_data_i(R_data_i),
    .w_full_o(R_w_full_lo),
    .r_clk_i(L_clk_i),
    .r_reset_i(L_reset_i),
    .r_deq_i(_1_net_),
    .r_data_o(L_data_o),
    .r_valid_o(L_v_o)
  );


  bsg_async_fifo_lg_size_p6_width_p50
  l2r_fifo
  (
    .w_clk_i(L_clk_i),
    .w_reset_i(L_reset_i),
    .w_enq_i(L_yumi_o),
    .w_data_i(L_data_i),
    .w_full_o(L_w_full_lo),
    .r_clk_i(R_clk_i),
    .r_reset_i(R_reset_i),
    .r_deq_i(R_yumi_i),
    .r_data_o(R_data_o),
    .r_valid_o(R_v_o)
  );


  bsg_sync_sync_width_p1
  fsb_en_sync
  (
    .oclk_i(L_clk_i),
    .iclk_data_i(R_en_i),
    .oclk_data_o(L_en_o)
  );

  assign R_ready_o = ~R_w_full_lo;
  assign _1_net_ = L_v_o & L_ready_i;
  assign _0_net_ = N0 & R_v_i;
  assign N0 = ~R_w_full_lo;
  assign L_yumi_o = N1 & L_v_i;
  assign N1 = ~L_w_full_lo;

endmodule

